-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b87fa",
          2049 => x"f80d0b0b",
          2050 => x"0b93e904",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b93",
          2121 => x"cd040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b93b0",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b83bd",
          2210 => x"e4738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"93b50400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b0bac",
          2219 => x"cc2d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b0bab",
          2227 => x"ab2d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"96040b0b",
          2317 => x"0b8ca604",
          2318 => x"0b0b0b8c",
          2319 => x"b6040b0b",
          2320 => x"0b8cc604",
          2321 => x"0b0b0b8c",
          2322 => x"d6040b0b",
          2323 => x"0b8ce604",
          2324 => x"0b0b0b8c",
          2325 => x"f6040b0b",
          2326 => x"0b8d8604",
          2327 => x"0b0b0b8d",
          2328 => x"96040b0b",
          2329 => x"0b8da604",
          2330 => x"0b0b0b8d",
          2331 => x"b6040b0b",
          2332 => x"0b8dc604",
          2333 => x"0b0b0b8d",
          2334 => x"d7040b0b",
          2335 => x"0b8de804",
          2336 => x"0b0b0b8d",
          2337 => x"f9040b0b",
          2338 => x"0b8e8a04",
          2339 => x"0b0b0b8e",
          2340 => x"9b040b0b",
          2341 => x"0b8eac04",
          2342 => x"0b0b0b8e",
          2343 => x"bd040b0b",
          2344 => x"0b8ece04",
          2345 => x"0b0b0b8e",
          2346 => x"df040b0b",
          2347 => x"0b8ef004",
          2348 => x"0b0b0b8f",
          2349 => x"81040b0b",
          2350 => x"0b8f9204",
          2351 => x"0b0b0b8f",
          2352 => x"a3040b0b",
          2353 => x"0b8fb404",
          2354 => x"0b0b0b8f",
          2355 => x"c5040b0b",
          2356 => x"0b8fd604",
          2357 => x"0b0b0b8f",
          2358 => x"e7040b0b",
          2359 => x"0b8ff804",
          2360 => x"0b0b0b90",
          2361 => x"89040b0b",
          2362 => x"0b909a04",
          2363 => x"0b0b0b90",
          2364 => x"ab040b0b",
          2365 => x"0b90bc04",
          2366 => x"0b0b0b90",
          2367 => x"cd040b0b",
          2368 => x"0b90de04",
          2369 => x"0b0b0b90",
          2370 => x"ef040b0b",
          2371 => x"0b918004",
          2372 => x"0b0b0b91",
          2373 => x"91040b0b",
          2374 => x"0b91a204",
          2375 => x"0b0b0b91",
          2376 => x"b3040b0b",
          2377 => x"0b91c404",
          2378 => x"0b0b0b91",
          2379 => x"d5040b0b",
          2380 => x"0b91e604",
          2381 => x"0b0b0b91",
          2382 => x"f7040b0b",
          2383 => x"0b928804",
          2384 => x"0b0b0b92",
          2385 => x"99040b0b",
          2386 => x"0b92aa04",
          2387 => x"0b0b0b92",
          2388 => x"bb040b0b",
          2389 => x"0b92cb04",
          2390 => x"0b0b0b92",
          2391 => x"dc040b0b",
          2392 => x"0b92ed04",
          2393 => x"0b0b0b92",
          2394 => x"fe04ffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0484b8f0",
          2434 => x"0c80d5ec",
          2435 => x"2d84b8f0",
          2436 => x"0880c080",
          2437 => x"900484b8",
          2438 => x"f00ca2ee",
          2439 => x"2d84b8f0",
          2440 => x"0880c080",
          2441 => x"900484b8",
          2442 => x"f00ca0f3",
          2443 => x"2d84b8f0",
          2444 => x"0880c080",
          2445 => x"900484b8",
          2446 => x"f00ca0e0",
          2447 => x"2d84b8f0",
          2448 => x"0880c080",
          2449 => x"900484b8",
          2450 => x"f00c94a3",
          2451 => x"2d84b8f0",
          2452 => x"0880c080",
          2453 => x"900484b8",
          2454 => x"f00ca1f6",
          2455 => x"2d84b8f0",
          2456 => x"0880c080",
          2457 => x"900484b8",
          2458 => x"f00caf86",
          2459 => x"2d84b8f0",
          2460 => x"0880c080",
          2461 => x"900484b8",
          2462 => x"f00cad82",
          2463 => x"2d84b8f0",
          2464 => x"0880c080",
          2465 => x"900484b8",
          2466 => x"f00c9488",
          2467 => x"2d84b8f0",
          2468 => x"0880c080",
          2469 => x"900484b8",
          2470 => x"f00c95a8",
          2471 => x"2d84b8f0",
          2472 => x"0880c080",
          2473 => x"900484b8",
          2474 => x"f00c95d1",
          2475 => x"2d84b8f0",
          2476 => x"0880c080",
          2477 => x"900484b8",
          2478 => x"f00cb18a",
          2479 => x"2d84b8f0",
          2480 => x"0880c080",
          2481 => x"900484b8",
          2482 => x"f00c80d4",
          2483 => x"d12d84b8",
          2484 => x"f00880c0",
          2485 => x"80900484",
          2486 => x"b8f00c80",
          2487 => x"d5b62d84",
          2488 => x"b8f00880",
          2489 => x"c0809004",
          2490 => x"84b8f00c",
          2491 => x"80d28d2d",
          2492 => x"84b8f008",
          2493 => x"80c08090",
          2494 => x"0484b8f0",
          2495 => x"0c80d3c0",
          2496 => x"2d84b8f0",
          2497 => x"0880c080",
          2498 => x"900484b8",
          2499 => x"f00c82c9",
          2500 => x"9d2d84b8",
          2501 => x"f00880c0",
          2502 => x"80900484",
          2503 => x"b8f00c82",
          2504 => x"e2ef2d84",
          2505 => x"b8f00880",
          2506 => x"c0809004",
          2507 => x"84b8f00c",
          2508 => x"82d28d2d",
          2509 => x"84b8f008",
          2510 => x"80c08090",
          2511 => x"0484b8f0",
          2512 => x"0c82d7af",
          2513 => x"2d84b8f0",
          2514 => x"0880c080",
          2515 => x"900484b8",
          2516 => x"f00c82ed",
          2517 => x"8c2d84b8",
          2518 => x"f00880c0",
          2519 => x"80900484",
          2520 => x"b8f00c82",
          2521 => x"fa942d84",
          2522 => x"b8f00880",
          2523 => x"c0809004",
          2524 => x"84b8f00c",
          2525 => x"82def62d",
          2526 => x"84b8f008",
          2527 => x"80c08090",
          2528 => x"0484b8f0",
          2529 => x"0c82f1ad",
          2530 => x"2d84b8f0",
          2531 => x"0880c080",
          2532 => x"900484b8",
          2533 => x"f00c82f2",
          2534 => x"fa2d84b8",
          2535 => x"f00880c0",
          2536 => x"80900484",
          2537 => x"b8f00c82",
          2538 => x"f3cf2d84",
          2539 => x"b8f00880",
          2540 => x"c0809004",
          2541 => x"84b8f00c",
          2542 => x"8384912d",
          2543 => x"84b8f008",
          2544 => x"80c08090",
          2545 => x"0484b8f0",
          2546 => x"0c82fed6",
          2547 => x"2d84b8f0",
          2548 => x"0880c080",
          2549 => x"900484b8",
          2550 => x"f00c838a",
          2551 => x"f52d84b8",
          2552 => x"f00880c0",
          2553 => x"80900484",
          2554 => x"b8f00c82",
          2555 => x"f5ac2d84",
          2556 => x"b8f00880",
          2557 => x"c0809004",
          2558 => x"84b8f00c",
          2559 => x"8393ec2d",
          2560 => x"84b8f008",
          2561 => x"80c08090",
          2562 => x"0484b8f0",
          2563 => x"0c8394f7",
          2564 => x"2d84b8f0",
          2565 => x"0880c080",
          2566 => x"900484b8",
          2567 => x"f00c82e5",
          2568 => x"bf2d84b8",
          2569 => x"f00880c0",
          2570 => x"80900484",
          2571 => x"b8f00c82",
          2572 => x"e3d62d84",
          2573 => x"b8f00880",
          2574 => x"c0809004",
          2575 => x"84b8f00c",
          2576 => x"82e6fd2d",
          2577 => x"84b8f008",
          2578 => x"80c08090",
          2579 => x"0484b8f0",
          2580 => x"0c82f696",
          2581 => x"2d84b8f0",
          2582 => x"0880c080",
          2583 => x"900484b8",
          2584 => x"f00c8396",
          2585 => x"892d84b8",
          2586 => x"f00880c0",
          2587 => x"80900484",
          2588 => x"b8f00c83",
          2589 => x"99e62d84",
          2590 => x"b8f00880",
          2591 => x"c0809004",
          2592 => x"84b8f00c",
          2593 => x"83a0d82d",
          2594 => x"84b8f008",
          2595 => x"80c08090",
          2596 => x"0484b8f0",
          2597 => x"0c82c6ee",
          2598 => x"2d84b8f0",
          2599 => x"0880c080",
          2600 => x"900484b8",
          2601 => x"f00c83a4",
          2602 => x"812d84b8",
          2603 => x"f00880c0",
          2604 => x"80900484",
          2605 => x"b8f00c83",
          2606 => x"b9822d84",
          2607 => x"b8f00880",
          2608 => x"c0809004",
          2609 => x"84b8f00c",
          2610 => x"83b7b42d",
          2611 => x"84b8f008",
          2612 => x"80c08090",
          2613 => x"0484b8f0",
          2614 => x"0c81f3d2",
          2615 => x"2d84b8f0",
          2616 => x"0880c080",
          2617 => x"900484b8",
          2618 => x"f00c81f4",
          2619 => x"d12d84b8",
          2620 => x"f00880c0",
          2621 => x"80900484",
          2622 => x"b8f00c81",
          2623 => x"f5d02d84",
          2624 => x"b8f00880",
          2625 => x"c0809004",
          2626 => x"84b8f00c",
          2627 => x"80d08f2d",
          2628 => x"84b8f008",
          2629 => x"80c08090",
          2630 => x"0484b8f0",
          2631 => x"0c80d1df",
          2632 => x"2d84b8f0",
          2633 => x"0880c080",
          2634 => x"900484b8",
          2635 => x"f00c80d7",
          2636 => x"8a2d84b8",
          2637 => x"f00880c0",
          2638 => x"80900484",
          2639 => x"b8f00cb1",
          2640 => x"9a2d84b8",
          2641 => x"f00880c0",
          2642 => x"80900484",
          2643 => x"b8f00c81",
          2644 => x"daf02d84",
          2645 => x"b8f00880",
          2646 => x"c0809004",
          2647 => x"84b8f00c",
          2648 => x"81dcab2d",
          2649 => x"84b8f008",
          2650 => x"80c08090",
          2651 => x"0484b8f0",
          2652 => x"0c81f1ac",
          2653 => x"2d84b8f0",
          2654 => x"0880c080",
          2655 => x"900484b8",
          2656 => x"f00c81d5",
          2657 => x"802d84b8",
          2658 => x"f00880c0",
          2659 => x"8090043c",
          2660 => x"04101010",
          2661 => x"10101010",
          2662 => x"10101010",
          2663 => x"10101010",
          2664 => x"10101010",
          2665 => x"10101010",
          2666 => x"10101010",
          2667 => x"10101010",
          2668 => x"53510400",
          2669 => x"007381ff",
          2670 => x"06738306",
          2671 => x"09810583",
          2672 => x"05101010",
          2673 => x"2b0772fc",
          2674 => x"060c5151",
          2675 => x"04727280",
          2676 => x"728106ff",
          2677 => x"05097206",
          2678 => x"05711052",
          2679 => x"720a100a",
          2680 => x"5372ed38",
          2681 => x"51515351",
          2682 => x"0484b8e4",
          2683 => x"7084d4d0",
          2684 => x"278e3880",
          2685 => x"71708405",
          2686 => x"530c0b0b",
          2687 => x"0b93ec04",
          2688 => x"8c815180",
          2689 => x"ceba0400",
          2690 => x"fc3d0d87",
          2691 => x"3d707084",
          2692 => x"05520856",
          2693 => x"53745284",
          2694 => x"d4c80851",
          2695 => x"81c53f86",
          2696 => x"3d0d04fa",
          2697 => x"3d0d787a",
          2698 => x"7c851133",
          2699 => x"81328106",
          2700 => x"80732507",
          2701 => x"56585557",
          2702 => x"80527272",
          2703 => x"2e098106",
          2704 => x"80d338ff",
          2705 => x"1477748a",
          2706 => x"32703070",
          2707 => x"72079f2a",
          2708 => x"51555556",
          2709 => x"54807425",
          2710 => x"b7387180",
          2711 => x"2eb23875",
          2712 => x"518efa3f",
          2713 => x"84b8e408",
          2714 => x"5384b8e4",
          2715 => x"08ff2eae",
          2716 => x"3884b8e4",
          2717 => x"08757081",
          2718 => x"055734ff",
          2719 => x"14738a32",
          2720 => x"70307072",
          2721 => x"079f2a51",
          2722 => x"54545473",
          2723 => x"8024cb38",
          2724 => x"80753476",
          2725 => x"527184b8",
          2726 => x"e40c883d",
          2727 => x"0d04800b",
          2728 => x"84b8e40c",
          2729 => x"883d0d04",
          2730 => x"f53d0d7d",
          2731 => x"54860284",
          2732 => x"05990534",
          2733 => x"7356fe0a",
          2734 => x"588e3d88",
          2735 => x"05537e52",
          2736 => x"8d3de405",
          2737 => x"519d3f73",
          2738 => x"19548074",
          2739 => x"348d3d0d",
          2740 => x"04fd3d0d",
          2741 => x"863d8805",
          2742 => x"53765275",
          2743 => x"51853f85",
          2744 => x"3d0d04f1",
          2745 => x"3d0d6163",
          2746 => x"65425d5d",
          2747 => x"80708c1f",
          2748 => x"0c851e33",
          2749 => x"70812a81",
          2750 => x"32810655",
          2751 => x"555bff54",
          2752 => x"727b2e09",
          2753 => x"810680d2",
          2754 => x"387b3357",
          2755 => x"767b2e80",
          2756 => x"c538811c",
          2757 => x"7b810654",
          2758 => x"5c72802e",
          2759 => x"818138d0",
          2760 => x"175f7e89",
          2761 => x"2681a338",
          2762 => x"76b03270",
          2763 => x"30708025",
          2764 => x"51545578",
          2765 => x"ae387280",
          2766 => x"2ea9387a",
          2767 => x"832a7081",
          2768 => x"32810640",
          2769 => x"547e802e",
          2770 => x"9e387a82",
          2771 => x"80075b7b",
          2772 => x"335776ff",
          2773 => x"bd388c1d",
          2774 => x"08547384",
          2775 => x"b8e40c91",
          2776 => x"3d0d047a",
          2777 => x"832a5478",
          2778 => x"10101079",
          2779 => x"10057098",
          2780 => x"2b70982c",
          2781 => x"19708180",
          2782 => x"0a298b0a",
          2783 => x"0570982c",
          2784 => x"525a5b56",
          2785 => x"5f807924",
          2786 => x"81863873",
          2787 => x"81065372",
          2788 => x"ffbd3878",
          2789 => x"7c335858",
          2790 => x"76fef738",
          2791 => x"ffb83976",
          2792 => x"a52e0981",
          2793 => x"06933881",
          2794 => x"73745a5a",
          2795 => x"5b8a7c33",
          2796 => x"585a76fe",
          2797 => x"dd38ff9e",
          2798 => x"397c5276",
          2799 => x"518baf3f",
          2800 => x"7b335776",
          2801 => x"fecc38ff",
          2802 => x"8d397a83",
          2803 => x"2a708106",
          2804 => x"5455788a",
          2805 => x"38817074",
          2806 => x"0640547e",
          2807 => x"9538e017",
          2808 => x"537280d8",
          2809 => x"26973872",
          2810 => x"101083c9",
          2811 => x"f4055473",
          2812 => x"080473e0",
          2813 => x"18545980",
          2814 => x"d87327eb",
          2815 => x"387c5276",
          2816 => x"518aeb3f",
          2817 => x"807c3358",
          2818 => x"5b76fe86",
          2819 => x"38fec739",
          2820 => x"80ff59fe",
          2821 => x"f639885a",
          2822 => x"7f608405",
          2823 => x"71087d83",
          2824 => x"ffcf065e",
          2825 => x"58415484",
          2826 => x"b8f45e79",
          2827 => x"52755193",
          2828 => x"9a3f84b8",
          2829 => x"e40881ff",
          2830 => x"0684b8e4",
          2831 => x"0818df05",
          2832 => x"56537289",
          2833 => x"26883884",
          2834 => x"b8e408b0",
          2835 => x"0555747e",
          2836 => x"70810540",
          2837 => x"34795275",
          2838 => x"5190ca3f",
          2839 => x"84b8e408",
          2840 => x"5684b8e4",
          2841 => x"08c5387d",
          2842 => x"84b8f431",
          2843 => x"982b7bb2",
          2844 => x"0640567e",
          2845 => x"802e8f38",
          2846 => x"77848080",
          2847 => x"29fc8080",
          2848 => x"0570902c",
          2849 => x"59557a86",
          2850 => x"2a708106",
          2851 => x"555f7380",
          2852 => x"2e9e3877",
          2853 => x"84808029",
          2854 => x"f8808005",
          2855 => x"5379902e",
          2856 => x"8b387784",
          2857 => x"808029fc",
          2858 => x"80800553",
          2859 => x"72902c58",
          2860 => x"7a832a70",
          2861 => x"81065455",
          2862 => x"72802e9e",
          2863 => x"3875982c",
          2864 => x"7081ff06",
          2865 => x"54547873",
          2866 => x"2486cc38",
          2867 => x"7a83fff7",
          2868 => x"0670832a",
          2869 => x"71862a41",
          2870 => x"565b7481",
          2871 => x"06547380",
          2872 => x"2e85f038",
          2873 => x"77793190",
          2874 => x"2b70902c",
          2875 => x"7c838006",
          2876 => x"56595373",
          2877 => x"802e8596",
          2878 => x"387a812a",
          2879 => x"81065473",
          2880 => x"85eb387a",
          2881 => x"842a8106",
          2882 => x"54738698",
          2883 => x"387a852a",
          2884 => x"81065473",
          2885 => x"8697387e",
          2886 => x"81065473",
          2887 => x"858f387a",
          2888 => x"882a8106",
          2889 => x"5f7e802e",
          2890 => x"b2387778",
          2891 => x"84808029",
          2892 => x"fc808005",
          2893 => x"70902c5a",
          2894 => x"40548074",
          2895 => x"259d387c",
          2896 => x"52b05188",
          2897 => x"a93f7778",
          2898 => x"84808029",
          2899 => x"fc808005",
          2900 => x"70902c5a",
          2901 => x"40547380",
          2902 => x"24e53874",
          2903 => x"81065372",
          2904 => x"802eb238",
          2905 => x"78798180",
          2906 => x"0a2981ff",
          2907 => x"0a057098",
          2908 => x"2c5b5555",
          2909 => x"8075259d",
          2910 => x"387c52b0",
          2911 => x"5187ef3f",
          2912 => x"78798180",
          2913 => x"0a2981ff",
          2914 => x"0a057098",
          2915 => x"2c5b5555",
          2916 => x"748024e5",
          2917 => x"387a872a",
          2918 => x"7081065c",
          2919 => x"557a802e",
          2920 => x"81b93876",
          2921 => x"80e32e84",
          2922 => x"d8387680",
          2923 => x"f32e81ca",
          2924 => x"387680d3",
          2925 => x"2e81e238",
          2926 => x"7d84b8f4",
          2927 => x"2e96387c",
          2928 => x"52ff1e70",
          2929 => x"33525e87",
          2930 => x"a53f7d84",
          2931 => x"b8f42e09",
          2932 => x"8106ec38",
          2933 => x"7481065b",
          2934 => x"7a802efc",
          2935 => x"a7387778",
          2936 => x"84808029",
          2937 => x"fc808005",
          2938 => x"70902c5a",
          2939 => x"40558075",
          2940 => x"25fc9138",
          2941 => x"7c52a051",
          2942 => x"86f43fe2",
          2943 => x"397a9007",
          2944 => x"5b7aa007",
          2945 => x"7c33585b",
          2946 => x"76fa8738",
          2947 => x"fac8397a",
          2948 => x"80c0075b",
          2949 => x"80f85790",
          2950 => x"60618405",
          2951 => x"71087e83",
          2952 => x"ffcf065f",
          2953 => x"5942555a",
          2954 => x"fbfd397f",
          2955 => x"60840577",
          2956 => x"fe800a06",
          2957 => x"83133370",
          2958 => x"982b7207",
          2959 => x"7c848080",
          2960 => x"29fc8080",
          2961 => x"0570902c",
          2962 => x"5e525a56",
          2963 => x"57415f7a",
          2964 => x"872a7081",
          2965 => x"065c557a",
          2966 => x"fec93877",
          2967 => x"78848080",
          2968 => x"29fc8080",
          2969 => x"0570902c",
          2970 => x"5a545f80",
          2971 => x"7f25feb3",
          2972 => x"387c52a0",
          2973 => x"5185f73f",
          2974 => x"e239ff1a",
          2975 => x"7083ffff",
          2976 => x"065b5779",
          2977 => x"83ffff2e",
          2978 => x"feca387c",
          2979 => x"52757081",
          2980 => x"05573351",
          2981 => x"85d83fe2",
          2982 => x"39ff1a70",
          2983 => x"83ffff06",
          2984 => x"5b547983",
          2985 => x"ffff2efe",
          2986 => x"ab387c52",
          2987 => x"75708105",
          2988 => x"57335185",
          2989 => x"b93fe239",
          2990 => x"75fc0a06",
          2991 => x"81fc0a07",
          2992 => x"78848080",
          2993 => x"29fc8080",
          2994 => x"0570902c",
          2995 => x"5a585680",
          2996 => x"e37b872a",
          2997 => x"7081065d",
          2998 => x"56577afd",
          2999 => x"c638fefb",
          3000 => x"397f6084",
          3001 => x"05710870",
          3002 => x"53404156",
          3003 => x"807e2482",
          3004 => x"df387a83",
          3005 => x"ffbf065b",
          3006 => x"84b8f45e",
          3007 => x"faad397a",
          3008 => x"84077c33",
          3009 => x"585b76f8",
          3010 => x"8938f8ca",
          3011 => x"397a8807",
          3012 => x"5b807c33",
          3013 => x"585976f7",
          3014 => x"f938f8ba",
          3015 => x"397f6084",
          3016 => x"05710877",
          3017 => x"81065658",
          3018 => x"415f7282",
          3019 => x"8a387551",
          3020 => x"87f63f84",
          3021 => x"b8e40883",
          3022 => x"ffff0678",
          3023 => x"7131902b",
          3024 => x"545a7290",
          3025 => x"2c58fe87",
          3026 => x"397a80c0",
          3027 => x"077c3358",
          3028 => x"5b76f7be",
          3029 => x"38f7ff39",
          3030 => x"7f608405",
          3031 => x"71087781",
          3032 => x"065d5841",
          3033 => x"547981cf",
          3034 => x"38755187",
          3035 => x"bb3f84b8",
          3036 => x"e40883ff",
          3037 => x"ff067871",
          3038 => x"31902b54",
          3039 => x"5ac4397a",
          3040 => x"8180077c",
          3041 => x"33585b76",
          3042 => x"f78838f7",
          3043 => x"c9397778",
          3044 => x"84808029",
          3045 => x"fc808005",
          3046 => x"70902c5a",
          3047 => x"54548074",
          3048 => x"25fad638",
          3049 => x"7c52a051",
          3050 => x"83c43fe2",
          3051 => x"397c52b0",
          3052 => x"5183bb3f",
          3053 => x"79902e09",
          3054 => x"8106fae3",
          3055 => x"387c5276",
          3056 => x"5183ab3f",
          3057 => x"7a882a81",
          3058 => x"065f7e80",
          3059 => x"2efb8c38",
          3060 => x"fad83975",
          3061 => x"982c7871",
          3062 => x"31902b70",
          3063 => x"902c7d83",
          3064 => x"8006575a",
          3065 => x"515373fa",
          3066 => x"9038ffa2",
          3067 => x"397c52ad",
          3068 => x"5182fb3f",
          3069 => x"7e810654",
          3070 => x"73802efa",
          3071 => x"a238ffad",
          3072 => x"397c5275",
          3073 => x"982a5182",
          3074 => x"e53f7481",
          3075 => x"065b7a80",
          3076 => x"2ef7f138",
          3077 => x"fbc83978",
          3078 => x"7431982b",
          3079 => x"70982c5a",
          3080 => x"53f9b739",
          3081 => x"7c52ab51",
          3082 => x"82c43fc8",
          3083 => x"397c52a0",
          3084 => x"5182bb3f",
          3085 => x"ffbe3978",
          3086 => x"52755188",
          3087 => x"8b3f84b8",
          3088 => x"e40883ff",
          3089 => x"ff067871",
          3090 => x"31902b54",
          3091 => x"5afdf339",
          3092 => x"7a82077e",
          3093 => x"307183ff",
          3094 => x"bf065257",
          3095 => x"5bfd9939",
          3096 => x"fe3d0d84",
          3097 => x"d4c40853",
          3098 => x"75527451",
          3099 => x"f3b53f84",
          3100 => x"3d0d04fa",
          3101 => x"3d0d7855",
          3102 => x"800b84d4",
          3103 => x"c8088511",
          3104 => x"3370812a",
          3105 => x"81327081",
          3106 => x"06515658",
          3107 => x"5557ff56",
          3108 => x"72772e09",
          3109 => x"810680d5",
          3110 => x"38747081",
          3111 => x"05563353",
          3112 => x"72772eb0",
          3113 => x"3884d4c8",
          3114 => x"08527251",
          3115 => x"90140853",
          3116 => x"722d84b8",
          3117 => x"e408802e",
          3118 => x"8338ff57",
          3119 => x"74708105",
          3120 => x"56335372",
          3121 => x"802e8838",
          3122 => x"84d4c808",
          3123 => x"54d73984",
          3124 => x"d4c80854",
          3125 => x"84d4c808",
          3126 => x"528a5190",
          3127 => x"14085574",
          3128 => x"2d84b8e4",
          3129 => x"08802e83",
          3130 => x"38ff5776",
          3131 => x"567584b8",
          3132 => x"e40c883d",
          3133 => x"0d04fa3d",
          3134 => x"0d787a56",
          3135 => x"54800b85",
          3136 => x"16337081",
          3137 => x"2a813270",
          3138 => x"81065155",
          3139 => x"5757ff56",
          3140 => x"72772e09",
          3141 => x"81069238",
          3142 => x"73708105",
          3143 => x"55335372",
          3144 => x"772e0981",
          3145 => x"06983876",
          3146 => x"567584b8",
          3147 => x"e40c883d",
          3148 => x"0d047370",
          3149 => x"81055533",
          3150 => x"5372802e",
          3151 => x"ea387452",
          3152 => x"72519015",
          3153 => x"0853722d",
          3154 => x"84b8e408",
          3155 => x"802ee338",
          3156 => x"ff747081",
          3157 => x"05563354",
          3158 => x"5772e338",
          3159 => x"ca39ff3d",
          3160 => x"0d84d4c8",
          3161 => x"08527351",
          3162 => x"853f833d",
          3163 => x"0d04fa3d",
          3164 => x"0d787a85",
          3165 => x"11337081",
          3166 => x"2a813281",
          3167 => x"06565656",
          3168 => x"57ff5672",
          3169 => x"ae387382",
          3170 => x"2a810654",
          3171 => x"73802eac",
          3172 => x"388c1508",
          3173 => x"53728816",
          3174 => x"08259138",
          3175 => x"74085676",
          3176 => x"76347408",
          3177 => x"8105750c",
          3178 => x"8c150853",
          3179 => x"81138c16",
          3180 => x"0c765675",
          3181 => x"84b8e40c",
          3182 => x"883d0d04",
          3183 => x"74527681",
          3184 => x"ff065190",
          3185 => x"15085473",
          3186 => x"2dff5684",
          3187 => x"b8e408e3",
          3188 => x"388c1508",
          3189 => x"81058c16",
          3190 => x"0c7656d7",
          3191 => x"39fb3d0d",
          3192 => x"77851133",
          3193 => x"7081ff06",
          3194 => x"70813281",
          3195 => x"06555556",
          3196 => x"56ff5471",
          3197 => x"b3387286",
          3198 => x"2a810652",
          3199 => x"71b33872",
          3200 => x"822a8106",
          3201 => x"5271802e",
          3202 => x"80c33875",
          3203 => x"08703353",
          3204 => x"5371802e",
          3205 => x"80f03881",
          3206 => x"13760c8c",
          3207 => x"16088105",
          3208 => x"8c170c71",
          3209 => x"81ff0654",
          3210 => x"7384b8e4",
          3211 => x"0c873d0d",
          3212 => x"0474ffbf",
          3213 => x"06537285",
          3214 => x"17348c16",
          3215 => x"0881058c",
          3216 => x"170c8416",
          3217 => x"3384b8e4",
          3218 => x"0c873d0d",
          3219 => x"04755194",
          3220 => x"16085574",
          3221 => x"2d84b8e4",
          3222 => x"085284b8",
          3223 => x"e4088025",
          3224 => x"ffb93885",
          3225 => x"16337090",
          3226 => x"07545284",
          3227 => x"b8e408ff",
          3228 => x"2e853871",
          3229 => x"a0075372",
          3230 => x"851734ff",
          3231 => x"547384b8",
          3232 => x"e40c873d",
          3233 => x"0d0474a0",
          3234 => x"07537285",
          3235 => x"1734ff54",
          3236 => x"ec39fd3d",
          3237 => x"0d757771",
          3238 => x"54545471",
          3239 => x"70810553",
          3240 => x"335170f7",
          3241 => x"38ff1252",
          3242 => x"72708105",
          3243 => x"54335170",
          3244 => x"72708105",
          3245 => x"543470f0",
          3246 => x"387384b8",
          3247 => x"e40c853d",
          3248 => x"0d04fc3d",
          3249 => x"0d767971",
          3250 => x"7a555552",
          3251 => x"5470802e",
          3252 => x"9d387372",
          3253 => x"27a13870",
          3254 => x"802e9338",
          3255 => x"71708105",
          3256 => x"53337370",
          3257 => x"81055534",
          3258 => x"ff115170",
          3259 => x"ef387384",
          3260 => x"b8e40c86",
          3261 => x"3d0d0470",
          3262 => x"12557375",
          3263 => x"27d93870",
          3264 => x"14755353",
          3265 => x"ff13ff13",
          3266 => x"53537133",
          3267 => x"7334ff11",
          3268 => x"5170802e",
          3269 => x"d938ff13",
          3270 => x"ff135353",
          3271 => x"71337334",
          3272 => x"ff115170",
          3273 => x"df38c739",
          3274 => x"fe3d0d74",
          3275 => x"70535371",
          3276 => x"70810553",
          3277 => x"335170f7",
          3278 => x"38ff1270",
          3279 => x"743184b8",
          3280 => x"e40c5184",
          3281 => x"3d0d04fd",
          3282 => x"3d0d7577",
          3283 => x"71545454",
          3284 => x"72708105",
          3285 => x"54335170",
          3286 => x"72708105",
          3287 => x"543470f0",
          3288 => x"387384b8",
          3289 => x"e40c853d",
          3290 => x"0d04fd3d",
          3291 => x"0d757871",
          3292 => x"79555552",
          3293 => x"5470802e",
          3294 => x"93387170",
          3295 => x"81055333",
          3296 => x"73708105",
          3297 => x"5534ff11",
          3298 => x"5170ef38",
          3299 => x"7384b8e4",
          3300 => x"0c853d0d",
          3301 => x"04fc3d0d",
          3302 => x"76787a55",
          3303 => x"56547280",
          3304 => x"2ea13873",
          3305 => x"33757081",
          3306 => x"05573352",
          3307 => x"5271712e",
          3308 => x"0981069a",
          3309 => x"38811454",
          3310 => x"71802eb7",
          3311 => x"38ff1353",
          3312 => x"72e13880",
          3313 => x"517084b8",
          3314 => x"e40c863d",
          3315 => x"0d047280",
          3316 => x"2ef13873",
          3317 => x"3353ff51",
          3318 => x"72802ee9",
          3319 => x"38ff1533",
          3320 => x"52815171",
          3321 => x"802ede38",
          3322 => x"72723184",
          3323 => x"b8e40c86",
          3324 => x"3d0d0471",
          3325 => x"84b8e40c",
          3326 => x"863d0d04",
          3327 => x"fb3d0d77",
          3328 => x"79537052",
          3329 => x"5680c13f",
          3330 => x"84b8e408",
          3331 => x"84b8e408",
          3332 => x"81055255",
          3333 => x"81b2d93f",
          3334 => x"84b8e408",
          3335 => x"5484b8e4",
          3336 => x"08802e9b",
          3337 => x"3884b8e4",
          3338 => x"08155480",
          3339 => x"74347453",
          3340 => x"755284b8",
          3341 => x"e40851fe",
          3342 => x"b13f84b8",
          3343 => x"e4085473",
          3344 => x"84b8e40c",
          3345 => x"873d0d04",
          3346 => x"fd3d0d75",
          3347 => x"77717154",
          3348 => x"55535471",
          3349 => x"802e9f38",
          3350 => x"72708105",
          3351 => x"54335170",
          3352 => x"802e8c38",
          3353 => x"ff125271",
          3354 => x"ff2e0981",
          3355 => x"06ea38ff",
          3356 => x"13707531",
          3357 => x"52527084",
          3358 => x"b8e40c85",
          3359 => x"3d0d04fd",
          3360 => x"3d0d7577",
          3361 => x"79725553",
          3362 => x"54547080",
          3363 => x"2e8e3872",
          3364 => x"72708105",
          3365 => x"5434ff11",
          3366 => x"5170f438",
          3367 => x"7384b8e4",
          3368 => x"0c853d0d",
          3369 => x"04fa3d0d",
          3370 => x"787a5854",
          3371 => x"a0527680",
          3372 => x"2e8b3876",
          3373 => x"5180f53f",
          3374 => x"84b8e408",
          3375 => x"52e01253",
          3376 => x"73802e8d",
          3377 => x"38735180",
          3378 => x"e33f7184",
          3379 => x"b8e40831",
          3380 => x"53805272",
          3381 => x"9f2680cb",
          3382 => x"38735272",
          3383 => x"9f2e80c3",
          3384 => x"38811374",
          3385 => x"712aa072",
          3386 => x"3176712b",
          3387 => x"57545455",
          3388 => x"80567476",
          3389 => x"2ea83872",
          3390 => x"10749f2a",
          3391 => x"07741077",
          3392 => x"07787231",
          3393 => x"ff119f2c",
          3394 => x"7081067b",
          3395 => x"72067571",
          3396 => x"31ff1c5c",
          3397 => x"56525255",
          3398 => x"58555374",
          3399 => x"da387310",
          3400 => x"76075271",
          3401 => x"84b8e40c",
          3402 => x"883d0d04",
          3403 => x"fc3d0d76",
          3404 => x"70fc8080",
          3405 => x"06703070",
          3406 => x"72078025",
          3407 => x"70842b90",
          3408 => x"71317571",
          3409 => x"2a7083fe",
          3410 => x"80067030",
          3411 => x"70802583",
          3412 => x"2b887131",
          3413 => x"74712a70",
          3414 => x"81f00670",
          3415 => x"30708025",
          3416 => x"822b8471",
          3417 => x"3174712a",
          3418 => x"5553751b",
          3419 => x"05738c06",
          3420 => x"70307080",
          3421 => x"25108271",
          3422 => x"3177712a",
          3423 => x"70812a81",
          3424 => x"32708106",
          3425 => x"70308274",
          3426 => x"31067519",
          3427 => x"0584b8e4",
          3428 => x"0c515254",
          3429 => x"55515456",
          3430 => x"5a535555",
          3431 => x"55515656",
          3432 => x"56565158",
          3433 => x"56545286",
          3434 => x"3d0d04fd",
          3435 => x"3d0d7577",
          3436 => x"70547153",
          3437 => x"54548194",
          3438 => x"3f84b8e4",
          3439 => x"08732974",
          3440 => x"713184b8",
          3441 => x"e40c5385",
          3442 => x"3d0d04fa",
          3443 => x"3d0d787a",
          3444 => x"5854a053",
          3445 => x"76802e8b",
          3446 => x"387651fe",
          3447 => x"cf3f84b8",
          3448 => x"e40853e0",
          3449 => x"13527380",
          3450 => x"2e8d3873",
          3451 => x"51febd3f",
          3452 => x"7284b8e4",
          3453 => x"08315273",
          3454 => x"53719f26",
          3455 => x"80c53880",
          3456 => x"53719f2e",
          3457 => x"be388112",
          3458 => x"74712aa0",
          3459 => x"72317671",
          3460 => x"2b575454",
          3461 => x"55805674",
          3462 => x"762ea838",
          3463 => x"7210749f",
          3464 => x"2a077410",
          3465 => x"77077872",
          3466 => x"31ff119f",
          3467 => x"2c708106",
          3468 => x"7b720675",
          3469 => x"7131ff1c",
          3470 => x"5c565252",
          3471 => x"55585553",
          3472 => x"74da3872",
          3473 => x"84b8e40c",
          3474 => x"883d0d04",
          3475 => x"fa3d0d78",
          3476 => x"9f2c7a9f",
          3477 => x"2c7a9f2c",
          3478 => x"7b327c9f",
          3479 => x"2c7d3273",
          3480 => x"73327174",
          3481 => x"31577275",
          3482 => x"31565956",
          3483 => x"595556fc",
          3484 => x"b43f84b8",
          3485 => x"e4087532",
          3486 => x"753184b8",
          3487 => x"e40c883d",
          3488 => x"0d04f73d",
          3489 => x"0d7b7d5b",
          3490 => x"5780707b",
          3491 => x"0c770870",
          3492 => x"33565659",
          3493 => x"73a02e09",
          3494 => x"81068f38",
          3495 => x"81157078",
          3496 => x"0c703355",
          3497 => x"5573a02e",
          3498 => x"f33873ad",
          3499 => x"2e80f538",
          3500 => x"73b02e81",
          3501 => x"8338d014",
          3502 => x"58805677",
          3503 => x"892680db",
          3504 => x"388a5880",
          3505 => x"56a07427",
          3506 => x"80c43880",
          3507 => x"e0742789",
          3508 => x"38e01470",
          3509 => x"81ff0655",
          3510 => x"53d01470",
          3511 => x"81ff0651",
          3512 => x"53907327",
          3513 => x"8f38f913",
          3514 => x"7081ff06",
          3515 => x"54548973",
          3516 => x"27818938",
          3517 => x"72782781",
          3518 => x"83387776",
          3519 => x"29138116",
          3520 => x"70790c70",
          3521 => x"33565656",
          3522 => x"73a026ff",
          3523 => x"be387880",
          3524 => x"2e843875",
          3525 => x"3056757a",
          3526 => x"0c815675",
          3527 => x"84b8e40c",
          3528 => x"8b3d0d04",
          3529 => x"81701670",
          3530 => x"790c7033",
          3531 => x"56565973",
          3532 => x"b02e0981",
          3533 => x"06feff38",
          3534 => x"81157078",
          3535 => x"0c703355",
          3536 => x"557380e2",
          3537 => x"2ea63890",
          3538 => x"587380f8",
          3539 => x"2ea03881",
          3540 => x"56a07427",
          3541 => x"c638d014",
          3542 => x"53805688",
          3543 => x"58897327",
          3544 => x"fee13875",
          3545 => x"84b8e40c",
          3546 => x"8b3d0d04",
          3547 => x"82588115",
          3548 => x"70780c70",
          3549 => x"33555580",
          3550 => x"56feca39",
          3551 => x"800b84b8",
          3552 => x"e40c8b3d",
          3553 => x"0d04f73d",
          3554 => x"0d7b7d5b",
          3555 => x"5780707b",
          3556 => x"0c770870",
          3557 => x"33565659",
          3558 => x"73a02e09",
          3559 => x"81068f38",
          3560 => x"81157078",
          3561 => x"0c703355",
          3562 => x"5573a02e",
          3563 => x"f33873ad",
          3564 => x"2e80f538",
          3565 => x"73b02e81",
          3566 => x"8338d014",
          3567 => x"58805677",
          3568 => x"892680db",
          3569 => x"388a5880",
          3570 => x"56a07427",
          3571 => x"80c43880",
          3572 => x"e0742789",
          3573 => x"38e01470",
          3574 => x"81ff0655",
          3575 => x"53d01470",
          3576 => x"81ff0651",
          3577 => x"53907327",
          3578 => x"8f38f913",
          3579 => x"7081ff06",
          3580 => x"54548973",
          3581 => x"27818938",
          3582 => x"72782781",
          3583 => x"83387776",
          3584 => x"29138116",
          3585 => x"70790c70",
          3586 => x"33565656",
          3587 => x"73a026ff",
          3588 => x"be387880",
          3589 => x"2e843875",
          3590 => x"3056757a",
          3591 => x"0c815675",
          3592 => x"84b8e40c",
          3593 => x"8b3d0d04",
          3594 => x"81701670",
          3595 => x"790c7033",
          3596 => x"56565973",
          3597 => x"b02e0981",
          3598 => x"06feff38",
          3599 => x"81157078",
          3600 => x"0c703355",
          3601 => x"557380e2",
          3602 => x"2ea63890",
          3603 => x"587380f8",
          3604 => x"2ea03881",
          3605 => x"56a07427",
          3606 => x"c638d014",
          3607 => x"53805688",
          3608 => x"58897327",
          3609 => x"fee13875",
          3610 => x"84b8e40c",
          3611 => x"8b3d0d04",
          3612 => x"82588115",
          3613 => x"70780c70",
          3614 => x"33555580",
          3615 => x"56feca39",
          3616 => x"800b84b8",
          3617 => x"e40c8b3d",
          3618 => x"0d0480d6",
          3619 => x"d13f84b8",
          3620 => x"e40881ff",
          3621 => x"0684b8e4",
          3622 => x"0c04ff3d",
          3623 => x"0d735271",
          3624 => x"93268c38",
          3625 => x"71101083",
          3626 => x"bdf40552",
          3627 => x"71080483",
          3628 => x"ce8c51ef",
          3629 => x"be3f833d",
          3630 => x"0d0483ce",
          3631 => x"9c51efb3",
          3632 => x"3f833d0d",
          3633 => x"0483ceb4",
          3634 => x"51efa83f",
          3635 => x"833d0d04",
          3636 => x"83cecc51",
          3637 => x"ef9d3f83",
          3638 => x"3d0d0483",
          3639 => x"cee451ef",
          3640 => x"923f833d",
          3641 => x"0d0483ce",
          3642 => x"f451ef87",
          3643 => x"3f833d0d",
          3644 => x"0483cf94",
          3645 => x"51eefc3f",
          3646 => x"833d0d04",
          3647 => x"83cfa451",
          3648 => x"eef13f83",
          3649 => x"3d0d0483",
          3650 => x"cfcc51ee",
          3651 => x"e63f833d",
          3652 => x"0d0483cf",
          3653 => x"e051eedb",
          3654 => x"3f833d0d",
          3655 => x"0483cffc",
          3656 => x"51eed03f",
          3657 => x"833d0d04",
          3658 => x"83d09451",
          3659 => x"eec53f83",
          3660 => x"3d0d0483",
          3661 => x"d0ac51ee",
          3662 => x"ba3f833d",
          3663 => x"0d0483d0",
          3664 => x"c451eeaf",
          3665 => x"3f833d0d",
          3666 => x"0483d0d4",
          3667 => x"51eea43f",
          3668 => x"833d0d04",
          3669 => x"83d0e851",
          3670 => x"ee993f83",
          3671 => x"3d0d0483",
          3672 => x"d0f851ee",
          3673 => x"8e3f833d",
          3674 => x"0d0483d1",
          3675 => x"8851ee83",
          3676 => x"3f833d0d",
          3677 => x"0483d198",
          3678 => x"51edf83f",
          3679 => x"833d0d04",
          3680 => x"83d1a851",
          3681 => x"eded3f83",
          3682 => x"3d0d0483",
          3683 => x"d1b451ed",
          3684 => x"e23f833d",
          3685 => x"0d04ec3d",
          3686 => x"0d660284",
          3687 => x"0580e305",
          3688 => x"335b5880",
          3689 => x"68793070",
          3690 => x"7b077325",
          3691 => x"51575759",
          3692 => x"78577587",
          3693 => x"ff268338",
          3694 => x"81577477",
          3695 => x"077081ff",
          3696 => x"06515593",
          3697 => x"577480e2",
          3698 => x"38815377",
          3699 => x"528c3d70",
          3700 => x"52588295",
          3701 => x"c83f84b8",
          3702 => x"e4085784",
          3703 => x"b8e40880",
          3704 => x"2e80d038",
          3705 => x"775182af",
          3706 => x"863f7630",
          3707 => x"70780780",
          3708 => x"257b3070",
          3709 => x"9f2a7206",
          3710 => x"53575758",
          3711 => x"77802eaa",
          3712 => x"3887c098",
          3713 => x"88085574",
          3714 => x"87e72680",
          3715 => x"e0387452",
          3716 => x"7887e829",
          3717 => x"51f58e3f",
          3718 => x"84b8e408",
          3719 => x"5483d1e4",
          3720 => x"53785283",
          3721 => x"d1c051df",
          3722 => x"df3f7684",
          3723 => x"b8e40c96",
          3724 => x"3d0d0484",
          3725 => x"b8e40887",
          3726 => x"c098880c",
          3727 => x"84b8e408",
          3728 => x"59963dd4",
          3729 => x"05548480",
          3730 => x"53755277",
          3731 => x"51829dbd",
          3732 => x"3f84b8e4",
          3733 => x"085784b8",
          3734 => x"e408ff88",
          3735 => x"387a5574",
          3736 => x"802eff80",
          3737 => x"38741975",
          3738 => x"175759d5",
          3739 => x"3987e852",
          3740 => x"7451f4b1",
          3741 => x"3f84b8e4",
          3742 => x"08527851",
          3743 => x"f4a73f84",
          3744 => x"b8e40854",
          3745 => x"83d1e453",
          3746 => x"785283d1",
          3747 => x"c051def8",
          3748 => x"3fff9739",
          3749 => x"f83d0d7c",
          3750 => x"028405b7",
          3751 => x"05335859",
          3752 => x"ff588053",
          3753 => x"7b527a51",
          3754 => x"fdec3f84",
          3755 => x"b8e4088b",
          3756 => x"3876802e",
          3757 => x"91387681",
          3758 => x"2e8a3877",
          3759 => x"84b8e40c",
          3760 => x"8a3d0d04",
          3761 => x"780484d4",
          3762 => x"c4566155",
          3763 => x"605484b8",
          3764 => x"e4537f52",
          3765 => x"7e51782d",
          3766 => x"84b8e408",
          3767 => x"84b8e40c",
          3768 => x"8a3d0d04",
          3769 => x"f33d0d7f",
          3770 => x"6163028c",
          3771 => x"0580cf05",
          3772 => x"33737315",
          3773 => x"68415f5c",
          3774 => x"5c5f5d5e",
          3775 => x"78802e83",
          3776 => x"82387a52",
          3777 => x"83d1ec51",
          3778 => x"ddfe3f83",
          3779 => x"d1f451dd",
          3780 => x"f73f8054",
          3781 => x"737927b2",
          3782 => x"387c902e",
          3783 => x"81ed387c",
          3784 => x"a02e82a8",
          3785 => x"38731853",
          3786 => x"727a2781",
          3787 => x"a7387233",
          3788 => x"5283d1f8",
          3789 => x"51ddd13f",
          3790 => x"811484d4",
          3791 => x"c8085354",
          3792 => x"a051ecaa",
          3793 => x"3f787426",
          3794 => x"dc3883d2",
          3795 => x"8051ddb8",
          3796 => x"3f805675",
          3797 => x"792780c0",
          3798 => x"38751870",
          3799 => x"33555380",
          3800 => x"55727a27",
          3801 => x"83388155",
          3802 => x"80539f74",
          3803 => x"27833881",
          3804 => x"53747306",
          3805 => x"7081ff06",
          3806 => x"56577480",
          3807 => x"2e883880",
          3808 => x"fe742781",
          3809 => x"ee3884d4",
          3810 => x"c80852a0",
          3811 => x"51ebdf3f",
          3812 => x"81165678",
          3813 => x"7626c238",
          3814 => x"83d28451",
          3815 => x"e9d53f78",
          3816 => x"18791c5c",
          3817 => x"5880519d",
          3818 => x"a83f84b8",
          3819 => x"e408982b",
          3820 => x"70982c58",
          3821 => x"5476a02e",
          3822 => x"81ee3876",
          3823 => x"9b2e82c3",
          3824 => x"387b1e57",
          3825 => x"767826fe",
          3826 => x"b938ff0b",
          3827 => x"84b8e40c",
          3828 => x"8f3d0d04",
          3829 => x"83d28851",
          3830 => x"dcae3f81",
          3831 => x"1484d4c8",
          3832 => x"085354a0",
          3833 => x"51eb873f",
          3834 => x"787426fe",
          3835 => x"b838feda",
          3836 => x"3983d298",
          3837 => x"51dc913f",
          3838 => x"821484d4",
          3839 => x"c8085354",
          3840 => x"a051eaea",
          3841 => x"3f737927",
          3842 => x"fec03873",
          3843 => x"1853727a",
          3844 => x"27df3872",
          3845 => x"225283d2",
          3846 => x"8c51dbec",
          3847 => x"3f821484",
          3848 => x"d4c80853",
          3849 => x"54a051ea",
          3850 => x"c53f7874",
          3851 => x"26dd38fe",
          3852 => x"993983d2",
          3853 => x"9451dbd0",
          3854 => x"3f841484",
          3855 => x"d4c80853",
          3856 => x"54a051ea",
          3857 => x"a93f7379",
          3858 => x"27fdff38",
          3859 => x"73185372",
          3860 => x"7a27df38",
          3861 => x"72085283",
          3862 => x"d1ec51db",
          3863 => x"ab3f8414",
          3864 => x"84d4c808",
          3865 => x"5354a051",
          3866 => x"ea843f78",
          3867 => x"7426dd38",
          3868 => x"fdd83984",
          3869 => x"d4c80852",
          3870 => x"7351e9f2",
          3871 => x"3f811656",
          3872 => x"fe913980",
          3873 => x"ced83f84",
          3874 => x"b8e40881",
          3875 => x"ff065388",
          3876 => x"5972a82e",
          3877 => x"fcec38a0",
          3878 => x"597280d0",
          3879 => x"2e098106",
          3880 => x"fce03890",
          3881 => x"59fcdb39",
          3882 => x"80519ba5",
          3883 => x"3f84b8e4",
          3884 => x"08982b70",
          3885 => x"982c70a0",
          3886 => x"32703072",
          3887 => x"9b327030",
          3888 => x"70720773",
          3889 => x"75070651",
          3890 => x"55585957",
          3891 => x"58537280",
          3892 => x"25fde838",
          3893 => x"80519af9",
          3894 => x"3f84b8e4",
          3895 => x"08982b70",
          3896 => x"982c70a0",
          3897 => x"32703072",
          3898 => x"9b327030",
          3899 => x"70720773",
          3900 => x"75070651",
          3901 => x"55585957",
          3902 => x"58538073",
          3903 => x"24ffa938",
          3904 => x"fdb93980",
          3905 => x"0b84b8e4",
          3906 => x"0c8f3d0d",
          3907 => x"04fe3d0d",
          3908 => x"87c09680",
          3909 => x"0853aac7",
          3910 => x"3f81519c",
          3911 => x"ed3f83d2",
          3912 => x"dc519cfe",
          3913 => x"3f80519c",
          3914 => x"e13f7281",
          3915 => x"2a708106",
          3916 => x"51527182",
          3917 => x"b7387282",
          3918 => x"2a708106",
          3919 => x"51527182",
          3920 => x"89387283",
          3921 => x"2a708106",
          3922 => x"51527181",
          3923 => x"db387284",
          3924 => x"2a708106",
          3925 => x"51527181",
          3926 => x"ad387285",
          3927 => x"2a708106",
          3928 => x"51527180",
          3929 => x"ff387286",
          3930 => x"2a708106",
          3931 => x"51527180",
          3932 => x"d2387287",
          3933 => x"2a708106",
          3934 => x"515271a9",
          3935 => x"3872882a",
          3936 => x"81065372",
          3937 => x"8838a9df",
          3938 => x"3f843d0d",
          3939 => x"0481519b",
          3940 => x"f93f83d2",
          3941 => x"f4519c8a",
          3942 => x"3f80519b",
          3943 => x"ed3fa9c7",
          3944 => x"3f843d0d",
          3945 => x"0481519b",
          3946 => x"e13f83d3",
          3947 => x"88519bf2",
          3948 => x"3f80519b",
          3949 => x"d53f7288",
          3950 => x"2a810653",
          3951 => x"72802ec6",
          3952 => x"38cb3981",
          3953 => x"519bc33f",
          3954 => x"83d39c51",
          3955 => x"9bd43f80",
          3956 => x"519bb73f",
          3957 => x"72872a70",
          3958 => x"81065152",
          3959 => x"71802eff",
          3960 => x"9c38c239",
          3961 => x"81519ba2",
          3962 => x"3f83d3b0",
          3963 => x"519bb33f",
          3964 => x"80519b96",
          3965 => x"3f72862a",
          3966 => x"70810651",
          3967 => x"5271802e",
          3968 => x"fef038ff",
          3969 => x"be398151",
          3970 => x"9b803f83",
          3971 => x"d3c4519b",
          3972 => x"913f8051",
          3973 => x"9af43f72",
          3974 => x"852a7081",
          3975 => x"06515271",
          3976 => x"802efec2",
          3977 => x"38ffbd39",
          3978 => x"81519ade",
          3979 => x"3f83d3d8",
          3980 => x"519aef3f",
          3981 => x"80519ad2",
          3982 => x"3f72842a",
          3983 => x"70810651",
          3984 => x"5271802e",
          3985 => x"fe9438ff",
          3986 => x"bd398151",
          3987 => x"9abc3f83",
          3988 => x"d3ec519a",
          3989 => x"cd3f8051",
          3990 => x"9ab03f72",
          3991 => x"832a7081",
          3992 => x"06515271",
          3993 => x"802efde6",
          3994 => x"38ffbd39",
          3995 => x"81519a9a",
          3996 => x"3f83d3fc",
          3997 => x"519aab3f",
          3998 => x"80519a8e",
          3999 => x"3f72822a",
          4000 => x"70810651",
          4001 => x"5271802e",
          4002 => x"fdb838ff",
          4003 => x"bd39ca3d",
          4004 => x"0d807041",
          4005 => x"41ff6184",
          4006 => x"cff00c42",
          4007 => x"81526051",
          4008 => x"81b5fb3f",
          4009 => x"84b8e408",
          4010 => x"81ff069b",
          4011 => x"3d405978",
          4012 => x"612e84b1",
          4013 => x"3883d4d0",
          4014 => x"51e3b83f",
          4015 => x"983d4383",
          4016 => x"d58851d6",
          4017 => x"c33f7e48",
          4018 => x"80f85380",
          4019 => x"527e51eb",
          4020 => x"ae3f0b0b",
          4021 => x"83edd833",
          4022 => x"7081ff06",
          4023 => x"5b597980",
          4024 => x"2e82f138",
          4025 => x"79812e83",
          4026 => x"88387881",
          4027 => x"ff065e7d",
          4028 => x"822e83c1",
          4029 => x"3867705a",
          4030 => x"5a79802e",
          4031 => x"83dc3879",
          4032 => x"335c7ba0",
          4033 => x"2e098106",
          4034 => x"8c38811a",
          4035 => x"70335d5a",
          4036 => x"7ba02ef6",
          4037 => x"38805c7b",
          4038 => x"9b26be38",
          4039 => x"7b902983",
          4040 => x"eddc0570",
          4041 => x"08525be7",
          4042 => x"ff3f84b8",
          4043 => x"e40884b8",
          4044 => x"e408547a",
          4045 => x"537b0852",
          4046 => x"5de8da3f",
          4047 => x"84b8e408",
          4048 => x"8b38841b",
          4049 => x"335e7d81",
          4050 => x"2e838038",
          4051 => x"811c7081",
          4052 => x"ff065d5b",
          4053 => x"9b7c27c4",
          4054 => x"389a3d33",
          4055 => x"5c7b802e",
          4056 => x"fedd3880",
          4057 => x"f8527e51",
          4058 => x"e9923f84",
          4059 => x"b8e4085e",
          4060 => x"84b8e408",
          4061 => x"802e8dc9",
          4062 => x"3884b8e4",
          4063 => x"0848b83d",
          4064 => x"ff800551",
          4065 => x"91893f84",
          4066 => x"b8e40860",
          4067 => x"62065c5c",
          4068 => x"7a802e81",
          4069 => x"843884b8",
          4070 => x"e40851e7",
          4071 => x"8b3f84b8",
          4072 => x"e4088f26",
          4073 => x"80f33881",
          4074 => x"0ba53d5e",
          4075 => x"5b7a822e",
          4076 => x"8d85387a",
          4077 => x"82248ce2",
          4078 => x"387a812e",
          4079 => x"82e4387b",
          4080 => x"54805383",
          4081 => x"d58c527c",
          4082 => x"51d5dd3f",
          4083 => x"83f1a058",
          4084 => x"84b99457",
          4085 => x"7d566755",
          4086 => x"80549080",
          4087 => x"0a539080",
          4088 => x"0a527c51",
          4089 => x"f5ae3f84",
          4090 => x"b8e40884",
          4091 => x"b8e40809",
          4092 => x"70307072",
          4093 => x"07802551",
          4094 => x"5b5b4280",
          4095 => x"5a7a8326",
          4096 => x"8338815a",
          4097 => x"787a0659",
          4098 => x"78802e8d",
          4099 => x"38811b70",
          4100 => x"81ff065c",
          4101 => x"5a7aff95",
          4102 => x"387f8132",
          4103 => x"61813207",
          4104 => x"5d7c81ee",
          4105 => x"3861ff2e",
          4106 => x"81e8387d",
          4107 => x"518194d0",
          4108 => x"3f83d588",
          4109 => x"51d3d13f",
          4110 => x"7e4880f8",
          4111 => x"5380527e",
          4112 => x"51e8bc3f",
          4113 => x"0b0b83ed",
          4114 => x"d8337081",
          4115 => x"ff065b59",
          4116 => x"79fd9138",
          4117 => x"815383d4",
          4118 => x"b45284cf",
          4119 => x"f4518288",
          4120 => x"bc3f84b8",
          4121 => x"e40880c5",
          4122 => x"38810b0b",
          4123 => x"0b83edd8",
          4124 => x"3484cff4",
          4125 => x"5380f852",
          4126 => x"7e5182f6",
          4127 => x"b73f84b8",
          4128 => x"e408802e",
          4129 => x"a03884b8",
          4130 => x"e40851df",
          4131 => x"e63f0b0b",
          4132 => x"83edd833",
          4133 => x"7081ff06",
          4134 => x"5f597d82",
          4135 => x"2e098106",
          4136 => x"fcd33891",
          4137 => x"3984cff4",
          4138 => x"5182a1c3",
          4139 => x"3f820b0b",
          4140 => x"0b83edd8",
          4141 => x"3483d4c4",
          4142 => x"5380f852",
          4143 => x"7e51a7c3",
          4144 => x"3f67705a",
          4145 => x"5a79fcb7",
          4146 => x"3890397c",
          4147 => x"1a630c85",
          4148 => x"1b335978",
          4149 => x"818926fd",
          4150 => x"80387810",
          4151 => x"1083bec4",
          4152 => x"055a7908",
          4153 => x"04835383",
          4154 => x"d594527e",
          4155 => x"51e4fb3f",
          4156 => x"60537e52",
          4157 => x"84ba9051",
          4158 => x"8284f33f",
          4159 => x"84b8e408",
          4160 => x"612e0981",
          4161 => x"06fbae38",
          4162 => x"81709a3d",
          4163 => x"454141fb",
          4164 => x"ae3983d5",
          4165 => x"9851dedb",
          4166 => x"3f7d5181",
          4167 => x"92e23ffe",
          4168 => x"903983d5",
          4169 => x"a8567b55",
          4170 => x"83d5ac54",
          4171 => x"805383d5",
          4172 => x"b0527c51",
          4173 => x"d2f23ffd",
          4174 => x"9339818c",
          4175 => x"9a3ffaff",
          4176 => x"399add3f",
          4177 => x"faf93981",
          4178 => x"528351bf",
          4179 => x"933ffaef",
          4180 => x"39818dc5",
          4181 => x"3ffae839",
          4182 => x"83d5c051",
          4183 => x"de953f80",
          4184 => x"59780483",
          4185 => x"d5d451de",
          4186 => x"8a3fd0fd",
          4187 => x"3ffad039",
          4188 => x"b83dff84",
          4189 => x"1153ff80",
          4190 => x"0551ec8a",
          4191 => x"3f84b8e4",
          4192 => x"08802efa",
          4193 => x"ba386852",
          4194 => x"83d5f051",
          4195 => x"d0fa3f68",
          4196 => x"5a792d84",
          4197 => x"b8e40880",
          4198 => x"2efaa438",
          4199 => x"84b8e408",
          4200 => x"5283d68c",
          4201 => x"51d0e13f",
          4202 => x"fa9539b8",
          4203 => x"3dff8411",
          4204 => x"53ff8005",
          4205 => x"51ebcf3f",
          4206 => x"84b8e408",
          4207 => x"802ef9ff",
          4208 => x"38685283",
          4209 => x"d6a851d0",
          4210 => x"bf3f6859",
          4211 => x"7804b83d",
          4212 => x"fef41153",
          4213 => x"ff800551",
          4214 => x"e9a83f84",
          4215 => x"b8e40880",
          4216 => x"2ef9dc38",
          4217 => x"b83dfef0",
          4218 => x"1153ff80",
          4219 => x"0551e992",
          4220 => x"3f84b8e4",
          4221 => x"0886d038",
          4222 => x"64597808",
          4223 => x"53785283",
          4224 => x"d6c451d0",
          4225 => x"833f84d4",
          4226 => x"c4085380",
          4227 => x"f8527e51",
          4228 => x"d0913f7e",
          4229 => x"487e3359",
          4230 => x"78ae2ef9",
          4231 => x"a238789f",
          4232 => x"2687d338",
          4233 => x"64840570",
          4234 => x"4659cf39",
          4235 => x"b83dfef4",
          4236 => x"1153ff80",
          4237 => x"0551e8ca",
          4238 => x"3f84b8e4",
          4239 => x"08802ef8",
          4240 => x"fe38b83d",
          4241 => x"fef01153",
          4242 => x"ff800551",
          4243 => x"e8b43f84",
          4244 => x"b8e40886",
          4245 => x"b0386459",
          4246 => x"78225378",
          4247 => x"5283d6d4",
          4248 => x"51cfa53f",
          4249 => x"84d4c408",
          4250 => x"5380f852",
          4251 => x"7e51cfb3",
          4252 => x"3f7e487e",
          4253 => x"335978ae",
          4254 => x"2ef8c438",
          4255 => x"789f2687",
          4256 => x"ca386482",
          4257 => x"05704659",
          4258 => x"cf39b83d",
          4259 => x"ff841153",
          4260 => x"ff800551",
          4261 => x"e9f03f84",
          4262 => x"b8e40880",
          4263 => x"2ef8a038",
          4264 => x"b83dfefc",
          4265 => x"1153ff80",
          4266 => x"0551e9da",
          4267 => x"3f84b8e4",
          4268 => x"08802ef8",
          4269 => x"8a38b83d",
          4270 => x"fef81153",
          4271 => x"ff800551",
          4272 => x"e9c43f84",
          4273 => x"b8e40880",
          4274 => x"2ef7f438",
          4275 => x"83d6e051",
          4276 => x"ceb63f68",
          4277 => x"675d5978",
          4278 => x"7c27838d",
          4279 => x"38657033",
          4280 => x"7a335f5c",
          4281 => x"5a7a7d2e",
          4282 => x"95387a55",
          4283 => x"79547833",
          4284 => x"53785283",
          4285 => x"d6f051ce",
          4286 => x"8f3f6666",
          4287 => x"5b5c8119",
          4288 => x"811b4759",
          4289 => x"d239b83d",
          4290 => x"ff841153",
          4291 => x"ff800551",
          4292 => x"e8f43f84",
          4293 => x"b8e40880",
          4294 => x"2ef7a438",
          4295 => x"b83dfefc",
          4296 => x"1153ff80",
          4297 => x"0551e8de",
          4298 => x"3f84b8e4",
          4299 => x"08802ef7",
          4300 => x"8e38b83d",
          4301 => x"fef81153",
          4302 => x"ff800551",
          4303 => x"e8c83f84",
          4304 => x"b8e40880",
          4305 => x"2ef6f838",
          4306 => x"83d78c51",
          4307 => x"cdba3f68",
          4308 => x"5a796727",
          4309 => x"82933865",
          4310 => x"5c797081",
          4311 => x"055b337c",
          4312 => x"34658105",
          4313 => x"46eb39b8",
          4314 => x"3dff8411",
          4315 => x"53ff8005",
          4316 => x"51e8933f",
          4317 => x"84b8e408",
          4318 => x"802ef6c3",
          4319 => x"38b83dfe",
          4320 => x"fc1153ff",
          4321 => x"800551e7",
          4322 => x"fd3f84b8",
          4323 => x"e408b138",
          4324 => x"68703354",
          4325 => x"5283d798",
          4326 => x"51cced3f",
          4327 => x"84d4c408",
          4328 => x"5380f852",
          4329 => x"7e51ccfb",
          4330 => x"3f7e487e",
          4331 => x"335978ae",
          4332 => x"2ef68c38",
          4333 => x"789f2684",
          4334 => x"97386881",
          4335 => x"0549d139",
          4336 => x"68590280",
          4337 => x"db053379",
          4338 => x"34688105",
          4339 => x"49b83dfe",
          4340 => x"fc1153ff",
          4341 => x"800551e7",
          4342 => x"ad3f84b8",
          4343 => x"e408802e",
          4344 => x"f5dd3868",
          4345 => x"590280db",
          4346 => x"05337934",
          4347 => x"68810549",
          4348 => x"b83dfefc",
          4349 => x"1153ff80",
          4350 => x"0551e78a",
          4351 => x"3f84b8e4",
          4352 => x"08ffbd38",
          4353 => x"f5b939b8",
          4354 => x"3dff8411",
          4355 => x"53ff8005",
          4356 => x"51e6f33f",
          4357 => x"84b8e408",
          4358 => x"802ef5a3",
          4359 => x"38b83dfe",
          4360 => x"fc1153ff",
          4361 => x"800551e6",
          4362 => x"dd3f84b8",
          4363 => x"e408802e",
          4364 => x"f58d38b8",
          4365 => x"3dfef811",
          4366 => x"53ff8005",
          4367 => x"51e6c73f",
          4368 => x"84b8e408",
          4369 => x"863884b8",
          4370 => x"e4084683",
          4371 => x"d7a451cb",
          4372 => x"b73f6867",
          4373 => x"5b59787a",
          4374 => x"278f3865",
          4375 => x"5b7a7970",
          4376 => x"84055b0c",
          4377 => x"797926f5",
          4378 => x"388a51d9",
          4379 => x"f13ff4cf",
          4380 => x"39b83dff",
          4381 => x"80055187",
          4382 => x"963f84b8",
          4383 => x"e408b93d",
          4384 => x"ff800552",
          4385 => x"5988d83f",
          4386 => x"815384b8",
          4387 => x"e4085278",
          4388 => x"51ea833f",
          4389 => x"84b8e408",
          4390 => x"802ef4a3",
          4391 => x"3884b8e4",
          4392 => x"0851e7f6",
          4393 => x"3ff49839",
          4394 => x"b83dff84",
          4395 => x"1153ff80",
          4396 => x"0551e5d2",
          4397 => x"3f84b8e4",
          4398 => x"08913883",
          4399 => x"f1e8335a",
          4400 => x"79802e83",
          4401 => x"c03883f1",
          4402 => x"a00849b8",
          4403 => x"3dfefc11",
          4404 => x"53ff8005",
          4405 => x"51e5af3f",
          4406 => x"84b8e408",
          4407 => x"913883f1",
          4408 => x"e8335a79",
          4409 => x"802e838a",
          4410 => x"3883f1a4",
          4411 => x"0847b83d",
          4412 => x"fef81153",
          4413 => x"ff800551",
          4414 => x"e58c3f84",
          4415 => x"b8e40880",
          4416 => x"2ea53880",
          4417 => x"665c5c7a",
          4418 => x"882e8338",
          4419 => x"815c7a90",
          4420 => x"32703070",
          4421 => x"72079f2a",
          4422 => x"7e065c5f",
          4423 => x"5d79802e",
          4424 => x"88387aa0",
          4425 => x"2e833888",
          4426 => x"4683d7b4",
          4427 => x"51d6c43f",
          4428 => x"80556854",
          4429 => x"65536652",
          4430 => x"6851eba8",
          4431 => x"3f83d7c0",
          4432 => x"51d6b03f",
          4433 => x"f2f93964",
          4434 => x"64710c59",
          4435 => x"64840545",
          4436 => x"b83dfef0",
          4437 => x"1153ff80",
          4438 => x"0551e2a6",
          4439 => x"3f84b8e4",
          4440 => x"08802ef2",
          4441 => x"da386464",
          4442 => x"710c5964",
          4443 => x"840545b8",
          4444 => x"3dfef011",
          4445 => x"53ff8005",
          4446 => x"51e2873f",
          4447 => x"84b8e408",
          4448 => x"c638f2bb",
          4449 => x"39645e02",
          4450 => x"80ce0522",
          4451 => x"7e708205",
          4452 => x"40237d45",
          4453 => x"b83dfef0",
          4454 => x"1153ff80",
          4455 => x"0551e1e2",
          4456 => x"3f84b8e4",
          4457 => x"08802ef2",
          4458 => x"9638645e",
          4459 => x"0280ce05",
          4460 => x"227e7082",
          4461 => x"0540237d",
          4462 => x"45b83dfe",
          4463 => x"f01153ff",
          4464 => x"800551e1",
          4465 => x"bd3f84b8",
          4466 => x"e408ffb9",
          4467 => x"38f1f039",
          4468 => x"b83dfefc",
          4469 => x"1153ff80",
          4470 => x"0551e3aa",
          4471 => x"3f84b8e4",
          4472 => x"08802e81",
          4473 => x"dc38685c",
          4474 => x"0280db05",
          4475 => x"337c3468",
          4476 => x"810549fb",
          4477 => x"9b39b83d",
          4478 => x"fef01153",
          4479 => x"ff800551",
          4480 => x"e1803f84",
          4481 => x"b8e40880",
          4482 => x"2e819838",
          4483 => x"6464710c",
          4484 => x"5d648405",
          4485 => x"704659f7",
          4486 => x"e1397a83",
          4487 => x"2e098106",
          4488 => x"f39d387b",
          4489 => x"5583d5ac",
          4490 => x"54805383",
          4491 => x"d7cc527c",
          4492 => x"51c8f53f",
          4493 => x"f396397b",
          4494 => x"527c51da",
          4495 => x"8a3ff38c",
          4496 => x"3983d7d8",
          4497 => x"51d4ac3f",
          4498 => x"f0f539b8",
          4499 => x"3dfef011",
          4500 => x"53ff8005",
          4501 => x"51e0ab3f",
          4502 => x"84b8e408",
          4503 => x"802eb838",
          4504 => x"64590280",
          4505 => x"ce052279",
          4506 => x"7082055b",
          4507 => x"237845f7",
          4508 => x"e73983f1",
          4509 => x"e9335c7b",
          4510 => x"802e80cf",
          4511 => x"3883f1ac",
          4512 => x"0847fcea",
          4513 => x"3983f1e9",
          4514 => x"335c7b80",
          4515 => x"2ea13883",
          4516 => x"f1a80849",
          4517 => x"fcb53983",
          4518 => x"d88451d3",
          4519 => x"d63f6459",
          4520 => x"f7b63983",
          4521 => x"d88451d3",
          4522 => x"ca3f6459",
          4523 => x"f6cc3983",
          4524 => x"f1ea3359",
          4525 => x"78802ea5",
          4526 => x"3883f1b0",
          4527 => x"0849fc8b",
          4528 => x"3983d884",
          4529 => x"51d3ac3f",
          4530 => x"f9c63983",
          4531 => x"f1ea3359",
          4532 => x"78802e9b",
          4533 => x"3883f1b4",
          4534 => x"0847fc92",
          4535 => x"3983f1eb",
          4536 => x"335e7d80",
          4537 => x"2e9b3883",
          4538 => x"f1b80849",
          4539 => x"fbdd3983",
          4540 => x"f1eb335e",
          4541 => x"7d802e9b",
          4542 => x"3883f1bc",
          4543 => x"0847fbee",
          4544 => x"3983f1e6",
          4545 => x"335d7c80",
          4546 => x"2e9b3883",
          4547 => x"f1c00849",
          4548 => x"fbb93983",
          4549 => x"f1e6335d",
          4550 => x"7c802e94",
          4551 => x"3883f1c4",
          4552 => x"0847fbca",
          4553 => x"3983f1d0",
          4554 => x"08fc8005",
          4555 => x"49fb9c39",
          4556 => x"83f1d008",
          4557 => x"880547fb",
          4558 => x"b539f33d",
          4559 => x"0d800b84",
          4560 => x"b9943487",
          4561 => x"c0948c70",
          4562 => x"08565787",
          4563 => x"84805274",
          4564 => x"51dad23f",
          4565 => x"84b8e408",
          4566 => x"902b7708",
          4567 => x"57558784",
          4568 => x"80527551",
          4569 => x"dabf3f74",
          4570 => x"84b8e408",
          4571 => x"07770c87",
          4572 => x"c0949c70",
          4573 => x"08565787",
          4574 => x"84805274",
          4575 => x"51daa63f",
          4576 => x"84b8e408",
          4577 => x"902b7708",
          4578 => x"57558784",
          4579 => x"80527551",
          4580 => x"da933f74",
          4581 => x"84b8e408",
          4582 => x"07770c8c",
          4583 => x"80830b87",
          4584 => x"c094840c",
          4585 => x"8c80830b",
          4586 => x"87c09494",
          4587 => x"0c81bce1",
          4588 => x"5c81c7e0",
          4589 => x"5d830284",
          4590 => x"05a10534",
          4591 => x"805e84d4",
          4592 => x"c40b893d",
          4593 => x"7088130c",
          4594 => x"70720c84",
          4595 => x"d4c80c56",
          4596 => x"b6f43f89",
          4597 => x"833f9587",
          4598 => x"3fba8d51",
          4599 => x"94fc3f83",
          4600 => x"d2a05283",
          4601 => x"d2a451c4",
          4602 => x"9f3f83f1",
          4603 => x"d4702252",
          4604 => x"5594873f",
          4605 => x"83d2ac54",
          4606 => x"83d2b853",
          4607 => x"81153352",
          4608 => x"83d2c051",
          4609 => x"c4823f8d",
          4610 => x"973fed82",
          4611 => x"3f8004fb",
          4612 => x"3d0d7770",
          4613 => x"08565680",
          4614 => x"75525374",
          4615 => x"732e8183",
          4616 => x"38743370",
          4617 => x"81ff0652",
          4618 => x"5270a02e",
          4619 => x"09810691",
          4620 => x"38811570",
          4621 => x"337081ff",
          4622 => x"06535355",
          4623 => x"70a02ef1",
          4624 => x"387181ff",
          4625 => x"065473a2",
          4626 => x"2e818238",
          4627 => x"74527281",
          4628 => x"2e80e738",
          4629 => x"80723370",
          4630 => x"81ff0653",
          4631 => x"545470a0",
          4632 => x"2e833881",
          4633 => x"5470802e",
          4634 => x"8b387380",
          4635 => x"2e863881",
          4636 => x"1252e139",
          4637 => x"807381ff",
          4638 => x"06525470",
          4639 => x"a02e0981",
          4640 => x"06833881",
          4641 => x"5470a232",
          4642 => x"70307080",
          4643 => x"25760752",
          4644 => x"52537280",
          4645 => x"2e883880",
          4646 => x"72708105",
          4647 => x"54347176",
          4648 => x"0c745170",
          4649 => x"84b8e40c",
          4650 => x"873d0d04",
          4651 => x"70802ec4",
          4652 => x"3873802e",
          4653 => x"ffbe3881",
          4654 => x"12528072",
          4655 => x"337081ff",
          4656 => x"06535454",
          4657 => x"70a22ee4",
          4658 => x"388154e0",
          4659 => x"39811555",
          4660 => x"81755353",
          4661 => x"72812e09",
          4662 => x"8106fef8",
          4663 => x"38dc39fc",
          4664 => x"3d0d7653",
          4665 => x"72088b38",
          4666 => x"800b84b8",
          4667 => x"e40c863d",
          4668 => x"0d04863d",
          4669 => x"fc055272",
          4670 => x"51db873f",
          4671 => x"84b8e408",
          4672 => x"802ee538",
          4673 => x"7484b8e4",
          4674 => x"0c863d0d",
          4675 => x"04fc3d0d",
          4676 => x"76821133",
          4677 => x"ff055253",
          4678 => x"8152708b",
          4679 => x"26819838",
          4680 => x"831333ff",
          4681 => x"05548252",
          4682 => x"739e2681",
          4683 => x"8a388413",
          4684 => x"33518352",
          4685 => x"70972680",
          4686 => x"fe388513",
          4687 => x"33548452",
          4688 => x"73bb2680",
          4689 => x"f2388613",
          4690 => x"33558552",
          4691 => x"74bb2680",
          4692 => x"e6388813",
          4693 => x"22558652",
          4694 => x"7487e726",
          4695 => x"80d9388a",
          4696 => x"13225487",
          4697 => x"527387e7",
          4698 => x"2680cc38",
          4699 => x"810b87c0",
          4700 => x"989c0c72",
          4701 => x"2287c098",
          4702 => x"bc0c8213",
          4703 => x"3387c098",
          4704 => x"b80c8313",
          4705 => x"3387c098",
          4706 => x"b40c8413",
          4707 => x"3387c098",
          4708 => x"b00c8513",
          4709 => x"3387c098",
          4710 => x"ac0c8613",
          4711 => x"3387c098",
          4712 => x"a80c7487",
          4713 => x"c098a40c",
          4714 => x"7387c098",
          4715 => x"a00c800b",
          4716 => x"87c0989c",
          4717 => x"0c805271",
          4718 => x"84b8e40c",
          4719 => x"863d0d04",
          4720 => x"f33d0d7f",
          4721 => x"5b87c098",
          4722 => x"9c5d817d",
          4723 => x"0c87c098",
          4724 => x"bc085e7d",
          4725 => x"7b2387c0",
          4726 => x"98b8085c",
          4727 => x"7b821c34",
          4728 => x"87c098b4",
          4729 => x"085a7983",
          4730 => x"1c3487c0",
          4731 => x"98b0085c",
          4732 => x"7b841c34",
          4733 => x"87c098ac",
          4734 => x"085a7985",
          4735 => x"1c3487c0",
          4736 => x"98a8085c",
          4737 => x"7b861c34",
          4738 => x"87c098a4",
          4739 => x"085c7b88",
          4740 => x"1c2387c0",
          4741 => x"98a0085a",
          4742 => x"798a1c23",
          4743 => x"807d0c79",
          4744 => x"83ffff06",
          4745 => x"597b83ff",
          4746 => x"ff065886",
          4747 => x"1b335785",
          4748 => x"1b335684",
          4749 => x"1b335583",
          4750 => x"1b335482",
          4751 => x"1b33537d",
          4752 => x"83ffff06",
          4753 => x"5283d888",
          4754 => x"51ffbfbc",
          4755 => x"3f8f3d0d",
          4756 => x"04fe3d0d",
          4757 => x"02930533",
          4758 => x"5372812e",
          4759 => x"a8387251",
          4760 => x"80e8b03f",
          4761 => x"84b8e408",
          4762 => x"982b7098",
          4763 => x"2c515271",
          4764 => x"ff2e0981",
          4765 => x"06863872",
          4766 => x"832ee338",
          4767 => x"7184b8e4",
          4768 => x"0c843d0d",
          4769 => x"04725180",
          4770 => x"e8893f84",
          4771 => x"b8e40898",
          4772 => x"2b70982c",
          4773 => x"515271ff",
          4774 => x"2e098106",
          4775 => x"df387251",
          4776 => x"80e7f03f",
          4777 => x"84b8e408",
          4778 => x"982b7098",
          4779 => x"2c515271",
          4780 => x"ff2ed238",
          4781 => x"c739fd3d",
          4782 => x"0d807054",
          4783 => x"5271882b",
          4784 => x"54815180",
          4785 => x"e7cd3f84",
          4786 => x"b8e40898",
          4787 => x"2b70982c",
          4788 => x"515271ff",
          4789 => x"2eeb3873",
          4790 => x"72078114",
          4791 => x"54528373",
          4792 => x"25db3871",
          4793 => x"84b8e40c",
          4794 => x"853d0d04",
          4795 => x"fc3d0d02",
          4796 => x"9b053383",
          4797 => x"f19c3370",
          4798 => x"81ff0653",
          4799 => x"55557080",
          4800 => x"2e80f438",
          4801 => x"87c09494",
          4802 => x"0870962a",
          4803 => x"70810653",
          4804 => x"54527080",
          4805 => x"2e8c3871",
          4806 => x"912a7081",
          4807 => x"06515170",
          4808 => x"e3387281",
          4809 => x"32810653",
          4810 => x"72802e8a",
          4811 => x"3871932a",
          4812 => x"81065271",
          4813 => x"cf387381",
          4814 => x"ff065187",
          4815 => x"c0948052",
          4816 => x"70802e86",
          4817 => x"3887c094",
          4818 => x"90527472",
          4819 => x"0c7484b8",
          4820 => x"e40c863d",
          4821 => x"0d047191",
          4822 => x"2a708106",
          4823 => x"51517097",
          4824 => x"38728132",
          4825 => x"81065372",
          4826 => x"802ecb38",
          4827 => x"71932a81",
          4828 => x"06527180",
          4829 => x"2ec03887",
          4830 => x"c0948408",
          4831 => x"70962a70",
          4832 => x"81065354",
          4833 => x"5270cf38",
          4834 => x"d839ff3d",
          4835 => x"0d028f05",
          4836 => x"33703070",
          4837 => x"9f2a5152",
          4838 => x"527083f1",
          4839 => x"9c34833d",
          4840 => x"0d04fa3d",
          4841 => x"0d785580",
          4842 => x"75337056",
          4843 => x"52577077",
          4844 => x"2e80e738",
          4845 => x"811583f1",
          4846 => x"9c337081",
          4847 => x"ff065457",
          4848 => x"5571802e",
          4849 => x"80ff3887",
          4850 => x"c0949408",
          4851 => x"70962a70",
          4852 => x"81065354",
          4853 => x"5270802e",
          4854 => x"8c387191",
          4855 => x"2a708106",
          4856 => x"515170e3",
          4857 => x"38728132",
          4858 => x"81065372",
          4859 => x"802e8a38",
          4860 => x"71932a81",
          4861 => x"065271cf",
          4862 => x"387581ff",
          4863 => x"065187c0",
          4864 => x"94805270",
          4865 => x"802e8638",
          4866 => x"87c09490",
          4867 => x"5273720c",
          4868 => x"81177533",
          4869 => x"555773ff",
          4870 => x"9b387684",
          4871 => x"b8e40c88",
          4872 => x"3d0d0471",
          4873 => x"912a7081",
          4874 => x"06515170",
          4875 => x"98387281",
          4876 => x"32810653",
          4877 => x"72802ec1",
          4878 => x"3871932a",
          4879 => x"81065271",
          4880 => x"802effb5",
          4881 => x"3887c094",
          4882 => x"84087096",
          4883 => x"2a708106",
          4884 => x"53545270",
          4885 => x"ce38d739",
          4886 => x"ff3d0d87",
          4887 => x"c09e8008",
          4888 => x"709c2a8a",
          4889 => x"06525270",
          4890 => x"802e84ab",
          4891 => x"3887c09e",
          4892 => x"a40883f1",
          4893 => x"a00c87c0",
          4894 => x"9ea80883",
          4895 => x"f1a40c87",
          4896 => x"c09e9408",
          4897 => x"83f1a80c",
          4898 => x"87c09e98",
          4899 => x"0883f1ac",
          4900 => x"0c87c09e",
          4901 => x"9c0883f1",
          4902 => x"b00c87c0",
          4903 => x"9ea00883",
          4904 => x"f1b40c87",
          4905 => x"c09eac08",
          4906 => x"83f1b80c",
          4907 => x"87c09eb0",
          4908 => x"0883f1bc",
          4909 => x"0c87c09e",
          4910 => x"b40883f1",
          4911 => x"c00c87c0",
          4912 => x"9eb80883",
          4913 => x"f1c40c87",
          4914 => x"c09ebc08",
          4915 => x"83f1c80c",
          4916 => x"87c09ec0",
          4917 => x"0883f1cc",
          4918 => x"0c87c09e",
          4919 => x"c40883f1",
          4920 => x"d00c87c0",
          4921 => x"9e800852",
          4922 => x"7183f1d4",
          4923 => x"2387c09e",
          4924 => x"840883f1",
          4925 => x"d80c87c0",
          4926 => x"9e880883",
          4927 => x"f1dc0c87",
          4928 => x"c09e8c08",
          4929 => x"83f1e00c",
          4930 => x"810b83f1",
          4931 => x"e434800b",
          4932 => x"87c09e90",
          4933 => x"08708480",
          4934 => x"0a065152",
          4935 => x"527082fb",
          4936 => x"387183f1",
          4937 => x"e534800b",
          4938 => x"87c09e90",
          4939 => x"08708880",
          4940 => x"0a065152",
          4941 => x"5270802e",
          4942 => x"83388152",
          4943 => x"7183f1e6",
          4944 => x"34800b87",
          4945 => x"c09e9008",
          4946 => x"7090800a",
          4947 => x"06515252",
          4948 => x"70802e83",
          4949 => x"38815271",
          4950 => x"83f1e734",
          4951 => x"800b87c0",
          4952 => x"9e900870",
          4953 => x"88808006",
          4954 => x"51525270",
          4955 => x"802e8338",
          4956 => x"81527183",
          4957 => x"f1e83480",
          4958 => x"0b87c09e",
          4959 => x"900870a0",
          4960 => x"80800651",
          4961 => x"52527080",
          4962 => x"2e833881",
          4963 => x"527183f1",
          4964 => x"e934800b",
          4965 => x"87c09e90",
          4966 => x"08709080",
          4967 => x"80065152",
          4968 => x"5270802e",
          4969 => x"83388152",
          4970 => x"7183f1ea",
          4971 => x"34800b87",
          4972 => x"c09e9008",
          4973 => x"70848080",
          4974 => x"06515252",
          4975 => x"70802e83",
          4976 => x"38815271",
          4977 => x"83f1eb34",
          4978 => x"800b87c0",
          4979 => x"9e900870",
          4980 => x"82808006",
          4981 => x"51525270",
          4982 => x"802e8338",
          4983 => x"81527183",
          4984 => x"f1ec3480",
          4985 => x"0b87c09e",
          4986 => x"90087081",
          4987 => x"80800651",
          4988 => x"52527080",
          4989 => x"2e833881",
          4990 => x"527183f1",
          4991 => x"ed34800b",
          4992 => x"87c09e90",
          4993 => x"087080c0",
          4994 => x"80065152",
          4995 => x"5270802e",
          4996 => x"83388152",
          4997 => x"7183f1ee",
          4998 => x"34800b87",
          4999 => x"c09e9008",
          5000 => x"70a08006",
          5001 => x"51525270",
          5002 => x"802e8338",
          5003 => x"81527183",
          5004 => x"f1ef3487",
          5005 => x"c09e9008",
          5006 => x"98800670",
          5007 => x"8a2a5351",
          5008 => x"7183f1f0",
          5009 => x"34800b87",
          5010 => x"c09e9008",
          5011 => x"70848006",
          5012 => x"51525270",
          5013 => x"802e8338",
          5014 => x"81527183",
          5015 => x"f1f13487",
          5016 => x"c09e9008",
          5017 => x"83f00670",
          5018 => x"842a5351",
          5019 => x"7183f1f2",
          5020 => x"34800b87",
          5021 => x"c09e9008",
          5022 => x"70880651",
          5023 => x"52527080",
          5024 => x"2e833881",
          5025 => x"527183f1",
          5026 => x"f33487c0",
          5027 => x"9e900887",
          5028 => x"06517083",
          5029 => x"f1f43483",
          5030 => x"3d0d0481",
          5031 => x"52fd8239",
          5032 => x"fb3d0d83",
          5033 => x"d8a051ff",
          5034 => x"b6de3f83",
          5035 => x"f1e43354",
          5036 => x"7386aa38",
          5037 => x"83d8b451",
          5038 => x"c3b93f83",
          5039 => x"f1e63355",
          5040 => x"7485fa38",
          5041 => x"83f1eb33",
          5042 => x"547385d1",
          5043 => x"3883f1e8",
          5044 => x"33567585",
          5045 => x"a83883f1",
          5046 => x"e9335574",
          5047 => x"84ff3883",
          5048 => x"f1ea3354",
          5049 => x"7384d638",
          5050 => x"83f1ef33",
          5051 => x"567584b3",
          5052 => x"3883f1f3",
          5053 => x"33547384",
          5054 => x"903883f1",
          5055 => x"f1335574",
          5056 => x"83ed3883",
          5057 => x"f1e53356",
          5058 => x"7583cf38",
          5059 => x"83f1e733",
          5060 => x"547383b1",
          5061 => x"3883f1ec",
          5062 => x"33557483",
          5063 => x"933883f1",
          5064 => x"ed335675",
          5065 => x"82f43883",
          5066 => x"f1ee3354",
          5067 => x"7381ec38",
          5068 => x"83d8cc51",
          5069 => x"c2bd3f83",
          5070 => x"f1c80852",
          5071 => x"83d8d851",
          5072 => x"ffb5c53f",
          5073 => x"83f1cc08",
          5074 => x"5283d980",
          5075 => x"51ffb5b8",
          5076 => x"3f83f1d0",
          5077 => x"085283d9",
          5078 => x"a851ffb5",
          5079 => x"ab3f83d9",
          5080 => x"d051c28f",
          5081 => x"3f83f1d4",
          5082 => x"225283d9",
          5083 => x"d851ffb5",
          5084 => x"973f83f1",
          5085 => x"d80856bd",
          5086 => x"84c05275",
          5087 => x"51caa63f",
          5088 => x"84b8e408",
          5089 => x"bd84c029",
          5090 => x"76713154",
          5091 => x"5484b8e4",
          5092 => x"085283da",
          5093 => x"8051ffb4",
          5094 => x"ef3f83f1",
          5095 => x"eb335574",
          5096 => x"80c33883",
          5097 => x"f1e63355",
          5098 => x"748a388a",
          5099 => x"51c3af3f",
          5100 => x"873d0d04",
          5101 => x"83f1e008",
          5102 => x"56bd84c0",
          5103 => x"527551c9",
          5104 => x"e43f84b8",
          5105 => x"e408bd84",
          5106 => x"c0297671",
          5107 => x"31545484",
          5108 => x"b8e40852",
          5109 => x"83daac51",
          5110 => x"ffb4ad3f",
          5111 => x"8a51c2fe",
          5112 => x"3f873d0d",
          5113 => x"0483f1dc",
          5114 => x"0856bd84",
          5115 => x"c0527551",
          5116 => x"c9b33f84",
          5117 => x"b8e408bd",
          5118 => x"84c02976",
          5119 => x"71315454",
          5120 => x"84b8e408",
          5121 => x"5283dad8",
          5122 => x"51ffb3fc",
          5123 => x"3f83f1e6",
          5124 => x"33557480",
          5125 => x"2eff9438",
          5126 => x"ff9a3983",
          5127 => x"db8451c0",
          5128 => x"d23f83d8",
          5129 => x"cc51c0cb",
          5130 => x"3f83f1c8",
          5131 => x"085283d8",
          5132 => x"d851ffb3",
          5133 => x"d33f83f1",
          5134 => x"cc085283",
          5135 => x"d98051ff",
          5136 => x"b3c63f83",
          5137 => x"f1d00852",
          5138 => x"83d9a851",
          5139 => x"ffb3b93f",
          5140 => x"83d9d051",
          5141 => x"c09d3f83",
          5142 => x"f1d42252",
          5143 => x"83d9d851",
          5144 => x"ffb3a53f",
          5145 => x"83f1d808",
          5146 => x"56bd84c0",
          5147 => x"527551c8",
          5148 => x"b43f84b8",
          5149 => x"e408bd84",
          5150 => x"c0297671",
          5151 => x"31545484",
          5152 => x"b8e40852",
          5153 => x"83da8051",
          5154 => x"ffb2fd3f",
          5155 => x"83f1eb33",
          5156 => x"5574802e",
          5157 => x"fe8d38fe",
          5158 => x"cc3983db",
          5159 => x"8c51ffbf",
          5160 => x"d23f83f1",
          5161 => x"ee335473",
          5162 => x"802efd84",
          5163 => x"38feec39",
          5164 => x"83db9451",
          5165 => x"ffbfbc3f",
          5166 => x"83f1ed33",
          5167 => x"5675802e",
          5168 => x"fce538d6",
          5169 => x"3983dba0",
          5170 => x"51ffbfa7",
          5171 => x"3f83f1ec",
          5172 => x"33557480",
          5173 => x"2efcc738",
          5174 => x"d73983db",
          5175 => x"ac51ffbf",
          5176 => x"923f83f1",
          5177 => x"e7335473",
          5178 => x"802efca9",
          5179 => x"38d73983",
          5180 => x"f1f23352",
          5181 => x"83dbc051",
          5182 => x"ffb28d3f",
          5183 => x"83f1e533",
          5184 => x"5675802e",
          5185 => x"fc8638d2",
          5186 => x"3983f1f4",
          5187 => x"335283db",
          5188 => x"e051ffb1",
          5189 => x"f33f83f1",
          5190 => x"f1335574",
          5191 => x"802efbe3",
          5192 => x"38cd3983",
          5193 => x"f1f03352",
          5194 => x"83dc8051",
          5195 => x"ffb1d93f",
          5196 => x"83f1f333",
          5197 => x"5473802e",
          5198 => x"fbc038cd",
          5199 => x"3983f1b0",
          5200 => x"0883f1b4",
          5201 => x"08115452",
          5202 => x"83dca051",
          5203 => x"ffb1b93f",
          5204 => x"83f1ef33",
          5205 => x"5675802e",
          5206 => x"fb9738c7",
          5207 => x"3983f1a8",
          5208 => x"0883f1ac",
          5209 => x"08115452",
          5210 => x"83dcbc51",
          5211 => x"ffb1993f",
          5212 => x"83f1ea33",
          5213 => x"5473802e",
          5214 => x"faee38c1",
          5215 => x"3983f1a0",
          5216 => x"0883f1a4",
          5217 => x"08115452",
          5218 => x"83dcd851",
          5219 => x"ffb0f93f",
          5220 => x"83f1e933",
          5221 => x"5574802e",
          5222 => x"fac538c1",
          5223 => x"3983f1b8",
          5224 => x"0883f1bc",
          5225 => x"08115452",
          5226 => x"83dcf451",
          5227 => x"ffb0d93f",
          5228 => x"83f1e833",
          5229 => x"5675802e",
          5230 => x"fa9c38c1",
          5231 => x"3983f1c0",
          5232 => x"0883f1c4",
          5233 => x"08115452",
          5234 => x"83dd9051",
          5235 => x"ffb0b93f",
          5236 => x"83f1eb33",
          5237 => x"5473802e",
          5238 => x"f9f338c1",
          5239 => x"3983ddac",
          5240 => x"51ffb0a4",
          5241 => x"3f83d8b4",
          5242 => x"51ffbd87",
          5243 => x"3f83f1e6",
          5244 => x"33557480",
          5245 => x"2ef9cd38",
          5246 => x"c439ff3d",
          5247 => x"0d028e05",
          5248 => x"33527185",
          5249 => x"268c3871",
          5250 => x"101083c2",
          5251 => x"ec055271",
          5252 => x"080483dd",
          5253 => x"c051ffaf",
          5254 => x"ef3f833d",
          5255 => x"0d0483dd",
          5256 => x"c851ffaf",
          5257 => x"e33f833d",
          5258 => x"0d0483dd",
          5259 => x"d051ffaf",
          5260 => x"d73f833d",
          5261 => x"0d0483dd",
          5262 => x"d851ffaf",
          5263 => x"cb3f833d",
          5264 => x"0d0483dd",
          5265 => x"e051ffaf",
          5266 => x"bf3f833d",
          5267 => x"0d0483dd",
          5268 => x"e851ffaf",
          5269 => x"b33f833d",
          5270 => x"0d047188",
          5271 => x"800c0480",
          5272 => x"0b87c096",
          5273 => x"840c0483",
          5274 => x"f1f80887",
          5275 => x"c096840c",
          5276 => x"04d93d0d",
          5277 => x"aa3d08ad",
          5278 => x"3d085a5a",
          5279 => x"81705758",
          5280 => x"805283f2",
          5281 => x"d0085182",
          5282 => x"88823f84",
          5283 => x"b8e40880",
          5284 => x"ed388b3d",
          5285 => x"57ff0b83",
          5286 => x"f2d00854",
          5287 => x"5580f852",
          5288 => x"765182d2",
          5289 => x"8f3f84b8",
          5290 => x"e408802e",
          5291 => x"a4387651",
          5292 => x"c0f63f84",
          5293 => x"b8e40881",
          5294 => x"17575580",
          5295 => x"0b84b8e4",
          5296 => x"08258e38",
          5297 => x"84b8e408",
          5298 => x"ff057018",
          5299 => x"55558074",
          5300 => x"34740970",
          5301 => x"30707207",
          5302 => x"9f2a5155",
          5303 => x"5578762e",
          5304 => x"853873ff",
          5305 => x"b03883f2",
          5306 => x"d0088c11",
          5307 => x"08535182",
          5308 => x"879a3f84",
          5309 => x"b8e4088f",
          5310 => x"3878762e",
          5311 => x"9a387784",
          5312 => x"b8e40ca9",
          5313 => x"3d0d0483",
          5314 => x"e19851ff",
          5315 => x"adfa3f78",
          5316 => x"762e0981",
          5317 => x"06e83876",
          5318 => x"527951c0",
          5319 => x"aa3f7951",
          5320 => x"c0863fab",
          5321 => x"3d085684",
          5322 => x"b8e40876",
          5323 => x"34765283",
          5324 => x"e1c451ff",
          5325 => x"add23f80",
          5326 => x"0b84b8e4",
          5327 => x"0ca93d0d",
          5328 => x"04d83d0d",
          5329 => x"ab3d08ad",
          5330 => x"3d087172",
          5331 => x"5d723357",
          5332 => x"575a5773",
          5333 => x"a02e8191",
          5334 => x"38800b8d",
          5335 => x"3d595675",
          5336 => x"10101083",
          5337 => x"f2d80570",
          5338 => x"085254ff",
          5339 => x"bfba3f84",
          5340 => x"b8e40853",
          5341 => x"79527308",
          5342 => x"51c09a3f",
          5343 => x"84b8e408",
          5344 => x"90388414",
          5345 => x"33547381",
          5346 => x"2e818838",
          5347 => x"73822e99",
          5348 => x"38811670",
          5349 => x"81ff0657",
          5350 => x"54827627",
          5351 => x"c2388054",
          5352 => x"7384b8e4",
          5353 => x"0caa3d0d",
          5354 => x"04811a5a",
          5355 => x"aa3dff84",
          5356 => x"1153ff80",
          5357 => x"0551c7ce",
          5358 => x"3f84b8e4",
          5359 => x"08802ed1",
          5360 => x"38ff1b53",
          5361 => x"78527651",
          5362 => x"fda73f84",
          5363 => x"b8e40881",
          5364 => x"ff065473",
          5365 => x"802ec938",
          5366 => x"81167081",
          5367 => x"ff065754",
          5368 => x"827627fe",
          5369 => x"fa38ffb6",
          5370 => x"39783377",
          5371 => x"05567676",
          5372 => x"27fee638",
          5373 => x"8115705b",
          5374 => x"70335555",
          5375 => x"73a02e09",
          5376 => x"8106fed5",
          5377 => x"38757526",
          5378 => x"eb38800b",
          5379 => x"8d3d5956",
          5380 => x"fecd3973",
          5381 => x"84b8e408",
          5382 => x"5383f2d0",
          5383 => x"08525682",
          5384 => x"84ea3f84",
          5385 => x"b8e40880",
          5386 => x"d03883f2",
          5387 => x"d0085380",
          5388 => x"f8527751",
          5389 => x"82cefd3f",
          5390 => x"84b8e408",
          5391 => x"802eba38",
          5392 => x"7751ffbd",
          5393 => x"e33f84b8",
          5394 => x"e4085580",
          5395 => x"0b84b8e4",
          5396 => x"08259d38",
          5397 => x"84b8e408",
          5398 => x"ff057019",
          5399 => x"58558077",
          5400 => x"34775375",
          5401 => x"52811683",
          5402 => x"e18c5256",
          5403 => x"ffab993f",
          5404 => x"74ff2e09",
          5405 => x"8106ffb2",
          5406 => x"38810b84",
          5407 => x"b8e40caa",
          5408 => x"3d0d04ce",
          5409 => x"3d0db53d",
          5410 => x"08b73d08",
          5411 => x"b93d085a",
          5412 => x"415c800b",
          5413 => x"b43d3483",
          5414 => x"f2d43383",
          5415 => x"f2d00856",
          5416 => x"5d749e38",
          5417 => x"7483f2cc",
          5418 => x"33565674",
          5419 => x"802e82cb",
          5420 => x"3877802e",
          5421 => x"918d3881",
          5422 => x"7077065a",
          5423 => x"577890a0",
          5424 => x"3877802e",
          5425 => x"90fd3893",
          5426 => x"3db43d5f",
          5427 => x"5f8051eb",
          5428 => x"803f84b8",
          5429 => x"e408982b",
          5430 => x"70982c5b",
          5431 => x"5679ff2e",
          5432 => x"ec387981",
          5433 => x"ff0684d0",
          5434 => x"a0337098",
          5435 => x"2b70982c",
          5436 => x"84d09c33",
          5437 => x"70982b70",
          5438 => x"972c7198",
          5439 => x"2c057010",
          5440 => x"1083ddec",
          5441 => x"05700815",
          5442 => x"70335253",
          5443 => x"5c5d4652",
          5444 => x"5b585c59",
          5445 => x"81577479",
          5446 => x"2e80cd38",
          5447 => x"78752781",
          5448 => x"87387581",
          5449 => x"800a2981",
          5450 => x"ff0a0570",
          5451 => x"982c5755",
          5452 => x"80762481",
          5453 => x"cb387510",
          5454 => x"1670822b",
          5455 => x"5657800b",
          5456 => x"83ddf016",
          5457 => x"33425777",
          5458 => x"61259138",
          5459 => x"83ddec15",
          5460 => x"08187033",
          5461 => x"56417875",
          5462 => x"2e819538",
          5463 => x"76802ec2",
          5464 => x"387584d0",
          5465 => x"9c348157",
          5466 => x"76802e81",
          5467 => x"9938811b",
          5468 => x"70982b70",
          5469 => x"982c84d0",
          5470 => x"9c337098",
          5471 => x"2b70972c",
          5472 => x"71982c05",
          5473 => x"70822b83",
          5474 => x"ddf01133",
          5475 => x"5f535f5d",
          5476 => x"585d5757",
          5477 => x"7a782e81",
          5478 => x"90387684",
          5479 => x"d0a034fe",
          5480 => x"ac398157",
          5481 => x"76ffba38",
          5482 => x"7581800a",
          5483 => x"2981800a",
          5484 => x"0570982c",
          5485 => x"7081ff06",
          5486 => x"59574176",
          5487 => x"952680c0",
          5488 => x"38751016",
          5489 => x"70822b51",
          5490 => x"55800b83",
          5491 => x"ddf01633",
          5492 => x"42577761",
          5493 => x"25ce3883",
          5494 => x"ddec1508",
          5495 => x"18703342",
          5496 => x"5578612e",
          5497 => x"ffbc3876",
          5498 => x"802effbc",
          5499 => x"38fef239",
          5500 => x"81577680",
          5501 => x"2efeab38",
          5502 => x"fee73981",
          5503 => x"56fdb239",
          5504 => x"805776fe",
          5505 => x"e9387684",
          5506 => x"d0a03476",
          5507 => x"84d09c34",
          5508 => x"797e3476",
          5509 => x"7f0c6255",
          5510 => x"749526fd",
          5511 => x"b0387410",
          5512 => x"1083c384",
          5513 => x"05577608",
          5514 => x"0483ddf4",
          5515 => x"15087f0c",
          5516 => x"800b84d0",
          5517 => x"a034800b",
          5518 => x"84d09c34",
          5519 => x"d93984d0",
          5520 => x"a8335675",
          5521 => x"802efd85",
          5522 => x"3884d4c8",
          5523 => x"08528851",
          5524 => x"ffb69b3f",
          5525 => x"84d0a833",
          5526 => x"ff055776",
          5527 => x"84d0a834",
          5528 => x"fceb3984",
          5529 => x"d0a83370",
          5530 => x"81ff0684",
          5531 => x"d0a4335b",
          5532 => x"57557579",
          5533 => x"27fcd638",
          5534 => x"84d4c808",
          5535 => x"52811558",
          5536 => x"7784d0a8",
          5537 => x"347b1670",
          5538 => x"335255ff",
          5539 => x"b5e03ffc",
          5540 => x"bc397c93",
          5541 => x"2e8bda38",
          5542 => x"7c101083",
          5543 => x"f2800570",
          5544 => x"08575975",
          5545 => x"8f833875",
          5546 => x"84d0a434",
          5547 => x"757c3484",
          5548 => x"d0a43384",
          5549 => x"d0a83356",
          5550 => x"5674802e",
          5551 => x"b63884d4",
          5552 => x"c8085288",
          5553 => x"51ffb5a6",
          5554 => x"3f84d4c8",
          5555 => x"0852a051",
          5556 => x"ffb59b3f",
          5557 => x"84d4c808",
          5558 => x"528851ff",
          5559 => x"b5903f84",
          5560 => x"d0a833ff",
          5561 => x"055b7a84",
          5562 => x"d0a8347a",
          5563 => x"81ff0655",
          5564 => x"74cc387b",
          5565 => x"51ffa690",
          5566 => x"3f7584d0",
          5567 => x"a834fbcd",
          5568 => x"397c8a38",
          5569 => x"83f2c808",
          5570 => x"56758d9e",
          5571 => x"387c1010",
          5572 => x"83f1fc05",
          5573 => x"fc110857",
          5574 => x"55758ef9",
          5575 => x"38740856",
          5576 => x"75802efb",
          5577 => x"a8387551",
          5578 => x"ffb7fd3f",
          5579 => x"84b8e408",
          5580 => x"84d0a434",
          5581 => x"84b8e408",
          5582 => x"81ff0681",
          5583 => x"05537552",
          5584 => x"7b51ffb8",
          5585 => x"a53f84d0",
          5586 => x"a43384d0",
          5587 => x"a8335656",
          5588 => x"74802eff",
          5589 => x"9e3884d4",
          5590 => x"c8085288",
          5591 => x"51ffb48e",
          5592 => x"3f84d4c8",
          5593 => x"0852a051",
          5594 => x"ffb4833f",
          5595 => x"84d4c808",
          5596 => x"528851ff",
          5597 => x"b3f83f84",
          5598 => x"d0a833ff",
          5599 => x"05557484",
          5600 => x"d0a83474",
          5601 => x"81ff0655",
          5602 => x"c73984d0",
          5603 => x"a8337081",
          5604 => x"ff0684d0",
          5605 => x"a4335b57",
          5606 => x"55757927",
          5607 => x"faaf3884",
          5608 => x"d4c80852",
          5609 => x"81155776",
          5610 => x"84d0a834",
          5611 => x"7b167033",
          5612 => x"5255ffb3",
          5613 => x"b93f84d0",
          5614 => x"a8337081",
          5615 => x"ff0684d0",
          5616 => x"a4335a57",
          5617 => x"55757827",
          5618 => x"fa833884",
          5619 => x"d4c80852",
          5620 => x"81155776",
          5621 => x"84d0a834",
          5622 => x"7b167033",
          5623 => x"5255ffb3",
          5624 => x"8d3f84d0",
          5625 => x"a8337081",
          5626 => x"ff0684d0",
          5627 => x"a4335a57",
          5628 => x"55777626",
          5629 => x"ffa938f9",
          5630 => x"d43984d0",
          5631 => x"a83384d0",
          5632 => x"a4335656",
          5633 => x"74762ef9",
          5634 => x"c438ff15",
          5635 => x"5b7a84d0",
          5636 => x"a4347598",
          5637 => x"2b70982c",
          5638 => x"7c81ff06",
          5639 => x"43575a60",
          5640 => x"762480ef",
          5641 => x"3884d4c8",
          5642 => x"0852a051",
          5643 => x"ffb2bf3f",
          5644 => x"84d0a833",
          5645 => x"70982b70",
          5646 => x"982c84d0",
          5647 => x"a4335a57",
          5648 => x"57417477",
          5649 => x"24f98638",
          5650 => x"84d4c808",
          5651 => x"528851ff",
          5652 => x"b29c3f74",
          5653 => x"81800a29",
          5654 => x"81800a05",
          5655 => x"70982c84",
          5656 => x"d0a4335d",
          5657 => x"565a747b",
          5658 => x"24f8e238",
          5659 => x"84d4c808",
          5660 => x"528851ff",
          5661 => x"b1f83f74",
          5662 => x"81800a29",
          5663 => x"81800a05",
          5664 => x"70982c84",
          5665 => x"d0a4335d",
          5666 => x"565a7a75",
          5667 => x"25ffb938",
          5668 => x"f8bb397b",
          5669 => x"16588118",
          5670 => x"33783484",
          5671 => x"d4c80852",
          5672 => x"773351ff",
          5673 => x"b1c83f75",
          5674 => x"81800a29",
          5675 => x"81800a05",
          5676 => x"70982c84",
          5677 => x"d0a4335b",
          5678 => x"57557579",
          5679 => x"25fee638",
          5680 => x"7b165881",
          5681 => x"18337834",
          5682 => x"84d4c808",
          5683 => x"52773351",
          5684 => x"ffb19b3f",
          5685 => x"7581800a",
          5686 => x"2981800a",
          5687 => x"0570982c",
          5688 => x"84d0a433",
          5689 => x"5b575578",
          5690 => x"7624ffa7",
          5691 => x"38feb639",
          5692 => x"84d0a833",
          5693 => x"5574802e",
          5694 => x"f7d33884",
          5695 => x"d4c80852",
          5696 => x"8851ffb0",
          5697 => x"e93f84d0",
          5698 => x"a833ff05",
          5699 => x"577684d0",
          5700 => x"a8347681",
          5701 => x"ff0655dd",
          5702 => x"3984d0a4",
          5703 => x"337c055f",
          5704 => x"807f3484",
          5705 => x"d4c80852",
          5706 => x"8a51ffb0",
          5707 => x"c13f84d0",
          5708 => x"a4527b51",
          5709 => x"f48b3f84",
          5710 => x"b8e40881",
          5711 => x"ff065877",
          5712 => x"89cf3884",
          5713 => x"d0a43357",
          5714 => x"76802e80",
          5715 => x"d83883f2",
          5716 => x"d4337010",
          5717 => x"1083f1fc",
          5718 => x"05700857",
          5719 => x"5e56748b",
          5720 => x"a0387582",
          5721 => x"2b87fc06",
          5722 => x"83f1fc05",
          5723 => x"81187053",
          5724 => x"575b80e7",
          5725 => x"fb3f84b8",
          5726 => x"e4087b0c",
          5727 => x"83f2d433",
          5728 => x"70101083",
          5729 => x"f1fc0570",
          5730 => x"08574141",
          5731 => x"748bad38",
          5732 => x"83f2d008",
          5733 => x"5675802e",
          5734 => x"8c3883f2",
          5735 => x"cc335877",
          5736 => x"802e8bbc",
          5737 => x"38800b84",
          5738 => x"d0a83480",
          5739 => x"0b84d0a4",
          5740 => x"347b84b8",
          5741 => x"e40cb43d",
          5742 => x"0d0484d0",
          5743 => x"a8335574",
          5744 => x"802eb638",
          5745 => x"84d4c808",
          5746 => x"528851ff",
          5747 => x"afa03f84",
          5748 => x"d4c80852",
          5749 => x"a051ffaf",
          5750 => x"953f84d4",
          5751 => x"c8085288",
          5752 => x"51ffaf8a",
          5753 => x"3f84d0a8",
          5754 => x"33ff0556",
          5755 => x"7584d0a8",
          5756 => x"347581ff",
          5757 => x"065574cc",
          5758 => x"3883d1e0",
          5759 => x"51ffa088",
          5760 => x"3f800b84",
          5761 => x"d0a83480",
          5762 => x"0b84d0a4",
          5763 => x"34f5be39",
          5764 => x"837c3480",
          5765 => x"0b811d34",
          5766 => x"84d0a833",
          5767 => x"5574802e",
          5768 => x"b63884d4",
          5769 => x"c8085288",
          5770 => x"51ffaec2",
          5771 => x"3f84d4c8",
          5772 => x"0852a051",
          5773 => x"ffaeb73f",
          5774 => x"84d4c808",
          5775 => x"528851ff",
          5776 => x"aeac3f84",
          5777 => x"d0a833ff",
          5778 => x"055d7c84",
          5779 => x"d0a8347c",
          5780 => x"81ff0655",
          5781 => x"74cc3883",
          5782 => x"d1e051ff",
          5783 => x"9faa3f80",
          5784 => x"0b84d0a8",
          5785 => x"34800b84",
          5786 => x"d0a4347b",
          5787 => x"84b8e40c",
          5788 => x"b43d0d04",
          5789 => x"84d0a833",
          5790 => x"7081ff06",
          5791 => x"5c567a80",
          5792 => x"2ef4ca38",
          5793 => x"84d0a433",
          5794 => x"ff055978",
          5795 => x"84d0a434",
          5796 => x"ff165877",
          5797 => x"84d0a834",
          5798 => x"84d4c808",
          5799 => x"528851ff",
          5800 => x"adcc3f84",
          5801 => x"d0a83370",
          5802 => x"982b7098",
          5803 => x"2c84d0a4",
          5804 => x"335a525b",
          5805 => x"56767624",
          5806 => x"80ef3884",
          5807 => x"d4c80852",
          5808 => x"a051ffad",
          5809 => x"a93f84d0",
          5810 => x"a8337098",
          5811 => x"2b70982c",
          5812 => x"84d0a433",
          5813 => x"5d575956",
          5814 => x"747a24f3",
          5815 => x"f03884d4",
          5816 => x"c8085288",
          5817 => x"51ffad86",
          5818 => x"3f748180",
          5819 => x"0a298180",
          5820 => x"0a057098",
          5821 => x"2c84d0a4",
          5822 => x"335b5155",
          5823 => x"747924f3",
          5824 => x"cc3884d4",
          5825 => x"c8085288",
          5826 => x"51fface2",
          5827 => x"3f748180",
          5828 => x"0a298180",
          5829 => x"0a057098",
          5830 => x"2c84d0a4",
          5831 => x"335b5155",
          5832 => x"787525ff",
          5833 => x"b938f3a5",
          5834 => x"397b1657",
          5835 => x"81173377",
          5836 => x"3484d4c8",
          5837 => x"08527633",
          5838 => x"51ffacb2",
          5839 => x"3f758180",
          5840 => x"0a298180",
          5841 => x"0a057098",
          5842 => x"2c84d0a4",
          5843 => x"3343575b",
          5844 => x"756125fe",
          5845 => x"e6387b16",
          5846 => x"57811733",
          5847 => x"773484d4",
          5848 => x"c8085276",
          5849 => x"3351ffac",
          5850 => x"853f7581",
          5851 => x"800a2981",
          5852 => x"800a0570",
          5853 => x"982c84d0",
          5854 => x"a4334357",
          5855 => x"5b607624",
          5856 => x"ffa738fe",
          5857 => x"b63984d0",
          5858 => x"a8337081",
          5859 => x"ff065858",
          5860 => x"76602ef2",
          5861 => x"b83884d0",
          5862 => x"a4335576",
          5863 => x"7527ae38",
          5864 => x"74982b70",
          5865 => x"982c5741",
          5866 => x"767624a1",
          5867 => x"387b165b",
          5868 => x"7a33811c",
          5869 => x"34758180",
          5870 => x"0a2981ff",
          5871 => x"0a057098",
          5872 => x"2c84d0a8",
          5873 => x"33525758",
          5874 => x"757825e1",
          5875 => x"38811855",
          5876 => x"7484d0a8",
          5877 => x"347781ff",
          5878 => x"067c055a",
          5879 => x"b33d337a",
          5880 => x"3484d0a4",
          5881 => x"33577660",
          5882 => x"258b3881",
          5883 => x"17567584",
          5884 => x"d0a43475",
          5885 => x"5784d0a8",
          5886 => x"33708180",
          5887 => x"0a2981ff",
          5888 => x"0a057098",
          5889 => x"2c7981ff",
          5890 => x"0644585c",
          5891 => x"58607624",
          5892 => x"81ef3877",
          5893 => x"982b7098",
          5894 => x"2c7881ff",
          5895 => x"065c5759",
          5896 => x"757a25f1",
          5897 => x"a83884d4",
          5898 => x"c8085288",
          5899 => x"51ffaabe",
          5900 => x"3f758180",
          5901 => x"0a298180",
          5902 => x"0a057098",
          5903 => x"2c84d0a4",
          5904 => x"33575741",
          5905 => x"757525f1",
          5906 => x"843884d4",
          5907 => x"c8085288",
          5908 => x"51ffaa9a",
          5909 => x"3f758180",
          5910 => x"0a298180",
          5911 => x"0a057098",
          5912 => x"2c84d0a4",
          5913 => x"33575741",
          5914 => x"747624ff",
          5915 => x"b938f0dd",
          5916 => x"3983f1fc",
          5917 => x"08567580",
          5918 => x"2ef49d38",
          5919 => x"7551ffad",
          5920 => x"a73f84b8",
          5921 => x"e40884d0",
          5922 => x"a43484b8",
          5923 => x"e40881ff",
          5924 => x"06810553",
          5925 => x"75527b51",
          5926 => x"ffadcf3f",
          5927 => x"84d0a433",
          5928 => x"84d0a833",
          5929 => x"56567480",
          5930 => x"2ef4c838",
          5931 => x"84d4c808",
          5932 => x"528851ff",
          5933 => x"a9b83f84",
          5934 => x"d4c80852",
          5935 => x"a051ffa9",
          5936 => x"ad3f84d4",
          5937 => x"c8085288",
          5938 => x"51ffa9a2",
          5939 => x"3f84d0a8",
          5940 => x"33ff055b",
          5941 => x"7a84d0a8",
          5942 => x"347a81ff",
          5943 => x"0655c739",
          5944 => x"a85180e1",
          5945 => x"8b3f84b8",
          5946 => x"e40883f2",
          5947 => x"d00c84b8",
          5948 => x"e40885a5",
          5949 => x"387683f2",
          5950 => x"cc3477ef",
          5951 => x"ca3880c3",
          5952 => x"3984d4c8",
          5953 => x"08527b16",
          5954 => x"70335258",
          5955 => x"ffa8df3f",
          5956 => x"7581800a",
          5957 => x"2981800a",
          5958 => x"0570982c",
          5959 => x"84d0a433",
          5960 => x"52575776",
          5961 => x"7624da38",
          5962 => x"84d0a833",
          5963 => x"70982b70",
          5964 => x"982c7981",
          5965 => x"ff065d58",
          5966 => x"5a58757a",
          5967 => x"25ef8e38",
          5968 => x"fde43983",
          5969 => x"f2d00880",
          5970 => x"2eeefc38",
          5971 => x"83f1fc57",
          5972 => x"93567608",
          5973 => x"5574bb38",
          5974 => x"ff168418",
          5975 => x"58567580",
          5976 => x"25f03880",
          5977 => x"0b83f2d4",
          5978 => x"3483f2d0",
          5979 => x"08557480",
          5980 => x"2eeed438",
          5981 => x"745181e7",
          5982 => x"f63f83f2",
          5983 => x"d0085180",
          5984 => x"d9fe3f80",
          5985 => x"0b83f2d0",
          5986 => x"0c933db4",
          5987 => x"3d5f5fee",
          5988 => x"bc397451",
          5989 => x"80d9e93f",
          5990 => x"80770cff",
          5991 => x"16841858",
          5992 => x"56758025",
          5993 => x"ffac38ff",
          5994 => x"ba397551",
          5995 => x"ffaaf93f",
          5996 => x"84b8e408",
          5997 => x"84d0a434",
          5998 => x"84b8e408",
          5999 => x"81ff0681",
          6000 => x"05537552",
          6001 => x"7b51ffab",
          6002 => x"a13f930b",
          6003 => x"84d0a433",
          6004 => x"84d0a833",
          6005 => x"57575d74",
          6006 => x"802ef297",
          6007 => x"3884d4c8",
          6008 => x"08528851",
          6009 => x"ffa7873f",
          6010 => x"84d4c808",
          6011 => x"52a051ff",
          6012 => x"a6fc3f84",
          6013 => x"d4c80852",
          6014 => x"8851ffa6",
          6015 => x"f13f84d0",
          6016 => x"a833ff05",
          6017 => x"5a7984d0",
          6018 => x"a8347981",
          6019 => x"ff0655c7",
          6020 => x"39807c34",
          6021 => x"800b84d0",
          6022 => x"a834800b",
          6023 => x"84d0a434",
          6024 => x"7b84b8e4",
          6025 => x"0cb43d0d",
          6026 => x"047551ff",
          6027 => x"a9fa3f84",
          6028 => x"b8e40884",
          6029 => x"d0a43484",
          6030 => x"b8e40881",
          6031 => x"ff068105",
          6032 => x"5375527b",
          6033 => x"51ffaaa2",
          6034 => x"3f811d70",
          6035 => x"81ff0684",
          6036 => x"d0a43384",
          6037 => x"d0a83358",
          6038 => x"525e5674",
          6039 => x"802ef193",
          6040 => x"3884d4c8",
          6041 => x"08528851",
          6042 => x"ffa6833f",
          6043 => x"84d4c808",
          6044 => x"52a051ff",
          6045 => x"a5f83f84",
          6046 => x"d4c80852",
          6047 => x"8851ffa5",
          6048 => x"ed3f84d0",
          6049 => x"a833ff05",
          6050 => x"577684d0",
          6051 => x"a8347681",
          6052 => x"ff0655c7",
          6053 => x"397551ff",
          6054 => x"a98e3f84",
          6055 => x"b8e40884",
          6056 => x"d0a43484",
          6057 => x"b8e40881",
          6058 => x"ff068105",
          6059 => x"5375527b",
          6060 => x"51ffa9b6",
          6061 => x"3fff1d70",
          6062 => x"81ff0684",
          6063 => x"d0a43384",
          6064 => x"d0a83358",
          6065 => x"585e5874",
          6066 => x"802ef0a7",
          6067 => x"3884d4c8",
          6068 => x"08528851",
          6069 => x"ffa5973f",
          6070 => x"84d4c808",
          6071 => x"52a051ff",
          6072 => x"a58c3f84",
          6073 => x"d4c80852",
          6074 => x"8851ffa5",
          6075 => x"813f84d0",
          6076 => x"a833ff05",
          6077 => x"416084d0",
          6078 => x"a8346081",
          6079 => x"ff0655c7",
          6080 => x"39745180",
          6081 => x"d6fa3f83",
          6082 => x"f2d43370",
          6083 => x"822b87fc",
          6084 => x"0683f1fc",
          6085 => x"05811970",
          6086 => x"54525c56",
          6087 => x"80dcd13f",
          6088 => x"84b8e408",
          6089 => x"7b0c83f2",
          6090 => x"d4337010",
          6091 => x"1083f1fc",
          6092 => x"05700857",
          6093 => x"41417480",
          6094 => x"2ef4d538",
          6095 => x"75537b52",
          6096 => x"7451ffa8",
          6097 => x"a53f83f2",
          6098 => x"d4338105",
          6099 => x"7081ff06",
          6100 => x"5a569379",
          6101 => x"2782f238",
          6102 => x"7783f2d4",
          6103 => x"34f4b139",
          6104 => x"b43dfef8",
          6105 => x"05547653",
          6106 => x"7b527551",
          6107 => x"81d8c03f",
          6108 => x"83f2d008",
          6109 => x"528a5182",
          6110 => x"ba883f83",
          6111 => x"f2d00851",
          6112 => x"81dff33f",
          6113 => x"800b84d0",
          6114 => x"a834800b",
          6115 => x"84d0a434",
          6116 => x"7b84b8e4",
          6117 => x"0cb43d0d",
          6118 => x"04935377",
          6119 => x"5284b8e4",
          6120 => x"085181c9",
          6121 => x"f83f84b8",
          6122 => x"e40882a5",
          6123 => x"3884b8e4",
          6124 => x"08963d5c",
          6125 => x"5d83f2d0",
          6126 => x"085380f8",
          6127 => x"527a5182",
          6128 => x"b7f23f84",
          6129 => x"b8e4085a",
          6130 => x"84b8e408",
          6131 => x"7b2e0981",
          6132 => x"06e9ee38",
          6133 => x"84b8e408",
          6134 => x"51ffa6cc",
          6135 => x"3f84b8e4",
          6136 => x"0856800b",
          6137 => x"84b8e408",
          6138 => x"2580e338",
          6139 => x"84b8e408",
          6140 => x"ff05701b",
          6141 => x"58568077",
          6142 => x"347581ff",
          6143 => x"0683f2d4",
          6144 => x"33701010",
          6145 => x"83f1fc05",
          6146 => x"70085840",
          6147 => x"58597480",
          6148 => x"f2387682",
          6149 => x"2b87fc06",
          6150 => x"83f1fc05",
          6151 => x"811a7053",
          6152 => x"585580da",
          6153 => x"cb3f84b8",
          6154 => x"e408750c",
          6155 => x"83f2d433",
          6156 => x"70101083",
          6157 => x"f1fc0570",
          6158 => x"08574041",
          6159 => x"74a03881",
          6160 => x"1d7081ff",
          6161 => x"065e5793",
          6162 => x"7d278338",
          6163 => x"805d75ff",
          6164 => x"2e098106",
          6165 => x"fedf3877",
          6166 => x"e8ed38f9",
          6167 => x"e6397653",
          6168 => x"79527451",
          6169 => x"ffa6833f",
          6170 => x"83f2d433",
          6171 => x"81057081",
          6172 => x"ff065b57",
          6173 => x"937a2780",
          6174 => x"c838800b",
          6175 => x"83f2d434",
          6176 => x"ffbd3974",
          6177 => x"5180d3f8",
          6178 => x"3f83f2d4",
          6179 => x"3370822b",
          6180 => x"87fc0683",
          6181 => x"f1fc0581",
          6182 => x"1b705452",
          6183 => x"565780d9",
          6184 => x"cf3f84b8",
          6185 => x"e408750c",
          6186 => x"83f2d433",
          6187 => x"70101083",
          6188 => x"f1fc0570",
          6189 => x"08574041",
          6190 => x"74802eff",
          6191 => x"8238ff9e",
          6192 => x"397683f2",
          6193 => x"d434fef7",
          6194 => x"397583f2",
          6195 => x"d434f1c0",
          6196 => x"3983e0cc",
          6197 => x"51ff9f9b",
          6198 => x"3f77e7eb",
          6199 => x"38f8e439",
          6200 => x"f23d0d02",
          6201 => x"80c30533",
          6202 => x"02840580",
          6203 => x"c705335b",
          6204 => x"53728326",
          6205 => x"818d3872",
          6206 => x"812e818b",
          6207 => x"38817325",
          6208 => x"839e3872",
          6209 => x"822e82a8",
          6210 => x"3886a7a0",
          6211 => x"805986a7",
          6212 => x"b080705e",
          6213 => x"5780569f",
          6214 => x"a0587976",
          6215 => x"2e903875",
          6216 => x"83f89434",
          6217 => x"7583f895",
          6218 => x"347583f8",
          6219 => x"922383f8",
          6220 => x"90337098",
          6221 => x"2b71902b",
          6222 => x"0771882b",
          6223 => x"0771077a",
          6224 => x"7f565656",
          6225 => x"5b787727",
          6226 => x"94388074",
          6227 => x"70840556",
          6228 => x"0c747370",
          6229 => x"8405550c",
          6230 => x"767426ee",
          6231 => x"38757827",
          6232 => x"a23883f8",
          6233 => x"90338497",
          6234 => x"b6177978",
          6235 => x"31555555",
          6236 => x"a00be0e0",
          6237 => x"15347474",
          6238 => x"70810556",
          6239 => x"34ff1353",
          6240 => x"72ee3890",
          6241 => x"3d0d0486",
          6242 => x"a7a0800b",
          6243 => x"83f89433",
          6244 => x"70101011",
          6245 => x"83f89533",
          6246 => x"71902911",
          6247 => x"74055b41",
          6248 => x"58405986",
          6249 => x"a7b0800b",
          6250 => x"84b6d833",
          6251 => x"7081ff06",
          6252 => x"84b6d733",
          6253 => x"7081ff06",
          6254 => x"83f89222",
          6255 => x"7083ffff",
          6256 => x"06707529",
          6257 => x"5d595d58",
          6258 => x"5e575b5d",
          6259 => x"73732687",
          6260 => x"38727431",
          6261 => x"75295679",
          6262 => x"81ff067e",
          6263 => x"81ff067c",
          6264 => x"81ff067a",
          6265 => x"83ffff06",
          6266 => x"6281ff06",
          6267 => x"70752914",
          6268 => x"5d425757",
          6269 => x"5b5c7474",
          6270 => x"268f3883",
          6271 => x"f8943374",
          6272 => x"76310570",
          6273 => x"7d291b59",
          6274 => x"5f768306",
          6275 => x"5c7b802e",
          6276 => x"fe9c3878",
          6277 => x"7d555372",
          6278 => x"7726fec1",
          6279 => x"38807370",
          6280 => x"81055534",
          6281 => x"83f89033",
          6282 => x"74708105",
          6283 => x"5634e839",
          6284 => x"86a7a080",
          6285 => x"5986a7b0",
          6286 => x"807084b6",
          6287 => x"d8337081",
          6288 => x"ff0684b6",
          6289 => x"d7337081",
          6290 => x"ff0683f8",
          6291 => x"92227074",
          6292 => x"295d5b5d",
          6293 => x"575e565e",
          6294 => x"57747827",
          6295 => x"81df3873",
          6296 => x"81ff0673",
          6297 => x"81ff0671",
          6298 => x"7129185a",
          6299 => x"54547980",
          6300 => x"2efdbb38",
          6301 => x"800b83f8",
          6302 => x"9434800b",
          6303 => x"83f89534",
          6304 => x"83f89033",
          6305 => x"70982b71",
          6306 => x"902b0771",
          6307 => x"882b0771",
          6308 => x"077a7f56",
          6309 => x"56565b76",
          6310 => x"7926fdae",
          6311 => x"38fdbe39",
          6312 => x"72fce638",
          6313 => x"83f89433",
          6314 => x"7081ff06",
          6315 => x"70101011",
          6316 => x"83f89533",
          6317 => x"71902911",
          6318 => x"86a7a080",
          6319 => x"115e575b",
          6320 => x"56565f86",
          6321 => x"a7b08070",
          6322 => x"1484b6d8",
          6323 => x"337081ff",
          6324 => x"0684b6d7",
          6325 => x"337081ff",
          6326 => x"0683f892",
          6327 => x"227083ff",
          6328 => x"ff067c75",
          6329 => x"2960055e",
          6330 => x"5a415f58",
          6331 => x"5f405e57",
          6332 => x"7973268b",
          6333 => x"38727a31",
          6334 => x"15707d29",
          6335 => x"1957537d",
          6336 => x"81ff0674",
          6337 => x"81ff0671",
          6338 => x"71297d83",
          6339 => x"ffff0662",
          6340 => x"81ff0670",
          6341 => x"7529585f",
          6342 => x"5b5c5d55",
          6343 => x"7b782685",
          6344 => x"38777529",
          6345 => x"53797331",
          6346 => x"16798306",
          6347 => x"5b5879fd",
          6348 => x"e2387683",
          6349 => x"065c7bfd",
          6350 => x"da38fbf2",
          6351 => x"39747831",
          6352 => x"7b2956fe",
          6353 => x"9a39fb3d",
          6354 => x"0d86ee80",
          6355 => x"8c53ff8a",
          6356 => x"73348773",
          6357 => x"34857334",
          6358 => x"81733486",
          6359 => x"ee809c55",
          6360 => x"80f47534",
          6361 => x"ffb07534",
          6362 => x"86ee8098",
          6363 => x"56807634",
          6364 => x"80763486",
          6365 => x"ee809454",
          6366 => x"8a743480",
          6367 => x"7434ff80",
          6368 => x"75348152",
          6369 => x"8351fad8",
          6370 => x"3f86a087",
          6371 => x"e0700854",
          6372 => x"5481f856",
          6373 => x"86a081f8",
          6374 => x"73770684",
          6375 => x"07545572",
          6376 => x"75347308",
          6377 => x"7080ff06",
          6378 => x"80c00751",
          6379 => x"53727534",
          6380 => x"86a087cc",
          6381 => x"08707706",
          6382 => x"81075153",
          6383 => x"7286a081",
          6384 => x"f3347308",
          6385 => x"81f70688",
          6386 => x"07537275",
          6387 => x"3480d00b",
          6388 => x"84b6d834",
          6389 => x"800b84b8",
          6390 => x"e40c873d",
          6391 => x"0d0484b6",
          6392 => x"d83384b8",
          6393 => x"e40c04f7",
          6394 => x"3d0d02af",
          6395 => x"05330284",
          6396 => x"05b30533",
          6397 => x"84b6d733",
          6398 => x"5b595681",
          6399 => x"53757926",
          6400 => x"82da3884",
          6401 => x"b6d83383",
          6402 => x"f8953383",
          6403 => x"f8943372",
          6404 => x"71291286",
          6405 => x"a7a08011",
          6406 => x"83f89222",
          6407 => x"5f515759",
          6408 => x"717c2905",
          6409 => x"7083ffff",
          6410 => x"0683f6ea",
          6411 => x"33535758",
          6412 => x"5372812e",
          6413 => x"83c43883",
          6414 => x"f8922276",
          6415 => x"05557483",
          6416 => x"f8922383",
          6417 => x"f8943376",
          6418 => x"057081ff",
          6419 => x"067a81ff",
          6420 => x"06555b55",
          6421 => x"727a2682",
          6422 => x"8c38ff19",
          6423 => x"537283f8",
          6424 => x"943483f8",
          6425 => x"92227083",
          6426 => x"ffff0684",
          6427 => x"b6d6335c",
          6428 => x"55577974",
          6429 => x"26828938",
          6430 => x"84b6d833",
          6431 => x"76712954",
          6432 => x"58805472",
          6433 => x"9f9f26ac",
          6434 => x"388497b6",
          6435 => x"70145455",
          6436 => x"e0e01333",
          6437 => x"e0e01634",
          6438 => x"72708105",
          6439 => x"54337570",
          6440 => x"81055734",
          6441 => x"81145484",
          6442 => x"b6d57327",
          6443 => x"e338739f",
          6444 => x"9f26a138",
          6445 => x"83f89033",
          6446 => x"8497b615",
          6447 => x"5455a00b",
          6448 => x"e0e01434",
          6449 => x"74737081",
          6450 => x"05553481",
          6451 => x"14549f9f",
          6452 => x"7427eb38",
          6453 => x"84b6d633",
          6454 => x"ff055675",
          6455 => x"83f89223",
          6456 => x"75577881",
          6457 => x"ff067783",
          6458 => x"ffff0654",
          6459 => x"54737326",
          6460 => x"81fd3872",
          6461 => x"74318105",
          6462 => x"84b6d833",
          6463 => x"71712958",
          6464 => x"55577555",
          6465 => x"86a7a080",
          6466 => x"5886a7b0",
          6467 => x"807981ff",
          6468 => x"067581ff",
          6469 => x"06717129",
          6470 => x"195c5c54",
          6471 => x"57757927",
          6472 => x"b9388497",
          6473 => x"b61654e0",
          6474 => x"e0143353",
          6475 => x"84b6e013",
          6476 => x"33787081",
          6477 => x"055a3473",
          6478 => x"70810555",
          6479 => x"33777081",
          6480 => x"05593481",
          6481 => x"1584b6d8",
          6482 => x"3384b6d7",
          6483 => x"33717129",
          6484 => x"19565c5a",
          6485 => x"55727526",
          6486 => x"ce388053",
          6487 => x"7284b8e4",
          6488 => x"0c8b3d0d",
          6489 => x"047483f8",
          6490 => x"943483f8",
          6491 => x"92227083",
          6492 => x"ffff0684",
          6493 => x"b6d6335c",
          6494 => x"5557737a",
          6495 => x"27fdf938",
          6496 => x"77802efe",
          6497 => x"dd387881",
          6498 => x"ff06ff05",
          6499 => x"83f89433",
          6500 => x"56537275",
          6501 => x"2e098106",
          6502 => x"fec83873",
          6503 => x"76318105",
          6504 => x"84b6d833",
          6505 => x"71712978",
          6506 => x"72291156",
          6507 => x"52595473",
          6508 => x"7327feae",
          6509 => x"3883f890",
          6510 => x"338497b6",
          6511 => x"15747631",
          6512 => x"555656a0",
          6513 => x"0be0e016",
          6514 => x"34757570",
          6515 => x"81055734",
          6516 => x"ff135372",
          6517 => x"802efe8a",
          6518 => x"38a00be0",
          6519 => x"e0163475",
          6520 => x"75708105",
          6521 => x"5734ff13",
          6522 => x"5372d838",
          6523 => x"fdf43980",
          6524 => x"0b84b6d8",
          6525 => x"335556fe",
          6526 => x"893983f8",
          6527 => x"96153359",
          6528 => x"84b6e019",
          6529 => x"33743484",
          6530 => x"b6d73359",
          6531 => x"fca939fc",
          6532 => x"3d0d7602",
          6533 => x"84059f05",
          6534 => x"33535170",
          6535 => x"86269b38",
          6536 => x"70101083",
          6537 => x"c3dc0551",
          6538 => x"70080484",
          6539 => x"b6d83351",
          6540 => x"71712786",
          6541 => x"387183f8",
          6542 => x"9534800b",
          6543 => x"84b8e40c",
          6544 => x"863d0d04",
          6545 => x"800b83f8",
          6546 => x"953483f8",
          6547 => x"94337081",
          6548 => x"ff065452",
          6549 => x"72802ee2",
          6550 => x"38ff1251",
          6551 => x"7083f894",
          6552 => x"34800b84",
          6553 => x"b8e40c86",
          6554 => x"3d0d0483",
          6555 => x"f8943370",
          6556 => x"73317009",
          6557 => x"709f2c72",
          6558 => x"06545553",
          6559 => x"547083f8",
          6560 => x"9434de39",
          6561 => x"83f89433",
          6562 => x"720584b6",
          6563 => x"d733ff11",
          6564 => x"55565170",
          6565 => x"75258338",
          6566 => x"70537283",
          6567 => x"f8943480",
          6568 => x"0b84b8e4",
          6569 => x"0c863d0d",
          6570 => x"0483f895",
          6571 => x"33707331",
          6572 => x"7009709f",
          6573 => x"2c720654",
          6574 => x"56535570",
          6575 => x"83f89534",
          6576 => x"800b84b8",
          6577 => x"e40c863d",
          6578 => x"0d0483f8",
          6579 => x"95337205",
          6580 => x"84b6d833",
          6581 => x"ff115555",
          6582 => x"51707425",
          6583 => x"83387053",
          6584 => x"7283f895",
          6585 => x"34800b84",
          6586 => x"b8e40c86",
          6587 => x"3d0d0480",
          6588 => x"0b83f895",
          6589 => x"3483f894",
          6590 => x"3384b6d7",
          6591 => x"33ff0556",
          6592 => x"52717525",
          6593 => x"feb43881",
          6594 => x"12517083",
          6595 => x"f89434fe",
          6596 => x"d039ff3d",
          6597 => x"0d028f05",
          6598 => x"335170b1",
          6599 => x"26b33870",
          6600 => x"101083c3",
          6601 => x"f8055170",
          6602 => x"080483f8",
          6603 => x"90337080",
          6604 => x"f0067184",
          6605 => x"2b80f006",
          6606 => x"7072842a",
          6607 => x"07515253",
          6608 => x"517180f0",
          6609 => x"2e098106",
          6610 => x"9c3880f2",
          6611 => x"0b83f890",
          6612 => x"34800b84",
          6613 => x"b8e40c83",
          6614 => x"3d0d0483",
          6615 => x"f8903381",
          6616 => x"9f069007",
          6617 => x"517083f8",
          6618 => x"9034800b",
          6619 => x"84b8e40c",
          6620 => x"833d0d04",
          6621 => x"83f89033",
          6622 => x"80f00751",
          6623 => x"7083f890",
          6624 => x"34e83983",
          6625 => x"f8903381",
          6626 => x"fe068607",
          6627 => x"517083f8",
          6628 => x"9034d739",
          6629 => x"80f10b83",
          6630 => x"f8903480",
          6631 => x"0b84b8e4",
          6632 => x"0c833d0d",
          6633 => x"0483f890",
          6634 => x"3381fc06",
          6635 => x"84075170",
          6636 => x"83f89034",
          6637 => x"ffb43983",
          6638 => x"f8903387",
          6639 => x"07517083",
          6640 => x"f89034ff",
          6641 => x"a53983f8",
          6642 => x"903381fd",
          6643 => x"06850751",
          6644 => x"7083f890",
          6645 => x"34ff9339",
          6646 => x"83f89033",
          6647 => x"81fb0683",
          6648 => x"07517083",
          6649 => x"f89034ff",
          6650 => x"813983f8",
          6651 => x"903381f9",
          6652 => x"06810751",
          6653 => x"7083f890",
          6654 => x"34feef39",
          6655 => x"83f89033",
          6656 => x"81f80651",
          6657 => x"7083f890",
          6658 => x"34fedf39",
          6659 => x"83f89033",
          6660 => x"81df0680",
          6661 => x"d0075170",
          6662 => x"83f89034",
          6663 => x"fecc3983",
          6664 => x"f8903381",
          6665 => x"bf06b007",
          6666 => x"517083f8",
          6667 => x"9034feba",
          6668 => x"3983f890",
          6669 => x"3381ef06",
          6670 => x"80e00751",
          6671 => x"7083f890",
          6672 => x"34fea739",
          6673 => x"83f89033",
          6674 => x"81cf0680",
          6675 => x"c0075170",
          6676 => x"83f89034",
          6677 => x"fe943983",
          6678 => x"f8903381",
          6679 => x"af06a007",
          6680 => x"517083f8",
          6681 => x"9034fe82",
          6682 => x"3983f890",
          6683 => x"33818f06",
          6684 => x"517083f8",
          6685 => x"9034fdf2",
          6686 => x"3983f890",
          6687 => x"3381fa06",
          6688 => x"82075170",
          6689 => x"83f89034",
          6690 => x"fde039f3",
          6691 => x"3d0d02bf",
          6692 => x"05330284",
          6693 => x"0580c305",
          6694 => x"3383f894",
          6695 => x"3383f893",
          6696 => x"3383f895",
          6697 => x"3384b6da",
          6698 => x"3343415f",
          6699 => x"5d5b5978",
          6700 => x"822e82a1",
          6701 => x"38788224",
          6702 => x"a5387881",
          6703 => x"2e818238",
          6704 => x"7d84b6da",
          6705 => x"34800b84",
          6706 => x"b6dc347a",
          6707 => x"83f89434",
          6708 => x"7b83f892",
          6709 => x"237c83f8",
          6710 => x"95348f3d",
          6711 => x"0d047883",
          6712 => x"2e098106",
          6713 => x"db38800b",
          6714 => x"84b6da34",
          6715 => x"810b84b6",
          6716 => x"dc34820b",
          6717 => x"83f89434",
          6718 => x"a80b83f8",
          6719 => x"9534820b",
          6720 => x"83f89223",
          6721 => x"795884b6",
          6722 => x"d8335784",
          6723 => x"b6d73356",
          6724 => x"84b6d633",
          6725 => x"557b547c",
          6726 => x"537a5283",
          6727 => x"e2d851ff",
          6728 => x"81e63f7d",
          6729 => x"84b6da34",
          6730 => x"800b84b6",
          6731 => x"dc347a83",
          6732 => x"f894347b",
          6733 => x"83f89223",
          6734 => x"7c83f895",
          6735 => x"348f3d0d",
          6736 => x"04800b84",
          6737 => x"b6da3481",
          6738 => x"0b84b6dc",
          6739 => x"34800b83",
          6740 => x"f89434a8",
          6741 => x"0b83f895",
          6742 => x"34800b83",
          6743 => x"f8922384",
          6744 => x"b7e73358",
          6745 => x"84b7e633",
          6746 => x"5784b7e5",
          6747 => x"33567955",
          6748 => x"7b547c53",
          6749 => x"7a5283e2",
          6750 => x"f451ff81",
          6751 => x"8b3f800b",
          6752 => x"84b7e533",
          6753 => x"5a5a7979",
          6754 => x"27a53879",
          6755 => x"1084b8b8",
          6756 => x"05702253",
          6757 => x"5983e38c",
          6758 => x"51ff80ec",
          6759 => x"3f811a70",
          6760 => x"81ff0684",
          6761 => x"b7e53352",
          6762 => x"5b59787a",
          6763 => x"26dd3883",
          6764 => x"d29451ff",
          6765 => x"80d23f7d",
          6766 => x"84b6da34",
          6767 => x"800b84b6",
          6768 => x"dc347a83",
          6769 => x"f894347b",
          6770 => x"83f89223",
          6771 => x"7c83f895",
          6772 => x"348f3d0d",
          6773 => x"04800b84",
          6774 => x"b6da3481",
          6775 => x"0b84b6dc",
          6776 => x"34810b83",
          6777 => x"f89434a8",
          6778 => x"0b83f895",
          6779 => x"34810b83",
          6780 => x"f8922383",
          6781 => x"f6c851ff",
          6782 => x"92ae3f84",
          6783 => x"b8e40852",
          6784 => x"83e39051",
          6785 => x"ff80813f",
          6786 => x"805983f6",
          6787 => x"c851ff92",
          6788 => x"973f7884",
          6789 => x"b8e40827",
          6790 => x"fda63883",
          6791 => x"f6c81933",
          6792 => x"5283e398",
          6793 => x"51feffe0",
          6794 => x"3f811970",
          6795 => x"81ff065a",
          6796 => x"5ad839f9",
          6797 => x"3d0d7a02",
          6798 => x"8405a705",
          6799 => x"3384b6d8",
          6800 => x"3383f895",
          6801 => x"3383f894",
          6802 => x"33727129",
          6803 => x"1286a7a0",
          6804 => x"801183f8",
          6805 => x"92225351",
          6806 => x"595c717c",
          6807 => x"29057083",
          6808 => x"ffff0683",
          6809 => x"f6ea3352",
          6810 => x"59515557",
          6811 => x"5772812e",
          6812 => x"81e93875",
          6813 => x"892e81f9",
          6814 => x"38758924",
          6815 => x"81b93875",
          6816 => x"812e8385",
          6817 => x"3875882e",
          6818 => x"82d53884",
          6819 => x"b6d83383",
          6820 => x"f8943383",
          6821 => x"f8953372",
          6822 => x"72290555",
          6823 => x"565484b6",
          6824 => x"e0163386",
          6825 => x"a7a08014",
          6826 => x"3484b6d8",
          6827 => x"3383f895",
          6828 => x"3383f892",
          6829 => x"22727129",
          6830 => x"125a5a56",
          6831 => x"537583f8",
          6832 => x"96183483",
          6833 => x"f8943373",
          6834 => x"71291658",
          6835 => x"5483f890",
          6836 => x"3386a7b0",
          6837 => x"80183484",
          6838 => x"b6d83370",
          6839 => x"81ff0683",
          6840 => x"f8922283",
          6841 => x"f8953372",
          6842 => x"72291157",
          6843 => x"5b575557",
          6844 => x"83f89033",
          6845 => x"8497b614",
          6846 => x"34811870",
          6847 => x"81ff0659",
          6848 => x"55737826",
          6849 => x"81993884",
          6850 => x"b6d93358",
          6851 => x"7781ea38",
          6852 => x"ff175372",
          6853 => x"83f89534",
          6854 => x"84b6db33",
          6855 => x"5372802e",
          6856 => x"8c3884b6",
          6857 => x"dc335776",
          6858 => x"802e80fb",
          6859 => x"38800b84",
          6860 => x"b8e40c89",
          6861 => x"3d0d0475",
          6862 => x"8d2e9738",
          6863 => x"758d2480",
          6864 => x"f738758a",
          6865 => x"2e098106",
          6866 => x"fec13881",
          6867 => x"528151f1",
          6868 => x"963f800b",
          6869 => x"83f89534",
          6870 => x"ffbe3983",
          6871 => x"f8961533",
          6872 => x"5384b6e0",
          6873 => x"13337434",
          6874 => x"75892e09",
          6875 => x"8106fe89",
          6876 => x"38805376",
          6877 => x"52a051fd",
          6878 => x"ba3f8113",
          6879 => x"7081ff06",
          6880 => x"54547283",
          6881 => x"26ff9138",
          6882 => x"7652a051",
          6883 => x"fda53f81",
          6884 => x"137081ff",
          6885 => x"06545483",
          6886 => x"7327d838",
          6887 => x"fefa3974",
          6888 => x"83f89534",
          6889 => x"fef23975",
          6890 => x"528351f9",
          6891 => x"de3f800b",
          6892 => x"84b8e40c",
          6893 => x"893d0d04",
          6894 => x"7580ff2e",
          6895 => x"098106fd",
          6896 => x"ca3883f8",
          6897 => x"95337081",
          6898 => x"ff0655ff",
          6899 => x"05537383",
          6900 => x"38735372",
          6901 => x"83f89534",
          6902 => x"7652a051",
          6903 => x"fcd53f83",
          6904 => x"f8953370",
          6905 => x"81ff0655",
          6906 => x"ff055373",
          6907 => x"fea53873",
          6908 => x"537283f8",
          6909 => x"9534fea0",
          6910 => x"39800b83",
          6911 => x"f8953481",
          6912 => x"528151ef",
          6913 => x"e23ffe90",
          6914 => x"39805275",
          6915 => x"51efd83f",
          6916 => x"fe8639e6",
          6917 => x"3d0d0280",
          6918 => x"f3053384",
          6919 => x"b7e00857",
          6920 => x"5975812e",
          6921 => x"81b83875",
          6922 => x"822e8382",
          6923 => x"38788a2e",
          6924 => x"84b53878",
          6925 => x"8a2482d1",
          6926 => x"3878882e",
          6927 => x"84b93878",
          6928 => x"892e888f",
          6929 => x"3884b6d8",
          6930 => x"3383f894",
          6931 => x"3383f895",
          6932 => x"33727229",
          6933 => x"05585e5c",
          6934 => x"84b6e019",
          6935 => x"3386a7a0",
          6936 => x"80173484",
          6937 => x"b6d83383",
          6938 => x"f8953383",
          6939 => x"f8922272",
          6940 => x"7129125a",
          6941 => x"5a424078",
          6942 => x"83f89618",
          6943 => x"3483f894",
          6944 => x"33607129",
          6945 => x"6205405a",
          6946 => x"83f89033",
          6947 => x"7f86a7b0",
          6948 => x"80053484",
          6949 => x"b6d83370",
          6950 => x"81ff0683",
          6951 => x"f8922283",
          6952 => x"f8953372",
          6953 => x"72291142",
          6954 => x"405d5859",
          6955 => x"83f89033",
          6956 => x"8497b61f",
          6957 => x"34811d70",
          6958 => x"81ff0642",
          6959 => x"58766126",
          6960 => x"81b83884",
          6961 => x"b6d9335a",
          6962 => x"7986f138",
          6963 => x"ff195675",
          6964 => x"83f89534",
          6965 => x"800b84b8",
          6966 => x"e40c9c3d",
          6967 => x"0d0478b7",
          6968 => x"2e848a38",
          6969 => x"b7792581",
          6970 => x"fd3878b8",
          6971 => x"2e9bb338",
          6972 => x"7880db2e",
          6973 => x"89cc3880",
          6974 => x"0b84b7e0",
          6975 => x"0c84b6d8",
          6976 => x"3383f894",
          6977 => x"3383f895",
          6978 => x"33727229",
          6979 => x"055e4040",
          6980 => x"84b6e019",
          6981 => x"3386a7a0",
          6982 => x"801d3484",
          6983 => x"b6d83383",
          6984 => x"f8953383",
          6985 => x"f8922272",
          6986 => x"71291241",
          6987 => x"5f595678",
          6988 => x"83f8961f",
          6989 => x"3483f894",
          6990 => x"33767129",
          6991 => x"195b5783",
          6992 => x"f8903386",
          6993 => x"a7b0801b",
          6994 => x"3484b6d8",
          6995 => x"337081ff",
          6996 => x"0683f892",
          6997 => x"2283f895",
          6998 => x"33727229",
          6999 => x"11444243",
          7000 => x"585983f8",
          7001 => x"90336084",
          7002 => x"97b60534",
          7003 => x"811f5877",
          7004 => x"81ff0641",
          7005 => x"607727fe",
          7006 => x"ca387783",
          7007 => x"f8953480",
          7008 => x"0b84b8e4",
          7009 => x"0c9c3d0d",
          7010 => x"04789b2e",
          7011 => x"82b73878",
          7012 => x"9b248381",
          7013 => x"38788d2e",
          7014 => x"098106fd",
          7015 => x"a838800b",
          7016 => x"83f89534",
          7017 => x"800b84b8",
          7018 => x"e40c9c3d",
          7019 => x"0d04789b",
          7020 => x"2e82aa38",
          7021 => x"d0195675",
          7022 => x"892684d0",
          7023 => x"3884b7e4",
          7024 => x"33811159",
          7025 => x"577784b7",
          7026 => x"e4347884",
          7027 => x"b7e81834",
          7028 => x"7781ff06",
          7029 => x"59800b84",
          7030 => x"b7e81a34",
          7031 => x"800b84b8",
          7032 => x"e40c9c3d",
          7033 => x"0d04789b",
          7034 => x"2efde938",
          7035 => x"800b84b7",
          7036 => x"e00c84b6",
          7037 => x"d83383f8",
          7038 => x"943383f8",
          7039 => x"95337272",
          7040 => x"29055e40",
          7041 => x"4084b6e0",
          7042 => x"193386a7",
          7043 => x"a0801d34",
          7044 => x"84b6d833",
          7045 => x"83f89533",
          7046 => x"83f89222",
          7047 => x"72712912",
          7048 => x"415f5956",
          7049 => x"7883f896",
          7050 => x"1f3483f8",
          7051 => x"94337671",
          7052 => x"29195b57",
          7053 => x"83f89033",
          7054 => x"86a7b080",
          7055 => x"1b3484b6",
          7056 => x"d8337081",
          7057 => x"ff0683f8",
          7058 => x"922283f8",
          7059 => x"95337272",
          7060 => x"29114442",
          7061 => x"43585983",
          7062 => x"f8903360",
          7063 => x"8497b605",
          7064 => x"34811f58",
          7065 => x"fe893981",
          7066 => x"528151ea",
          7067 => x"fa3f800b",
          7068 => x"83f89534",
          7069 => x"feae3984",
          7070 => x"b6d83383",
          7071 => x"f8953370",
          7072 => x"81ff0683",
          7073 => x"f8943373",
          7074 => x"71291286",
          7075 => x"a7a08005",
          7076 => x"83f89222",
          7077 => x"40515d72",
          7078 => x"7e290570",
          7079 => x"83ffff06",
          7080 => x"83f6ea33",
          7081 => x"5a51595a",
          7082 => x"5c75812e",
          7083 => x"86a43878",
          7084 => x"81ff06ff",
          7085 => x"1a575776",
          7086 => x"fc953876",
          7087 => x"567583f8",
          7088 => x"9534fc90",
          7089 => x"39800b84",
          7090 => x"b7e43480",
          7091 => x"0b84b7e5",
          7092 => x"34800b84",
          7093 => x"b7e63480",
          7094 => x"0b84b7e7",
          7095 => x"34810b84",
          7096 => x"b7e00c80",
          7097 => x"0b84b8e4",
          7098 => x"0c9c3d0d",
          7099 => x"0483f894",
          7100 => x"3384b8cc",
          7101 => x"3483f895",
          7102 => x"3384b8cd",
          7103 => x"3483f893",
          7104 => x"3384b8ce",
          7105 => x"34800b84",
          7106 => x"b7e00c80",
          7107 => x"0b84b8e4",
          7108 => x"0c9c3d0d",
          7109 => x"047880ff",
          7110 => x"2e098106",
          7111 => x"faa73883",
          7112 => x"f8943384",
          7113 => x"b6d83370",
          7114 => x"81ff0683",
          7115 => x"f8953370",
          7116 => x"81ff0672",
          7117 => x"75291186",
          7118 => x"a7a08005",
          7119 => x"83f89222",
          7120 => x"5c40727b",
          7121 => x"29057083",
          7122 => x"ffff0683",
          7123 => x"f6ea3344",
          7124 => x"5c435c42",
          7125 => x"5b5c7d81",
          7126 => x"2e85fe38",
          7127 => x"7881ff06",
          7128 => x"ff1a5856",
          7129 => x"75833875",
          7130 => x"577683f8",
          7131 => x"95347b81",
          7132 => x"ff067a81",
          7133 => x"ff067881",
          7134 => x"ff067272",
          7135 => x"29055f40",
          7136 => x"5b84b780",
          7137 => x"3386a7a0",
          7138 => x"801e3484",
          7139 => x"b6d83383",
          7140 => x"f8953383",
          7141 => x"f8922272",
          7142 => x"7129125a",
          7143 => x"5e4240a0",
          7144 => x"0b83f896",
          7145 => x"183483f8",
          7146 => x"94336071",
          7147 => x"2962055a",
          7148 => x"5683f890",
          7149 => x"3386a7b0",
          7150 => x"801a3484",
          7151 => x"b6d83370",
          7152 => x"81ff0683",
          7153 => x"f8922283",
          7154 => x"f8953372",
          7155 => x"72291143",
          7156 => x"5d5a5e59",
          7157 => x"83f89033",
          7158 => x"7f8497b6",
          7159 => x"0534811a",
          7160 => x"7081ff06",
          7161 => x"5c587c7b",
          7162 => x"2695ea38",
          7163 => x"84b6d933",
          7164 => x"5a7996d0",
          7165 => x"38ff1958",
          7166 => x"7783f895",
          7167 => x"3483f895",
          7168 => x"337081ff",
          7169 => x"0658ff05",
          7170 => x"56fdac39",
          7171 => x"78bb2e95",
          7172 => x"d83878bd",
          7173 => x"2e83d738",
          7174 => x"78bf2e95",
          7175 => x"a83884b7",
          7176 => x"e4335f7e",
          7177 => x"83f938ff",
          7178 => x"bf195675",
          7179 => x"b42684c8",
          7180 => x"38751010",
          7181 => x"83c5c005",
          7182 => x"58770804",
          7183 => x"800b83f8",
          7184 => x"95348052",
          7185 => x"8151e79f",
          7186 => x"3f800b84",
          7187 => x"b8e40c9c",
          7188 => x"3d0d0483",
          7189 => x"f8943384",
          7190 => x"b6d83370",
          7191 => x"81ff0683",
          7192 => x"f8953370",
          7193 => x"81ff0672",
          7194 => x"75291186",
          7195 => x"a7a08005",
          7196 => x"83f89222",
          7197 => x"5c41727b",
          7198 => x"29057083",
          7199 => x"ffff0683",
          7200 => x"f6ea3346",
          7201 => x"53455c59",
          7202 => x"5b5b7f81",
          7203 => x"2e82ef38",
          7204 => x"805c7a81",
          7205 => x"ff067a81",
          7206 => x"ff067a81",
          7207 => x"ff067272",
          7208 => x"29055c58",
          7209 => x"4084b780",
          7210 => x"3386a7a0",
          7211 => x"801b3484",
          7212 => x"b6d83383",
          7213 => x"f8953383",
          7214 => x"f8922272",
          7215 => x"7129125e",
          7216 => x"415e56a0",
          7217 => x"0b83f896",
          7218 => x"1c3483f8",
          7219 => x"94337671",
          7220 => x"291e5a5e",
          7221 => x"83f89033",
          7222 => x"86a7b080",
          7223 => x"1a3484b6",
          7224 => x"d8337081",
          7225 => x"ff0683f8",
          7226 => x"922283f8",
          7227 => x"95337272",
          7228 => x"29115b44",
          7229 => x"5a405983",
          7230 => x"f8903384",
          7231 => x"97b61834",
          7232 => x"60810570",
          7233 => x"81ff065b",
          7234 => x"587e7a26",
          7235 => x"81ac3884",
          7236 => x"b6d93358",
          7237 => x"7792fb38",
          7238 => x"ff195675",
          7239 => x"83f89534",
          7240 => x"811c7081",
          7241 => x"ff065d59",
          7242 => x"7b8326f7",
          7243 => x"a73883f8",
          7244 => x"943384b6",
          7245 => x"d83383f8",
          7246 => x"95337281",
          7247 => x"ff067281",
          7248 => x"ff067281",
          7249 => x"ff067272",
          7250 => x"2905545b",
          7251 => x"435b5b5b",
          7252 => x"84b78033",
          7253 => x"86a7a080",
          7254 => x"1b3484b6",
          7255 => x"d83383f8",
          7256 => x"953383f8",
          7257 => x"92227271",
          7258 => x"29125e41",
          7259 => x"5e56a00b",
          7260 => x"83f8961c",
          7261 => x"3483f894",
          7262 => x"33767129",
          7263 => x"1e5a5e83",
          7264 => x"f8903386",
          7265 => x"a7b0801a",
          7266 => x"3484b6d8",
          7267 => x"337081ff",
          7268 => x"0683f892",
          7269 => x"2283f895",
          7270 => x"33727229",
          7271 => x"115b445a",
          7272 => x"405983f8",
          7273 => x"90338497",
          7274 => x"b6183460",
          7275 => x"81057081",
          7276 => x"ff065b58",
          7277 => x"797f27fe",
          7278 => x"d6387783",
          7279 => x"f89534fe",
          7280 => x"df39820b",
          7281 => x"84b7e00c",
          7282 => x"800b84b8",
          7283 => x"e40c9c3d",
          7284 => x"0d0483f8",
          7285 => x"96173359",
          7286 => x"84b6e019",
          7287 => x"337a3483",
          7288 => x"f8953370",
          7289 => x"81ff0658",
          7290 => x"ff0556f9",
          7291 => x"ca39810b",
          7292 => x"84b7e634",
          7293 => x"800b84b8",
          7294 => x"e40c9c3d",
          7295 => x"0d0483f8",
          7296 => x"9617335b",
          7297 => x"84b6e01b",
          7298 => x"337c3483",
          7299 => x"f8943384",
          7300 => x"b6d83383",
          7301 => x"f895335b",
          7302 => x"5b5b805c",
          7303 => x"fcf43984",
          7304 => x"b7e8429c",
          7305 => x"3ddc1153",
          7306 => x"d80551ff",
          7307 => x"8ad83f84",
          7308 => x"b8e40880",
          7309 => x"2efbf038",
          7310 => x"84b7e533",
          7311 => x"8111575a",
          7312 => x"7584b7e5",
          7313 => x"34791083",
          7314 => x"fe064102",
          7315 => x"80ca0522",
          7316 => x"6184b8b8",
          7317 => x"0523fbcf",
          7318 => x"3983f896",
          7319 => x"17335c84",
          7320 => x"b6e01c33",
          7321 => x"7b3483f8",
          7322 => x"943384b6",
          7323 => x"d83383f8",
          7324 => x"95335b5b",
          7325 => x"5cf9e539",
          7326 => x"84b6d833",
          7327 => x"83f89433",
          7328 => x"83f89533",
          7329 => x"72722905",
          7330 => x"415d5b84",
          7331 => x"b6e01933",
          7332 => x"7f86a7a0",
          7333 => x"80053484",
          7334 => x"b6d83383",
          7335 => x"f8953383",
          7336 => x"f8922272",
          7337 => x"7129125a",
          7338 => x"435b5678",
          7339 => x"83f89618",
          7340 => x"3483f894",
          7341 => x"33767129",
          7342 => x"1b415e83",
          7343 => x"f8903360",
          7344 => x"86a7b080",
          7345 => x"053484b6",
          7346 => x"d8337081",
          7347 => x"ff0683f8",
          7348 => x"922283f8",
          7349 => x"95337272",
          7350 => x"2911415f",
          7351 => x"5a425a83",
          7352 => x"f8903384",
          7353 => x"97b61e34",
          7354 => x"811c7081",
          7355 => x"ff065c58",
          7356 => x"607b2690",
          7357 => x"a23884b6",
          7358 => x"d9335877",
          7359 => x"90e238ff",
          7360 => x"1a567583",
          7361 => x"f8953480",
          7362 => x"0b84b7e0",
          7363 => x"0c84b6db",
          7364 => x"33407f80",
          7365 => x"2ef3bd38",
          7366 => x"84b6dc33",
          7367 => x"5675f3b4",
          7368 => x"38785281",
          7369 => x"51eae43f",
          7370 => x"800b84b8",
          7371 => x"e40c9c3d",
          7372 => x"0d0484b8",
          7373 => x"cc3383f8",
          7374 => x"943484b8",
          7375 => x"cd3383f8",
          7376 => x"953484b8",
          7377 => x"ce335776",
          7378 => x"83f89223",
          7379 => x"ffb93983",
          7380 => x"f8943384",
          7381 => x"b8cc3483",
          7382 => x"f8953384",
          7383 => x"b8cd3483",
          7384 => x"f8933384",
          7385 => x"b8ce34ff",
          7386 => x"9e3984b7",
          7387 => x"e5335b7a",
          7388 => x"802eff93",
          7389 => x"3884b8b8",
          7390 => x"225d7c86",
          7391 => x"2e098106",
          7392 => x"ff853883",
          7393 => x"f8953381",
          7394 => x"055583f8",
          7395 => x"94338105",
          7396 => x"549b5383",
          7397 => x"e3a05294",
          7398 => x"3d705257",
          7399 => x"feee893f",
          7400 => x"7651feff",
          7401 => x"833f84b8",
          7402 => x"e40881ff",
          7403 => x"0683f6e8",
          7404 => x"33577605",
          7405 => x"4160a024",
          7406 => x"fecd3876",
          7407 => x"5283f6c8",
          7408 => x"51fefdce",
          7409 => x"3ffec039",
          7410 => x"800b84b7",
          7411 => x"e5335b58",
          7412 => x"7981ff06",
          7413 => x"5b777b27",
          7414 => x"fead3877",
          7415 => x"1084b8b8",
          7416 => x"05811133",
          7417 => x"574175b1",
          7418 => x"268aa538",
          7419 => x"75101083",
          7420 => x"c794055f",
          7421 => x"7e080484",
          7422 => x"b7e5335e",
          7423 => x"7d802e8f",
          7424 => x"a43883f8",
          7425 => x"943384b8",
          7426 => x"b9337171",
          7427 => x"31700970",
          7428 => x"9f2c7206",
          7429 => x"5a42595e",
          7430 => x"5c7583f8",
          7431 => x"9434fde7",
          7432 => x"3984b7e5",
          7433 => x"33567580",
          7434 => x"2e8ee738",
          7435 => x"84b8b933",
          7436 => x"ff057081",
          7437 => x"ff0684b6",
          7438 => x"d8335d57",
          7439 => x"5f757b27",
          7440 => x"fdc53875",
          7441 => x"83f89534",
          7442 => x"fdbd3980",
          7443 => x"0b83f895",
          7444 => x"3483f894",
          7445 => x"337081ff",
          7446 => x"065d577b",
          7447 => x"802efda7",
          7448 => x"38ff1756",
          7449 => x"7583f894",
          7450 => x"34fd9c39",
          7451 => x"800b83f8",
          7452 => x"953483f8",
          7453 => x"943384b6",
          7454 => x"d733ff05",
          7455 => x"57577676",
          7456 => x"25fd8438",
          7457 => x"81175675",
          7458 => x"83f89434",
          7459 => x"fcf93984",
          7460 => x"b7e53340",
          7461 => x"7f802e8d",
          7462 => x"e03883f8",
          7463 => x"953384b8",
          7464 => x"b9337171",
          7465 => x"31700970",
          7466 => x"9f2c7206",
          7467 => x"5a415942",
          7468 => x"5a7583f8",
          7469 => x"9534fccf",
          7470 => x"3984b7e5",
          7471 => x"335b7a80",
          7472 => x"2efcc438",
          7473 => x"84b8b822",
          7474 => x"4160992e",
          7475 => x"098106fc",
          7476 => x"b63884b6",
          7477 => x"d83383f8",
          7478 => x"953383f8",
          7479 => x"94337271",
          7480 => x"291286a7",
          7481 => x"a0801183",
          7482 => x"f8922243",
          7483 => x"515a5871",
          7484 => x"60290570",
          7485 => x"83ffff06",
          7486 => x"83f6e808",
          7487 => x"87fffe80",
          7488 => x"06425a5d",
          7489 => x"5d7e8482",
          7490 => x"802e92bf",
          7491 => x"38800b83",
          7492 => x"f6e934fb",
          7493 => x"f23984b7",
          7494 => x"e5335a79",
          7495 => x"802efbe7",
          7496 => x"3884b8b8",
          7497 => x"22587799",
          7498 => x"2e098106",
          7499 => x"fbd93881",
          7500 => x"0b83f6e9",
          7501 => x"34fbd039",
          7502 => x"84b7e533",
          7503 => x"5675802e",
          7504 => x"90be3884",
          7505 => x"b8b93383",
          7506 => x"f895335d",
          7507 => x"7c0584b6",
          7508 => x"d833ff11",
          7509 => x"595e5675",
          7510 => x"7d258338",
          7511 => x"75577683",
          7512 => x"f89534fb",
          7513 => x"a23984b7",
          7514 => x"e5335776",
          7515 => x"802e8cc8",
          7516 => x"3884b8b9",
          7517 => x"3383f894",
          7518 => x"33426105",
          7519 => x"84b6d733",
          7520 => x"ff115941",
          7521 => x"56756025",
          7522 => x"83387557",
          7523 => x"7683f894",
          7524 => x"34faf439",
          7525 => x"83e3ac51",
          7526 => x"fee8ed3f",
          7527 => x"800b84b7",
          7528 => x"e5335757",
          7529 => x"7676278b",
          7530 => x"c7387610",
          7531 => x"84b8b805",
          7532 => x"7022535a",
          7533 => x"83e38c51",
          7534 => x"fee8cd3f",
          7535 => x"81177081",
          7536 => x"ff0684b7",
          7537 => x"e5335858",
          7538 => x"58da3982",
          7539 => x"0b84b7e5",
          7540 => x"335f577d",
          7541 => x"802e8d38",
          7542 => x"84b8b822",
          7543 => x"56758326",
          7544 => x"83387557",
          7545 => x"81527681",
          7546 => x"ff0651d5",
          7547 => x"f33ffa97",
          7548 => x"3984b7e5",
          7549 => x"33578177",
          7550 => x"278eb738",
          7551 => x"84b8bb33",
          7552 => x"ff057081",
          7553 => x"ff0684b8",
          7554 => x"b933ff05",
          7555 => x"7081ff06",
          7556 => x"84b6d733",
          7557 => x"7081ff06",
          7558 => x"ff114043",
          7559 => x"525b595c",
          7560 => x"5c777e27",
          7561 => x"8338775a",
          7562 => x"7983f892",
          7563 => x"237681ff",
          7564 => x"06ff1858",
          7565 => x"5f777f27",
          7566 => x"83387757",
          7567 => x"7683f894",
          7568 => x"3484b6d8",
          7569 => x"33ff1157",
          7570 => x"407a6027",
          7571 => x"f9b4387a",
          7572 => x"567583f8",
          7573 => x"9534f9af",
          7574 => x"3984b7e5",
          7575 => x"335f7e80",
          7576 => x"2e8aef38",
          7577 => x"84b8b933",
          7578 => x"84b6d733",
          7579 => x"405b7a7f",
          7580 => x"26f99438",
          7581 => x"83f89433",
          7582 => x"84b6d833",
          7583 => x"7081ff06",
          7584 => x"83f89533",
          7585 => x"71742911",
          7586 => x"86a7a080",
          7587 => x"0583f892",
          7588 => x"225f4071",
          7589 => x"7e290570",
          7590 => x"83ffff06",
          7591 => x"83f6ea33",
          7592 => x"46525959",
          7593 => x"5f5d6081",
          7594 => x"2e84f038",
          7595 => x"7983ffff",
          7596 => x"06707c31",
          7597 => x"5d57807c",
          7598 => x"248efe38",
          7599 => x"84b6d733",
          7600 => x"56767627",
          7601 => x"8ed638ff",
          7602 => x"16567583",
          7603 => x"f892237c",
          7604 => x"81ff0670",
          7605 => x"7c314157",
          7606 => x"8060248e",
          7607 => x"e53884b6",
          7608 => x"d7335676",
          7609 => x"76278dee",
          7610 => x"38ff1656",
          7611 => x"7583f894",
          7612 => x"347e81ff",
          7613 => x"0683f892",
          7614 => x"22575780",
          7615 => x"5a767626",
          7616 => x"90387577",
          7617 => x"3181057e",
          7618 => x"81ff0671",
          7619 => x"71295c5e",
          7620 => x"5b795886",
          7621 => x"a7a0805b",
          7622 => x"86a7b080",
          7623 => x"7f81ff06",
          7624 => x"7f81ff06",
          7625 => x"7171291d",
          7626 => x"4258425c",
          7627 => x"797f27f7",
          7628 => x"d6388497",
          7629 => x"b61a57e0",
          7630 => x"e017335f",
          7631 => x"84b6e01f",
          7632 => x"337b7081",
          7633 => x"055d3476",
          7634 => x"70810558",
          7635 => x"337c7081",
          7636 => x"055e3481",
          7637 => x"1884b6d8",
          7638 => x"3384b6d7",
          7639 => x"33717129",
          7640 => x"1d43405e",
          7641 => x"58776027",
          7642 => x"f79d38e0",
          7643 => x"e017335f",
          7644 => x"84b6e01f",
          7645 => x"337b7081",
          7646 => x"055d3476",
          7647 => x"70810558",
          7648 => x"337c7081",
          7649 => x"055e3481",
          7650 => x"1884b6d8",
          7651 => x"3384b6d7",
          7652 => x"33717129",
          7653 => x"1d43405e",
          7654 => x"587f7826",
          7655 => x"ff9938f6",
          7656 => x"e63984b7",
          7657 => x"e5335675",
          7658 => x"802e87e0",
          7659 => x"38805284",
          7660 => x"b8b93351",
          7661 => x"d8b13ff6",
          7662 => x"ce39800b",
          7663 => x"84b6d833",
          7664 => x"ff1184b7",
          7665 => x"e5335d59",
          7666 => x"40587978",
          7667 => x"2e943884",
          7668 => x"b8b82256",
          7669 => x"75782e09",
          7670 => x"81068bbe",
          7671 => x"3883f895",
          7672 => x"33587681",
          7673 => x"ff0683f8",
          7674 => x"94337943",
          7675 => x"5c5c76ff",
          7676 => x"2e81ed38",
          7677 => x"84b6d733",
          7678 => x"407a6026",
          7679 => x"f689387e",
          7680 => x"81ff0656",
          7681 => x"607626f5",
          7682 => x"fe387b76",
          7683 => x"26617d27",
          7684 => x"075776f5",
          7685 => x"f2387a10",
          7686 => x"101b7090",
          7687 => x"29620586",
          7688 => x"a7a08011",
          7689 => x"701f5d5a",
          7690 => x"86a7b080",
          7691 => x"05798306",
          7692 => x"58515d75",
          7693 => x"8bac3879",
          7694 => x"83065776",
          7695 => x"8ba43883",
          7696 => x"f8903370",
          7697 => x"982b7190",
          7698 => x"2b077188",
          7699 => x"2b077107",
          7700 => x"797f5952",
          7701 => x"5f57777a",
          7702 => x"279e3880",
          7703 => x"77708405",
          7704 => x"590c7d76",
          7705 => x"70840558",
          7706 => x"0c797726",
          7707 => x"ee3884b6",
          7708 => x"d83384b6",
          7709 => x"d733415f",
          7710 => x"7e81ff06",
          7711 => x"6081ff06",
          7712 => x"83f89222",
          7713 => x"7d732964",
          7714 => x"05595959",
          7715 => x"5a777726",
          7716 => x"8c387678",
          7717 => x"311b707b",
          7718 => x"29620557",
          7719 => x"4075761d",
          7720 => x"57577676",
          7721 => x"26f4e038",
          7722 => x"83f89033",
          7723 => x"8497b618",
          7724 => x"595aa00b",
          7725 => x"e0e01934",
          7726 => x"79787081",
          7727 => x"055a3481",
          7728 => x"17577676",
          7729 => x"26f4c038",
          7730 => x"a00be0e0",
          7731 => x"19347978",
          7732 => x"7081055a",
          7733 => x"34811757",
          7734 => x"757727d6",
          7735 => x"38f4a839",
          7736 => x"ff1f7081",
          7737 => x"ff065d58",
          7738 => x"fe8a3983",
          7739 => x"f8903370",
          7740 => x"80f00671",
          7741 => x"842b80f0",
          7742 => x"0671842a",
          7743 => x"07585d57",
          7744 => x"7b80f02e",
          7745 => x"098106be",
          7746 => x"3880f20b",
          7747 => x"83f89034",
          7748 => x"81187081",
          7749 => x"ff065956",
          7750 => x"f5b63983",
          7751 => x"f8961733",
          7752 => x"5e84b6e0",
          7753 => x"1e337c34",
          7754 => x"83f89433",
          7755 => x"84b6d833",
          7756 => x"83f89222",
          7757 => x"84b6d733",
          7758 => x"425c5f5d",
          7759 => x"faee3983",
          7760 => x"f8903387",
          7761 => x"07567583",
          7762 => x"f8903481",
          7763 => x"187081ff",
          7764 => x"065956f4",
          7765 => x"fb3983f8",
          7766 => x"903381fd",
          7767 => x"06850756",
          7768 => x"7583f890",
          7769 => x"34e53983",
          7770 => x"f8903381",
          7771 => x"fb068307",
          7772 => x"567583f8",
          7773 => x"9034d439",
          7774 => x"83f89033",
          7775 => x"81f90681",
          7776 => x"07567583",
          7777 => x"f89034c3",
          7778 => x"3983f890",
          7779 => x"33819f06",
          7780 => x"90075675",
          7781 => x"83f89034",
          7782 => x"ffb13980",
          7783 => x"f10b83f8",
          7784 => x"90348118",
          7785 => x"7081ff06",
          7786 => x"5956f4a4",
          7787 => x"3983f890",
          7788 => x"33818f06",
          7789 => x"567583f8",
          7790 => x"9034ff8f",
          7791 => x"3983f890",
          7792 => x"33819f06",
          7793 => x"90075675",
          7794 => x"83f89034",
          7795 => x"fefd3983",
          7796 => x"f8903381",
          7797 => x"ef0680e0",
          7798 => x"07567583",
          7799 => x"f89034fe",
          7800 => x"ea3983f8",
          7801 => x"903381cf",
          7802 => x"0680c007",
          7803 => x"567583f8",
          7804 => x"9034fed7",
          7805 => x"3983f890",
          7806 => x"3381af06",
          7807 => x"a0075675",
          7808 => x"83f89034",
          7809 => x"fec53983",
          7810 => x"f8903381",
          7811 => x"fe068607",
          7812 => x"567583f8",
          7813 => x"9034feb3",
          7814 => x"3983f890",
          7815 => x"3381fc06",
          7816 => x"84075675",
          7817 => x"83f89034",
          7818 => x"fea13983",
          7819 => x"f8903381",
          7820 => x"fa068207",
          7821 => x"567583f8",
          7822 => x"9034fe8f",
          7823 => x"3983f890",
          7824 => x"3381f806",
          7825 => x"567583f8",
          7826 => x"9034fdff",
          7827 => x"3983f890",
          7828 => x"3380f007",
          7829 => x"567583f8",
          7830 => x"9034fdef",
          7831 => x"3983f890",
          7832 => x"3380f007",
          7833 => x"567583f8",
          7834 => x"9034fddf",
          7835 => x"3983f890",
          7836 => x"3381df06",
          7837 => x"80d00756",
          7838 => x"7583f890",
          7839 => x"34fdcc39",
          7840 => x"83f89033",
          7841 => x"81bf06b0",
          7842 => x"07567583",
          7843 => x"f89034fd",
          7844 => x"ba39800b",
          7845 => x"83f89534",
          7846 => x"80528151",
          7847 => x"d2c93fec",
          7848 => x"ff3984b8",
          7849 => x"cc3383f8",
          7850 => x"943484b8",
          7851 => x"cd3383f8",
          7852 => x"953484b8",
          7853 => x"ce335978",
          7854 => x"83f89223",
          7855 => x"800b84b7",
          7856 => x"e00ce8c7",
          7857 => x"39810b84",
          7858 => x"b7e73480",
          7859 => x"0b84b8e4",
          7860 => x"0c9c3d0d",
          7861 => x"047783f8",
          7862 => x"953483f8",
          7863 => x"95337081",
          7864 => x"ff0658ff",
          7865 => x"0556e7cf",
          7866 => x"3984b7e8",
          7867 => x"429c3ddc",
          7868 => x"1153d805",
          7869 => x"51fef98e",
          7870 => x"3f84b8e4",
          7871 => x"08a13884",
          7872 => x"b8e40884",
          7873 => x"b7e00c80",
          7874 => x"0b84b7e4",
          7875 => x"34800b84",
          7876 => x"b8e40c9c",
          7877 => x"3d0d0477",
          7878 => x"83f89534",
          7879 => x"efe93984",
          7880 => x"b7e53381",
          7881 => x"115c5c7a",
          7882 => x"84b7e534",
          7883 => x"7b1083fe",
          7884 => x"065d0280",
          7885 => x"ca052284",
          7886 => x"b8b81e23",
          7887 => x"800b84b7",
          7888 => x"e434ca39",
          7889 => x"800b83f8",
          7890 => x"95348052",
          7891 => x"8151d197",
          7892 => x"3f83f895",
          7893 => x"337081ff",
          7894 => x"0658ff05",
          7895 => x"56e6d839",
          7896 => x"800b83f8",
          7897 => x"95348052",
          7898 => x"8151d0fb",
          7899 => x"3fef9839",
          7900 => x"8a51feeb",
          7901 => x"e93fef8f",
          7902 => x"3983f895",
          7903 => x"33ff0570",
          7904 => x"09709f2c",
          7905 => x"7206585f",
          7906 => x"57f2a639",
          7907 => x"75528151",
          7908 => x"d93984b6",
          7909 => x"d8334075",
          7910 => x"6027eeeb",
          7911 => x"387583f8",
          7912 => x"9534eee3",
          7913 => x"3983f894",
          7914 => x"33ff0570",
          7915 => x"09709f2c",
          7916 => x"72065840",
          7917 => x"57f0e239",
          7918 => x"83f89433",
          7919 => x"810584b6",
          7920 => x"d733ff11",
          7921 => x"59595675",
          7922 => x"7825f3c0",
          7923 => x"387557f3",
          7924 => x"bb3984b6",
          7925 => x"d7337081",
          7926 => x"ff06585c",
          7927 => x"817726ee",
          7928 => x"a63883f8",
          7929 => x"943384b6",
          7930 => x"d8337081",
          7931 => x"ff0683f8",
          7932 => x"95337174",
          7933 => x"291186a7",
          7934 => x"a0800583",
          7935 => x"f892225f",
          7936 => x"5f717e29",
          7937 => x"057083ff",
          7938 => x"ff0683f6",
          7939 => x"ea335d5b",
          7940 => x"44425f5d",
          7941 => x"77812e81",
          7942 => x"f5387983",
          7943 => x"ffff06ff",
          7944 => x"115c5780",
          7945 => x"7b248489",
          7946 => x"3884b6d7",
          7947 => x"33567676",
          7948 => x"27839838",
          7949 => x"ff165675",
          7950 => x"83f89223",
          7951 => x"7c81ff06",
          7952 => x"ff115757",
          7953 => x"80762483",
          7954 => x"df3884b6",
          7955 => x"d7335676",
          7956 => x"762782ec",
          7957 => x"38ff1656",
          7958 => x"7583f894",
          7959 => x"347b81ff",
          7960 => x"0683f892",
          7961 => x"22575780",
          7962 => x"5a767626",
          7963 => x"90387577",
          7964 => x"3181057e",
          7965 => x"81ff0671",
          7966 => x"71295c5e",
          7967 => x"5f795886",
          7968 => x"a7a0805b",
          7969 => x"86a7b080",
          7970 => x"7c81ff06",
          7971 => x"7f81ff06",
          7972 => x"7171291d",
          7973 => x"4142425d",
          7974 => x"797e27ec",
          7975 => x"ea388497",
          7976 => x"b61a57e0",
          7977 => x"e017335e",
          7978 => x"84b6e01e",
          7979 => x"337b7081",
          7980 => x"055d3476",
          7981 => x"70810558",
          7982 => x"337d7081",
          7983 => x"055f3481",
          7984 => x"1884b6d8",
          7985 => x"3384b6d7",
          7986 => x"33717129",
          7987 => x"1d59415d",
          7988 => x"58777627",
          7989 => x"ecb138e0",
          7990 => x"e017335e",
          7991 => x"84b6e01e",
          7992 => x"337b7081",
          7993 => x"055d3476",
          7994 => x"70810558",
          7995 => x"337d7081",
          7996 => x"055f3481",
          7997 => x"1884b6d8",
          7998 => x"3384b6d7",
          7999 => x"33717129",
          8000 => x"1d59415d",
          8001 => x"58757826",
          8002 => x"ff9938eb",
          8003 => x"fa3983f8",
          8004 => x"9617335c",
          8005 => x"84b6e01c",
          8006 => x"337b3483",
          8007 => x"f8943384",
          8008 => x"b6d83383",
          8009 => x"f8922284",
          8010 => x"b6d7335f",
          8011 => x"5c5f5dfd",
          8012 => x"e93976eb",
          8013 => x"d23884b6",
          8014 => x"d7337081",
          8015 => x"ff06ff11",
          8016 => x"5c425876",
          8017 => x"61278338",
          8018 => x"765a7983",
          8019 => x"f8922377",
          8020 => x"81ff06ff",
          8021 => x"19585a80",
          8022 => x"7a278338",
          8023 => x"80577683",
          8024 => x"f8943484",
          8025 => x"b6d83370",
          8026 => x"81ff06ff",
          8027 => x"12525956",
          8028 => x"807827eb",
          8029 => x"8d388056",
          8030 => x"7583f895",
          8031 => x"34eb8839",
          8032 => x"83f89533",
          8033 => x"810584b6",
          8034 => x"d833ff11",
          8035 => x"59405675",
          8036 => x"7f25efca",
          8037 => x"387557ef",
          8038 => x"c5397581",
          8039 => x"2e098106",
          8040 => x"f4c03883",
          8041 => x"f8953370",
          8042 => x"81ff0683",
          8043 => x"f894337a",
          8044 => x"445d5d57",
          8045 => x"76ff2e09",
          8046 => x"8106f4b8",
          8047 => x"38f6a139",
          8048 => x"ff1d5675",
          8049 => x"83f89434",
          8050 => x"fd9339ff",
          8051 => x"1a567583",
          8052 => x"f89223fc",
          8053 => x"e7397c7b",
          8054 => x"31567583",
          8055 => x"f89434f2",
          8056 => x"9039777d",
          8057 => x"5856777a",
          8058 => x"26f58d38",
          8059 => x"80767081",
          8060 => x"05583483",
          8061 => x"f8903377",
          8062 => x"70810559",
          8063 => x"34757a26",
          8064 => x"f4ec3880",
          8065 => x"76708105",
          8066 => x"583483f8",
          8067 => x"90337770",
          8068 => x"81055934",
          8069 => x"797627d4",
          8070 => x"38f4d339",
          8071 => x"797b3156",
          8072 => x"7583f892",
          8073 => x"23f1a839",
          8074 => x"800b83f8",
          8075 => x"9434fcad",
          8076 => x"397e83f8",
          8077 => x"9223fc84",
          8078 => x"39800b83",
          8079 => x"f89223f1",
          8080 => x"8e39800b",
          8081 => x"83f89434",
          8082 => x"f1a73983",
          8083 => x"f8961833",
          8084 => x"5a84b6e0",
          8085 => x"1a337734",
          8086 => x"800b83f6",
          8087 => x"e934e9a7",
          8088 => x"39fd3d0d",
          8089 => x"02970533",
          8090 => x"84b6da33",
          8091 => x"54547280",
          8092 => x"2e903873",
          8093 => x"51db9c3f",
          8094 => x"800b84b8",
          8095 => x"e40c853d",
          8096 => x"0d047652",
          8097 => x"7351d7ab",
          8098 => x"3f800b84",
          8099 => x"b8e40c85",
          8100 => x"3d0d04f3",
          8101 => x"3d0d02bf",
          8102 => x"05335cff",
          8103 => x"0b83f6e8",
          8104 => x"337081ff",
          8105 => x"0683f6c8",
          8106 => x"11335855",
          8107 => x"55597480",
          8108 => x"2e80d638",
          8109 => x"81145675",
          8110 => x"83f6e834",
          8111 => x"74597884",
          8112 => x"b8e40c8f",
          8113 => x"3d0d0483",
          8114 => x"f6c40854",
          8115 => x"82537380",
          8116 => x"2e913873",
          8117 => x"73327030",
          8118 => x"71077009",
          8119 => x"709f2a56",
          8120 => x"5d5e5872",
          8121 => x"83f6c40c",
          8122 => x"ff598054",
          8123 => x"7b812e09",
          8124 => x"81068338",
          8125 => x"7b547b83",
          8126 => x"32703070",
          8127 => x"80257607",
          8128 => x"5c5c5d79",
          8129 => x"802e85c4",
          8130 => x"3884b6d8",
          8131 => x"3383f895",
          8132 => x"3383f894",
          8133 => x"33727129",
          8134 => x"1286a7a0",
          8135 => x"800583f8",
          8136 => x"92225b59",
          8137 => x"5d717929",
          8138 => x"057083ff",
          8139 => x"ff0683f6",
          8140 => x"e9335859",
          8141 => x"55587481",
          8142 => x"2e838c38",
          8143 => x"81f05473",
          8144 => x"86ee8080",
          8145 => x"34800b87",
          8146 => x"c098880c",
          8147 => x"87c09888",
          8148 => x"08567580",
          8149 => x"2ef63886",
          8150 => x"ee808408",
          8151 => x"577683f4",
          8152 => x"94153481",
          8153 => x"147081ff",
          8154 => x"06555581",
          8155 => x"f97427cf",
          8156 => x"38805483",
          8157 => x"f6841433",
          8158 => x"7081ff06",
          8159 => x"83f68e16",
          8160 => x"33585455",
          8161 => x"72762e85",
          8162 => x"c1387281",
          8163 => x"ff2e86b4",
          8164 => x"387483f6",
          8165 => x"98153475",
          8166 => x"81ff065a",
          8167 => x"7981ff2e",
          8168 => x"85cd3875",
          8169 => x"83f6a215",
          8170 => x"3483f684",
          8171 => x"143383f6",
          8172 => x"8e153481",
          8173 => x"147081ff",
          8174 => x"06555e89",
          8175 => x"7427ffb3",
          8176 => x"3883f68c",
          8177 => x"3370982b",
          8178 => x"70802558",
          8179 => x"56547583",
          8180 => x"f6bc3473",
          8181 => x"81ff0670",
          8182 => x"862a8132",
          8183 => x"70810651",
          8184 => x"54587280",
          8185 => x"2e85e738",
          8186 => x"810b83f6",
          8187 => x"bd347309",
          8188 => x"81065372",
          8189 => x"802e85e4",
          8190 => x"38810b83",
          8191 => x"f6be3480",
          8192 => x"0b83f6bd",
          8193 => x"3383f6c4",
          8194 => x"0883f6be",
          8195 => x"337083f6",
          8196 => x"c03383f6",
          8197 => x"bf335d5d",
          8198 => x"425e5c5e",
          8199 => x"5683f698",
          8200 => x"16335574",
          8201 => x"81ff2e8d",
          8202 => x"3883f6ac",
          8203 => x"16335473",
          8204 => x"802e8282",
          8205 => x"3883f6a2",
          8206 => x"16335372",
          8207 => x"81ff2e8b",
          8208 => x"3883f6ac",
          8209 => x"16335473",
          8210 => x"81ec3874",
          8211 => x"81ff0654",
          8212 => x"7381ff2e",
          8213 => x"8d3883f6",
          8214 => x"ac163353",
          8215 => x"72812e81",
          8216 => x"da387481",
          8217 => x"ff065372",
          8218 => x"81ff2e84",
          8219 => x"8c3883f6",
          8220 => x"ac163354",
          8221 => x"81742784",
          8222 => x"803883f6",
          8223 => x"b80887e8",
          8224 => x"0587c098",
          8225 => x"9c085454",
          8226 => x"73732783",
          8227 => x"ec38810b",
          8228 => x"87c0989c",
          8229 => x"0883f6b8",
          8230 => x"0c588116",
          8231 => x"7081ff06",
          8232 => x"57548976",
          8233 => x"27fef638",
          8234 => x"7683f6bf",
          8235 => x"347783f6",
          8236 => x"c034fe9e",
          8237 => x"1953729c",
          8238 => x"26828b38",
          8239 => x"72101083",
          8240 => x"c8dc055a",
          8241 => x"79080483",
          8242 => x"f6ec0854",
          8243 => x"73802e91",
          8244 => x"3883f414",
          8245 => x"87c0989c",
          8246 => x"085e5e7d",
          8247 => x"7d27fcdc",
          8248 => x"38800b83",
          8249 => x"f6ea3354",
          8250 => x"5472812e",
          8251 => x"83387454",
          8252 => x"7383f6ea",
          8253 => x"3487c098",
          8254 => x"9c0883f6",
          8255 => x"ec0c7381",
          8256 => x"ff065877",
          8257 => x"812e9438",
          8258 => x"83f89617",
          8259 => x"335484b6",
          8260 => x"e0143376",
          8261 => x"3481f054",
          8262 => x"fca53983",
          8263 => x"f6c40853",
          8264 => x"72802e82",
          8265 => x"9c387281",
          8266 => x"2e83f438",
          8267 => x"80c37634",
          8268 => x"81f054fc",
          8269 => x"8a398058",
          8270 => x"fee03980",
          8271 => x"74565783",
          8272 => x"597c812e",
          8273 => x"9b387977",
          8274 => x"2e098106",
          8275 => x"83b4387d",
          8276 => x"812e80ed",
          8277 => x"3879812e",
          8278 => x"80d73879",
          8279 => x"81ff0659",
          8280 => x"87772775",
          8281 => x"982b5454",
          8282 => x"728025a1",
          8283 => x"3873802e",
          8284 => x"9c388117",
          8285 => x"7081ff06",
          8286 => x"761081fe",
          8287 => x"06877227",
          8288 => x"71982b57",
          8289 => x"53575854",
          8290 => x"807324e1",
          8291 => x"38781010",
          8292 => x"10791005",
          8293 => x"7611832b",
          8294 => x"780583f2",
          8295 => x"f4057033",
          8296 => x"5b565478",
          8297 => x"87c0989c",
          8298 => x"0883f6b8",
          8299 => x"0c57fdea",
          8300 => x"3980597d",
          8301 => x"812effa8",
          8302 => x"387981ff",
          8303 => x"0659ffa0",
          8304 => x"398259ff",
          8305 => x"9b3978ff",
          8306 => x"2efa9f38",
          8307 => x"800b84b6",
          8308 => x"da335454",
          8309 => x"72812e83",
          8310 => x"e8387b82",
          8311 => x"32703070",
          8312 => x"80257607",
          8313 => x"4059567d",
          8314 => x"8a387b83",
          8315 => x"2e098106",
          8316 => x"f9cc3878",
          8317 => x"ff2ef9c6",
          8318 => x"38805372",
          8319 => x"10101083",
          8320 => x"f6f00570",
          8321 => x"335d5478",
          8322 => x"7c2e83ba",
          8323 => x"38811370",
          8324 => x"81ff0654",
          8325 => x"57937327",
          8326 => x"e23884b6",
          8327 => x"db335372",
          8328 => x"802ef99a",
          8329 => x"3884b6dc",
          8330 => x"335574f9",
          8331 => x"91387881",
          8332 => x"ff065282",
          8333 => x"51ccd43f",
          8334 => x"7884b8e4",
          8335 => x"0c8f3d0d",
          8336 => x"04be7634",
          8337 => x"81f054f9",
          8338 => x"f6397281",
          8339 => x"ff2e9238",
          8340 => x"83f6ac14",
          8341 => x"3381055b",
          8342 => x"7a83f6ac",
          8343 => x"1534fac9",
          8344 => x"39800b83",
          8345 => x"f6ac1534",
          8346 => x"ff0b83f6",
          8347 => x"981534ff",
          8348 => x"0b83f6a2",
          8349 => x"1534fab1",
          8350 => x"397481ff",
          8351 => x"06537281",
          8352 => x"ff2efc96",
          8353 => x"3883f6ac",
          8354 => x"16335581",
          8355 => x"7527fc8a",
          8356 => x"387781ff",
          8357 => x"06547381",
          8358 => x"2e098106",
          8359 => x"fbfc3883",
          8360 => x"f6b80881",
          8361 => x"fa0587c0",
          8362 => x"989c0854",
          8363 => x"55747327",
          8364 => x"fbe83887",
          8365 => x"c0989c08",
          8366 => x"83f6b80c",
          8367 => x"7681ff06",
          8368 => x"59fbd739",
          8369 => x"ff0b83f6",
          8370 => x"981534f9",
          8371 => x"ca397283",
          8372 => x"f6bd3473",
          8373 => x"09810653",
          8374 => x"72fa9e38",
          8375 => x"7283f6be",
          8376 => x"34800b83",
          8377 => x"f6bd3383",
          8378 => x"f6c40883",
          8379 => x"f6be3370",
          8380 => x"83f6c033",
          8381 => x"83f6bf33",
          8382 => x"5d5d425e",
          8383 => x"5c5e56fa",
          8384 => x"9c397982",
          8385 => x"2e098106",
          8386 => x"fccb387a",
          8387 => x"597a812e",
          8388 => x"fcce3879",
          8389 => x"812e0981",
          8390 => x"06fcc038",
          8391 => x"fd9339ef",
          8392 => x"763481f0",
          8393 => x"54f89839",
          8394 => x"800b84b6",
          8395 => x"db335754",
          8396 => x"75833881",
          8397 => x"547384b6",
          8398 => x"db34ff59",
          8399 => x"f7ac3980",
          8400 => x"0b84b6da",
          8401 => x"33585476",
          8402 => x"83388154",
          8403 => x"7384b6da",
          8404 => x"34ff59f7",
          8405 => x"95398153",
          8406 => x"83f6c408",
          8407 => x"842ef783",
          8408 => x"38840b83",
          8409 => x"f6c40cf6",
          8410 => x"ff3984b6",
          8411 => x"d7337081",
          8412 => x"ff06ff11",
          8413 => x"575a5480",
          8414 => x"79278338",
          8415 => x"80557483",
          8416 => x"f8922373",
          8417 => x"81ff06ff",
          8418 => x"15555380",
          8419 => x"73278338",
          8420 => x"80547383",
          8421 => x"f8943484",
          8422 => x"b6d83370",
          8423 => x"81ff0656",
          8424 => x"ff055380",
          8425 => x"75278338",
          8426 => x"80537283",
          8427 => x"f89534ff",
          8428 => x"59f6b739",
          8429 => x"81528351",
          8430 => x"ffbaa53f",
          8431 => x"ff59f6aa",
          8432 => x"397254fc",
          8433 => x"95398414",
          8434 => x"085283f6",
          8435 => x"c851fede",
          8436 => x"f63f810b",
          8437 => x"83f6e834",
          8438 => x"83f6c833",
          8439 => x"59fcbb39",
          8440 => x"803d0d81",
          8441 => x"51f5ac3f",
          8442 => x"823d0d04",
          8443 => x"fa3d0d80",
          8444 => x"0b83f2f0",
          8445 => x"08535702",
          8446 => x"a3053382",
          8447 => x"133483f2",
          8448 => x"f0085180",
          8449 => x"e0713485",
          8450 => x"0b83f2f0",
          8451 => x"085556fe",
          8452 => x"0b811534",
          8453 => x"800b86f0",
          8454 => x"80e83487",
          8455 => x"c0989c08",
          8456 => x"83f2f008",
          8457 => x"5580ce90",
          8458 => x"055387c0",
          8459 => x"989c0852",
          8460 => x"87c0989c",
          8461 => x"08517072",
          8462 => x"2ef63881",
          8463 => x"143387c0",
          8464 => x"989c0856",
          8465 => x"52747327",
          8466 => x"87387181",
          8467 => x"fe2edb38",
          8468 => x"87c098a4",
          8469 => x"0851ff55",
          8470 => x"70732780",
          8471 => x"c8387155",
          8472 => x"71ff2e80",
          8473 => x"c03887c0",
          8474 => x"989c0880",
          8475 => x"ce900553",
          8476 => x"87c0989c",
          8477 => x"085287c0",
          8478 => x"989c0855",
          8479 => x"74722ef6",
          8480 => x"38811433",
          8481 => x"87c0989c",
          8482 => x"08525270",
          8483 => x"73278738",
          8484 => x"7181ff2e",
          8485 => x"db3887c0",
          8486 => x"98a40855",
          8487 => x"72752683",
          8488 => x"38ff5271",
          8489 => x"55ff1670",
          8490 => x"81ff0657",
          8491 => x"5375802e",
          8492 => x"98387481",
          8493 => x"ff065271",
          8494 => x"fed53874",
          8495 => x"ff2e8a38",
          8496 => x"7684b8e4",
          8497 => x"0c883d0d",
          8498 => x"04810b84",
          8499 => x"b8e40c88",
          8500 => x"3d0d04fa",
          8501 => x"3d0d7902",
          8502 => x"8405a305",
          8503 => x"33565280",
          8504 => x"0b83f2f0",
          8505 => x"0873882b",
          8506 => x"87fc8080",
          8507 => x"06707598",
          8508 => x"2a075155",
          8509 => x"55577183",
          8510 => x"15347290",
          8511 => x"2a517084",
          8512 => x"15347190",
          8513 => x"2a567585",
          8514 => x"15347286",
          8515 => x"153483f2",
          8516 => x"f0085274",
          8517 => x"82133483",
          8518 => x"f2f00851",
          8519 => x"80e17134",
          8520 => x"850b83f2",
          8521 => x"f0085556",
          8522 => x"fe0b8115",
          8523 => x"34800b86",
          8524 => x"f080e834",
          8525 => x"87c0989c",
          8526 => x"0883f2f0",
          8527 => x"085580ce",
          8528 => x"90055387",
          8529 => x"c0989c08",
          8530 => x"5287c098",
          8531 => x"9c085170",
          8532 => x"722ef638",
          8533 => x"81143387",
          8534 => x"c0989c08",
          8535 => x"56527473",
          8536 => x"27873871",
          8537 => x"81fe2edb",
          8538 => x"3887c098",
          8539 => x"a40851ff",
          8540 => x"55707327",
          8541 => x"80c83871",
          8542 => x"5571ff2e",
          8543 => x"80c03887",
          8544 => x"c0989c08",
          8545 => x"80ce9005",
          8546 => x"5387c098",
          8547 => x"9c085287",
          8548 => x"c0989c08",
          8549 => x"5574722e",
          8550 => x"f6388114",
          8551 => x"3387c098",
          8552 => x"9c085252",
          8553 => x"70732787",
          8554 => x"387181ff",
          8555 => x"2edb3887",
          8556 => x"c098a408",
          8557 => x"55727526",
          8558 => x"8338ff52",
          8559 => x"7155ff16",
          8560 => x"7081ff06",
          8561 => x"57537580",
          8562 => x"2e80c738",
          8563 => x"7481ff06",
          8564 => x"5271fed4",
          8565 => x"38745170",
          8566 => x"81ff0656",
          8567 => x"75aa3880",
          8568 => x"c6147b84",
          8569 => x"80115552",
          8570 => x"52707327",
          8571 => x"92387170",
          8572 => x"81055333",
          8573 => x"71708105",
          8574 => x"53347271",
          8575 => x"26f03876",
          8576 => x"84b8e40c",
          8577 => x"883d0d04",
          8578 => x"810b84b8",
          8579 => x"e40c883d",
          8580 => x"0d04ff51",
          8581 => x"c239fa3d",
          8582 => x"0d790284",
          8583 => x"05a30533",
          8584 => x"5656800b",
          8585 => x"83f2f008",
          8586 => x"77882b87",
          8587 => x"fc808006",
          8588 => x"7079982a",
          8589 => x"07515555",
          8590 => x"57758315",
          8591 => x"3472902a",
          8592 => x"51708415",
          8593 => x"3475902a",
          8594 => x"52718515",
          8595 => x"34728615",
          8596 => x"347a83f2",
          8597 => x"f00880c6",
          8598 => x"11848013",
          8599 => x"56545551",
          8600 => x"70732797",
          8601 => x"38707081",
          8602 => x"05523372",
          8603 => x"70810554",
          8604 => x"34727126",
          8605 => x"f03883f2",
          8606 => x"f0085474",
          8607 => x"82153483",
          8608 => x"f2f00855",
          8609 => x"80e27534",
          8610 => x"850b83f2",
          8611 => x"f0085556",
          8612 => x"fe0b8115",
          8613 => x"34800b86",
          8614 => x"f080e834",
          8615 => x"87c0989c",
          8616 => x"0883f2f0",
          8617 => x"085580ce",
          8618 => x"90055387",
          8619 => x"c0989c08",
          8620 => x"5287c098",
          8621 => x"9c085170",
          8622 => x"722ef638",
          8623 => x"81143387",
          8624 => x"c0989c08",
          8625 => x"56527473",
          8626 => x"27873871",
          8627 => x"81fe2edb",
          8628 => x"3887c098",
          8629 => x"a40851ff",
          8630 => x"55707327",
          8631 => x"80c83871",
          8632 => x"5571ff2e",
          8633 => x"80c03887",
          8634 => x"c0989c08",
          8635 => x"80ce9005",
          8636 => x"5387c098",
          8637 => x"9c085287",
          8638 => x"c0989c08",
          8639 => x"5574722e",
          8640 => x"f6388114",
          8641 => x"3387c098",
          8642 => x"9c085252",
          8643 => x"70732787",
          8644 => x"387181ff",
          8645 => x"2edb3887",
          8646 => x"c098a408",
          8647 => x"55727526",
          8648 => x"8338ff52",
          8649 => x"7155ff16",
          8650 => x"7081ff06",
          8651 => x"57537580",
          8652 => x"2ea13874",
          8653 => x"81ff0652",
          8654 => x"71fed538",
          8655 => x"74517081",
          8656 => x"ff065473",
          8657 => x"802e8338",
          8658 => x"81577684",
          8659 => x"b8e40c88",
          8660 => x"3d0d04ff",
          8661 => x"51e839fb",
          8662 => x"3d0d83f2",
          8663 => x"f0085180",
          8664 => x"d0713485",
          8665 => x"0b83f2f0",
          8666 => x"085656fe",
          8667 => x"0b811634",
          8668 => x"800b86f0",
          8669 => x"80e83487",
          8670 => x"c0989c08",
          8671 => x"83f2f008",
          8672 => x"5680ce90",
          8673 => x"055487c0",
          8674 => x"989c0852",
          8675 => x"87c0989c",
          8676 => x"08537272",
          8677 => x"2ef63881",
          8678 => x"153387c0",
          8679 => x"989c0852",
          8680 => x"52707427",
          8681 => x"87387181",
          8682 => x"fe2edb38",
          8683 => x"87c098a4",
          8684 => x"0851ff53",
          8685 => x"70742780",
          8686 => x"c8387153",
          8687 => x"71ff2e80",
          8688 => x"c03887c0",
          8689 => x"989c0880",
          8690 => x"ce900553",
          8691 => x"87c0989c",
          8692 => x"085287c0",
          8693 => x"989c0851",
          8694 => x"70722ef6",
          8695 => x"38811533",
          8696 => x"87c0989c",
          8697 => x"08555273",
          8698 => x"73278738",
          8699 => x"7181ff2e",
          8700 => x"db3887c0",
          8701 => x"98a40851",
          8702 => x"72712683",
          8703 => x"38ff5271",
          8704 => x"53ff1670",
          8705 => x"81ff0657",
          8706 => x"5275802e",
          8707 => x"8a387281",
          8708 => x"ff065473",
          8709 => x"fed538ff",
          8710 => x"39803d0d",
          8711 => x"83e3e851",
          8712 => x"fed0d03f",
          8713 => x"823d0d04",
          8714 => x"f93d0d84",
          8715 => x"b8d4087a",
          8716 => x"7131832a",
          8717 => x"7083ffff",
          8718 => x"0670832b",
          8719 => x"73117033",
          8720 => x"81123371",
          8721 => x"8b2b7183",
          8722 => x"2b077711",
          8723 => x"70338112",
          8724 => x"3371982b",
          8725 => x"71902b07",
          8726 => x"5c544153",
          8727 => x"535d5759",
          8728 => x"52565753",
          8729 => x"80712481",
          8730 => x"af387216",
          8731 => x"82113383",
          8732 => x"1233718b",
          8733 => x"2b71832b",
          8734 => x"07760570",
          8735 => x"33811233",
          8736 => x"71982b71",
          8737 => x"902b0757",
          8738 => x"535c5259",
          8739 => x"56528071",
          8740 => x"24839e38",
          8741 => x"84133385",
          8742 => x"1433718b",
          8743 => x"2b71832b",
          8744 => x"07750576",
          8745 => x"882a5254",
          8746 => x"56577486",
          8747 => x"13347381",
          8748 => x"ff065473",
          8749 => x"87133484",
          8750 => x"b8d40870",
          8751 => x"17841233",
          8752 => x"85133371",
          8753 => x"882b0770",
          8754 => x"882a5c55",
          8755 => x"59545177",
          8756 => x"84143471",
          8757 => x"85143484",
          8758 => x"b8d40816",
          8759 => x"52800b86",
          8760 => x"1334800b",
          8761 => x"87133484",
          8762 => x"b8d40853",
          8763 => x"74841434",
          8764 => x"73851434",
          8765 => x"84b8d408",
          8766 => x"16703381",
          8767 => x"12337188",
          8768 => x"2b078280",
          8769 => x"80077088",
          8770 => x"2a585852",
          8771 => x"52747234",
          8772 => x"75811334",
          8773 => x"893d0d04",
          8774 => x"86123387",
          8775 => x"1333718b",
          8776 => x"2b71832b",
          8777 => x"07751184",
          8778 => x"16338517",
          8779 => x"3371882b",
          8780 => x"0770882a",
          8781 => x"58585451",
          8782 => x"53585871",
          8783 => x"84123472",
          8784 => x"85123484",
          8785 => x"b8d40870",
          8786 => x"16841133",
          8787 => x"85123371",
          8788 => x"8b2b7183",
          8789 => x"2b07565a",
          8790 => x"5a527205",
          8791 => x"86123387",
          8792 => x"13337188",
          8793 => x"2b077088",
          8794 => x"2a525559",
          8795 => x"52778613",
          8796 => x"34728713",
          8797 => x"3484b8d4",
          8798 => x"08157033",
          8799 => x"81123371",
          8800 => x"882b0781",
          8801 => x"ffff0670",
          8802 => x"882a5a5a",
          8803 => x"54527672",
          8804 => x"34778113",
          8805 => x"3484b8d4",
          8806 => x"08701770",
          8807 => x"33811233",
          8808 => x"718b2b71",
          8809 => x"832b0774",
          8810 => x"05703381",
          8811 => x"12337188",
          8812 => x"2b077083",
          8813 => x"2b8ffff8",
          8814 => x"0677057b",
          8815 => x"882a5452",
          8816 => x"53545c5a",
          8817 => x"57545277",
          8818 => x"82143473",
          8819 => x"83143484",
          8820 => x"b8d40870",
          8821 => x"17703381",
          8822 => x"1233718b",
          8823 => x"2b71832b",
          8824 => x"07740570",
          8825 => x"33811233",
          8826 => x"71882b07",
          8827 => x"81ffff06",
          8828 => x"70882a5f",
          8829 => x"5253555a",
          8830 => x"57545277",
          8831 => x"73347081",
          8832 => x"143484b8",
          8833 => x"d4087017",
          8834 => x"82113383",
          8835 => x"1233718b",
          8836 => x"2b71832b",
          8837 => x"07740570",
          8838 => x"33811233",
          8839 => x"71982b71",
          8840 => x"902b0758",
          8841 => x"535d525a",
          8842 => x"57535370",
          8843 => x"8025fce4",
          8844 => x"38713381",
          8845 => x"13337188",
          8846 => x"2b078280",
          8847 => x"80077088",
          8848 => x"2a595954",
          8849 => x"76753477",
          8850 => x"81163484",
          8851 => x"b8d40870",
          8852 => x"17703381",
          8853 => x"1233718b",
          8854 => x"2b71832b",
          8855 => x"07740582",
          8856 => x"14338315",
          8857 => x"3371882b",
          8858 => x"0770882a",
          8859 => x"575c5c52",
          8860 => x"58565253",
          8861 => x"72821534",
          8862 => x"75831534",
          8863 => x"893d0d04",
          8864 => x"f93d0d79",
          8865 => x"84b8d408",
          8866 => x"58587680",
          8867 => x"2e8f3877",
          8868 => x"802e8638",
          8869 => x"7751fb90",
          8870 => x"3f893d0d",
          8871 => x"0484fff4",
          8872 => x"0b84b8d4",
          8873 => x"0ca0800b",
          8874 => x"84b8d023",
          8875 => x"82808053",
          8876 => x"765284ff",
          8877 => x"f451fed3",
          8878 => x"c63f84b8",
          8879 => x"d4085576",
          8880 => x"7534810b",
          8881 => x"81163484",
          8882 => x"b8d40854",
          8883 => x"76841534",
          8884 => x"810b8515",
          8885 => x"3484b8d4",
          8886 => x"08567686",
          8887 => x"1734810b",
          8888 => x"87173484",
          8889 => x"b8d40884",
          8890 => x"b8d022ff",
          8891 => x"05fe8080",
          8892 => x"077083ff",
          8893 => x"ff067088",
          8894 => x"2a585155",
          8895 => x"56748817",
          8896 => x"34738917",
          8897 => x"3484b8d0",
          8898 => x"22701010",
          8899 => x"1084b8d4",
          8900 => x"0805f805",
          8901 => x"55557682",
          8902 => x"1534810b",
          8903 => x"831534fe",
          8904 => x"ee39f73d",
          8905 => x"0d7b5280",
          8906 => x"53815184",
          8907 => x"72278e38",
          8908 => x"fb12832a",
          8909 => x"82057083",
          8910 => x"ffff0651",
          8911 => x"517083ff",
          8912 => x"ff0684b8",
          8913 => x"d4088411",
          8914 => x"33851233",
          8915 => x"71882b07",
          8916 => x"7052595a",
          8917 => x"585581ff",
          8918 => x"ff547580",
          8919 => x"2e80cc38",
          8920 => x"75101010",
          8921 => x"17703381",
          8922 => x"12337188",
          8923 => x"2b077081",
          8924 => x"ffff0679",
          8925 => x"317083ff",
          8926 => x"ff06707a",
          8927 => x"2756535c",
          8928 => x"5c545272",
          8929 => x"74278a38",
          8930 => x"70802e85",
          8931 => x"38757355",
          8932 => x"58841233",
          8933 => x"85133371",
          8934 => x"882b0757",
          8935 => x"5a75c138",
          8936 => x"7381ffff",
          8937 => x"2e853877",
          8938 => x"74545680",
          8939 => x"76832b78",
          8940 => x"11703381",
          8941 => x"12337188",
          8942 => x"2b077081",
          8943 => x"ffff0656",
          8944 => x"565d5659",
          8945 => x"5970792e",
          8946 => x"83388159",
          8947 => x"80517473",
          8948 => x"26828d38",
          8949 => x"78517880",
          8950 => x"2e828538",
          8951 => x"72752e82",
          8952 => x"88387416",
          8953 => x"70832b78",
          8954 => x"11748280",
          8955 => x"80077088",
          8956 => x"2a5b5c56",
          8957 => x"565a7674",
          8958 => x"34788115",
          8959 => x"3484b8d4",
          8960 => x"08157688",
          8961 => x"2a535371",
          8962 => x"82143475",
          8963 => x"83143484",
          8964 => x"b8d40870",
          8965 => x"19703381",
          8966 => x"12337188",
          8967 => x"2b077083",
          8968 => x"2b8ffff8",
          8969 => x"0674057e",
          8970 => x"83ffff06",
          8971 => x"70882a5c",
          8972 => x"58535759",
          8973 => x"52527582",
          8974 => x"12347281",
          8975 => x"ff065372",
          8976 => x"83123484",
          8977 => x"b8d40818",
          8978 => x"54757434",
          8979 => x"72811534",
          8980 => x"84b8d408",
          8981 => x"70198611",
          8982 => x"33871233",
          8983 => x"718b2b71",
          8984 => x"832b0774",
          8985 => x"05585c5c",
          8986 => x"53577584",
          8987 => x"15347285",
          8988 => x"153484b8",
          8989 => x"d4087016",
          8990 => x"55780586",
          8991 => x"11338712",
          8992 => x"3371882b",
          8993 => x"0770882a",
          8994 => x"54545859",
          8995 => x"70861534",
          8996 => x"71871534",
          8997 => x"84b8d408",
          8998 => x"70198411",
          8999 => x"33851233",
          9000 => x"718b2b71",
          9001 => x"832b0774",
          9002 => x"05585a5c",
          9003 => x"5a527586",
          9004 => x"15347287",
          9005 => x"153484b8",
          9006 => x"d4087016",
          9007 => x"55780584",
          9008 => x"11338512",
          9009 => x"3371882b",
          9010 => x"0770882a",
          9011 => x"545c5759",
          9012 => x"70841534",
          9013 => x"79851534",
          9014 => x"84b8d408",
          9015 => x"18840551",
          9016 => x"7084b8e4",
          9017 => x"0c8b3d0d",
          9018 => x"04861433",
          9019 => x"87153371",
          9020 => x"8b2b7183",
          9021 => x"2b077905",
          9022 => x"84173385",
          9023 => x"18337188",
          9024 => x"2b077088",
          9025 => x"2a5a5b59",
          9026 => x"53545274",
          9027 => x"84123476",
          9028 => x"85123484",
          9029 => x"b8d40870",
          9030 => x"19841133",
          9031 => x"85123371",
          9032 => x"8b2b7183",
          9033 => x"2b077405",
          9034 => x"86143387",
          9035 => x"15337188",
          9036 => x"2b077088",
          9037 => x"2a585d5f",
          9038 => x"52565b57",
          9039 => x"5270861a",
          9040 => x"3476871a",
          9041 => x"3484b8d4",
          9042 => x"08187033",
          9043 => x"81123371",
          9044 => x"882b0781",
          9045 => x"ffff0670",
          9046 => x"882a5957",
          9047 => x"54577577",
          9048 => x"34748118",
          9049 => x"3484b8d4",
          9050 => x"08188405",
          9051 => x"51fef139",
          9052 => x"f93d0d79",
          9053 => x"84b8d408",
          9054 => x"58587680",
          9055 => x"2ea03877",
          9056 => x"54778a38",
          9057 => x"7384b8e4",
          9058 => x"0c893d0d",
          9059 => x"047751fb",
          9060 => x"913f84b8",
          9061 => x"e40884b8",
          9062 => x"e40c893d",
          9063 => x"0d0484ff",
          9064 => x"f40b84b8",
          9065 => x"d40ca080",
          9066 => x"0b84b8d0",
          9067 => x"23828080",
          9068 => x"53765284",
          9069 => x"fff451fe",
          9070 => x"cdc53f84",
          9071 => x"b8d40855",
          9072 => x"76753481",
          9073 => x"0b811634",
          9074 => x"84b8d408",
          9075 => x"54768415",
          9076 => x"34810b85",
          9077 => x"153484b8",
          9078 => x"d4085676",
          9079 => x"86173481",
          9080 => x"0b871734",
          9081 => x"84b8d408",
          9082 => x"84b8d022",
          9083 => x"ff05fe80",
          9084 => x"80077083",
          9085 => x"ffff0670",
          9086 => x"882a5851",
          9087 => x"55567488",
          9088 => x"17347389",
          9089 => x"173484b8",
          9090 => x"d0227010",
          9091 => x"101084b8",
          9092 => x"d40805f8",
          9093 => x"05555576",
          9094 => x"82153481",
          9095 => x"0b831534",
          9096 => x"77547780",
          9097 => x"2efedd38",
          9098 => x"fee339ed",
          9099 => x"3d0d6567",
          9100 => x"415f8070",
          9101 => x"84b8d408",
          9102 => x"59454176",
          9103 => x"612e84aa",
          9104 => x"387e802e",
          9105 => x"85af387f",
          9106 => x"802e88d7",
          9107 => x"38815484",
          9108 => x"60278f38",
          9109 => x"7ffb0583",
          9110 => x"2a820570",
          9111 => x"83ffff06",
          9112 => x"55587383",
          9113 => x"ffff067f",
          9114 => x"7831832a",
          9115 => x"7083ffff",
          9116 => x"0670832b",
          9117 => x"7a117033",
          9118 => x"81123371",
          9119 => x"882b0770",
          9120 => x"75317083",
          9121 => x"ffff0670",
          9122 => x"101010fc",
          9123 => x"0573832b",
          9124 => x"61117033",
          9125 => x"81123371",
          9126 => x"882b0770",
          9127 => x"902b7090",
          9128 => x"2c534245",
          9129 => x"46445354",
          9130 => x"43445c48",
          9131 => x"59525e5f",
          9132 => x"42807a24",
          9133 => x"85fd3882",
          9134 => x"15338316",
          9135 => x"3371882b",
          9136 => x"07701010",
          9137 => x"10197033",
          9138 => x"81123371",
          9139 => x"982b7190",
          9140 => x"2b07535c",
          9141 => x"53565656",
          9142 => x"80742485",
          9143 => x"c9387a62",
          9144 => x"2782f638",
          9145 => x"631b5877",
          9146 => x"622e87a2",
          9147 => x"3860802e",
          9148 => x"85f93860",
          9149 => x"1b587762",
          9150 => x"2587be38",
          9151 => x"63185961",
          9152 => x"792492f7",
          9153 => x"38761e70",
          9154 => x"33811233",
          9155 => x"718b2b71",
          9156 => x"832b077a",
          9157 => x"11703381",
          9158 => x"12337198",
          9159 => x"2b71902b",
          9160 => x"07474359",
          9161 => x"5253575b",
          9162 => x"58806024",
          9163 => x"8cba3876",
          9164 => x"1e821133",
          9165 => x"83123371",
          9166 => x"8b2b7183",
          9167 => x"2b077a11",
          9168 => x"86113387",
          9169 => x"1233718b",
          9170 => x"2b71832b",
          9171 => x"077e0584",
          9172 => x"14338515",
          9173 => x"3371882b",
          9174 => x"0770882a",
          9175 => x"59574852",
          9176 => x"5b415853",
          9177 => x"5c595677",
          9178 => x"841d3479",
          9179 => x"851d3484",
          9180 => x"b8d40870",
          9181 => x"17841133",
          9182 => x"85123371",
          9183 => x"8b2b7183",
          9184 => x"2b077405",
          9185 => x"86143387",
          9186 => x"15337188",
          9187 => x"2b077088",
          9188 => x"2a5f425e",
          9189 => x"52405741",
          9190 => x"57778616",
          9191 => x"347b8716",
          9192 => x"3484b8d4",
          9193 => x"08167033",
          9194 => x"81123371",
          9195 => x"882b0781",
          9196 => x"ffff0670",
          9197 => x"882a5a5c",
          9198 => x"5e597679",
          9199 => x"3479811a",
          9200 => x"3484b8d4",
          9201 => x"08701f82",
          9202 => x"11338312",
          9203 => x"33718b2b",
          9204 => x"71832b07",
          9205 => x"74057333",
          9206 => x"81153371",
          9207 => x"882b0770",
          9208 => x"882a415c",
          9209 => x"455d5f5a",
          9210 => x"55557979",
          9211 => x"3475811a",
          9212 => x"3484b8d4",
          9213 => x"08701f70",
          9214 => x"33811233",
          9215 => x"718b2b71",
          9216 => x"832b0774",
          9217 => x"05821433",
          9218 => x"83153371",
          9219 => x"882b0770",
          9220 => x"882a415c",
          9221 => x"455d5f5a",
          9222 => x"55557982",
          9223 => x"1a347583",
          9224 => x"1a3484b8",
          9225 => x"d408701f",
          9226 => x"82113383",
          9227 => x"12337188",
          9228 => x"2b076657",
          9229 => x"62567083",
          9230 => x"2b42525a",
          9231 => x"5d7e0584",
          9232 => x"0551fec4",
          9233 => x"fd3f84b8",
          9234 => x"d4081e84",
          9235 => x"05616505",
          9236 => x"1c7083ff",
          9237 => x"ff065d44",
          9238 => x"5f7a6226",
          9239 => x"81b6387e",
          9240 => x"547384b8",
          9241 => x"e40c953d",
          9242 => x"0d0484ff",
          9243 => x"f40b84b8",
          9244 => x"d40ca080",
          9245 => x"0b84b8d0",
          9246 => x"23828080",
          9247 => x"53605284",
          9248 => x"fff451fe",
          9249 => x"c7f93f84",
          9250 => x"b8d4085e",
          9251 => x"607e3481",
          9252 => x"0b811f34",
          9253 => x"84b8d408",
          9254 => x"5d60841e",
          9255 => x"34810b85",
          9256 => x"1e3484b8",
          9257 => x"d4085c60",
          9258 => x"861d3481",
          9259 => x"0b871d34",
          9260 => x"84b8d408",
          9261 => x"84b8d022",
          9262 => x"ff05fe80",
          9263 => x"80077083",
          9264 => x"ffff0670",
          9265 => x"882a5c5a",
          9266 => x"5b577888",
          9267 => x"18347789",
          9268 => x"183484b8",
          9269 => x"d0227010",
          9270 => x"101084b8",
          9271 => x"d40805f8",
          9272 => x"05555660",
          9273 => x"82153481",
          9274 => x"0b831534",
          9275 => x"84b8d408",
          9276 => x"577efad3",
          9277 => x"3876802e",
          9278 => x"828c387e",
          9279 => x"547f802e",
          9280 => x"fedf387f",
          9281 => x"51f49b3f",
          9282 => x"84b8e408",
          9283 => x"84b8e40c",
          9284 => x"953d0d04",
          9285 => x"611c84b8",
          9286 => x"d4087183",
          9287 => x"2b71115e",
          9288 => x"447f0570",
          9289 => x"33811233",
          9290 => x"71882b07",
          9291 => x"81ffff06",
          9292 => x"70882a48",
          9293 => x"445b5e40",
          9294 => x"637b3460",
          9295 => x"811c3461",
          9296 => x"84b8d408",
          9297 => x"057c882a",
          9298 => x"57587582",
          9299 => x"19347b83",
          9300 => x"193484b8",
          9301 => x"d408701f",
          9302 => x"70338112",
          9303 => x"3371882b",
          9304 => x"0770832b",
          9305 => x"8ffff806",
          9306 => x"74056483",
          9307 => x"ffff0670",
          9308 => x"882a4a5c",
          9309 => x"47575e5b",
          9310 => x"5d636382",
          9311 => x"05347681",
          9312 => x"ff064160",
          9313 => x"63830534",
          9314 => x"84b8d408",
          9315 => x"1e5b637b",
          9316 => x"3460811c",
          9317 => x"346184b8",
          9318 => x"d4080584",
          9319 => x"0551ed88",
          9320 => x"3f7e54fd",
          9321 => x"bc397b75",
          9322 => x"317083ff",
          9323 => x"ff064254",
          9324 => x"faac3977",
          9325 => x"81ffff06",
          9326 => x"76317083",
          9327 => x"ffff0682",
          9328 => x"17338318",
          9329 => x"3371882b",
          9330 => x"07701010",
          9331 => x"101b7033",
          9332 => x"81123371",
          9333 => x"982b7190",
          9334 => x"2b07535e",
          9335 => x"53545858",
          9336 => x"45547380",
          9337 => x"25f9f738",
          9338 => x"ffbc3961",
          9339 => x"7824fa83",
          9340 => x"38807a24",
          9341 => x"8b8f3877",
          9342 => x"83ffff06",
          9343 => x"5b617b27",
          9344 => x"fcdd38fe",
          9345 => x"8f3984ff",
          9346 => x"f40b84b8",
          9347 => x"d40ca080",
          9348 => x"0b84b8d0",
          9349 => x"23828080",
          9350 => x"537e5284",
          9351 => x"fff451fe",
          9352 => x"c4dd3f84",
          9353 => x"b8d4085a",
          9354 => x"7e7a3481",
          9355 => x"0b811b34",
          9356 => x"84b8d408",
          9357 => x"597e841a",
          9358 => x"34810b85",
          9359 => x"1a3484b8",
          9360 => x"d408587e",
          9361 => x"86193481",
          9362 => x"0b871934",
          9363 => x"84b8d408",
          9364 => x"84b8d022",
          9365 => x"ff05fe80",
          9366 => x"80077083",
          9367 => x"ffff0670",
          9368 => x"882a5856",
          9369 => x"57447464",
          9370 => x"88053473",
          9371 => x"64890534",
          9372 => x"84b8d022",
          9373 => x"70101010",
          9374 => x"84b8d408",
          9375 => x"05f80542",
          9376 => x"437e6182",
          9377 => x"05348161",
          9378 => x"830534fc",
          9379 => x"ee39807a",
          9380 => x"2483de38",
          9381 => x"6183ffff",
          9382 => x"065b617b",
          9383 => x"27fbc038",
          9384 => x"fcf23976",
          9385 => x"802e82bd",
          9386 => x"387e51ea",
          9387 => x"fb3f7f54",
          9388 => x"7384b8e4",
          9389 => x"0c953d0d",
          9390 => x"04761e82",
          9391 => x"11338312",
          9392 => x"33718b2b",
          9393 => x"71832b07",
          9394 => x"7a118611",
          9395 => x"33871233",
          9396 => x"718b2b71",
          9397 => x"832b077e",
          9398 => x"05841433",
          9399 => x"85153371",
          9400 => x"882b0770",
          9401 => x"882a4344",
          9402 => x"45565b46",
          9403 => x"58535c45",
          9404 => x"56786484",
          9405 => x"05347a64",
          9406 => x"85053484",
          9407 => x"b8d40870",
          9408 => x"17841133",
          9409 => x"85123371",
          9410 => x"8b2b7183",
          9411 => x"2b077405",
          9412 => x"86143387",
          9413 => x"15337188",
          9414 => x"2b077088",
          9415 => x"2a5b4142",
          9416 => x"485d595d",
          9417 => x"41736486",
          9418 => x"05347a64",
          9419 => x"87053484",
          9420 => x"b8d40816",
          9421 => x"70338112",
          9422 => x"3371882b",
          9423 => x"0781ffff",
          9424 => x"0670882a",
          9425 => x"5f5c5a5d",
          9426 => x"7b7d3479",
          9427 => x"811e3484",
          9428 => x"b8d40870",
          9429 => x"1f821133",
          9430 => x"83123371",
          9431 => x"8b2b7183",
          9432 => x"2b077405",
          9433 => x"73338115",
          9434 => x"3371882b",
          9435 => x"0770882a",
          9436 => x"5e5c5e40",
          9437 => x"43574554",
          9438 => x"767c3475",
          9439 => x"811d3484",
          9440 => x"b8d40870",
          9441 => x"1f703381",
          9442 => x"1233718b",
          9443 => x"2b71832b",
          9444 => x"07740582",
          9445 => x"14338315",
          9446 => x"3371882b",
          9447 => x"0770882a",
          9448 => x"4047405b",
          9449 => x"405c5555",
          9450 => x"78821834",
          9451 => x"60831834",
          9452 => x"84b8d408",
          9453 => x"701f8211",
          9454 => x"33831233",
          9455 => x"71882b07",
          9456 => x"66576256",
          9457 => x"70832b42",
          9458 => x"52585d7e",
          9459 => x"05840551",
          9460 => x"febdef3f",
          9461 => x"84b8d408",
          9462 => x"1e840578",
          9463 => x"83ffff06",
          9464 => x"5c5ffc99",
          9465 => x"3984fff4",
          9466 => x"0b84b8d4",
          9467 => x"0ca0800b",
          9468 => x"84b8d023",
          9469 => x"82808053",
          9470 => x"7f5284ff",
          9471 => x"f451fec0",
          9472 => x"fe3f84b8",
          9473 => x"d408567f",
          9474 => x"7634810b",
          9475 => x"81173484",
          9476 => x"b8d40855",
          9477 => x"7f841634",
          9478 => x"810b8516",
          9479 => x"3484b8d4",
          9480 => x"08547f86",
          9481 => x"1534810b",
          9482 => x"87153484",
          9483 => x"b8d40884",
          9484 => x"b8d022ff",
          9485 => x"05fe8080",
          9486 => x"077083ff",
          9487 => x"ff067088",
          9488 => x"2a454344",
          9489 => x"5e61881f",
          9490 => x"3460891f",
          9491 => x"3484b8d0",
          9492 => x"22701010",
          9493 => x"1084b8d4",
          9494 => x"0805f805",
          9495 => x"5c5d7f82",
          9496 => x"1c34810b",
          9497 => x"831c347e",
          9498 => x"51e7bd3f",
          9499 => x"7f54fcc0",
          9500 => x"39861933",
          9501 => x"871a3371",
          9502 => x"8b2b7183",
          9503 => x"2b077905",
          9504 => x"841c3385",
          9505 => x"1d337188",
          9506 => x"2b077088",
          9507 => x"2a5c485e",
          9508 => x"43595576",
          9509 => x"61840534",
          9510 => x"63618505",
          9511 => x"3484b8d4",
          9512 => x"08701e84",
          9513 => x"11338512",
          9514 => x"33718b2b",
          9515 => x"71832b07",
          9516 => x"74058614",
          9517 => x"33871533",
          9518 => x"71882b07",
          9519 => x"70882a41",
          9520 => x"5f484859",
          9521 => x"56594079",
          9522 => x"64860534",
          9523 => x"78648705",
          9524 => x"3484b8d4",
          9525 => x"081d7033",
          9526 => x"81123371",
          9527 => x"882b0781",
          9528 => x"ffff0670",
          9529 => x"882a5942",
          9530 => x"58587578",
          9531 => x"347f8119",
          9532 => x"3484b8d4",
          9533 => x"08701f70",
          9534 => x"33811233",
          9535 => x"718b2b71",
          9536 => x"832b0774",
          9537 => x"05703381",
          9538 => x"12337188",
          9539 => x"2b077083",
          9540 => x"2b8ffff8",
          9541 => x"06770563",
          9542 => x"882a485d",
          9543 => x"5d5a5d40",
          9544 => x"5d44417f",
          9545 => x"8217347b",
          9546 => x"83173484",
          9547 => x"b8d40870",
          9548 => x"1f703381",
          9549 => x"1233718b",
          9550 => x"2b71832b",
          9551 => x"07740570",
          9552 => x"33811233",
          9553 => x"71882b07",
          9554 => x"81ffff06",
          9555 => x"70882a48",
          9556 => x"5d5e5e46",
          9557 => x"5a415b60",
          9558 => x"60347660",
          9559 => x"81053461",
          9560 => x"83ffff06",
          9561 => x"5bfab339",
          9562 => x"86153387",
          9563 => x"1633718b",
          9564 => x"2b71832b",
          9565 => x"07790584",
          9566 => x"18338519",
          9567 => x"3371882b",
          9568 => x"0770882a",
          9569 => x"5e5e5a52",
          9570 => x"415d7884",
          9571 => x"1e347985",
          9572 => x"1e3484b8",
          9573 => x"d4087019",
          9574 => x"84113385",
          9575 => x"1233718b",
          9576 => x"2b71832b",
          9577 => x"07740586",
          9578 => x"14338715",
          9579 => x"3371882b",
          9580 => x"0770882a",
          9581 => x"44565e52",
          9582 => x"5a425556",
          9583 => x"7c608605",
          9584 => x"34756087",
          9585 => x"053484b8",
          9586 => x"d4081870",
          9587 => x"33811233",
          9588 => x"71882b07",
          9589 => x"81ffff06",
          9590 => x"70882a5b",
          9591 => x"5b585577",
          9592 => x"75347881",
          9593 => x"163484b8",
          9594 => x"d408701f",
          9595 => x"70338112",
          9596 => x"33718b2b",
          9597 => x"71832b07",
          9598 => x"74057033",
          9599 => x"81123371",
          9600 => x"882b0770",
          9601 => x"832b8fff",
          9602 => x"f8067705",
          9603 => x"63882a56",
          9604 => x"545f5f58",
          9605 => x"59425e55",
          9606 => x"7f821734",
          9607 => x"7b831734",
          9608 => x"84b8d408",
          9609 => x"701f7033",
          9610 => x"81123371",
          9611 => x"8b2b7183",
          9612 => x"2b077405",
          9613 => x"70338112",
          9614 => x"3371882b",
          9615 => x"0781ffff",
          9616 => x"0670882a",
          9617 => x"5d545e58",
          9618 => x"5b595d55",
          9619 => x"757c3476",
          9620 => x"811d3484",
          9621 => x"b8d40870",
          9622 => x"1f821133",
          9623 => x"83123371",
          9624 => x"8b2b7183",
          9625 => x"2b077411",
          9626 => x"86113387",
          9627 => x"1233718b",
          9628 => x"2b71832b",
          9629 => x"07780584",
          9630 => x"14338515",
          9631 => x"3371882b",
          9632 => x"0770882a",
          9633 => x"59574952",
          9634 => x"5c425953",
          9635 => x"5d5a5757",
          9636 => x"77841d34",
          9637 => x"79851d34",
          9638 => x"84b8d408",
          9639 => x"70178411",
          9640 => x"33851233",
          9641 => x"718b2b71",
          9642 => x"832b0774",
          9643 => x"05861433",
          9644 => x"87153371",
          9645 => x"882b0770",
          9646 => x"882a5f42",
          9647 => x"5e524057",
          9648 => x"41577786",
          9649 => x"16347b87",
          9650 => x"163484b8",
          9651 => x"d4081670",
          9652 => x"33811233",
          9653 => x"71882b07",
          9654 => x"81ffff06",
          9655 => x"70882a5a",
          9656 => x"5c5e5976",
          9657 => x"79347981",
          9658 => x"1a3484b8",
          9659 => x"d408701f",
          9660 => x"82113383",
          9661 => x"1233718b",
          9662 => x"2b71832b",
          9663 => x"07740573",
          9664 => x"33811533",
          9665 => x"71882b07",
          9666 => x"70882a41",
          9667 => x"5c455d5f",
          9668 => x"5a555579",
          9669 => x"79347581",
          9670 => x"1a3484b8",
          9671 => x"d408701f",
          9672 => x"70338112",
          9673 => x"33718b2b",
          9674 => x"71832b07",
          9675 => x"74058214",
          9676 => x"33831533",
          9677 => x"71882b07",
          9678 => x"70882a41",
          9679 => x"5c455d5f",
          9680 => x"5a555579",
          9681 => x"821a3475",
          9682 => x"831a3484",
          9683 => x"b8d40870",
          9684 => x"1f821133",
          9685 => x"83123371",
          9686 => x"882b0766",
          9687 => x"57625670",
          9688 => x"832b4252",
          9689 => x"5a5d7e05",
          9690 => x"840551fe",
          9691 => x"b6d43f84",
          9692 => x"b8d4081e",
          9693 => x"84056165",
          9694 => x"051c7083",
          9695 => x"ffff065d",
          9696 => x"445ff1d5",
          9697 => x"39861933",
          9698 => x"871a3371",
          9699 => x"8b2b7183",
          9700 => x"2b077905",
          9701 => x"841c3385",
          9702 => x"1d337188",
          9703 => x"2b077088",
          9704 => x"2a40485d",
          9705 => x"4341557a",
          9706 => x"61840534",
          9707 => x"63618505",
          9708 => x"3484b8d4",
          9709 => x"08701e84",
          9710 => x"11338512",
          9711 => x"33718b2b",
          9712 => x"71832b07",
          9713 => x"74058614",
          9714 => x"33871533",
          9715 => x"71882b07",
          9716 => x"70882a5b",
          9717 => x"415f485c",
          9718 => x"59415673",
          9719 => x"64860534",
          9720 => x"7a648705",
          9721 => x"3484b8d4",
          9722 => x"081d7033",
          9723 => x"81123371",
          9724 => x"882b0781",
          9725 => x"ffff0670",
          9726 => x"882a5c5f",
          9727 => x"42557875",
          9728 => x"347c8116",
          9729 => x"3484b8d4",
          9730 => x"08701f70",
          9731 => x"33811233",
          9732 => x"718b2b71",
          9733 => x"832b0774",
          9734 => x"05703381",
          9735 => x"12337188",
          9736 => x"2b077083",
          9737 => x"2b8ffff8",
          9738 => x"06770563",
          9739 => x"882a5d44",
          9740 => x"5c49585e",
          9741 => x"45584074",
          9742 => x"821e347b",
          9743 => x"831e3484",
          9744 => x"b8d40870",
          9745 => x"1f703381",
          9746 => x"1233718b",
          9747 => x"2b71832b",
          9748 => x"07740570",
          9749 => x"33811233",
          9750 => x"71882b07",
          9751 => x"81ffff06",
          9752 => x"70882a47",
          9753 => x"5f495846",
          9754 => x"595e5b7f",
          9755 => x"7d347881",
          9756 => x"1e347783",
          9757 => x"ffff065b",
          9758 => x"f383397e",
          9759 => x"605254e5",
          9760 => x"a13f84b8",
          9761 => x"e4085f84",
          9762 => x"b8e40880",
          9763 => x"2e933862",
          9764 => x"53735284",
          9765 => x"b8e40851",
          9766 => x"feb5cf3f",
          9767 => x"7351df88",
          9768 => x"3f615b61",
          9769 => x"7b27efb7",
          9770 => x"38f0e939",
          9771 => x"f93d0d7a",
          9772 => x"7a2984b8",
          9773 => x"d4085858",
          9774 => x"76802eb7",
          9775 => x"38775477",
          9776 => x"8a387384",
          9777 => x"b8e40c89",
          9778 => x"3d0d0477",
          9779 => x"51e4d33f",
          9780 => x"84b8e408",
          9781 => x"5484b8e4",
          9782 => x"08802ee6",
          9783 => x"38775380",
          9784 => x"5284b8e4",
          9785 => x"0851feb7",
          9786 => x"963f7384",
          9787 => x"b8e40c89",
          9788 => x"3d0d0484",
          9789 => x"fff40b84",
          9790 => x"b8d40ca0",
          9791 => x"800b84b8",
          9792 => x"d0238280",
          9793 => x"80537652",
          9794 => x"84fff451",
          9795 => x"feb6f03f",
          9796 => x"84b8d408",
          9797 => x"55767534",
          9798 => x"810b8116",
          9799 => x"3484b8d4",
          9800 => x"08547684",
          9801 => x"1534810b",
          9802 => x"85153484",
          9803 => x"b8d40856",
          9804 => x"76861734",
          9805 => x"810b8717",
          9806 => x"3484b8d4",
          9807 => x"0884b8d0",
          9808 => x"22ff05fe",
          9809 => x"80800770",
          9810 => x"83ffff06",
          9811 => x"70882a58",
          9812 => x"51555674",
          9813 => x"88173473",
          9814 => x"89173484",
          9815 => x"b8d02270",
          9816 => x"10101084",
          9817 => x"b8d40805",
          9818 => x"f8055555",
          9819 => x"76821534",
          9820 => x"810b8315",
          9821 => x"34775477",
          9822 => x"802efec6",
          9823 => x"38fecc39",
          9824 => x"ff3d0d02",
          9825 => x"8f053351",
          9826 => x"81527072",
          9827 => x"26873884",
          9828 => x"b8e01133",
          9829 => x"527184b8",
          9830 => x"e40c833d",
          9831 => x"0d04fe3d",
          9832 => x"0d029305",
          9833 => x"33528353",
          9834 => x"7181269d",
          9835 => x"387151d4",
          9836 => x"bb3f84b8",
          9837 => x"e40881ff",
          9838 => x"06537287",
          9839 => x"387284b8",
          9840 => x"e0133484",
          9841 => x"b8e01233",
          9842 => x"537284b8",
          9843 => x"e40c843d",
          9844 => x"0d04f73d",
          9845 => x"0d7c7e60",
          9846 => x"028c05af",
          9847 => x"05335a5c",
          9848 => x"57598154",
          9849 => x"76742687",
          9850 => x"3884b8e0",
          9851 => x"17335473",
          9852 => x"81065483",
          9853 => x"5573bd38",
          9854 => x"7358850b",
          9855 => x"87c0988c",
          9856 => x"0c785375",
          9857 => x"527651d5",
          9858 => x"ca3f84b8",
          9859 => x"e40881ff",
          9860 => x"06557480",
          9861 => x"2ea73887",
          9862 => x"c0988c08",
          9863 => x"5473e238",
          9864 => x"797826d6",
          9865 => x"3874fc80",
          9866 => x"80065473",
          9867 => x"802e8338",
          9868 => x"81547355",
          9869 => x"7484b8e4",
          9870 => x"0c8b3d0d",
          9871 => x"04848016",
          9872 => x"81197081",
          9873 => x"ff065a55",
          9874 => x"56797826",
          9875 => x"ffac38d5",
          9876 => x"39f73d0d",
          9877 => x"7c7e6002",
          9878 => x"8c05af05",
          9879 => x"335a5c57",
          9880 => x"59815476",
          9881 => x"74268738",
          9882 => x"84b8e017",
          9883 => x"33547381",
          9884 => x"06548355",
          9885 => x"73bd3873",
          9886 => x"58850b87",
          9887 => x"c0988c0c",
          9888 => x"78537552",
          9889 => x"7651d78e",
          9890 => x"3f84b8e4",
          9891 => x"0881ff06",
          9892 => x"5574802e",
          9893 => x"a73887c0",
          9894 => x"988c0854",
          9895 => x"73e23879",
          9896 => x"7826d638",
          9897 => x"74fc8080",
          9898 => x"06547380",
          9899 => x"2e833881",
          9900 => x"54735574",
          9901 => x"84b8e40c",
          9902 => x"8b3d0d04",
          9903 => x"84801681",
          9904 => x"197081ff",
          9905 => x"065a5556",
          9906 => x"797826ff",
          9907 => x"ac38d539",
          9908 => x"fc3d0d78",
          9909 => x"0284059b",
          9910 => x"05330288",
          9911 => x"059f0533",
          9912 => x"53535581",
          9913 => x"53717326",
          9914 => x"873884b8",
          9915 => x"e0123353",
          9916 => x"72810654",
          9917 => x"8353739b",
          9918 => x"38850b87",
          9919 => x"c0988c0c",
          9920 => x"81537073",
          9921 => x"2e963872",
          9922 => x"7125ad38",
          9923 => x"70832e9a",
          9924 => x"38845372",
          9925 => x"84b8e40c",
          9926 => x"863d0d04",
          9927 => x"88800a75",
          9928 => x"0c7384b8",
          9929 => x"e40c863d",
          9930 => x"0d048180",
          9931 => x"750c800b",
          9932 => x"84b8e40c",
          9933 => x"863d0d04",
          9934 => x"71842b87",
          9935 => x"c0928c11",
          9936 => x"535470cd",
          9937 => x"38710870",
          9938 => x"812a8106",
          9939 => x"51517080",
          9940 => x"2e8a3887",
          9941 => x"c0988c08",
          9942 => x"5574ea38",
          9943 => x"87c0988c",
          9944 => x"085170ca",
          9945 => x"3881720c",
          9946 => x"87c0928c",
          9947 => x"14527108",
          9948 => x"82065473",
          9949 => x"802eff9b",
          9950 => x"38710882",
          9951 => x"065473ee",
          9952 => x"38ff9039",
          9953 => x"f63d0d7c",
          9954 => x"58800b83",
          9955 => x"1933715b",
          9956 => x"56577477",
          9957 => x"2e098106",
          9958 => x"a8387733",
          9959 => x"5675832e",
          9960 => x"81873880",
          9961 => x"53805281",
          9962 => x"183351fe",
          9963 => x"a33f84b8",
          9964 => x"e408802e",
          9965 => x"83388159",
          9966 => x"7884b8e4",
          9967 => x"0c8c3d0d",
          9968 => x"048154b4",
          9969 => x"180853b8",
          9970 => x"18705381",
          9971 => x"1933525a",
          9972 => x"fcff3f81",
          9973 => x"5984b8e4",
          9974 => x"08772e09",
          9975 => x"8106d938",
          9976 => x"84b8e408",
          9977 => x"831934b4",
          9978 => x"180870a8",
          9979 => x"1a0831a0",
          9980 => x"1a0884b8",
          9981 => x"e4085c58",
          9982 => x"565b7476",
          9983 => x"27ff9b38",
          9984 => x"82183355",
          9985 => x"74822e09",
          9986 => x"8106ff8e",
          9987 => x"38815475",
          9988 => x"1b537952",
          9989 => x"81183351",
          9990 => x"fcb73f76",
          9991 => x"78335759",
          9992 => x"75832e09",
          9993 => x"8106fefb",
          9994 => x"38841833",
          9995 => x"5776812e",
          9996 => x"098106fe",
          9997 => x"ee38b818",
          9998 => x"5a84807a",
          9999 => x"56578075",
         10000 => x"70810557",
         10001 => x"34ff1757",
         10002 => x"76f43880",
         10003 => x"d50b84b6",
         10004 => x"1934ffaa",
         10005 => x"0b84b719",
         10006 => x"3480d27a",
         10007 => x"3480d20b",
         10008 => x"b9193480",
         10009 => x"e10bba19",
         10010 => x"3480c10b",
         10011 => x"bb193480",
         10012 => x"f20b849c",
         10013 => x"193480f2",
         10014 => x"0b849d19",
         10015 => x"3480c10b",
         10016 => x"849e1934",
         10017 => x"80e10b84",
         10018 => x"9f193494",
         10019 => x"18085574",
         10020 => x"84a01934",
         10021 => x"74882a5b",
         10022 => x"7a84a119",
         10023 => x"3474902a",
         10024 => x"567584a2",
         10025 => x"19347498",
         10026 => x"2a5b7a84",
         10027 => x"a3193490",
         10028 => x"18085b7a",
         10029 => x"84a41934",
         10030 => x"7a882a55",
         10031 => x"7484a519",
         10032 => x"347a902a",
         10033 => x"567584a6",
         10034 => x"19347a98",
         10035 => x"2a557484",
         10036 => x"a71934a4",
         10037 => x"18088105",
         10038 => x"70b41a0c",
         10039 => x"5b81547a",
         10040 => x"53795281",
         10041 => x"183351fa",
         10042 => x"e83f7684",
         10043 => x"19348053",
         10044 => x"80528118",
         10045 => x"3351fbd8",
         10046 => x"3f84b8e4",
         10047 => x"08802efd",
         10048 => x"b738fdb2",
         10049 => x"39f33d0d",
         10050 => x"60607008",
         10051 => x"59565681",
         10052 => x"76278838",
         10053 => x"9c170876",
         10054 => x"268c3881",
         10055 => x"587784b8",
         10056 => x"e40c8f3d",
         10057 => x"0d04ff77",
         10058 => x"33565874",
         10059 => x"822e81cc",
         10060 => x"38748224",
         10061 => x"82a53874",
         10062 => x"812e0981",
         10063 => x"06dd3875",
         10064 => x"812a1670",
         10065 => x"892aa819",
         10066 => x"08055a5a",
         10067 => x"805bb417",
         10068 => x"08792eb0",
         10069 => x"38831733",
         10070 => x"5c7b7b2e",
         10071 => x"09810683",
         10072 => x"de388154",
         10073 => x"7853b817",
         10074 => x"52811733",
         10075 => x"51f8e33f",
         10076 => x"84b8e408",
         10077 => x"802e8538",
         10078 => x"ff59815b",
         10079 => x"78b4180c",
         10080 => x"7aff9a38",
         10081 => x"7983ff06",
         10082 => x"17b81133",
         10083 => x"811c7089",
         10084 => x"2aa81b08",
         10085 => x"05535d5d",
         10086 => x"59b41708",
         10087 => x"792eb538",
         10088 => x"800b8318",
         10089 => x"33715c56",
         10090 => x"5d747d2e",
         10091 => x"09810684",
         10092 => x"b5388154",
         10093 => x"7853b817",
         10094 => x"52811733",
         10095 => x"51f8933f",
         10096 => x"84b8e408",
         10097 => x"802e8538",
         10098 => x"ff59815a",
         10099 => x"78b4180c",
         10100 => x"79feca38",
         10101 => x"7a83ff06",
         10102 => x"17b81133",
         10103 => x"70882b7e",
         10104 => x"07788106",
         10105 => x"71842a53",
         10106 => x"5d59595d",
         10107 => x"79feae38",
         10108 => x"769fff06",
         10109 => x"84b8e40c",
         10110 => x"8f3d0d04",
         10111 => x"75882aa8",
         10112 => x"18080559",
         10113 => x"b4170879",
         10114 => x"2eb53880",
         10115 => x"0b831833",
         10116 => x"715c5d5b",
         10117 => x"7b7b2e09",
         10118 => x"810681c2",
         10119 => x"38815478",
         10120 => x"53b81752",
         10121 => x"81173351",
         10122 => x"f7a83f84",
         10123 => x"b8e40880",
         10124 => x"2e8538ff",
         10125 => x"59815a78",
         10126 => x"b4180c79",
         10127 => x"fddf3875",
         10128 => x"1083fe06",
         10129 => x"7705b805",
         10130 => x"81113371",
         10131 => x"3371882b",
         10132 => x"0784b8e4",
         10133 => x"0c575b8f",
         10134 => x"3d0d0474",
         10135 => x"832e0981",
         10136 => x"06fdb838",
         10137 => x"75872aa8",
         10138 => x"18080559",
         10139 => x"b4170879",
         10140 => x"2eb53880",
         10141 => x"0b831833",
         10142 => x"715c5e5b",
         10143 => x"7c7b2e09",
         10144 => x"81068281",
         10145 => x"38815478",
         10146 => x"53b81752",
         10147 => x"81173351",
         10148 => x"f6c03f84",
         10149 => x"b8e40880",
         10150 => x"2e8538ff",
         10151 => x"59815a78",
         10152 => x"b4180c79",
         10153 => x"fcf73875",
         10154 => x"822b83fc",
         10155 => x"067705b8",
         10156 => x"05831133",
         10157 => x"82123371",
         10158 => x"902b7188",
         10159 => x"2b078114",
         10160 => x"33707207",
         10161 => x"882b7533",
         10162 => x"7180ffff",
         10163 => x"fe800607",
         10164 => x"84b8e40c",
         10165 => x"415c5e59",
         10166 => x"5a568f3d",
         10167 => x"0d048154",
         10168 => x"b4170853",
         10169 => x"b8177053",
         10170 => x"81183352",
         10171 => x"5cf6e23f",
         10172 => x"815a84b8",
         10173 => x"e4087b2e",
         10174 => x"098106fe",
         10175 => x"be3884b8",
         10176 => x"e4088318",
         10177 => x"34b41708",
         10178 => x"a8180831",
         10179 => x"84b8e408",
         10180 => x"5b5e7da0",
         10181 => x"180827fe",
         10182 => x"84388217",
         10183 => x"33557482",
         10184 => x"2e098106",
         10185 => x"fdf73881",
         10186 => x"54b41708",
         10187 => x"a0180805",
         10188 => x"537b5281",
         10189 => x"173351f6",
         10190 => x"983f7a5a",
         10191 => x"fddf3981",
         10192 => x"54b41708",
         10193 => x"53b81770",
         10194 => x"53811833",
         10195 => x"525cf681",
         10196 => x"3f84b8e4",
         10197 => x"087b2e09",
         10198 => x"81068281",
         10199 => x"3884b8e4",
         10200 => x"08831834",
         10201 => x"b41708a8",
         10202 => x"1808315d",
         10203 => x"7ca01808",
         10204 => x"278b3882",
         10205 => x"17335e7d",
         10206 => x"822e81cb",
         10207 => x"3884b8e4",
         10208 => x"085bfbde",
         10209 => x"398154b4",
         10210 => x"170853b8",
         10211 => x"17705381",
         10212 => x"1833525c",
         10213 => x"f5bb3f81",
         10214 => x"5a84b8e4",
         10215 => x"087b2e09",
         10216 => x"8106fdff",
         10217 => x"3884b8e4",
         10218 => x"08831834",
         10219 => x"b41708a8",
         10220 => x"18083184",
         10221 => x"b8e4085b",
         10222 => x"5e7da018",
         10223 => x"0827fdc5",
         10224 => x"38821733",
         10225 => x"5574822e",
         10226 => x"098106fd",
         10227 => x"b8388154",
         10228 => x"b41708a0",
         10229 => x"18080553",
         10230 => x"7b528117",
         10231 => x"3351f4f1",
         10232 => x"3f7a5afd",
         10233 => x"a0398154",
         10234 => x"b4170853",
         10235 => x"b8177053",
         10236 => x"81183352",
         10237 => x"5ef4da3f",
         10238 => x"815a84b8",
         10239 => x"e4087d2e",
         10240 => x"098106fb",
         10241 => x"cb3884b8",
         10242 => x"e4088318",
         10243 => x"34b41708",
         10244 => x"a8180831",
         10245 => x"84b8e408",
         10246 => x"5b5574a0",
         10247 => x"180827fb",
         10248 => x"91388217",
         10249 => x"33557482",
         10250 => x"2e098106",
         10251 => x"fb843881",
         10252 => x"54b41708",
         10253 => x"a0180805",
         10254 => x"537d5281",
         10255 => x"173351f4",
         10256 => x"903f7c5a",
         10257 => x"faec3981",
         10258 => x"54b41708",
         10259 => x"a0180805",
         10260 => x"537b5281",
         10261 => x"173351f3",
         10262 => x"f83ffa86",
         10263 => x"39815b7a",
         10264 => x"f9bb38fa",
         10265 => x"9f39f23d",
         10266 => x"0d606264",
         10267 => x"5d575982",
         10268 => x"58817627",
         10269 => x"9c38759c",
         10270 => x"1a082795",
         10271 => x"38783355",
         10272 => x"74782e96",
         10273 => x"38747824",
         10274 => x"81803874",
         10275 => x"812e828a",
         10276 => x"387784b8",
         10277 => x"e40c903d",
         10278 => x"0d047588",
         10279 => x"2aa81a08",
         10280 => x"0558800b",
         10281 => x"b41a0858",
         10282 => x"5c76782e",
         10283 => x"86b63883",
         10284 => x"19337c5b",
         10285 => x"5d7c7c2e",
         10286 => x"09810683",
         10287 => x"fa388154",
         10288 => x"7753b819",
         10289 => x"52811933",
         10290 => x"51f2873f",
         10291 => x"84b8e408",
         10292 => x"802e8538",
         10293 => x"ff58815a",
         10294 => x"77b41a0c",
         10295 => x"795879ff",
         10296 => x"b0387510",
         10297 => x"83fe0679",
         10298 => x"057b83ff",
         10299 => x"ff06585e",
         10300 => x"76b81f34",
         10301 => x"76882a5a",
         10302 => x"79b91f34",
         10303 => x"810b831a",
         10304 => x"347784b8",
         10305 => x"e40c903d",
         10306 => x"0d047483",
         10307 => x"2e098106",
         10308 => x"feff3875",
         10309 => x"872aa81a",
         10310 => x"08055880",
         10311 => x"0bb41a08",
         10312 => x"585c7678",
         10313 => x"2e85e138",
         10314 => x"8319337c",
         10315 => x"5b5d7c7c",
         10316 => x"2e098106",
         10317 => x"84bd3881",
         10318 => x"547753b8",
         10319 => x"19528119",
         10320 => x"3351f18e",
         10321 => x"3f84b8e4",
         10322 => x"08802e85",
         10323 => x"38ff5881",
         10324 => x"5a77b41a",
         10325 => x"0c795879",
         10326 => x"feb73875",
         10327 => x"822b83fc",
         10328 => x"067905b8",
         10329 => x"11831133",
         10330 => x"70982b8f",
         10331 => x"0a067ef0",
         10332 => x"0a060741",
         10333 => x"575e5c7d",
         10334 => x"7d347d88",
         10335 => x"2a5675b9",
         10336 => x"1d347d90",
         10337 => x"2a5a79ba",
         10338 => x"1d347d98",
         10339 => x"2a5b7abb",
         10340 => x"1d34810b",
         10341 => x"831a34fe",
         10342 => x"e8397581",
         10343 => x"2a167089",
         10344 => x"2aa81b08",
         10345 => x"05b41b08",
         10346 => x"59595a76",
         10347 => x"782eb738",
         10348 => x"800b831a",
         10349 => x"33715e56",
         10350 => x"5d747d2e",
         10351 => x"09810682",
         10352 => x"d4388154",
         10353 => x"7753b819",
         10354 => x"52811933",
         10355 => x"51f0833f",
         10356 => x"84b8e408",
         10357 => x"802e8538",
         10358 => x"ff58815c",
         10359 => x"77b41a0c",
         10360 => x"7b587bfd",
         10361 => x"ac387983",
         10362 => x"ff0619b8",
         10363 => x"05811b77",
         10364 => x"81065f5f",
         10365 => x"577a557c",
         10366 => x"802e8f38",
         10367 => x"7a842b9f",
         10368 => x"f0067733",
         10369 => x"8f067107",
         10370 => x"565a7477",
         10371 => x"34810b83",
         10372 => x"1a347d89",
         10373 => x"2aa81a08",
         10374 => x"0556800b",
         10375 => x"b41a0856",
         10376 => x"5f74762e",
         10377 => x"83dd3881",
         10378 => x"547453b8",
         10379 => x"19705381",
         10380 => x"1a335257",
         10381 => x"f09b3f81",
         10382 => x"5884b8e4",
         10383 => x"087f2e09",
         10384 => x"810680c7",
         10385 => x"3884b8e4",
         10386 => x"08831a34",
         10387 => x"b4190870",
         10388 => x"a81b0831",
         10389 => x"a01b0884",
         10390 => x"b8e4085b",
         10391 => x"5c565c74",
         10392 => x"7a278b38",
         10393 => x"82193355",
         10394 => x"74822e82",
         10395 => x"e4388154",
         10396 => x"75537652",
         10397 => x"81193351",
         10398 => x"eed83f84",
         10399 => x"b8e40880",
         10400 => x"2e8538ff",
         10401 => x"56815875",
         10402 => x"b41a0c77",
         10403 => x"fc83387d",
         10404 => x"83ff0619",
         10405 => x"b8057b84",
         10406 => x"2a56567c",
         10407 => x"8f387a88",
         10408 => x"2a763381",
         10409 => x"f006718f",
         10410 => x"0607565c",
         10411 => x"74763481",
         10412 => x"0b831a34",
         10413 => x"fccb3981",
         10414 => x"547653b8",
         10415 => x"19705381",
         10416 => x"1a33525d",
         10417 => x"ef8b3f81",
         10418 => x"5a84b8e4",
         10419 => x"087c2e09",
         10420 => x"8106fc88",
         10421 => x"3884b8e4",
         10422 => x"08831a34",
         10423 => x"b4190870",
         10424 => x"a81b0831",
         10425 => x"a01b0884",
         10426 => x"b8e4085d",
         10427 => x"59405e7e",
         10428 => x"7727fbca",
         10429 => x"38821933",
         10430 => x"5574822e",
         10431 => x"098106fb",
         10432 => x"bd388154",
         10433 => x"761e537c",
         10434 => x"52811933",
         10435 => x"51eec23f",
         10436 => x"7b5afbaa",
         10437 => x"39815476",
         10438 => x"53b81970",
         10439 => x"53811a33",
         10440 => x"5257eead",
         10441 => x"3f815c84",
         10442 => x"b8e4087d",
         10443 => x"2e098106",
         10444 => x"fdae3884",
         10445 => x"b8e40883",
         10446 => x"1a34b419",
         10447 => x"0870a81b",
         10448 => x"0831a01b",
         10449 => x"0884b8e4",
         10450 => x"085f4056",
         10451 => x"5f747e27",
         10452 => x"fcf03882",
         10453 => x"19335574",
         10454 => x"822e0981",
         10455 => x"06fce338",
         10456 => x"81547d1f",
         10457 => x"53765281",
         10458 => x"193351ed",
         10459 => x"e43f7c5c",
         10460 => x"fcd03981",
         10461 => x"547653b8",
         10462 => x"19705381",
         10463 => x"1a335257",
         10464 => x"edcf3f81",
         10465 => x"5a84b8e4",
         10466 => x"087c2e09",
         10467 => x"8106fbc5",
         10468 => x"3884b8e4",
         10469 => x"08831a34",
         10470 => x"b4190870",
         10471 => x"a81b0831",
         10472 => x"a01b0884",
         10473 => x"b8e4085d",
         10474 => x"5f405e7e",
         10475 => x"7d27fb87",
         10476 => x"38821933",
         10477 => x"5574822e",
         10478 => x"098106fa",
         10479 => x"fa388154",
         10480 => x"7c1e5376",
         10481 => x"52811933",
         10482 => x"51ed863f",
         10483 => x"7b5afae7",
         10484 => x"39815479",
         10485 => x"1c537652",
         10486 => x"81193351",
         10487 => x"ecf33f7e",
         10488 => x"58fd8b39",
         10489 => x"7b761083",
         10490 => x"fe067a05",
         10491 => x"7c83ffff",
         10492 => x"06595f58",
         10493 => x"76b81f34",
         10494 => x"76882a5a",
         10495 => x"79b91f34",
         10496 => x"f9fa397e",
         10497 => x"58fd8839",
         10498 => x"7b76822b",
         10499 => x"83fc067a",
         10500 => x"05b81183",
         10501 => x"11337098",
         10502 => x"2b8f0a06",
         10503 => x"7ff00a06",
         10504 => x"0742585f",
         10505 => x"5d587d7d",
         10506 => x"347d882a",
         10507 => x"5675b91d",
         10508 => x"347d902a",
         10509 => x"5a79ba1d",
         10510 => x"347d982a",
         10511 => x"5b7abb1d",
         10512 => x"34facf39",
         10513 => x"f63d0d7c",
         10514 => x"7e71085b",
         10515 => x"5c5a7a81",
         10516 => x"8a389019",
         10517 => x"08577680",
         10518 => x"2e80f438",
         10519 => x"769c1a08",
         10520 => x"2780ec38",
         10521 => x"94190870",
         10522 => x"56547380",
         10523 => x"2e80d738",
         10524 => x"767b2e81",
         10525 => x"93387656",
         10526 => x"8116569c",
         10527 => x"19087626",
         10528 => x"89388256",
         10529 => x"75772682",
         10530 => x"b2387552",
         10531 => x"7951f0f5",
         10532 => x"3f84b8e4",
         10533 => x"08802e81",
         10534 => x"d0388058",
         10535 => x"84b8e408",
         10536 => x"812eb138",
         10537 => x"84b8e408",
         10538 => x"09703070",
         10539 => x"72078025",
         10540 => x"707b0751",
         10541 => x"51555573",
         10542 => x"82aa3875",
         10543 => x"772e0981",
         10544 => x"06ffb538",
         10545 => x"73557484",
         10546 => x"b8e40c8c",
         10547 => x"3d0d0481",
         10548 => x"57ff9139",
         10549 => x"84b8e408",
         10550 => x"58ca397a",
         10551 => x"527951f0",
         10552 => x"a43f8155",
         10553 => x"7484b8e4",
         10554 => x"0827db38",
         10555 => x"84b8e408",
         10556 => x"5584b8e4",
         10557 => x"08ff2ece",
         10558 => x"389c1908",
         10559 => x"84b8e408",
         10560 => x"26c4387a",
         10561 => x"57fedd39",
         10562 => x"811b569c",
         10563 => x"19087626",
         10564 => x"83388256",
         10565 => x"75527951",
         10566 => x"efeb3f80",
         10567 => x"5884b8e4",
         10568 => x"08812e81",
         10569 => x"a03884b8",
         10570 => x"e4080970",
         10571 => x"30707207",
         10572 => x"8025707b",
         10573 => x"0784b8e4",
         10574 => x"08545151",
         10575 => x"555573ff",
         10576 => x"853884b8",
         10577 => x"e408802e",
         10578 => x"9a389019",
         10579 => x"08548174",
         10580 => x"27fea338",
         10581 => x"739c1a08",
         10582 => x"27fe9b38",
         10583 => x"73705757",
         10584 => x"fe963975",
         10585 => x"802efe8e",
         10586 => x"38ff5375",
         10587 => x"527851f5",
         10588 => x"f53f84b8",
         10589 => x"e40884b8",
         10590 => x"e4083070",
         10591 => x"84b8e408",
         10592 => x"07802556",
         10593 => x"58557a80",
         10594 => x"c4387480",
         10595 => x"e3387590",
         10596 => x"1a0c9c19",
         10597 => x"08fe0594",
         10598 => x"1a085658",
         10599 => x"74782686",
         10600 => x"38ff1594",
         10601 => x"1a0c8419",
         10602 => x"3381075a",
         10603 => x"79841a34",
         10604 => x"75557484",
         10605 => x"b8e40c8c",
         10606 => x"3d0d0480",
         10607 => x"0b84b8e4",
         10608 => x"0c8c3d0d",
         10609 => x"0484b8e4",
         10610 => x"0858feda",
         10611 => x"3973802e",
         10612 => x"ffb83875",
         10613 => x"537a5278",
         10614 => x"51f58b3f",
         10615 => x"84b8e408",
         10616 => x"55ffa739",
         10617 => x"84b8e408",
         10618 => x"84b8e40c",
         10619 => x"8c3d0d04",
         10620 => x"ff567481",
         10621 => x"2effb938",
         10622 => x"8155ffb6",
         10623 => x"39f83d0d",
         10624 => x"7a7c7108",
         10625 => x"59555873",
         10626 => x"f0800a26",
         10627 => x"80df3873",
         10628 => x"9f065372",
         10629 => x"80d73873",
         10630 => x"90190c88",
         10631 => x"18085574",
         10632 => x"80df3876",
         10633 => x"33567582",
         10634 => x"2680cc38",
         10635 => x"73852a53",
         10636 => x"820b8818",
         10637 => x"225a5672",
         10638 => x"7927a938",
         10639 => x"ac170898",
         10640 => x"190c7494",
         10641 => x"190c9818",
         10642 => x"08538256",
         10643 => x"72802e94",
         10644 => x"3873892a",
         10645 => x"1398190c",
         10646 => x"7383ff06",
         10647 => x"17b8059c",
         10648 => x"190c8056",
         10649 => x"7584b8e4",
         10650 => x"0c8a3d0d",
         10651 => x"04820b84",
         10652 => x"b8e40c8a",
         10653 => x"3d0d04ac",
         10654 => x"17085574",
         10655 => x"802effac",
         10656 => x"388a1722",
         10657 => x"70892b57",
         10658 => x"59737627",
         10659 => x"a5389c17",
         10660 => x"0853fe15",
         10661 => x"fe145456",
         10662 => x"80597573",
         10663 => x"278d388a",
         10664 => x"17227671",
         10665 => x"29b01908",
         10666 => x"055a5378",
         10667 => x"98190cff",
         10668 => x"91397452",
         10669 => x"7751eccd",
         10670 => x"3f84b8e4",
         10671 => x"085584b8",
         10672 => x"e408ff2e",
         10673 => x"a438810b",
         10674 => x"84b8e408",
         10675 => x"27ff9e38",
         10676 => x"9c170853",
         10677 => x"84b8e408",
         10678 => x"7327ff91",
         10679 => x"38737631",
         10680 => x"54737627",
         10681 => x"cd38ffaa",
         10682 => x"39810b84",
         10683 => x"b8e40c8a",
         10684 => x"3d0d04f3",
         10685 => x"3d0d7f70",
         10686 => x"08901208",
         10687 => x"a0055c5a",
         10688 => x"57f0800a",
         10689 => x"7a278638",
         10690 => x"800b9818",
         10691 => x"0c981708",
         10692 => x"55845674",
         10693 => x"802eb238",
         10694 => x"7983ff06",
         10695 => x"5b7a9d38",
         10696 => x"81159418",
         10697 => x"08575875",
         10698 => x"a9387985",
         10699 => x"2a881a22",
         10700 => x"57557476",
         10701 => x"2781f538",
         10702 => x"7798180c",
         10703 => x"7990180c",
         10704 => x"781bb805",
         10705 => x"9c180c80",
         10706 => x"567584b8",
         10707 => x"e40c8f3d",
         10708 => x"0d047798",
         10709 => x"180c8a19",
         10710 => x"22ff057a",
         10711 => x"892a065c",
         10712 => x"7bda3875",
         10713 => x"527651eb",
         10714 => x"9c3f84b8",
         10715 => x"e4085d82",
         10716 => x"56810b84",
         10717 => x"b8e40827",
         10718 => x"d0388156",
         10719 => x"84b8e408",
         10720 => x"ff2ec638",
         10721 => x"9c190884",
         10722 => x"b8e40826",
         10723 => x"82913860",
         10724 => x"802e8198",
         10725 => x"38941708",
         10726 => x"527651f9",
         10727 => x"a73f84b8",
         10728 => x"e4085d87",
         10729 => x"5684b8e4",
         10730 => x"08802eff",
         10731 => x"9c388256",
         10732 => x"84b8e408",
         10733 => x"812eff91",
         10734 => x"38815684",
         10735 => x"b8e408ff",
         10736 => x"2eff8638",
         10737 => x"84b8e408",
         10738 => x"831a335f",
         10739 => x"587d80ea",
         10740 => x"38fe189c",
         10741 => x"1a08fe05",
         10742 => x"5956805c",
         10743 => x"7578278d",
         10744 => x"388a1922",
         10745 => x"767129b0",
         10746 => x"1b08055d",
         10747 => x"5e7bb41a",
         10748 => x"0cb81958",
         10749 => x"84807857",
         10750 => x"55807670",
         10751 => x"81055834",
         10752 => x"ff155574",
         10753 => x"f4387456",
         10754 => x"8a192255",
         10755 => x"75752781",
         10756 => x"80388154",
         10757 => x"751c5377",
         10758 => x"52811933",
         10759 => x"51e4b23f",
         10760 => x"84b8e408",
         10761 => x"80e73881",
         10762 => x"1656dd39",
         10763 => x"7a98180c",
         10764 => x"840b84b8",
         10765 => x"e40c8f3d",
         10766 => x"0d047554",
         10767 => x"b4190853",
         10768 => x"b8197053",
         10769 => x"811a3352",
         10770 => x"56e4863f",
         10771 => x"84b8e408",
         10772 => x"80f33884",
         10773 => x"b8e40883",
         10774 => x"1a34b419",
         10775 => x"08a81a08",
         10776 => x"315574a0",
         10777 => x"1a0827fe",
         10778 => x"e8388219",
         10779 => x"335c7b82",
         10780 => x"2e098106",
         10781 => x"fedb3881",
         10782 => x"54b41908",
         10783 => x"a01a0805",
         10784 => x"53755281",
         10785 => x"193351e3",
         10786 => x"c83ffec5",
         10787 => x"398a1922",
         10788 => x"557483ff",
         10789 => x"ff065574",
         10790 => x"762e0981",
         10791 => x"06a7387c",
         10792 => x"94180cfe",
         10793 => x"1d9c1a08",
         10794 => x"fe055e56",
         10795 => x"8058757d",
         10796 => x"27fd8538",
         10797 => x"8a192276",
         10798 => x"7129b01b",
         10799 => x"08059819",
         10800 => x"0c5cfcf8",
         10801 => x"39810b84",
         10802 => x"b8e40c8f",
         10803 => x"3d0d04ee",
         10804 => x"3d0d6466",
         10805 => x"415c847c",
         10806 => x"085a5b81",
         10807 => x"ff70981e",
         10808 => x"08585e5e",
         10809 => x"75802e82",
         10810 => x"d238b819",
         10811 => x"5f755a80",
         10812 => x"58b41908",
         10813 => x"762e82d1",
         10814 => x"38831933",
         10815 => x"78585574",
         10816 => x"782e0981",
         10817 => x"06819438",
         10818 => x"81547553",
         10819 => x"b8195281",
         10820 => x"193351e1",
         10821 => x"bd3f84b8",
         10822 => x"e408802e",
         10823 => x"8538ff5a",
         10824 => x"815779b4",
         10825 => x"1a0c765b",
         10826 => x"76829038",
         10827 => x"9c1c0870",
         10828 => x"33585876",
         10829 => x"802e8281",
         10830 => x"388b1833",
         10831 => x"bf067081",
         10832 => x"ff065b41",
         10833 => x"60861d34",
         10834 => x"7681e532",
         10835 => x"703078ae",
         10836 => x"32703072",
         10837 => x"80257180",
         10838 => x"25075445",
         10839 => x"45575574",
         10840 => x"9338747a",
         10841 => x"df064356",
         10842 => x"61882e81",
         10843 => x"bf387560",
         10844 => x"2e818638",
         10845 => x"81ff5d80",
         10846 => x"527b51fa",
         10847 => x"f63f84b8",
         10848 => x"e4085b84",
         10849 => x"b8e40881",
         10850 => x"b238981c",
         10851 => x"085675fe",
         10852 => x"dc387a84",
         10853 => x"b8e40c94",
         10854 => x"3d0d0481",
         10855 => x"54b41908",
         10856 => x"537e5281",
         10857 => x"193351e1",
         10858 => x"a83f8157",
         10859 => x"84b8e408",
         10860 => x"782e0981",
         10861 => x"06feef38",
         10862 => x"84b8e408",
         10863 => x"831a34b4",
         10864 => x"1908a81a",
         10865 => x"083184b8",
         10866 => x"e408585b",
         10867 => x"7aa01a08",
         10868 => x"27feb538",
         10869 => x"82193341",
         10870 => x"60822e09",
         10871 => x"8106fea8",
         10872 => x"388154b4",
         10873 => x"1908a01a",
         10874 => x"0805537e",
         10875 => x"52811933",
         10876 => x"51e0de3f",
         10877 => x"7757fe90",
         10878 => x"39798f2e",
         10879 => x"09810681",
         10880 => x"e7387686",
         10881 => x"2a81065b",
         10882 => x"7a802e93",
         10883 => x"388d1833",
         10884 => x"7781bf06",
         10885 => x"70901f08",
         10886 => x"7fac050c",
         10887 => x"595e5e76",
         10888 => x"7d2eab38",
         10889 => x"81ff5574",
         10890 => x"5dfecc39",
         10891 => x"81567560",
         10892 => x"2e098106",
         10893 => x"febe38c1",
         10894 => x"39845b80",
         10895 => x"0b981d0c",
         10896 => x"7a84b8e4",
         10897 => x"0c943d0d",
         10898 => x"04775bfd",
         10899 => x"df398d18",
         10900 => x"33577d77",
         10901 => x"2e098106",
         10902 => x"cb388c19",
         10903 => x"089b1933",
         10904 => x"9a1a3371",
         10905 => x"882b0758",
         10906 => x"564175ff",
         10907 => x"b7387733",
         10908 => x"7081bf06",
         10909 => x"8d29f305",
         10910 => x"515a8176",
         10911 => x"585b83e4",
         10912 => x"e4173378",
         10913 => x"05811133",
         10914 => x"71337188",
         10915 => x"2b075244",
         10916 => x"567a802e",
         10917 => x"80c53879",
         10918 => x"81fe26ff",
         10919 => x"87387910",
         10920 => x"6105765c",
         10921 => x"42756223",
         10922 => x"811a5a81",
         10923 => x"17578c77",
         10924 => x"27cc3877",
         10925 => x"3370862a",
         10926 => x"81065957",
         10927 => x"77802e90",
         10928 => x"387981fe",
         10929 => x"26fedd38",
         10930 => x"79106105",
         10931 => x"43806323",
         10932 => x"ff1d7081",
         10933 => x"ff065e41",
         10934 => x"fd9d3975",
         10935 => x"83ffff2e",
         10936 => x"ca3881ff",
         10937 => x"55fec039",
         10938 => x"7ca8387c",
         10939 => x"558b5774",
         10940 => x"812a7581",
         10941 => x"80290578",
         10942 => x"7081055a",
         10943 => x"33407f05",
         10944 => x"7081ff06",
         10945 => x"ff195956",
         10946 => x"5976e438",
         10947 => x"747e2efd",
         10948 => x"8138ff0b",
         10949 => x"ac1d0c7a",
         10950 => x"84b8e40c",
         10951 => x"943d0d04",
         10952 => x"ef3d0d63",
         10953 => x"70085c5c",
         10954 => x"80527b51",
         10955 => x"f5cf3f84",
         10956 => x"b8e4085a",
         10957 => x"84b8e408",
         10958 => x"82803881",
         10959 => x"ff70405d",
         10960 => x"ff0bac1d",
         10961 => x"0cb81b5e",
         10962 => x"981c0856",
         10963 => x"8058b41b",
         10964 => x"08762e82",
         10965 => x"cc38831b",
         10966 => x"33785855",
         10967 => x"74782e09",
         10968 => x"810681df",
         10969 => x"38815475",
         10970 => x"53b81b52",
         10971 => x"811b3351",
         10972 => x"dce03f84",
         10973 => x"b8e40880",
         10974 => x"2e8538ff",
         10975 => x"56815775",
         10976 => x"b41c0c76",
         10977 => x"5a7681b2",
         10978 => x"389c1c08",
         10979 => x"70335859",
         10980 => x"76802e84",
         10981 => x"99388b19",
         10982 => x"33bf0670",
         10983 => x"81ff0657",
         10984 => x"5877861d",
         10985 => x"347681e5",
         10986 => x"2e80f238",
         10987 => x"75832a81",
         10988 => x"0655758f",
         10989 => x"2e81ef38",
         10990 => x"7480e238",
         10991 => x"758f2e81",
         10992 => x"e5387caa",
         10993 => x"38787d56",
         10994 => x"588b5774",
         10995 => x"812a7581",
         10996 => x"80290578",
         10997 => x"7081055a",
         10998 => x"33577605",
         10999 => x"7081ff06",
         11000 => x"ff195956",
         11001 => x"5d76e438",
         11002 => x"747f2e80",
         11003 => x"cd38ab1c",
         11004 => x"33810657",
         11005 => x"76a7388b",
         11006 => x"0ba01d59",
         11007 => x"57787081",
         11008 => x"055a3378",
         11009 => x"7081055a",
         11010 => x"33717131",
         11011 => x"ff1a5a58",
         11012 => x"42407680",
         11013 => x"2e81dc38",
         11014 => x"75802ee1",
         11015 => x"3881ff5d",
         11016 => x"ff0bac1d",
         11017 => x"0c80527b",
         11018 => x"51f5c83f",
         11019 => x"84b8e408",
         11020 => x"5a84b8e4",
         11021 => x"08802efe",
         11022 => x"8f387984",
         11023 => x"b8e40c93",
         11024 => x"3d0d0481",
         11025 => x"54b41b08",
         11026 => x"537d5281",
         11027 => x"1b3351dc",
         11028 => x"803f8157",
         11029 => x"84b8e408",
         11030 => x"782e0981",
         11031 => x"06fea438",
         11032 => x"84b8e408",
         11033 => x"831c34b4",
         11034 => x"1b08a81c",
         11035 => x"083184b8",
         11036 => x"e4085859",
         11037 => x"78a01c08",
         11038 => x"27fdea38",
         11039 => x"821b335a",
         11040 => x"79822e09",
         11041 => x"8106fddd",
         11042 => x"388154b4",
         11043 => x"1b08a01c",
         11044 => x"0805537d",
         11045 => x"52811b33",
         11046 => x"51dbb63f",
         11047 => x"7757fdc5",
         11048 => x"39775afd",
         11049 => x"e439ab1c",
         11050 => x"3370862a",
         11051 => x"81064255",
         11052 => x"60fef238",
         11053 => x"76862a81",
         11054 => x"065a7980",
         11055 => x"2e93388d",
         11056 => x"19337781",
         11057 => x"bf067090",
         11058 => x"1f087fac",
         11059 => x"050c595e",
         11060 => x"5f767d2e",
         11061 => x"af3881ff",
         11062 => x"55745d80",
         11063 => x"527b51f4",
         11064 => x"923f84b8",
         11065 => x"e4085a84",
         11066 => x"b8e40880",
         11067 => x"2efcd938",
         11068 => x"fec83975",
         11069 => x"802efec2",
         11070 => x"3881ff5d",
         11071 => x"ff0bac1d",
         11072 => x"0cfea239",
         11073 => x"8d193357",
         11074 => x"7e772e09",
         11075 => x"8106c738",
         11076 => x"8c1b089b",
         11077 => x"1a339a1b",
         11078 => x"3371882b",
         11079 => x"07594240",
         11080 => x"76ffb338",
         11081 => x"783370bf",
         11082 => x"068d29f3",
         11083 => x"055b5581",
         11084 => x"77595683",
         11085 => x"e4e41833",
         11086 => x"79058111",
         11087 => x"33713371",
         11088 => x"882b0752",
         11089 => x"42577580",
         11090 => x"2e80ed38",
         11091 => x"7981fe26",
         11092 => x"ff843876",
         11093 => x"5181a18a",
         11094 => x"3f84b8e4",
         11095 => x"087a1061",
         11096 => x"05702253",
         11097 => x"43811b5b",
         11098 => x"5681a0f6",
         11099 => x"3f7584b8",
         11100 => x"e4082e09",
         11101 => x"8106fede",
         11102 => x"38765681",
         11103 => x"18588c78",
         11104 => x"27ffb038",
         11105 => x"78337086",
         11106 => x"2a810656",
         11107 => x"5975802e",
         11108 => x"92387480",
         11109 => x"2e8d3879",
         11110 => x"10600570",
         11111 => x"2241417f",
         11112 => x"feb438ff",
         11113 => x"1d7081ff",
         11114 => x"065e5afe",
         11115 => x"ae39840b",
         11116 => x"84b8e40c",
         11117 => x"933d0d04",
         11118 => x"7683ffff",
         11119 => x"2effbc38",
         11120 => x"81ff55fe",
         11121 => x"9439ea3d",
         11122 => x"0d687008",
         11123 => x"70ab1333",
         11124 => x"81a00658",
         11125 => x"5a5d5e86",
         11126 => x"567485b5",
         11127 => x"38748c1d",
         11128 => x"08702257",
         11129 => x"575d7480",
         11130 => x"2e8e3881",
         11131 => x"1d701017",
         11132 => x"70225156",
         11133 => x"5d74f438",
         11134 => x"953da01f",
         11135 => x"5b408c60",
         11136 => x"7b585855",
         11137 => x"75708105",
         11138 => x"57337770",
         11139 => x"81055934",
         11140 => x"ff155574",
         11141 => x"ef380280",
         11142 => x"db053370",
         11143 => x"81065856",
         11144 => x"76802e82",
         11145 => x"aa3880c0",
         11146 => x"0bab1f34",
         11147 => x"810b943d",
         11148 => x"405b8c1c",
         11149 => x"087b5859",
         11150 => x"8b7a615a",
         11151 => x"57557770",
         11152 => x"81055933",
         11153 => x"76708105",
         11154 => x"5834ff15",
         11155 => x"5574ef38",
         11156 => x"857b2780",
         11157 => x"c2387a79",
         11158 => x"22565774",
         11159 => x"802eb838",
         11160 => x"74821a5a",
         11161 => x"568f5875",
         11162 => x"81067710",
         11163 => x"0776812a",
         11164 => x"7083ffff",
         11165 => x"0672902a",
         11166 => x"81064458",
         11167 => x"56576080",
         11168 => x"2e873876",
         11169 => x"84a0a132",
         11170 => x"57ff1858",
         11171 => x"778025d7",
         11172 => x"38782255",
         11173 => x"74ca3887",
         11174 => x"02840580",
         11175 => x"cf055758",
         11176 => x"76b007bf",
         11177 => x"0655b975",
         11178 => x"27843887",
         11179 => x"15557476",
         11180 => x"34ff16ff",
         11181 => x"1978842a",
         11182 => x"59595676",
         11183 => x"e338771f",
         11184 => x"5980fe79",
         11185 => x"34767a58",
         11186 => x"56807827",
         11187 => x"a0387933",
         11188 => x"5574a02e",
         11189 => x"98388116",
         11190 => x"56757827",
         11191 => x"88a23875",
         11192 => x"1a703356",
         11193 => x"5774a02e",
         11194 => x"098106ea",
         11195 => x"38811656",
         11196 => x"a0557787",
         11197 => x"268e3898",
         11198 => x"3d7805ec",
         11199 => x"05811971",
         11200 => x"33575941",
         11201 => x"74773487",
         11202 => x"762787f4",
         11203 => x"387d51f8",
         11204 => x"8f3f84b8",
         11205 => x"e4088b38",
         11206 => x"811b5b80",
         11207 => x"e37b27fe",
         11208 => x"91388756",
         11209 => x"7a80e42e",
         11210 => x"82e73884",
         11211 => x"b8e40856",
         11212 => x"84b8e408",
         11213 => x"842e0981",
         11214 => x"0682d638",
         11215 => x"0280db05",
         11216 => x"33ab1f34",
         11217 => x"7d080284",
         11218 => x"0580db05",
         11219 => x"33575875",
         11220 => x"812a8106",
         11221 => x"5f815b7e",
         11222 => x"802e9038",
         11223 => x"8d528c1d",
         11224 => x"51fe8ac1",
         11225 => x"3f84b8e4",
         11226 => x"081b5b80",
         11227 => x"527d51ed",
         11228 => x"8c3f84b8",
         11229 => x"e4085684",
         11230 => x"b8e40881",
         11231 => x"823884b8",
         11232 => x"e408b819",
         11233 => x"5e59981e",
         11234 => x"08568057",
         11235 => x"b4180876",
         11236 => x"2e85f338",
         11237 => x"83183340",
         11238 => x"7f772e09",
         11239 => x"810682a3",
         11240 => x"38815475",
         11241 => x"53b81852",
         11242 => x"81183351",
         11243 => x"d4a43f84",
         11244 => x"b8e40880",
         11245 => x"2e8538ff",
         11246 => x"56815775",
         11247 => x"b4190c76",
         11248 => x"5676bc38",
         11249 => x"9c1e0870",
         11250 => x"33564274",
         11251 => x"81e52e81",
         11252 => x"c9387430",
         11253 => x"70802578",
         11254 => x"07565f74",
         11255 => x"802e81c9",
         11256 => x"38811959",
         11257 => x"787b2e86",
         11258 => x"89388152",
         11259 => x"7d51ee83",
         11260 => x"3f84b8e4",
         11261 => x"085684b8",
         11262 => x"e408802e",
         11263 => x"ff883887",
         11264 => x"5875842e",
         11265 => x"81893875",
         11266 => x"58758183",
         11267 => x"38ff1b40",
         11268 => x"7f81f338",
         11269 => x"981e0857",
         11270 => x"b41c0877",
         11271 => x"2eaf3883",
         11272 => x"1c337857",
         11273 => x"407f8482",
         11274 => x"38815476",
         11275 => x"53b81c52",
         11276 => x"811c3351",
         11277 => x"d39c3f84",
         11278 => x"b8e40880",
         11279 => x"2e8538ff",
         11280 => x"57815676",
         11281 => x"b41d0c75",
         11282 => x"587580c3",
         11283 => x"38a00b9c",
         11284 => x"1f085755",
         11285 => x"80767081",
         11286 => x"055834ff",
         11287 => x"155574f4",
         11288 => x"388b0b9c",
         11289 => x"1f087b58",
         11290 => x"58557570",
         11291 => x"81055733",
         11292 => x"77708105",
         11293 => x"5934ff15",
         11294 => x"5574ef38",
         11295 => x"9c1e08ab",
         11296 => x"1f339806",
         11297 => x"5e5a7c8c",
         11298 => x"1b34810b",
         11299 => x"831d3477",
         11300 => x"567584b8",
         11301 => x"e40c983d",
         11302 => x"0d048175",
         11303 => x"30708025",
         11304 => x"72075740",
         11305 => x"5774feb9",
         11306 => x"38745981",
         11307 => x"527d51ec",
         11308 => x"c23f84b8",
         11309 => x"e4085684",
         11310 => x"b8e40880",
         11311 => x"2efdc738",
         11312 => x"febd3981",
         11313 => x"54b41808",
         11314 => x"537c5281",
         11315 => x"183351d3",
         11316 => x"803f84b8",
         11317 => x"e408772e",
         11318 => x"09810683",
         11319 => x"bf3884b8",
         11320 => x"e4088319",
         11321 => x"34b41808",
         11322 => x"a8190831",
         11323 => x"5574a019",
         11324 => x"08278b38",
         11325 => x"82183341",
         11326 => x"60822e84",
         11327 => x"ac3884b8",
         11328 => x"e40857fd",
         11329 => x"9c397f85",
         11330 => x"2b901f08",
         11331 => x"71315358",
         11332 => x"7d51e9e9",
         11333 => x"3f84b8e4",
         11334 => x"085884b8",
         11335 => x"e408feef",
         11336 => x"387984b8",
         11337 => x"e4085658",
         11338 => x"8b577481",
         11339 => x"2a758180",
         11340 => x"29057870",
         11341 => x"81055a33",
         11342 => x"57760570",
         11343 => x"81ff06ff",
         11344 => x"1959565d",
         11345 => x"76e43874",
         11346 => x"81ff06b8",
         11347 => x"1d434198",
         11348 => x"1e085780",
         11349 => x"56b41c08",
         11350 => x"772eb238",
         11351 => x"831c335b",
         11352 => x"7a762e09",
         11353 => x"810682c9",
         11354 => x"38815476",
         11355 => x"53b81c52",
         11356 => x"811c3351",
         11357 => x"d0dc3f84",
         11358 => x"b8e40880",
         11359 => x"2e8538ff",
         11360 => x"57815676",
         11361 => x"b41d0c75",
         11362 => x"5875fe83",
         11363 => x"388c1c08",
         11364 => x"9c1f0861",
         11365 => x"81ff065f",
         11366 => x"5c5f608d",
         11367 => x"1c348f0b",
         11368 => x"8b1c3475",
         11369 => x"8c1c3475",
         11370 => x"9a1c3475",
         11371 => x"9b1c347c",
         11372 => x"8d29f305",
         11373 => x"76775a58",
         11374 => x"597683ff",
         11375 => x"ff2e8b38",
         11376 => x"78101f70",
         11377 => x"22811b5b",
         11378 => x"585683e4",
         11379 => x"e418337b",
         11380 => x"05557675",
         11381 => x"70810557",
         11382 => x"3476882a",
         11383 => x"56757534",
         11384 => x"76853883",
         11385 => x"ffff5781",
         11386 => x"18588c78",
         11387 => x"27cb3876",
         11388 => x"83ffff2e",
         11389 => x"81b33878",
         11390 => x"101f7022",
         11391 => x"58587680",
         11392 => x"2e81a638",
         11393 => x"7c7b3481",
         11394 => x"0b831d34",
         11395 => x"80527d51",
         11396 => x"e9e13f84",
         11397 => x"b8e40858",
         11398 => x"84b8e408",
         11399 => x"fcf1387f",
         11400 => x"ff05407f",
         11401 => x"fea938fb",
         11402 => x"eb398154",
         11403 => x"b41c0853",
         11404 => x"b81c7053",
         11405 => x"811d3352",
         11406 => x"59d0963f",
         11407 => x"815684b8",
         11408 => x"e408fc83",
         11409 => x"3884b8e4",
         11410 => x"08831d34",
         11411 => x"b41c08a8",
         11412 => x"1d083184",
         11413 => x"b8e40857",
         11414 => x"4160a01d",
         11415 => x"0827fbc9",
         11416 => x"38821c33",
         11417 => x"4261822e",
         11418 => x"098106fb",
         11419 => x"bc388154",
         11420 => x"b41c08a0",
         11421 => x"1d080553",
         11422 => x"7852811c",
         11423 => x"3351cfd1",
         11424 => x"3f7756fb",
         11425 => x"a439769c",
         11426 => x"1f087033",
         11427 => x"57435674",
         11428 => x"81e52e09",
         11429 => x"8106faba",
         11430 => x"38fbff39",
         11431 => x"81705757",
         11432 => x"76802efa",
         11433 => x"9f38fad7",
         11434 => x"397c80c0",
         11435 => x"075dfed4",
         11436 => x"398154b4",
         11437 => x"1c085361",
         11438 => x"52811c33",
         11439 => x"51cf923f",
         11440 => x"84b8e408",
         11441 => x"762e0981",
         11442 => x"06bc3884",
         11443 => x"b8e40883",
         11444 => x"1d34b41c",
         11445 => x"08a81d08",
         11446 => x"315574a0",
         11447 => x"1d08278a",
         11448 => x"38821c33",
         11449 => x"5f7e822e",
         11450 => x"aa3884b8",
         11451 => x"e40856fc",
         11452 => x"f83975ff",
         11453 => x"1c41587f",
         11454 => x"802efa98",
         11455 => x"38fc8739",
         11456 => x"751a57f7",
         11457 => x"e8398170",
         11458 => x"59567580",
         11459 => x"2efcfe38",
         11460 => x"fafd3981",
         11461 => x"54b41c08",
         11462 => x"a01d0805",
         11463 => x"53615281",
         11464 => x"1c3351ce",
         11465 => x"ac3ffcc1",
         11466 => x"398154b4",
         11467 => x"1808a019",
         11468 => x"0805537c",
         11469 => x"52811833",
         11470 => x"51ce963f",
         11471 => x"f8e339f3",
         11472 => x"3d0d7f61",
         11473 => x"7108405e",
         11474 => x"5c800b96",
         11475 => x"1e34981c",
         11476 => x"08802e82",
         11477 => x"b538ac1c",
         11478 => x"08ff2e80",
         11479 => x"d9388070",
         11480 => x"71608c05",
         11481 => x"08702257",
         11482 => x"585b5c58",
         11483 => x"72782ebc",
         11484 => x"38775474",
         11485 => x"14702281",
         11486 => x"1b5b5556",
         11487 => x"7a829538",
         11488 => x"80d08014",
         11489 => x"7083ffff",
         11490 => x"06585a76",
         11491 => x"8fff2682",
         11492 => x"83387379",
         11493 => x"1a761170",
         11494 => x"225d5855",
         11495 => x"5b79d438",
         11496 => x"7a307080",
         11497 => x"2570307a",
         11498 => x"065a5c5e",
         11499 => x"7c189405",
         11500 => x"57800b82",
         11501 => x"18348070",
         11502 => x"891f5957",
         11503 => x"589c1c08",
         11504 => x"16703381",
         11505 => x"18585653",
         11506 => x"74a02eb2",
         11507 => x"3874852e",
         11508 => x"81bc3875",
         11509 => x"89327030",
         11510 => x"70720780",
         11511 => x"25555b54",
         11512 => x"778b2690",
         11513 => x"3872802e",
         11514 => x"8b38ae77",
         11515 => x"70810559",
         11516 => x"34811858",
         11517 => x"74777081",
         11518 => x"05593481",
         11519 => x"18588a76",
         11520 => x"27ffba38",
         11521 => x"7c188805",
         11522 => x"55800b81",
         11523 => x"1634961d",
         11524 => x"335372a5",
         11525 => x"387781f3",
         11526 => x"38bf0b96",
         11527 => x"1e348157",
         11528 => x"7c179405",
         11529 => x"56800b82",
         11530 => x"17349c1c",
         11531 => x"088c1133",
         11532 => x"55537389",
         11533 => x"3873891e",
         11534 => x"349c1c08",
         11535 => x"538b1333",
         11536 => x"881e349c",
         11537 => x"1c089c11",
         11538 => x"83113382",
         11539 => x"12337190",
         11540 => x"2b71882b",
         11541 => x"07811433",
         11542 => x"70720788",
         11543 => x"2b753371",
         11544 => x"07640c59",
         11545 => x"97163396",
         11546 => x"17337188",
         11547 => x"2b075f41",
         11548 => x"5b405a56",
         11549 => x"5b557786",
         11550 => x"1e239915",
         11551 => x"33981633",
         11552 => x"71882b07",
         11553 => x"5d547b84",
         11554 => x"1e238f3d",
         11555 => x"0d0481e5",
         11556 => x"55fec039",
         11557 => x"771d9611",
         11558 => x"81ff7a31",
         11559 => x"585b5783",
         11560 => x"b5527a90",
         11561 => x"2b740751",
         11562 => x"8191893f",
         11563 => x"84b8e408",
         11564 => x"83ffff06",
         11565 => x"5581ff75",
         11566 => x"27ad3881",
         11567 => x"762781b3",
         11568 => x"3874882a",
         11569 => x"54737a34",
         11570 => x"74971834",
         11571 => x"82780558",
         11572 => x"800b8c1f",
         11573 => x"08565b78",
         11574 => x"19751170",
         11575 => x"225c5754",
         11576 => x"79fd9038",
         11577 => x"fdba3974",
         11578 => x"30763070",
         11579 => x"78078025",
         11580 => x"72802507",
         11581 => x"58555775",
         11582 => x"80f93874",
         11583 => x"7a348178",
         11584 => x"0558800b",
         11585 => x"8c1f0856",
         11586 => x"5bcd3972",
         11587 => x"73891f33",
         11588 => x"5a575777",
         11589 => x"802efe88",
         11590 => x"387c961e",
         11591 => x"7e575954",
         11592 => x"891433ff",
         11593 => x"bf115a54",
         11594 => x"789926a4",
         11595 => x"389c1c08",
         11596 => x"8c113354",
         11597 => x"5b887627",
         11598 => x"b4387284",
         11599 => x"2a537281",
         11600 => x"065e7d80",
         11601 => x"2e8a38a0",
         11602 => x"147083ff",
         11603 => x"ff065553",
         11604 => x"73787081",
         11605 => x"055a3481",
         11606 => x"16811681",
         11607 => x"19718913",
         11608 => x"335e5759",
         11609 => x"565679ff",
         11610 => x"b738fdb4",
         11611 => x"3972832a",
         11612 => x"53cc3980",
         11613 => x"7b307080",
         11614 => x"25703073",
         11615 => x"06535d5f",
         11616 => x"58fca939",
         11617 => x"ef3d0d63",
         11618 => x"70087042",
         11619 => x"575c8065",
         11620 => x"70335755",
         11621 => x"5374af2e",
         11622 => x"83388153",
         11623 => x"7480dc2e",
         11624 => x"81df3872",
         11625 => x"802e81d9",
         11626 => x"38981608",
         11627 => x"881d0c73",
         11628 => x"33963d94",
         11629 => x"3d414255",
         11630 => x"9f752782",
         11631 => x"a7387342",
         11632 => x"8c160858",
         11633 => x"80576170",
         11634 => x"70810552",
         11635 => x"33555373",
         11636 => x"81df3872",
         11637 => x"7f0c73ff",
         11638 => x"2e81ec38",
         11639 => x"83ffff74",
         11640 => x"278b3876",
         11641 => x"10185680",
         11642 => x"76238117",
         11643 => x"577383ff",
         11644 => x"ff0670af",
         11645 => x"3270309f",
         11646 => x"73277180",
         11647 => x"2507575b",
         11648 => x"5b557382",
         11649 => x"90387480",
         11650 => x"dc2e8289",
         11651 => x"387480ff",
         11652 => x"26b23883",
         11653 => x"e4800b83",
         11654 => x"e4803370",
         11655 => x"81ff0656",
         11656 => x"54567380",
         11657 => x"2e81ab38",
         11658 => x"73752e8f",
         11659 => x"38811670",
         11660 => x"337081ff",
         11661 => x"06565456",
         11662 => x"73ee3872",
         11663 => x"81ff065b",
         11664 => x"7a818438",
         11665 => x"7681fe26",
         11666 => x"80fd3876",
         11667 => x"10185d74",
         11668 => x"7d238117",
         11669 => x"62707081",
         11670 => x"05523356",
         11671 => x"54577380",
         11672 => x"2efef038",
         11673 => x"80cb3981",
         11674 => x"7380dc32",
         11675 => x"70307080",
         11676 => x"25730751",
         11677 => x"55585572",
         11678 => x"802ea138",
         11679 => x"81147046",
         11680 => x"54807433",
         11681 => x"545572af",
         11682 => x"2edd3872",
         11683 => x"80dc3270",
         11684 => x"30708025",
         11685 => x"77075154",
         11686 => x"5772e138",
         11687 => x"72881d0c",
         11688 => x"7333963d",
         11689 => x"943d4142",
         11690 => x"55749f26",
         11691 => x"fe9038b4",
         11692 => x"3983b552",
         11693 => x"7351818d",
         11694 => x"e73f84b8",
         11695 => x"e40883ff",
         11696 => x"ff065473",
         11697 => x"fe8d3886",
         11698 => x"547384b8",
         11699 => x"e40c933d",
         11700 => x"0d0483e4",
         11701 => x"80337081",
         11702 => x"ff065c53",
         11703 => x"7a802efe",
         11704 => x"e338e439",
         11705 => x"ff800bab",
         11706 => x"1d348052",
         11707 => x"7b51de8d",
         11708 => x"3f84b8e4",
         11709 => x"0884b8e4",
         11710 => x"0c933d0d",
         11711 => x"04817380",
         11712 => x"dc327030",
         11713 => x"70802573",
         11714 => x"0741555a",
         11715 => x"567d802e",
         11716 => x"a1388114",
         11717 => x"42806270",
         11718 => x"33555556",
         11719 => x"72af2edd",
         11720 => x"387280dc",
         11721 => x"32703070",
         11722 => x"80257807",
         11723 => x"4054597d",
         11724 => x"e1387361",
         11725 => x"0c9f7527",
         11726 => x"822b5a76",
         11727 => x"812e84f8",
         11728 => x"3876822e",
         11729 => x"83d13876",
         11730 => x"17597680",
         11731 => x"2ea73876",
         11732 => x"177811fe",
         11733 => x"05702270",
         11734 => x"a0327030",
         11735 => x"709f2a52",
         11736 => x"42565f56",
         11737 => x"597cae2e",
         11738 => x"84387289",
         11739 => x"38ff1757",
         11740 => x"76dd3876",
         11741 => x"59771956",
         11742 => x"80762376",
         11743 => x"802efec7",
         11744 => x"38807822",
         11745 => x"7083ffff",
         11746 => x"0672585d",
         11747 => x"55567aa0",
         11748 => x"2e82e638",
         11749 => x"7383ffff",
         11750 => x"065372ae",
         11751 => x"2e82f138",
         11752 => x"76802eaa",
         11753 => x"387719fe",
         11754 => x"0570225a",
         11755 => x"5478ae2e",
         11756 => x"9d387610",
         11757 => x"18fe0554",
         11758 => x"ff175776",
         11759 => x"802e8f38",
         11760 => x"fe147022",
         11761 => x"5e547cae",
         11762 => x"2e098106",
         11763 => x"eb388b0b",
         11764 => x"a01d5553",
         11765 => x"a0747081",
         11766 => x"055634ff",
         11767 => x"135372f4",
         11768 => x"3872735c",
         11769 => x"5e887816",
         11770 => x"70228119",
         11771 => x"5957545d",
         11772 => x"74802e80",
         11773 => x"ed3874a0",
         11774 => x"2e83d038",
         11775 => x"74ae3270",
         11776 => x"30708025",
         11777 => x"555a5475",
         11778 => x"772e85ce",
         11779 => x"387283bb",
         11780 => x"3872597c",
         11781 => x"7b268338",
         11782 => x"81597577",
         11783 => x"32703070",
         11784 => x"72078025",
         11785 => x"707c0751",
         11786 => x"51545472",
         11787 => x"802e83e0",
         11788 => x"387c8b2e",
         11789 => x"86833875",
         11790 => x"772e8a38",
         11791 => x"7983075a",
         11792 => x"7577269e",
         11793 => x"38765688",
         11794 => x"5b8b7e82",
         11795 => x"2b81fc06",
         11796 => x"7718575f",
         11797 => x"5d771570",
         11798 => x"22811858",
         11799 => x"565374ff",
         11800 => x"9538a01c",
         11801 => x"33577681",
         11802 => x"e52e8384",
         11803 => x"387c882e",
         11804 => x"82e3387d",
         11805 => x"8c065877",
         11806 => x"8c2e82ed",
         11807 => x"387d8306",
         11808 => x"5574832e",
         11809 => x"82e33879",
         11810 => x"812a8106",
         11811 => x"56759d38",
         11812 => x"7d81065d",
         11813 => x"7c802e85",
         11814 => x"38799007",
         11815 => x"5a7d822a",
         11816 => x"81065e7d",
         11817 => x"802e8538",
         11818 => x"7988075a",
         11819 => x"79ab1d34",
         11820 => x"7b51e4ec",
         11821 => x"3f84b8e4",
         11822 => x"08ab1d33",
         11823 => x"565484b8",
         11824 => x"e408802e",
         11825 => x"81ac3884",
         11826 => x"b8e40884",
         11827 => x"2e098106",
         11828 => x"fbf73874",
         11829 => x"852a8106",
         11830 => x"5a79802e",
         11831 => x"84f03874",
         11832 => x"822a8106",
         11833 => x"59788298",
         11834 => x"387b0865",
         11835 => x"55567342",
         11836 => x"8c160858",
         11837 => x"8057f9ce",
         11838 => x"39811670",
         11839 => x"11791170",
         11840 => x"22404056",
         11841 => x"567ca02e",
         11842 => x"f0387580",
         11843 => x"2efd8538",
         11844 => x"7983075a",
         11845 => x"fd8a3982",
         11846 => x"18225675",
         11847 => x"ae2e0981",
         11848 => x"06fcac38",
         11849 => x"77225473",
         11850 => x"ae2e0981",
         11851 => x"06fca038",
         11852 => x"7610185b",
         11853 => x"807b2380",
         11854 => x"0ba01d56",
         11855 => x"53ae5476",
         11856 => x"73268338",
         11857 => x"a0547375",
         11858 => x"70810557",
         11859 => x"34811353",
         11860 => x"8a7327e9",
         11861 => x"3879a007",
         11862 => x"5877ab1d",
         11863 => x"347b51e3",
         11864 => x"bf3f84b8",
         11865 => x"e408ab1d",
         11866 => x"33565484",
         11867 => x"b8e408fe",
         11868 => x"d6387482",
         11869 => x"2a810658",
         11870 => x"77face38",
         11871 => x"861c3370",
         11872 => x"842a8106",
         11873 => x"565d7480",
         11874 => x"2e83cd38",
         11875 => x"901c0883",
         11876 => x"ff066005",
         11877 => x"80d31133",
         11878 => x"80d21233",
         11879 => x"71882b07",
         11880 => x"62334157",
         11881 => x"54547d83",
         11882 => x"2e82d838",
         11883 => x"74881d0c",
         11884 => x"7b086555",
         11885 => x"56feb739",
         11886 => x"77225574",
         11887 => x"ae2efef0",
         11888 => x"38761759",
         11889 => x"76fb8838",
         11890 => x"fbab3979",
         11891 => x"83077617",
         11892 => x"565afd81",
         11893 => x"397d822b",
         11894 => x"81fc0670",
         11895 => x"8c06595e",
         11896 => x"778c2e09",
         11897 => x"8106fd95",
         11898 => x"38798207",
         11899 => x"5afd9839",
         11900 => x"850ba01d",
         11901 => x"347c882e",
         11902 => x"098106fc",
         11903 => x"f638d639",
         11904 => x"ff800bab",
         11905 => x"1d34800b",
         11906 => x"84b8e40c",
         11907 => x"933d0d04",
         11908 => x"7480ff26",
         11909 => x"9d3881ff",
         11910 => x"752780c9",
         11911 => x"38ff1d59",
         11912 => x"787b2681",
         11913 => x"f7387983",
         11914 => x"077d7718",
         11915 => x"575c5afc",
         11916 => x"a4397982",
         11917 => x"075a83b5",
         11918 => x"52745181",
         11919 => x"85f63f84",
         11920 => x"b8e40883",
         11921 => x"ffff0670",
         11922 => x"872a8106",
         11923 => x"5a557880",
         11924 => x"2ec43874",
         11925 => x"80ff0683",
         11926 => x"e4f41133",
         11927 => x"56547481",
         11928 => x"ff26ffb9",
         11929 => x"3874802e",
         11930 => x"81853883",
         11931 => x"e48c0b83",
         11932 => x"e48c3370",
         11933 => x"81ff0656",
         11934 => x"54597380",
         11935 => x"2e80e038",
         11936 => x"73752e8f",
         11937 => x"38811970",
         11938 => x"337081ff",
         11939 => x"06565459",
         11940 => x"73ee3872",
         11941 => x"81ff0659",
         11942 => x"7880d438",
         11943 => x"ffbf1554",
         11944 => x"7399268a",
         11945 => x"387d8207",
         11946 => x"7081ff06",
         11947 => x"5f53ff9f",
         11948 => x"15597899",
         11949 => x"2693387d",
         11950 => x"81077081",
         11951 => x"ff06e017",
         11952 => x"7083ffff",
         11953 => x"0658565f",
         11954 => x"537b1ba0",
         11955 => x"05597479",
         11956 => x"34811b5b",
         11957 => x"751655fa",
         11958 => x"fc398053",
         11959 => x"fab33983",
         11960 => x"e48c3370",
         11961 => x"81ff065a",
         11962 => x"5378802e",
         11963 => x"ffae3880",
         11964 => x"df7a8307",
         11965 => x"7d1da005",
         11966 => x"5b5b5574",
         11967 => x"7934811b",
         11968 => x"5bd23980",
         11969 => x"cd143380",
         11970 => x"cc153371",
         11971 => x"982b7190",
         11972 => x"2b077707",
         11973 => x"881f0c5a",
         11974 => x"57fd9539",
         11975 => x"7b1ba005",
         11976 => x"75882a54",
         11977 => x"54727434",
         11978 => x"811b7c11",
         11979 => x"a0055a5b",
         11980 => x"74793481",
         11981 => x"1b5bff9c",
         11982 => x"39798307",
         11983 => x"a01d3358",
         11984 => x"5a7681e5",
         11985 => x"2e098106",
         11986 => x"faa338fd",
         11987 => x"a3397482",
         11988 => x"2a81065c",
         11989 => x"7bf6f238",
         11990 => x"850b84b8",
         11991 => x"e40c933d",
         11992 => x"0d04eb3d",
         11993 => x"0d676902",
         11994 => x"880580e7",
         11995 => x"05334242",
         11996 => x"5e80610c",
         11997 => x"ff7e0870",
         11998 => x"595b4279",
         11999 => x"802e85d7",
         12000 => x"38797081",
         12001 => x"055b3370",
         12002 => x"9f265656",
         12003 => x"75ba2e85",
         12004 => x"d03874ed",
         12005 => x"3875ba2e",
         12006 => x"85c73884",
         12007 => x"d0c03356",
         12008 => x"80762485",
         12009 => x"b2387510",
         12010 => x"1084d0ac",
         12011 => x"05700858",
         12012 => x"5a8c5876",
         12013 => x"802e8596",
         12014 => x"3876610c",
         12015 => x"7f81fe06",
         12016 => x"77335d59",
         12017 => x"7b802e9b",
         12018 => x"38811733",
         12019 => x"51ffbbb0",
         12020 => x"3f84b8e4",
         12021 => x"0881ff06",
         12022 => x"7081065e",
         12023 => x"587c802e",
         12024 => x"86963880",
         12025 => x"77347516",
         12026 => x"5d84b8d8",
         12027 => x"1d338118",
         12028 => x"34815281",
         12029 => x"173351ff",
         12030 => x"bba43f84",
         12031 => x"b8e40881",
         12032 => x"ff067081",
         12033 => x"06415683",
         12034 => x"587f84c2",
         12035 => x"3878802e",
         12036 => x"8d387582",
         12037 => x"2a810641",
         12038 => x"8a586084",
         12039 => x"b138805b",
         12040 => x"7a831834",
         12041 => x"ff0bb418",
         12042 => x"0c7a7b5a",
         12043 => x"5581547a",
         12044 => x"53b81770",
         12045 => x"53811833",
         12046 => x"5258ffbb",
         12047 => x"953f84b8",
         12048 => x"e4087b2e",
         12049 => x"8538ff55",
         12050 => x"815974b4",
         12051 => x"180c8456",
         12052 => x"78993884",
         12053 => x"b7173384",
         12054 => x"b6183371",
         12055 => x"882b0756",
         12056 => x"56835674",
         12057 => x"82d4d52e",
         12058 => x"85a53875",
         12059 => x"81268b38",
         12060 => x"84b8d91d",
         12061 => x"33426185",
         12062 => x"bf388158",
         12063 => x"75842e83",
         12064 => x"cd388d58",
         12065 => x"75812683",
         12066 => x"c53880c4",
         12067 => x"173380c3",
         12068 => x"18337188",
         12069 => x"2b075e59",
         12070 => x"7c84802e",
         12071 => x"09810683",
         12072 => x"ad3880cf",
         12073 => x"173380ce",
         12074 => x"18337188",
         12075 => x"2b07575a",
         12076 => x"75a43880",
         12077 => x"dc178311",
         12078 => x"33821233",
         12079 => x"71902b71",
         12080 => x"882b0781",
         12081 => x"14337072",
         12082 => x"07882b75",
         12083 => x"33710756",
         12084 => x"5a45435e",
         12085 => x"5f5675a0",
         12086 => x"180c80c8",
         12087 => x"17338218",
         12088 => x"3480c817",
         12089 => x"33ff1170",
         12090 => x"81ff065f",
         12091 => x"40598d58",
         12092 => x"7c812682",
         12093 => x"d9387881",
         12094 => x"ff067671",
         12095 => x"2980c519",
         12096 => x"335a5f5a",
         12097 => x"778a1823",
         12098 => x"77597780",
         12099 => x"2e87c438",
         12100 => x"ff187806",
         12101 => x"426187bb",
         12102 => x"3880ca17",
         12103 => x"3380c918",
         12104 => x"3371882b",
         12105 => x"07564074",
         12106 => x"88182374",
         12107 => x"758f065e",
         12108 => x"5a8d587c",
         12109 => x"82983880",
         12110 => x"cc173380",
         12111 => x"cb183371",
         12112 => x"882b0756",
         12113 => x"5c74a438",
         12114 => x"80d81783",
         12115 => x"11338212",
         12116 => x"3371902b",
         12117 => x"71882b07",
         12118 => x"81143370",
         12119 => x"7207882b",
         12120 => x"75337107",
         12121 => x"53445a58",
         12122 => x"42424280",
         12123 => x"c7173380",
         12124 => x"c6183371",
         12125 => x"882b075d",
         12126 => x"588d587b",
         12127 => x"802e81ce",
         12128 => x"387d1c7a",
         12129 => x"842a055a",
         12130 => x"79752681",
         12131 => x"c1387852",
         12132 => x"747a3151",
         12133 => x"fdee8e3f",
         12134 => x"84b8e408",
         12135 => x"5684b8e4",
         12136 => x"08802e81",
         12137 => x"a93884b8",
         12138 => x"e40880ff",
         12139 => x"fffff526",
         12140 => x"8338835d",
         12141 => x"7583fff5",
         12142 => x"26833882",
         12143 => x"5d759ff5",
         12144 => x"2685eb38",
         12145 => x"815d8216",
         12146 => x"709c190c",
         12147 => x"7ba4190c",
         12148 => x"7b1d70a8",
         12149 => x"1a0c7b1d",
         12150 => x"b01a0c57",
         12151 => x"597c832e",
         12152 => x"8a873888",
         12153 => x"17225c8d",
         12154 => x"587b802e",
         12155 => x"80e0387d",
         12156 => x"16ac180c",
         12157 => x"7819557c",
         12158 => x"822e8d38",
         12159 => x"78101970",
         12160 => x"812a7a81",
         12161 => x"0605565a",
         12162 => x"83ff1589",
         12163 => x"2a598d58",
         12164 => x"78a01808",
         12165 => x"26b838ff",
         12166 => x"0b94180c",
         12167 => x"ff0b9018",
         12168 => x"0cff800b",
         12169 => x"8418347c",
         12170 => x"832e8696",
         12171 => x"387c7734",
         12172 => x"84d0bc22",
         12173 => x"81055d7c",
         12174 => x"84d0bc23",
         12175 => x"7c861823",
         12176 => x"84d0c40b",
         12177 => x"8c180c80",
         12178 => x"0b98180c",
         12179 => x"80587784",
         12180 => x"b8e40c97",
         12181 => x"3d0d048b",
         12182 => x"0b84b8e4",
         12183 => x"0c973d0d",
         12184 => x"047633d0",
         12185 => x"117081ff",
         12186 => x"06575758",
         12187 => x"74892691",
         12188 => x"38821778",
         12189 => x"81ff06d0",
         12190 => x"055d5978",
         12191 => x"7a2e87fe",
         12192 => x"38807e08",
         12193 => x"83e4d45f",
         12194 => x"405c7c08",
         12195 => x"7f5a5b7a",
         12196 => x"7081055c",
         12197 => x"33797081",
         12198 => x"055b33ff",
         12199 => x"9f125a58",
         12200 => x"56779926",
         12201 => x"8938e016",
         12202 => x"7081ff06",
         12203 => x"5755ff9f",
         12204 => x"17587799",
         12205 => x"268938e0",
         12206 => x"177081ff",
         12207 => x"06585575",
         12208 => x"30709f2a",
         12209 => x"59557577",
         12210 => x"2e098106",
         12211 => x"853877ff",
         12212 => x"be38787a",
         12213 => x"32703070",
         12214 => x"72079f2a",
         12215 => x"7a075d58",
         12216 => x"557a802e",
         12217 => x"87983881",
         12218 => x"1c841e5e",
         12219 => x"5c837c25",
         12220 => x"ff983861",
         12221 => x"56f9a939",
         12222 => x"78802efe",
         12223 => x"cf387782",
         12224 => x"2a81065e",
         12225 => x"8a587dfe",
         12226 => x"c5388058",
         12227 => x"fec0397a",
         12228 => x"78335759",
         12229 => x"7581e92e",
         12230 => x"09810683",
         12231 => x"38815975",
         12232 => x"81eb3270",
         12233 => x"30708025",
         12234 => x"7b075a5b",
         12235 => x"5c7783ad",
         12236 => x"387581e8",
         12237 => x"2e83a638",
         12238 => x"933d7757",
         12239 => x"5a835983",
         12240 => x"fa163370",
         12241 => x"595b7a80",
         12242 => x"2ea53884",
         12243 => x"81163384",
         12244 => x"80173371",
         12245 => x"902b7188",
         12246 => x"2b0783ff",
         12247 => x"19337072",
         12248 => x"07882b83",
         12249 => x"fe1b3371",
         12250 => x"0752595b",
         12251 => x"40404077",
         12252 => x"7a708405",
         12253 => x"5c0cff19",
         12254 => x"90175759",
         12255 => x"788025ff",
         12256 => x"be3884b8",
         12257 => x"d91d3370",
         12258 => x"30709f2a",
         12259 => x"7271319b",
         12260 => x"3d711010",
         12261 => x"05f00584",
         12262 => x"b61c445d",
         12263 => x"52435b42",
         12264 => x"78085b83",
         12265 => x"567a802e",
         12266 => x"80fb3880",
         12267 => x"0b831834",
         12268 => x"ff0bb418",
         12269 => x"0c7a5580",
         12270 => x"567aff2e",
         12271 => x"a5388154",
         12272 => x"7a53b817",
         12273 => x"52811733",
         12274 => x"51ffb486",
         12275 => x"3f84b8e4",
         12276 => x"08762e85",
         12277 => x"38ff5581",
         12278 => x"5674b418",
         12279 => x"0c845875",
         12280 => x"bf38811f",
         12281 => x"337f3371",
         12282 => x"882b075d",
         12283 => x"5e83587b",
         12284 => x"82d4d52e",
         12285 => x"098106a8",
         12286 => x"38800bb8",
         12287 => x"18335758",
         12288 => x"7581e92e",
         12289 => x"82b73875",
         12290 => x"81eb3270",
         12291 => x"30708025",
         12292 => x"7a074242",
         12293 => x"427fbc38",
         12294 => x"7581e82e",
         12295 => x"b6388258",
         12296 => x"7781ff06",
         12297 => x"56800b84",
         12298 => x"b8d91e33",
         12299 => x"5d587b78",
         12300 => x"2e098106",
         12301 => x"83388158",
         12302 => x"817627f8",
         12303 => x"bd387780",
         12304 => x"2ef8b738",
         12305 => x"811a841a",
         12306 => x"5a5a837a",
         12307 => x"27fed138",
         12308 => x"f8a83983",
         12309 => x"0b80ee18",
         12310 => x"83e49440",
         12311 => x"5d587b70",
         12312 => x"81055d33",
         12313 => x"7e708105",
         12314 => x"40337171",
         12315 => x"31ff1b5b",
         12316 => x"52565677",
         12317 => x"802e80c5",
         12318 => x"3875802e",
         12319 => x"e138850b",
         12320 => x"818a1883",
         12321 => x"e498405d",
         12322 => x"587b7081",
         12323 => x"055d337e",
         12324 => x"70810540",
         12325 => x"33717131",
         12326 => x"ff1b5b58",
         12327 => x"42407780",
         12328 => x"2e858e38",
         12329 => x"75802ee1",
         12330 => x"388258fe",
         12331 => x"f3398d58",
         12332 => x"7cfa9338",
         12333 => x"7784b8e4",
         12334 => x"0c973d0d",
         12335 => x"04755875",
         12336 => x"802efedc",
         12337 => x"38850b81",
         12338 => x"8a1883e4",
         12339 => x"98405d58",
         12340 => x"ffb7398d",
         12341 => x"0b84b8e4",
         12342 => x"0c973d0d",
         12343 => x"04830b80",
         12344 => x"ee1883e4",
         12345 => x"945c5a58",
         12346 => x"78708105",
         12347 => x"5a337a70",
         12348 => x"81055c33",
         12349 => x"717131ff",
         12350 => x"1b5b575f",
         12351 => x"5f77802e",
         12352 => x"83d13874",
         12353 => x"802ee138",
         12354 => x"850b818a",
         12355 => x"1883e498",
         12356 => x"5c5a5878",
         12357 => x"7081055a",
         12358 => x"337a7081",
         12359 => x"055c3371",
         12360 => x"7131ff1b",
         12361 => x"5b584240",
         12362 => x"77802e84",
         12363 => x"91387580",
         12364 => x"2ee13893",
         12365 => x"3d77575a",
         12366 => x"8359fc83",
         12367 => x"398158fd",
         12368 => x"c63980e9",
         12369 => x"173380e8",
         12370 => x"18337188",
         12371 => x"2b075755",
         12372 => x"75812e09",
         12373 => x"8106f9d5",
         12374 => x"38811b58",
         12375 => x"805ab417",
         12376 => x"08782eb1",
         12377 => x"38831733",
         12378 => x"5b7a7a2e",
         12379 => x"09810682",
         12380 => x"9b388154",
         12381 => x"7753b817",
         12382 => x"52811733",
         12383 => x"51ffb0d2",
         12384 => x"3f84b8e4",
         12385 => x"08802e85",
         12386 => x"38ff5881",
         12387 => x"5a77b418",
         12388 => x"0c79f999",
         12389 => x"38798418",
         12390 => x"3484b717",
         12391 => x"3384b618",
         12392 => x"3371882b",
         12393 => x"07575e75",
         12394 => x"82d4d52e",
         12395 => x"098106f8",
         12396 => x"fc38b817",
         12397 => x"83113382",
         12398 => x"12337190",
         12399 => x"2b71882b",
         12400 => x"07811433",
         12401 => x"70720788",
         12402 => x"2b753371",
         12403 => x"075e4159",
         12404 => x"45425c59",
         12405 => x"77848b85",
         12406 => x"a4d22e09",
         12407 => x"8106f8cd",
         12408 => x"38849c17",
         12409 => x"83113382",
         12410 => x"12337190",
         12411 => x"2b71882b",
         12412 => x"07811433",
         12413 => x"70720788",
         12414 => x"2b753371",
         12415 => x"07474440",
         12416 => x"5b5c5a5e",
         12417 => x"60868a85",
         12418 => x"e4f22e09",
         12419 => x"8106f89d",
         12420 => x"3884a017",
         12421 => x"83113382",
         12422 => x"12337190",
         12423 => x"2b71882b",
         12424 => x"07811433",
         12425 => x"70720788",
         12426 => x"2b753371",
         12427 => x"07941e0c",
         12428 => x"5d84a41c",
         12429 => x"83113382",
         12430 => x"12337190",
         12431 => x"2b71882b",
         12432 => x"07811433",
         12433 => x"70720788",
         12434 => x"2b753371",
         12435 => x"07629005",
         12436 => x"0c594449",
         12437 => x"465c4540",
         12438 => x"455b565a",
         12439 => x"7c773484",
         12440 => x"d0bc2281",
         12441 => x"055d7c84",
         12442 => x"d0bc237c",
         12443 => x"86182384",
         12444 => x"d0c40b8c",
         12445 => x"180c800b",
         12446 => x"98180cf7",
         12447 => x"cf397b83",
         12448 => x"24f8f038",
         12449 => x"7b7a7f0c",
         12450 => x"56f29539",
         12451 => x"7554b417",
         12452 => x"0853b817",
         12453 => x"70538118",
         12454 => x"335259ff",
         12455 => x"afb33f84",
         12456 => x"b8e4087a",
         12457 => x"2e098106",
         12458 => x"81a43884",
         12459 => x"b8e40883",
         12460 => x"1834b417",
         12461 => x"08a81808",
         12462 => x"31407fa0",
         12463 => x"1808278b",
         12464 => x"38821733",
         12465 => x"4160822e",
         12466 => x"818d3884",
         12467 => x"b8e4085a",
         12468 => x"fda03974",
         12469 => x"5674802e",
         12470 => x"f3913885",
         12471 => x"0b818a18",
         12472 => x"83e4985c",
         12473 => x"5a58fcab",
         12474 => x"3980e317",
         12475 => x"3380e218",
         12476 => x"3371882b",
         12477 => x"075f5a8d",
         12478 => x"587df6d2",
         12479 => x"38881722",
         12480 => x"4261f6ca",
         12481 => x"3880e417",
         12482 => x"83113382",
         12483 => x"12337190",
         12484 => x"2b71882b",
         12485 => x"07811433",
         12486 => x"70720788",
         12487 => x"2b753371",
         12488 => x"07ac1e0c",
         12489 => x"5a7d822b",
         12490 => x"5a434440",
         12491 => x"5940f5d8",
         12492 => x"39755875",
         12493 => x"802ef9e8",
         12494 => x"388258f9",
         12495 => x"e3397580",
         12496 => x"2ef2a838",
         12497 => x"933d7757",
         12498 => x"5a8359f7",
         12499 => x"f239755a",
         12500 => x"79f5da38",
         12501 => x"fcbf3975",
         12502 => x"54b41708",
         12503 => x"a0180805",
         12504 => x"53785281",
         12505 => x"173351ff",
         12506 => x"ade73ffc",
         12507 => x"8539f03d",
         12508 => x"0d0280d3",
         12509 => x"05336470",
         12510 => x"43933d41",
         12511 => x"575dff76",
         12512 => x"5a407580",
         12513 => x"2e80e938",
         12514 => x"78708105",
         12515 => x"5a33709f",
         12516 => x"26555574",
         12517 => x"ba2e80e2",
         12518 => x"3873ed38",
         12519 => x"74ba2e80",
         12520 => x"d93884d0",
         12521 => x"c0335480",
         12522 => x"742480c4",
         12523 => x"38731010",
         12524 => x"84d0ac05",
         12525 => x"70085555",
         12526 => x"73802e84",
         12527 => x"38807434",
         12528 => x"62547380",
         12529 => x"2e863880",
         12530 => x"74346254",
         12531 => x"73750c7c",
         12532 => x"547c802e",
         12533 => x"92388053",
         12534 => x"933d7053",
         12535 => x"840551ef",
         12536 => x"813f84b8",
         12537 => x"e4085473",
         12538 => x"84b8e40c",
         12539 => x"923d0d04",
         12540 => x"8b0b84b8",
         12541 => x"e40c923d",
         12542 => x"0d047533",
         12543 => x"d0117081",
         12544 => x"ff065656",
         12545 => x"57738926",
         12546 => x"91388216",
         12547 => x"7781ff06",
         12548 => x"d0055c58",
         12549 => x"77792e80",
         12550 => x"f738807f",
         12551 => x"0883e4d4",
         12552 => x"5e5f5b7b",
         12553 => x"087e595a",
         12554 => x"79708105",
         12555 => x"5b337870",
         12556 => x"81055a33",
         12557 => x"ff9f1259",
         12558 => x"57557699",
         12559 => x"268938e0",
         12560 => x"157081ff",
         12561 => x"065654ff",
         12562 => x"9f165776",
         12563 => x"99268938",
         12564 => x"e0167081",
         12565 => x"ff065754",
         12566 => x"7430709f",
         12567 => x"2a585474",
         12568 => x"762e0981",
         12569 => x"06853876",
         12570 => x"ffbe3877",
         12571 => x"79327030",
         12572 => x"7072079f",
         12573 => x"2a79075c",
         12574 => x"57547980",
         12575 => x"2e923881",
         12576 => x"1b841d5d",
         12577 => x"5b837b25",
         12578 => x"ff99387f",
         12579 => x"54fe9839",
         12580 => x"7a8324f7",
         12581 => x"387a7960",
         12582 => x"0c54fe8b",
         12583 => x"39e63d0d",
         12584 => x"6c028405",
         12585 => x"80fb0533",
         12586 => x"56598956",
         12587 => x"78802ea6",
         12588 => x"3874bf06",
         12589 => x"70549d3d",
         12590 => x"cc05539e",
         12591 => x"3d840552",
         12592 => x"58ed9f3f",
         12593 => x"84b8e408",
         12594 => x"5784b8e4",
         12595 => x"08802e8f",
         12596 => x"3880790c",
         12597 => x"76567584",
         12598 => x"b8e40c9c",
         12599 => x"3d0d047e",
         12600 => x"406d5290",
         12601 => x"3d70525a",
         12602 => x"e19a3f84",
         12603 => x"b8e40857",
         12604 => x"84b8e408",
         12605 => x"802e81ba",
         12606 => x"38779c06",
         12607 => x"5d7c802e",
         12608 => x"81ca3876",
         12609 => x"802e83c1",
         12610 => x"3876842e",
         12611 => x"83ea3877",
         12612 => x"88075876",
         12613 => x"ffbb3877",
         12614 => x"832a8106",
         12615 => x"5b7a802e",
         12616 => x"81d13866",
         12617 => x"9b11339a",
         12618 => x"12337188",
         12619 => x"2b076170",
         12620 => x"3342585e",
         12621 => x"5e567d83",
         12622 => x"2e84e938",
         12623 => x"800b8e17",
         12624 => x"34800b8f",
         12625 => x"1734a10b",
         12626 => x"90173480",
         12627 => x"cc0b9117",
         12628 => x"346656a0",
         12629 => x"0b8b1734",
         12630 => x"7e67575e",
         12631 => x"800b9a17",
         12632 => x"34800b9b",
         12633 => x"17347d33",
         12634 => x"5d7c832e",
         12635 => x"84a93866",
         12636 => x"5b800b9c",
         12637 => x"1c34800b",
         12638 => x"9d1c3480",
         12639 => x"0b9e1c34",
         12640 => x"800b9f1c",
         12641 => x"347e5581",
         12642 => x"0b831634",
         12643 => x"7b802e80",
         12644 => x"e2387eb4",
         12645 => x"11087d7c",
         12646 => x"0853575f",
         12647 => x"57817c27",
         12648 => x"89389c17",
         12649 => x"087c2683",
         12650 => x"8a388257",
         12651 => x"80790cfe",
         12652 => x"a3390280",
         12653 => x"e7053370",
         12654 => x"982b5d5b",
         12655 => x"7b8025fe",
         12656 => x"b8388678",
         12657 => x"9c065e57",
         12658 => x"7cfeb838",
         12659 => x"76fe8238",
         12660 => x"0280c205",
         12661 => x"3370842a",
         12662 => x"81065d56",
         12663 => x"7b829138",
         12664 => x"77812a81",
         12665 => x"065e7d80",
         12666 => x"2e893875",
         12667 => x"81065a79",
         12668 => x"81f63877",
         12669 => x"832a8106",
         12670 => x"5675802e",
         12671 => x"86387780",
         12672 => x"c007587e",
         12673 => x"b41108a0",
         12674 => x"1b0c67a4",
         12675 => x"1b0c679b",
         12676 => x"11339a12",
         12677 => x"3371882b",
         12678 => x"07733340",
         12679 => x"5e40575a",
         12680 => x"7b832e81",
         12681 => x"f1387a88",
         12682 => x"1a0c9c16",
         12683 => x"83113382",
         12684 => x"12337190",
         12685 => x"2b71882b",
         12686 => x"07811433",
         12687 => x"70720788",
         12688 => x"2b753371",
         12689 => x"0770608c",
         12690 => x"050c6060",
         12691 => x"0c515241",
         12692 => x"59575d5e",
         12693 => x"861a2284",
         12694 => x"1a237790",
         12695 => x"1a34800b",
         12696 => x"911a3480",
         12697 => x"0b9c1a0c",
         12698 => x"77852a81",
         12699 => x"06557480",
         12700 => x"2e84ac38",
         12701 => x"75802e84",
         12702 => x"f1387594",
         12703 => x"1a0c8a1a",
         12704 => x"2270892b",
         12705 => x"7c525b58",
         12706 => x"76307078",
         12707 => x"07802556",
         12708 => x"5b797627",
         12709 => x"84923881",
         12710 => x"7076065f",
         12711 => x"5b7d802e",
         12712 => x"84863877",
         12713 => x"527851ff",
         12714 => x"acdb3f84",
         12715 => x"b8e40858",
         12716 => x"84b8e408",
         12717 => x"81268338",
         12718 => x"825784b8",
         12719 => x"e408ff2e",
         12720 => x"80cb3875",
         12721 => x"7a3156c0",
         12722 => x"390280c2",
         12723 => x"05339106",
         12724 => x"5e7d9538",
         12725 => x"77822a81",
         12726 => x"06557480",
         12727 => x"2efcb838",
         12728 => x"88578079",
         12729 => x"0cfbed39",
         12730 => x"87578079",
         12731 => x"0cfbe539",
         12732 => x"84578079",
         12733 => x"0cfbdd39",
         12734 => x"7951cdca",
         12735 => x"3f84b8e4",
         12736 => x"08788807",
         12737 => x"595776fb",
         12738 => x"c838fc8b",
         12739 => x"397a767b",
         12740 => x"315757fe",
         12741 => x"f3399516",
         12742 => x"33941733",
         12743 => x"71982b71",
         12744 => x"902b077d",
         12745 => x"075d5e5c",
         12746 => x"fdfc397c",
         12747 => x"557c7b27",
         12748 => x"81bd3874",
         12749 => x"527951ff",
         12750 => x"abcb3f84",
         12751 => x"b8e4085d",
         12752 => x"84b8e408",
         12753 => x"802e81a7",
         12754 => x"3884b8e4",
         12755 => x"08812efc",
         12756 => x"d93884b8",
         12757 => x"e408ff2e",
         12758 => x"83993880",
         12759 => x"53745276",
         12760 => x"51ffb282",
         12761 => x"3f84b8e4",
         12762 => x"08839038",
         12763 => x"9c1708fe",
         12764 => x"11941908",
         12765 => x"58565b75",
         12766 => x"7527ffaf",
         12767 => x"38811694",
         12768 => x"180c8417",
         12769 => x"33810755",
         12770 => x"74841834",
         12771 => x"7c557a7d",
         12772 => x"26ffa038",
         12773 => x"80d93980",
         12774 => x"0b941734",
         12775 => x"800b9517",
         12776 => x"34fbcc39",
         12777 => x"95163394",
         12778 => x"17337198",
         12779 => x"2b71902b",
         12780 => x"077e075e",
         12781 => x"565b800b",
         12782 => x"8e173480",
         12783 => x"0b8f1734",
         12784 => x"a10b9017",
         12785 => x"3480cc0b",
         12786 => x"91173466",
         12787 => x"56a00b8b",
         12788 => x"17347e67",
         12789 => x"575e800b",
         12790 => x"9a173480",
         12791 => x"0b9b1734",
         12792 => x"7d335d7c",
         12793 => x"832e0981",
         12794 => x"06fb8438",
         12795 => x"ffa93980",
         12796 => x"7f7f725e",
         12797 => x"59575db4",
         12798 => x"16087e2e",
         12799 => x"ae388316",
         12800 => x"335a797d",
         12801 => x"2e098106",
         12802 => x"b5388154",
         12803 => x"7d53b816",
         12804 => x"52811633",
         12805 => x"51ffa3ba",
         12806 => x"3f84b8e4",
         12807 => x"08802e85",
         12808 => x"38ff5781",
         12809 => x"5b76b417",
         12810 => x"0c7e567a",
         12811 => x"ff1d9018",
         12812 => x"0c577a80",
         12813 => x"2efbbc38",
         12814 => x"80790cf9",
         12815 => x"97398154",
         12816 => x"b4160853",
         12817 => x"b8167053",
         12818 => x"81173352",
         12819 => x"5affa481",
         12820 => x"3f84b8e4",
         12821 => x"087d2e09",
         12822 => x"810681aa",
         12823 => x"3884b8e4",
         12824 => x"08831734",
         12825 => x"b41608a8",
         12826 => x"17083184",
         12827 => x"b8e4085c",
         12828 => x"5574a017",
         12829 => x"0827ff92",
         12830 => x"38821633",
         12831 => x"5574822e",
         12832 => x"098106ff",
         12833 => x"85388154",
         12834 => x"b41608a0",
         12835 => x"17080553",
         12836 => x"79528116",
         12837 => x"3351ffa3",
         12838 => x"b83f7c5b",
         12839 => x"feec3974",
         12840 => x"941a0c76",
         12841 => x"56f8af39",
         12842 => x"77981a0c",
         12843 => x"76f8a238",
         12844 => x"7583ff06",
         12845 => x"5a79802e",
         12846 => x"f89a387e",
         12847 => x"fe199c12",
         12848 => x"08fe055f",
         12849 => x"595a777d",
         12850 => x"27f9df38",
         12851 => x"8a1a2278",
         12852 => x"7129b01c",
         12853 => x"0805565c",
         12854 => x"74802ef9",
         12855 => x"cd387589",
         12856 => x"2a159c1a",
         12857 => x"0c7656f7",
         12858 => x"ed397594",
         12859 => x"1a0c7656",
         12860 => x"f7e43981",
         12861 => x"5780790c",
         12862 => x"f7da3984",
         12863 => x"b8e40857",
         12864 => x"80790cf7",
         12865 => x"cf39817f",
         12866 => x"575bfe9f",
         12867 => x"39f03d0d",
         12868 => x"62656766",
         12869 => x"40405d5a",
         12870 => x"807e0c89",
         12871 => x"5779802e",
         12872 => x"9f387908",
         12873 => x"5675802e",
         12874 => x"97387533",
         12875 => x"5574802e",
         12876 => x"8f388616",
         12877 => x"22841b22",
         12878 => x"59597878",
         12879 => x"2e84b738",
         12880 => x"80557441",
         12881 => x"76557682",
         12882 => x"8c38911a",
         12883 => x"33557482",
         12884 => x"8438901a",
         12885 => x"33810657",
         12886 => x"87567680",
         12887 => x"2e81ed38",
         12888 => x"941a088c",
         12889 => x"1b087131",
         12890 => x"56567b75",
         12891 => x"2681ef38",
         12892 => x"7b802e81",
         12893 => x"d5386059",
         12894 => x"7583ff06",
         12895 => x"5b7a81e3",
         12896 => x"388a1922",
         12897 => x"ff057689",
         12898 => x"2a065b7a",
         12899 => x"9b387583",
         12900 => x"d338881a",
         12901 => x"08558175",
         12902 => x"27848538",
         12903 => x"74ff2e83",
         12904 => x"f0387498",
         12905 => x"1b0c6059",
         12906 => x"981a08fe",
         12907 => x"059c1a08",
         12908 => x"fe054157",
         12909 => x"76602783",
         12910 => x"e7388a19",
         12911 => x"22707829",
         12912 => x"b01b0805",
         12913 => x"56567480",
         12914 => x"2e83d538",
         12915 => x"7a157c89",
         12916 => x"2a595777",
         12917 => x"802e8381",
         12918 => x"38771b55",
         12919 => x"75752785",
         12920 => x"38757b31",
         12921 => x"58775476",
         12922 => x"537c5281",
         12923 => x"193351ff",
         12924 => x"9fe03f84",
         12925 => x"b8e40883",
         12926 => x"98386083",
         12927 => x"11335759",
         12928 => x"75802ea9",
         12929 => x"38b41908",
         12930 => x"77315675",
         12931 => x"78279e38",
         12932 => x"84807671",
         12933 => x"291eb81b",
         12934 => x"58585575",
         12935 => x"70810557",
         12936 => x"33777081",
         12937 => x"055934ff",
         12938 => x"155574ef",
         12939 => x"3877892b",
         12940 => x"587b7831",
         12941 => x"7e08197f",
         12942 => x"0c781e94",
         12943 => x"1c081a70",
         12944 => x"59941d0c",
         12945 => x"5e5c7bfe",
         12946 => x"af388056",
         12947 => x"7584b8e4",
         12948 => x"0c923d0d",
         12949 => x"047484b8",
         12950 => x"e40c923d",
         12951 => x"0d04745c",
         12952 => x"fe8e399c",
         12953 => x"1a085775",
         12954 => x"83ff0684",
         12955 => x"80713159",
         12956 => x"5b7b7827",
         12957 => x"83387b58",
         12958 => x"7656b419",
         12959 => x"08772eb6",
         12960 => x"38800b83",
         12961 => x"1a33715d",
         12962 => x"415f7f7f",
         12963 => x"2e098106",
         12964 => x"80e43881",
         12965 => x"547653b8",
         12966 => x"19528119",
         12967 => x"3351ff9e",
         12968 => x"b13f84b8",
         12969 => x"e408802e",
         12970 => x"8538ff56",
         12971 => x"815b75b4",
         12972 => x"1a0c7a81",
         12973 => x"dc386094",
         12974 => x"1b0883ff",
         12975 => x"0611797f",
         12976 => x"5a58b805",
         12977 => x"56597780",
         12978 => x"2efee638",
         12979 => x"74708105",
         12980 => x"56337770",
         12981 => x"81055934",
         12982 => x"ff165675",
         12983 => x"802efed1",
         12984 => x"38747081",
         12985 => x"05563377",
         12986 => x"70810559",
         12987 => x"34ff1656",
         12988 => x"75da38fe",
         12989 => x"bc398154",
         12990 => x"b4190853",
         12991 => x"b8197053",
         12992 => x"811a3352",
         12993 => x"40ff9ec9",
         12994 => x"3f815b84",
         12995 => x"b8e4087f",
         12996 => x"2e098106",
         12997 => x"ff9c3884",
         12998 => x"b8e40883",
         12999 => x"1a34b419",
         13000 => x"08a81a08",
         13001 => x"3184b8e4",
         13002 => x"085c5574",
         13003 => x"a01a0827",
         13004 => x"fee13882",
         13005 => x"19335574",
         13006 => x"822e0981",
         13007 => x"06fed438",
         13008 => x"8154b419",
         13009 => x"08a01a08",
         13010 => x"05537f52",
         13011 => x"81193351",
         13012 => x"ff9dfe3f",
         13013 => x"7e5bfebb",
         13014 => x"39769c1b",
         13015 => x"0c941a08",
         13016 => x"56fe8439",
         13017 => x"981a0852",
         13018 => x"7951ffa3",
         13019 => x"983f84b8",
         13020 => x"e40855fc",
         13021 => x"a1398116",
         13022 => x"3351ff9c",
         13023 => x"833f84b8",
         13024 => x"e4088106",
         13025 => x"5574fbb8",
         13026 => x"38747a08",
         13027 => x"5657fbb2",
         13028 => x"39810b91",
         13029 => x"1b34810b",
         13030 => x"84b8e40c",
         13031 => x"923d0d04",
         13032 => x"820b911b",
         13033 => x"34820b84",
         13034 => x"b8e40c92",
         13035 => x"3d0d04f0",
         13036 => x"3d0d6265",
         13037 => x"67664040",
         13038 => x"5c5a807e",
         13039 => x"0c895779",
         13040 => x"802e9f38",
         13041 => x"79085675",
         13042 => x"802e9738",
         13043 => x"75335574",
         13044 => x"802e8f38",
         13045 => x"86162284",
         13046 => x"1b225959",
         13047 => x"78782e85",
         13048 => x"fd388055",
         13049 => x"74417655",
         13050 => x"7682c438",
         13051 => x"911a3355",
         13052 => x"7482bc38",
         13053 => x"901a3370",
         13054 => x"812a8106",
         13055 => x"58588756",
         13056 => x"76802e82",
         13057 => x"a138941a",
         13058 => x"087b115d",
         13059 => x"577b7727",
         13060 => x"84387609",
         13061 => x"5b7a802e",
         13062 => x"82813876",
         13063 => x"83ff065f",
         13064 => x"7e82a238",
         13065 => x"608a1122",
         13066 => x"ff057889",
         13067 => x"2a065a56",
         13068 => x"78aa3876",
         13069 => x"849e3888",
         13070 => x"1a085574",
         13071 => x"802e84b1",
         13072 => x"3874812e",
         13073 => x"86a13874",
         13074 => x"ff2e868c",
         13075 => x"3874981b",
         13076 => x"0c881a08",
         13077 => x"85387488",
         13078 => x"1b0c6056",
         13079 => x"b416089c",
         13080 => x"1b082e81",
         13081 => x"d338981a",
         13082 => x"08fe059c",
         13083 => x"1708fe05",
         13084 => x"58587777",
         13085 => x"2785f038",
         13086 => x"8a162270",
         13087 => x"7929b018",
         13088 => x"08055657",
         13089 => x"74802e85",
         13090 => x"de387815",
         13091 => x"7b892a59",
         13092 => x"5c77802e",
         13093 => x"83983877",
         13094 => x"195f767f",
         13095 => x"27853876",
         13096 => x"79315877",
         13097 => x"547b537c",
         13098 => x"52811633",
         13099 => x"51ff9ba1",
         13100 => x"3f84b8e4",
         13101 => x"0885a138",
         13102 => x"60b41108",
         13103 => x"7d315657",
         13104 => x"747827a5",
         13105 => x"3884800b",
         13106 => x"b8187672",
         13107 => x"291f5758",
         13108 => x"56747081",
         13109 => x"05563377",
         13110 => x"70810559",
         13111 => x"34ff1656",
         13112 => x"75ef3860",
         13113 => x"5975831a",
         13114 => x"3477892b",
         13115 => x"597a7931",
         13116 => x"7e081a7f",
         13117 => x"0c791e94",
         13118 => x"1c081b70",
         13119 => x"71941f0c",
         13120 => x"8c1e085a",
         13121 => x"5a575e5b",
         13122 => x"75752783",
         13123 => x"38745675",
         13124 => x"8c1b0c7a",
         13125 => x"fe853890",
         13126 => x"1a335877",
         13127 => x"80c0075b",
         13128 => x"7a901b34",
         13129 => x"80567584",
         13130 => x"b8e40c92",
         13131 => x"3d0d0474",
         13132 => x"84b8e40c",
         13133 => x"923d0d04",
         13134 => x"83163355",
         13135 => x"7482c838",
         13136 => x"6056fea2",
         13137 => x"39609c1b",
         13138 => x"08595676",
         13139 => x"83ff0684",
         13140 => x"8071315a",
         13141 => x"5c7a7927",
         13142 => x"83387a59",
         13143 => x"7757b416",
         13144 => x"08782eb6",
         13145 => x"38800b83",
         13146 => x"1733715e",
         13147 => x"415f7f7f",
         13148 => x"2e098106",
         13149 => x"80d53881",
         13150 => x"547753b8",
         13151 => x"16528116",
         13152 => x"3351ff98",
         13153 => x"cd3f84b8",
         13154 => x"e408802e",
         13155 => x"8538ff57",
         13156 => x"815c76b4",
         13157 => x"170c7b83",
         13158 => x"bf386094",
         13159 => x"1b0883ff",
         13160 => x"06117a58",
         13161 => x"b8057e59",
         13162 => x"56587880",
         13163 => x"2e953876",
         13164 => x"70810558",
         13165 => x"33757081",
         13166 => x"055734ff",
         13167 => x"165675ef",
         13168 => x"38605881",
         13169 => x"0b831934",
         13170 => x"fea33981",
         13171 => x"54b41608",
         13172 => x"53b81670",
         13173 => x"53811733",
         13174 => x"5240ff98",
         13175 => x"f43f815c",
         13176 => x"84b8e408",
         13177 => x"7f2e0981",
         13178 => x"06ffab38",
         13179 => x"84b8e408",
         13180 => x"831734b4",
         13181 => x"1608a817",
         13182 => x"083184b8",
         13183 => x"e4085d55",
         13184 => x"74a01708",
         13185 => x"27fef038",
         13186 => x"82163355",
         13187 => x"74822e09",
         13188 => x"8106fee3",
         13189 => x"388154b4",
         13190 => x"1608a017",
         13191 => x"0805537f",
         13192 => x"52811633",
         13193 => x"51ff98a9",
         13194 => x"3f7e5cfe",
         13195 => x"ca39941a",
         13196 => x"08578c1a",
         13197 => x"08772693",
         13198 => x"38831633",
         13199 => x"407f81b9",
         13200 => x"38607cb4",
         13201 => x"120c941b",
         13202 => x"0858567b",
         13203 => x"7c9c1c0c",
         13204 => x"58fdf839",
         13205 => x"981a0852",
         13206 => x"7951ffab",
         13207 => x"e73f84b8",
         13208 => x"e4085584",
         13209 => x"b8e408fb",
         13210 => x"d838901a",
         13211 => x"3358fdab",
         13212 => x"39765279",
         13213 => x"51ffabcc",
         13214 => x"3f84b8e4",
         13215 => x"085584b8",
         13216 => x"e408fbbd",
         13217 => x"38e43981",
         13218 => x"54b41608",
         13219 => x"53b81670",
         13220 => x"53811733",
         13221 => x"5257ff97",
         13222 => x"b83f84b8",
         13223 => x"e40881b8",
         13224 => x"3884b8e4",
         13225 => x"08831734",
         13226 => x"b41608a8",
         13227 => x"17083158",
         13228 => x"77a01708",
         13229 => x"27fd8938",
         13230 => x"8216335c",
         13231 => x"7b822e09",
         13232 => x"8106fcfc",
         13233 => x"388154b4",
         13234 => x"1608a017",
         13235 => x"08055376",
         13236 => x"52811633",
         13237 => x"51ff96f9",
         13238 => x"3f6056fb",
         13239 => x"89398116",
         13240 => x"3351ff95",
         13241 => x"9b3f84b8",
         13242 => x"e4088106",
         13243 => x"5574f9f2",
         13244 => x"38747a08",
         13245 => x"5657f9ec",
         13246 => x"398154b4",
         13247 => x"160853b8",
         13248 => x"16705381",
         13249 => x"17335257",
         13250 => x"ff96c63f",
         13251 => x"84b8e408",
         13252 => x"80c63884",
         13253 => x"b8e40883",
         13254 => x"1734b416",
         13255 => x"08a81708",
         13256 => x"315574a0",
         13257 => x"170827fe",
         13258 => x"98388216",
         13259 => x"33587782",
         13260 => x"2e098106",
         13261 => x"fe8b3881",
         13262 => x"54b41608",
         13263 => x"a0170805",
         13264 => x"53765281",
         13265 => x"163351ff",
         13266 => x"96873f60",
         13267 => x"7cb4120c",
         13268 => x"941b0858",
         13269 => x"56fdf439",
         13270 => x"810b911b",
         13271 => x"34810b84",
         13272 => x"b8e40c92",
         13273 => x"3d0d0482",
         13274 => x"0b911b34",
         13275 => x"820b84b8",
         13276 => x"e40c923d",
         13277 => x"0d04f53d",
         13278 => x"0d7d5889",
         13279 => x"5a77802e",
         13280 => x"9f387708",
         13281 => x"5675802e",
         13282 => x"97387533",
         13283 => x"5574802e",
         13284 => x"8f388616",
         13285 => x"22841922",
         13286 => x"58597877",
         13287 => x"2e83b538",
         13288 => x"8055745c",
         13289 => x"79567981",
         13290 => x"d8389018",
         13291 => x"3370862a",
         13292 => x"81065c57",
         13293 => x"7a802e81",
         13294 => x"c8387ba0",
         13295 => x"19085a57",
         13296 => x"b4170879",
         13297 => x"2eac3883",
         13298 => x"17335b7a",
         13299 => x"81bc3881",
         13300 => x"547853b8",
         13301 => x"17528117",
         13302 => x"3351ff93",
         13303 => x"f53f84b8",
         13304 => x"e408802e",
         13305 => x"8538ff59",
         13306 => x"815678b4",
         13307 => x"180c7581",
         13308 => x"9038a418",
         13309 => x"088b1133",
         13310 => x"a0075a57",
         13311 => x"788b1834",
         13312 => x"77088819",
         13313 => x"087083ff",
         13314 => x"ff065d5a",
         13315 => x"567a9a18",
         13316 => x"347a882a",
         13317 => x"5a799b18",
         13318 => x"349c1776",
         13319 => x"3396195c",
         13320 => x"565b7483",
         13321 => x"2e81c138",
         13322 => x"8c180855",
         13323 => x"747b3474",
         13324 => x"882a5b7a",
         13325 => x"9d183474",
         13326 => x"902a5675",
         13327 => x"9e183474",
         13328 => x"982a5978",
         13329 => x"9f183480",
         13330 => x"7a34800b",
         13331 => x"971834a1",
         13332 => x"0b981834",
         13333 => x"80cc0b99",
         13334 => x"1834800b",
         13335 => x"92183480",
         13336 => x"0b931834",
         13337 => x"7b5b810b",
         13338 => x"831c347b",
         13339 => x"51ff9694",
         13340 => x"3f84b8e4",
         13341 => x"08901933",
         13342 => x"81bf065b",
         13343 => x"56799019",
         13344 => x"347584b8",
         13345 => x"e40c8d3d",
         13346 => x"0d048154",
         13347 => x"b4170853",
         13348 => x"b8177053",
         13349 => x"81183352",
         13350 => x"5bff93b5",
         13351 => x"3f815684",
         13352 => x"b8e408fe",
         13353 => x"c93884b8",
         13354 => x"e4088318",
         13355 => x"34b41708",
         13356 => x"a8180831",
         13357 => x"84b8e408",
         13358 => x"575574a0",
         13359 => x"180827fe",
         13360 => x"8e388217",
         13361 => x"33557482",
         13362 => x"2e098106",
         13363 => x"fe813881",
         13364 => x"54b41708",
         13365 => x"a0180805",
         13366 => x"537a5281",
         13367 => x"173351ff",
         13368 => x"92ef3f79",
         13369 => x"56fde839",
         13370 => x"78902a55",
         13371 => x"74941834",
         13372 => x"74882a56",
         13373 => x"75951834",
         13374 => x"8c180855",
         13375 => x"747b3474",
         13376 => x"882a5b7a",
         13377 => x"9d183474",
         13378 => x"902a5675",
         13379 => x"9e183474",
         13380 => x"982a5978",
         13381 => x"9f183480",
         13382 => x"7a34800b",
         13383 => x"971834a1",
         13384 => x"0b981834",
         13385 => x"80cc0b99",
         13386 => x"1834800b",
         13387 => x"92183480",
         13388 => x"0b931834",
         13389 => x"7b5b810b",
         13390 => x"831c347b",
         13391 => x"51ff94c4",
         13392 => x"3f84b8e4",
         13393 => x"08901933",
         13394 => x"81bf065b",
         13395 => x"56799019",
         13396 => x"34feae39",
         13397 => x"81163351",
         13398 => x"ff90a53f",
         13399 => x"84b8e408",
         13400 => x"81065574",
         13401 => x"fcba3874",
         13402 => x"7808565a",
         13403 => x"fcb439f9",
         13404 => x"3d0d7970",
         13405 => x"5255fbfe",
         13406 => x"3f84b8e4",
         13407 => x"085484b8",
         13408 => x"e408b138",
         13409 => x"89567480",
         13410 => x"2e9e3874",
         13411 => x"08537280",
         13412 => x"2e963872",
         13413 => x"33527180",
         13414 => x"2e8e3886",
         13415 => x"13228416",
         13416 => x"22585271",
         13417 => x"772e9638",
         13418 => x"80527158",
         13419 => x"75547584",
         13420 => x"3875750c",
         13421 => x"7384b8e4",
         13422 => x"0c893d0d",
         13423 => x"04811333",
         13424 => x"51ff8fbc",
         13425 => x"3f84b8e4",
         13426 => x"08810653",
         13427 => x"72da3873",
         13428 => x"75085356",
         13429 => x"d539f63d",
         13430 => x"0dff7d70",
         13431 => x"5b575b75",
         13432 => x"802eb238",
         13433 => x"75708105",
         13434 => x"5733709f",
         13435 => x"26525271",
         13436 => x"ba2eac38",
         13437 => x"70ee3871",
         13438 => x"ba2ea438",
         13439 => x"84d0c033",
         13440 => x"51807124",
         13441 => x"90387084",
         13442 => x"d0c03480",
         13443 => x"0b84b8e4",
         13444 => x"0c8c3d0d",
         13445 => x"048b0b84",
         13446 => x"b8e40c8c",
         13447 => x"3d0d0478",
         13448 => x"33d01170",
         13449 => x"81ff0653",
         13450 => x"53537089",
         13451 => x"26913882",
         13452 => x"197381ff",
         13453 => x"06d00559",
         13454 => x"5473762e",
         13455 => x"80f53880",
         13456 => x"0b83e4d4",
         13457 => x"5b587908",
         13458 => x"79565776",
         13459 => x"70810558",
         13460 => x"33757081",
         13461 => x"055733ff",
         13462 => x"9f125354",
         13463 => x"52709926",
         13464 => x"8938e012",
         13465 => x"7081ff06",
         13466 => x"5354ff9f",
         13467 => x"13517099",
         13468 => x"268938e0",
         13469 => x"137081ff",
         13470 => x"06545471",
         13471 => x"30709f2a",
         13472 => x"55517173",
         13473 => x"2e098106",
         13474 => x"853873ff",
         13475 => x"be387476",
         13476 => x"32703070",
         13477 => x"72079f2a",
         13478 => x"76075952",
         13479 => x"5276802e",
         13480 => x"92388118",
         13481 => x"841b5b58",
         13482 => x"837825ff",
         13483 => x"99387a51",
         13484 => x"fecf3977",
         13485 => x"8324f738",
         13486 => x"77765e51",
         13487 => x"fec339ea",
         13488 => x"3d0d8053",
         13489 => x"983dcc05",
         13490 => x"52993d51",
         13491 => x"d1943f84",
         13492 => x"b8e40855",
         13493 => x"84b8e408",
         13494 => x"802e8a38",
         13495 => x"7484b8e4",
         13496 => x"0c983d0d",
         13497 => x"047a5c68",
         13498 => x"52983dd0",
         13499 => x"0551c594",
         13500 => x"3f84b8e4",
         13501 => x"085584b8",
         13502 => x"e40880c6",
         13503 => x"380280d7",
         13504 => x"05337098",
         13505 => x"2b585a80",
         13506 => x"772480e2",
         13507 => x"3802b205",
         13508 => x"3370842a",
         13509 => x"81065759",
         13510 => x"75802eb2",
         13511 => x"387a639b",
         13512 => x"11339a12",
         13513 => x"3371882b",
         13514 => x"0773335e",
         13515 => x"5a5b5758",
         13516 => x"79832ea4",
         13517 => x"38769819",
         13518 => x"0c7484b8",
         13519 => x"e40c983d",
         13520 => x"0d0484b8",
         13521 => x"e408842e",
         13522 => x"098106ff",
         13523 => x"8f38850b",
         13524 => x"84b8e40c",
         13525 => x"983d0d04",
         13526 => x"95163394",
         13527 => x"17337198",
         13528 => x"2b71902b",
         13529 => x"07790798",
         13530 => x"1b0c5b54",
         13531 => x"cc397a7e",
         13532 => x"98120c58",
         13533 => x"7484b8e4",
         13534 => x"0c983d0d",
         13535 => x"04ff9e3d",
         13536 => x"0d80e63d",
         13537 => x"0880e63d",
         13538 => x"085d4080",
         13539 => x"7c348053",
         13540 => x"80e43dfd",
         13541 => x"b4055280",
         13542 => x"e53d51cf",
         13543 => x"c53f84b8",
         13544 => x"e4085984",
         13545 => x"b8e40883",
         13546 => x"c8386080",
         13547 => x"d93d0c7f",
         13548 => x"61981108",
         13549 => x"80dd3d0c",
         13550 => x"5880db3d",
         13551 => x"085b5879",
         13552 => x"802e82cc",
         13553 => x"3880d83d",
         13554 => x"983d405b",
         13555 => x"a0527a51",
         13556 => x"ffa4aa3f",
         13557 => x"84b8e408",
         13558 => x"5984b8e4",
         13559 => x"08839238",
         13560 => x"6080df3d",
         13561 => x"085856b4",
         13562 => x"1608772e",
         13563 => x"b13884b8",
         13564 => x"e4088317",
         13565 => x"335f5d7d",
         13566 => x"83c73881",
         13567 => x"547653b8",
         13568 => x"16528116",
         13569 => x"3351ff8b",
         13570 => x"c93f84b8",
         13571 => x"e408802e",
         13572 => x"8538ff57",
         13573 => x"815976b4",
         13574 => x"170c7882",
         13575 => x"d43880df",
         13576 => x"3d089b11",
         13577 => x"339a1233",
         13578 => x"71882b07",
         13579 => x"6370335d",
         13580 => x"40595656",
         13581 => x"78832e82",
         13582 => x"da387680",
         13583 => x"db3d0c80",
         13584 => x"527a51ff",
         13585 => x"a3b73f84",
         13586 => x"b8e40859",
         13587 => x"84b8e408",
         13588 => x"829f3880",
         13589 => x"527a51ff",
         13590 => x"a8f53f84",
         13591 => x"b8e40859",
         13592 => x"84b8e408",
         13593 => x"bb3880df",
         13594 => x"3d089b11",
         13595 => x"339a1233",
         13596 => x"71882b07",
         13597 => x"63703342",
         13598 => x"58595e56",
         13599 => x"7d832e81",
         13600 => x"fd38767a",
         13601 => x"2ea43884",
         13602 => x"b8e40852",
         13603 => x"7a51ffa4",
         13604 => x"e23f84b8",
         13605 => x"e4085984",
         13606 => x"b8e40880",
         13607 => x"2effb438",
         13608 => x"78842e83",
         13609 => x"d8387881",
         13610 => x"c83880e4",
         13611 => x"3dfdb805",
         13612 => x"527a51ff",
         13613 => x"bd893f78",
         13614 => x"7f820533",
         13615 => x"5b577980",
         13616 => x"2e903882",
         13617 => x"1f568117",
         13618 => x"81177033",
         13619 => x"5f57577c",
         13620 => x"f5388117",
         13621 => x"56757826",
         13622 => x"81953876",
         13623 => x"802e9c38",
         13624 => x"7e178205",
         13625 => x"56ff1880",
         13626 => x"e63d0811",
         13627 => x"ff19ff19",
         13628 => x"59595658",
         13629 => x"75337534",
         13630 => x"76eb38ff",
         13631 => x"1880e63d",
         13632 => x"08115f58",
         13633 => x"af7e3480",
         13634 => x"da3d085a",
         13635 => x"79fdbd38",
         13636 => x"77602e82",
         13637 => x"8a38800b",
         13638 => x"84d0c033",
         13639 => x"70101083",
         13640 => x"e4d40570",
         13641 => x"08703343",
         13642 => x"59595e5a",
         13643 => x"7e7a2e8d",
         13644 => x"38811a70",
         13645 => x"17703357",
         13646 => x"5f5a74f5",
         13647 => x"38821a5b",
         13648 => x"7a7826ab",
         13649 => x"38805776",
         13650 => x"7a279438",
         13651 => x"76165f7e",
         13652 => x"337c7081",
         13653 => x"055e3481",
         13654 => x"17577977",
         13655 => x"26ee38ba",
         13656 => x"7c708105",
         13657 => x"5e3476ff",
         13658 => x"2e098106",
         13659 => x"81df3891",
         13660 => x"59807c34",
         13661 => x"7884b8e4",
         13662 => x"0c80e43d",
         13663 => x"0d049516",
         13664 => x"33941733",
         13665 => x"71982b71",
         13666 => x"902b0779",
         13667 => x"0759565e",
         13668 => x"fdf03995",
         13669 => x"16339417",
         13670 => x"3371982b",
         13671 => x"71902b07",
         13672 => x"790780dd",
         13673 => x"3d0c5a5d",
         13674 => x"80527a51",
         13675 => x"ffa0ce3f",
         13676 => x"84b8e408",
         13677 => x"5984b8e4",
         13678 => x"08802efd",
         13679 => x"9638ffb1",
         13680 => x"398154b4",
         13681 => x"160853b8",
         13682 => x"16705381",
         13683 => x"1733525e",
         13684 => x"ff88fe3f",
         13685 => x"815984b8",
         13686 => x"e408fcbe",
         13687 => x"3884b8e4",
         13688 => x"08831734",
         13689 => x"b41608a8",
         13690 => x"17083184",
         13691 => x"b8e4085a",
         13692 => x"5574a017",
         13693 => x"0827fc83",
         13694 => x"38821633",
         13695 => x"5574822e",
         13696 => x"098106fb",
         13697 => x"f6388154",
         13698 => x"b41608a0",
         13699 => x"17080553",
         13700 => x"7d528116",
         13701 => x"3351ff88",
         13702 => x"b83f7c59",
         13703 => x"fbdd39ff",
         13704 => x"1880e63d",
         13705 => x"08115c58",
         13706 => x"af7b3480",
         13707 => x"0b84d0c0",
         13708 => x"33701010",
         13709 => x"83e4d405",
         13710 => x"70087033",
         13711 => x"4359595e",
         13712 => x"5a7e7a2e",
         13713 => x"098106fd",
         13714 => x"e838fdf1",
         13715 => x"3980e53d",
         13716 => x"08188119",
         13717 => x"595a7933",
         13718 => x"7c708105",
         13719 => x"5e347760",
         13720 => x"27fe8e38",
         13721 => x"80e53d08",
         13722 => x"18811959",
         13723 => x"5a79337c",
         13724 => x"7081055e",
         13725 => x"347f7826",
         13726 => x"d438fdf5",
         13727 => x"39825980",
         13728 => x"7c347884",
         13729 => x"b8e40c80",
         13730 => x"e43d0d04",
         13731 => x"f73d0d7b",
         13732 => x"7d585589",
         13733 => x"5674802e",
         13734 => x"9f387408",
         13735 => x"5473802e",
         13736 => x"97387333",
         13737 => x"5372802e",
         13738 => x"8f388614",
         13739 => x"22841622",
         13740 => x"59597878",
         13741 => x"2e83a038",
         13742 => x"8053725a",
         13743 => x"75537581",
         13744 => x"c2389115",
         13745 => x"33537281",
         13746 => x"ba388c15",
         13747 => x"08567676",
         13748 => x"2681b938",
         13749 => x"94150854",
         13750 => x"80587678",
         13751 => x"2e81cc38",
         13752 => x"798a1122",
         13753 => x"70892b52",
         13754 => x"5a567378",
         13755 => x"2e81f738",
         13756 => x"7552ff17",
         13757 => x"51fdbbad",
         13758 => x"3f84b8e4",
         13759 => x"08ff1577",
         13760 => x"54705355",
         13761 => x"53fdbb9d",
         13762 => x"3f84b8e4",
         13763 => x"08732681",
         13764 => x"d5387530",
         13765 => x"74067094",
         13766 => x"170c7771",
         13767 => x"31981708",
         13768 => x"56585973",
         13769 => x"802e8298",
         13770 => x"38757727",
         13771 => x"81d93876",
         13772 => x"76319416",
         13773 => x"08179417",
         13774 => x"0c901633",
         13775 => x"70812a81",
         13776 => x"06515a57",
         13777 => x"78802e81",
         13778 => x"fe387352",
         13779 => x"7451ff99",
         13780 => x"f33f84b8",
         13781 => x"e4085484",
         13782 => x"b8e40880",
         13783 => x"2e81a338",
         13784 => x"73ff2e98",
         13785 => x"38817427",
         13786 => x"82b43879",
         13787 => x"53739c14",
         13788 => x"082782aa",
         13789 => x"38739816",
         13790 => x"0cffae39",
         13791 => x"810b9116",
         13792 => x"34815372",
         13793 => x"84b8e40c",
         13794 => x"8b3d0d04",
         13795 => x"90153370",
         13796 => x"812a8106",
         13797 => x"555873fe",
         13798 => x"bb387594",
         13799 => x"16085557",
         13800 => x"80587678",
         13801 => x"2e098106",
         13802 => x"feb63877",
         13803 => x"94160c94",
         13804 => x"15085475",
         13805 => x"74279038",
         13806 => x"738c160c",
         13807 => x"90153380",
         13808 => x"c0075776",
         13809 => x"90163473",
         13810 => x"83ff0659",
         13811 => x"78802e8c",
         13812 => x"389c1508",
         13813 => x"782e8538",
         13814 => x"779c160c",
         13815 => x"800b84b8",
         13816 => x"e40c8b3d",
         13817 => x"0d04800b",
         13818 => x"94160c88",
         13819 => x"15085473",
         13820 => x"802e80fe",
         13821 => x"38739816",
         13822 => x"0c73802e",
         13823 => x"80c238fe",
         13824 => x"a83984b8",
         13825 => x"e4085794",
         13826 => x"15081794",
         13827 => x"160c7683",
         13828 => x"ff065675",
         13829 => x"802ea938",
         13830 => x"79fe159c",
         13831 => x"1208fe05",
         13832 => x"5a555673",
         13833 => x"782780f6",
         13834 => x"388a1622",
         13835 => x"747129b0",
         13836 => x"18080578",
         13837 => x"892a115a",
         13838 => x"5a537880",
         13839 => x"2e80df38",
         13840 => x"8c150856",
         13841 => x"fee93973",
         13842 => x"527451ff",
         13843 => x"89b73f84",
         13844 => x"b8e40854",
         13845 => x"fe8a3981",
         13846 => x"143351ff",
         13847 => x"82a23f84",
         13848 => x"b8e40881",
         13849 => x"065372fc",
         13850 => x"cf387275",
         13851 => x"085456fc",
         13852 => x"c9397352",
         13853 => x"7451ff97",
         13854 => x"cb3f84b8",
         13855 => x"e4085484",
         13856 => x"b8e40881",
         13857 => x"2e983884",
         13858 => x"b8e408ff",
         13859 => x"2efded38",
         13860 => x"84b8e408",
         13861 => x"88160c73",
         13862 => x"98160cfe",
         13863 => x"dc39820b",
         13864 => x"91163482",
         13865 => x"0b84b8e4",
         13866 => x"0c8b3d0d",
         13867 => x"04f63d0d",
         13868 => x"7c568954",
         13869 => x"75802ea2",
         13870 => x"3880538c",
         13871 => x"3dfc0552",
         13872 => x"8d3d8405",
         13873 => x"51c59b3f",
         13874 => x"84b8e408",
         13875 => x"5584b8e4",
         13876 => x"08802e8f",
         13877 => x"3880760c",
         13878 => x"74547384",
         13879 => x"b8e40c8c",
         13880 => x"3d0d047a",
         13881 => x"760c7d52",
         13882 => x"7551ffb9",
         13883 => x"973f84b8",
         13884 => x"e4085584",
         13885 => x"b8e40880",
         13886 => x"d138ab16",
         13887 => x"3370982b",
         13888 => x"59598078",
         13889 => x"24af3886",
         13890 => x"16337084",
         13891 => x"2a81065b",
         13892 => x"5479802e",
         13893 => x"80c5389c",
         13894 => x"16089b11",
         13895 => x"339a1233",
         13896 => x"71882b07",
         13897 => x"7d70335d",
         13898 => x"5d5a5557",
         13899 => x"78832eb3",
         13900 => x"38778817",
         13901 => x"0c7a5886",
         13902 => x"18228417",
         13903 => x"23745275",
         13904 => x"51ff99b9",
         13905 => x"3f84b8e4",
         13906 => x"08557484",
         13907 => x"2e8d3874",
         13908 => x"802eff84",
         13909 => x"3880760c",
         13910 => x"fefe3985",
         13911 => x"5580760c",
         13912 => x"fef63995",
         13913 => x"17339418",
         13914 => x"3371982b",
         13915 => x"71902b07",
         13916 => x"7a078819",
         13917 => x"0c5a5aff",
         13918 => x"bc39fa3d",
         13919 => x"0d785589",
         13920 => x"5474802e",
         13921 => x"9e387408",
         13922 => x"5372802e",
         13923 => x"96387233",
         13924 => x"5271802e",
         13925 => x"8e388613",
         13926 => x"22841622",
         13927 => x"57527176",
         13928 => x"2e943880",
         13929 => x"52715773",
         13930 => x"84387375",
         13931 => x"0c7384b8",
         13932 => x"e40c883d",
         13933 => x"0d048113",
         13934 => x"3351feff",
         13935 => x"c33f84b8",
         13936 => x"e4088106",
         13937 => x"5271dc38",
         13938 => x"71750853",
         13939 => x"54d739f8",
         13940 => x"3d0d7a7c",
         13941 => x"58558956",
         13942 => x"74802e9f",
         13943 => x"38740854",
         13944 => x"73802e97",
         13945 => x"38733353",
         13946 => x"72802e8f",
         13947 => x"38861422",
         13948 => x"84162259",
         13949 => x"5372782e",
         13950 => x"81973880",
         13951 => x"53725975",
         13952 => x"537580c7",
         13953 => x"3876802e",
         13954 => x"80f33875",
         13955 => x"527451ff",
         13956 => x"9dbd3f84",
         13957 => x"b8e40853",
         13958 => x"84b8e408",
         13959 => x"842eb538",
         13960 => x"84b8e408",
         13961 => x"a6387652",
         13962 => x"7451ffb2",
         13963 => x"923f7252",
         13964 => x"7451ff99",
         13965 => x"be3f84b8",
         13966 => x"e4088432",
         13967 => x"70307072",
         13968 => x"079f2c84",
         13969 => x"b8e40806",
         13970 => x"55575472",
         13971 => x"84b8e40c",
         13972 => x"8a3d0d04",
         13973 => x"75775375",
         13974 => x"5253ffb1",
         13975 => x"e23f7252",
         13976 => x"7451ff99",
         13977 => x"8e3f84b8",
         13978 => x"e4088432",
         13979 => x"70307072",
         13980 => x"079f2c84",
         13981 => x"b8e40806",
         13982 => x"555754cf",
         13983 => x"39755274",
         13984 => x"51ff96f9",
         13985 => x"3f84b8e4",
         13986 => x"0884b8e4",
         13987 => x"0c8a3d0d",
         13988 => x"04811433",
         13989 => x"51fefde8",
         13990 => x"3f84b8e4",
         13991 => x"08810653",
         13992 => x"72fed838",
         13993 => x"72750854",
         13994 => x"56fed239",
         13995 => x"ed3d0d66",
         13996 => x"57805389",
         13997 => x"3d705397",
         13998 => x"3d5256c1",
         13999 => x"a53f84b8",
         14000 => x"e4085584",
         14001 => x"b8e40880",
         14002 => x"2e8a3874",
         14003 => x"84b8e40c",
         14004 => x"953d0d04",
         14005 => x"65527551",
         14006 => x"ffb5a93f",
         14007 => x"84b8e408",
         14008 => x"5584b8e4",
         14009 => x"08e53802",
         14010 => x"80cb0533",
         14011 => x"70982b55",
         14012 => x"58807424",
         14013 => x"97387680",
         14014 => x"2ed13876",
         14015 => x"527551ff",
         14016 => x"b0bd3f74",
         14017 => x"84b8e40c",
         14018 => x"953d0d04",
         14019 => x"860b84b8",
         14020 => x"e40c953d",
         14021 => x"0d04ed3d",
         14022 => x"0d666856",
         14023 => x"5f805395",
         14024 => x"3dec0552",
         14025 => x"963d51c0",
         14026 => x"b93f84b8",
         14027 => x"e4085a84",
         14028 => x"b8e4089a",
         14029 => x"387f750c",
         14030 => x"74089c11",
         14031 => x"08fe1194",
         14032 => x"13085957",
         14033 => x"59577575",
         14034 => x"268d3875",
         14035 => x"7f0c7984",
         14036 => x"b8e40c95",
         14037 => x"3d0d0484",
         14038 => x"b8e40877",
         14039 => x"335a5b78",
         14040 => x"812e8293",
         14041 => x"3877a818",
         14042 => x"0884b8e4",
         14043 => x"085a5d59",
         14044 => x"7780c138",
         14045 => x"7b811d71",
         14046 => x"5c5d56b4",
         14047 => x"1708762e",
         14048 => x"82ef3883",
         14049 => x"1733785f",
         14050 => x"5d7c818d",
         14051 => x"38815475",
         14052 => x"53b81752",
         14053 => x"81173351",
         14054 => x"fefcb73f",
         14055 => x"84b8e408",
         14056 => x"802e8538",
         14057 => x"ff5a815e",
         14058 => x"79b4180c",
         14059 => x"7f7e5b57",
         14060 => x"7d80cc38",
         14061 => x"76335e7d",
         14062 => x"822e828d",
         14063 => x"387717b8",
         14064 => x"05831133",
         14065 => x"82123371",
         14066 => x"902b7188",
         14067 => x"2b078114",
         14068 => x"33707207",
         14069 => x"882b7533",
         14070 => x"7180ffff",
         14071 => x"fe800607",
         14072 => x"70307080",
         14073 => x"25630560",
         14074 => x"840583ff",
         14075 => x"0662ff05",
         14076 => x"43414353",
         14077 => x"54525358",
         14078 => x"405e5678",
         14079 => x"fef2387a",
         14080 => x"7f0c7a94",
         14081 => x"180c8417",
         14082 => x"33810758",
         14083 => x"77841834",
         14084 => x"7984b8e4",
         14085 => x"0c953d0d",
         14086 => x"048154b4",
         14087 => x"170853b8",
         14088 => x"17705381",
         14089 => x"1833525d",
         14090 => x"fefca63f",
         14091 => x"815e84b8",
         14092 => x"e408fef8",
         14093 => x"3884b8e4",
         14094 => x"08831834",
         14095 => x"b41708a8",
         14096 => x"18083184",
         14097 => x"b8e4085f",
         14098 => x"5574a018",
         14099 => x"0827febd",
         14100 => x"38821733",
         14101 => x"5574822e",
         14102 => x"098106fe",
         14103 => x"b0388154",
         14104 => x"b41708a0",
         14105 => x"18080553",
         14106 => x"7c528117",
         14107 => x"3351fefb",
         14108 => x"e03f775e",
         14109 => x"fe973982",
         14110 => x"7742923d",
         14111 => x"59567552",
         14112 => x"7751ff81",
         14113 => x"803f84b8",
         14114 => x"e408ff2e",
         14115 => x"80e83884",
         14116 => x"b8e40881",
         14117 => x"2e80f738",
         14118 => x"84b8e408",
         14119 => x"307084b8",
         14120 => x"e4080780",
         14121 => x"257c0581",
         14122 => x"18625a58",
         14123 => x"5c5c9c17",
         14124 => x"087626ca",
         14125 => x"387a7f0c",
         14126 => x"7a94180c",
         14127 => x"84173381",
         14128 => x"07587784",
         14129 => x"1834fec8",
         14130 => x"397717b8",
         14131 => x"05811133",
         14132 => x"71337188",
         14133 => x"2b077030",
         14134 => x"7080251f",
         14135 => x"821d83ff",
         14136 => x"06ff1f5f",
         14137 => x"5d5f595f",
         14138 => x"5f5578fd",
         14139 => x"8338fe8f",
         14140 => x"39775afd",
         14141 => x"bf398160",
         14142 => x"585a7a7f",
         14143 => x"0c7a9418",
         14144 => x"0c841733",
         14145 => x"81075877",
         14146 => x"841834fe",
         14147 => x"83398260",
         14148 => x"585ae739",
         14149 => x"f73d0d7b",
         14150 => x"57895676",
         14151 => x"802e9f38",
         14152 => x"76085574",
         14153 => x"802e9738",
         14154 => x"74335473",
         14155 => x"802e8f38",
         14156 => x"86152284",
         14157 => x"18225959",
         14158 => x"78782e81",
         14159 => x"da388054",
         14160 => x"735a7580",
         14161 => x"dc389117",
         14162 => x"33567580",
         14163 => x"d4389017",
         14164 => x"3370812a",
         14165 => x"81065558",
         14166 => x"87557380",
         14167 => x"2e80c438",
         14168 => x"94170854",
         14169 => x"738c1808",
         14170 => x"27b73873",
         14171 => x"81d53888",
         14172 => x"17087708",
         14173 => x"57548174",
         14174 => x"2788389c",
         14175 => x"16087426",
         14176 => x"b3388256",
         14177 => x"800b8818",
         14178 => x"0c941708",
         14179 => x"8c180c77",
         14180 => x"80c00759",
         14181 => x"78901834",
         14182 => x"75802e85",
         14183 => x"38759118",
         14184 => x"34755574",
         14185 => x"84b8e40c",
         14186 => x"8b3d0d04",
         14187 => x"78547878",
         14188 => x"2780ff38",
         14189 => x"73527651",
         14190 => x"fefeca3f",
         14191 => x"84b8e408",
         14192 => x"5984b8e4",
         14193 => x"08802e80",
         14194 => x"e93884b8",
         14195 => x"e408812e",
         14196 => x"82d83884",
         14197 => x"b8e408ff",
         14198 => x"2e82e538",
         14199 => x"80537352",
         14200 => x"7551ff85",
         14201 => x"813f84b8",
         14202 => x"e40882c8",
         14203 => x"389c1608",
         14204 => x"fe119418",
         14205 => x"08575558",
         14206 => x"747427ff",
         14207 => x"af388115",
         14208 => x"94170c84",
         14209 => x"16338107",
         14210 => x"54738417",
         14211 => x"34785477",
         14212 => x"7926ffa0",
         14213 => x"389c3981",
         14214 => x"153351fe",
         14215 => x"f6e23f84",
         14216 => x"b8e40881",
         14217 => x"065473fe",
         14218 => x"95387377",
         14219 => x"085556fe",
         14220 => x"8f39800b",
         14221 => x"90183359",
         14222 => x"54735680",
         14223 => x"0b88180c",
         14224 => x"fec73998",
         14225 => x"17085276",
         14226 => x"51fefdb9",
         14227 => x"3f84b8e4",
         14228 => x"08ff2e81",
         14229 => x"c23884b8",
         14230 => x"e408812e",
         14231 => x"81be3875",
         14232 => x"81ae3879",
         14233 => x"5884b8e4",
         14234 => x"089c1908",
         14235 => x"2781a138",
         14236 => x"84b8e408",
         14237 => x"98180878",
         14238 => x"08585654",
         14239 => x"810b84b8",
         14240 => x"e4082781",
         14241 => x"a13884b8",
         14242 => x"e4089c17",
         14243 => x"08278196",
         14244 => x"3874802e",
         14245 => x"9738ff53",
         14246 => x"74527551",
         14247 => x"ff83c73f",
         14248 => x"84b8e408",
         14249 => x"5584b8e4",
         14250 => x"0880e338",
         14251 => x"73527651",
         14252 => x"fefcd23f",
         14253 => x"84b8e408",
         14254 => x"5984b8e4",
         14255 => x"08802e80",
         14256 => x"cb3884b8",
         14257 => x"e408812e",
         14258 => x"80dc3884",
         14259 => x"b8e408ff",
         14260 => x"2e80fe38",
         14261 => x"80537352",
         14262 => x"7551ff83",
         14263 => x"893f84b8",
         14264 => x"e40880e6",
         14265 => x"389c1608",
         14266 => x"fe119418",
         14267 => x"08575558",
         14268 => x"74742790",
         14269 => x"38811594",
         14270 => x"170c8416",
         14271 => x"33810754",
         14272 => x"73841734",
         14273 => x"78547779",
         14274 => x"26ffa138",
         14275 => x"80557456",
         14276 => x"90173358",
         14277 => x"fcf33981",
         14278 => x"56febb39",
         14279 => x"820b9018",
         14280 => x"335956fc",
         14281 => x"e4398256",
         14282 => x"e739820b",
         14283 => x"90183359",
         14284 => x"54fe8639",
         14285 => x"84b8e408",
         14286 => x"90183359",
         14287 => x"54fdfa39",
         14288 => x"810b9018",
         14289 => x"335954fd",
         14290 => x"f03984b8",
         14291 => x"e40856c0",
         14292 => x"398156ff",
         14293 => x"bb39db3d",
         14294 => x"0d8253a7",
         14295 => x"3dff9c05",
         14296 => x"52a83d51",
         14297 => x"ffb7fb3f",
         14298 => x"84b8e408",
         14299 => x"5684b8e4",
         14300 => x"08802e8a",
         14301 => x"387584b8",
         14302 => x"e40ca73d",
         14303 => x"0d047d4b",
         14304 => x"a83d0852",
         14305 => x"9b3d7052",
         14306 => x"59ffabf8",
         14307 => x"3f84b8e4",
         14308 => x"085684b8",
         14309 => x"e408de38",
         14310 => x"02819305",
         14311 => x"3370852a",
         14312 => x"81065957",
         14313 => x"865677cd",
         14314 => x"3876982b",
         14315 => x"5b807b24",
         14316 => x"c4380280",
         14317 => x"ee053370",
         14318 => x"81065d57",
         14319 => x"87567bff",
         14320 => x"b4387da3",
         14321 => x"3d089b11",
         14322 => x"339a1233",
         14323 => x"71882b07",
         14324 => x"7333415e",
         14325 => x"5c57587c",
         14326 => x"832e80d5",
         14327 => x"3876842a",
         14328 => x"81065776",
         14329 => x"802e80ed",
         14330 => x"38875698",
         14331 => x"18087b2e",
         14332 => x"ff833877",
         14333 => x"5f7a4184",
         14334 => x"b8e40852",
         14335 => x"8f3d7052",
         14336 => x"55ff8bf9",
         14337 => x"3f84b8e4",
         14338 => x"085684b8",
         14339 => x"e408fee5",
         14340 => x"3884b8e4",
         14341 => x"08527451",
         14342 => x"ff91b43f",
         14343 => x"84b8e408",
         14344 => x"5684b8e4",
         14345 => x"08a03887",
         14346 => x"0b84b8e4",
         14347 => x"0ca73d0d",
         14348 => x"04951633",
         14349 => x"94173371",
         14350 => x"982b7190",
         14351 => x"2b077d07",
         14352 => x"5d5d5dff",
         14353 => x"983984b8",
         14354 => x"e408842e",
         14355 => x"883884b8",
         14356 => x"e408fea1",
         14357 => x"3878086f",
         14358 => x"a83d0857",
         14359 => x"5d5774ff",
         14360 => x"2e80d338",
         14361 => x"74527851",
         14362 => x"ff8b923f",
         14363 => x"84b8e408",
         14364 => x"5684b8e4",
         14365 => x"08802ebe",
         14366 => x"38753070",
         14367 => x"77078025",
         14368 => x"565a7a80",
         14369 => x"2e9a3874",
         14370 => x"802e9538",
         14371 => x"7a790858",
         14372 => x"55817b27",
         14373 => x"89389c17",
         14374 => x"087b2681",
         14375 => x"fd388256",
         14376 => x"75fdd238",
         14377 => x"7d51fef5",
         14378 => x"db3f84b8",
         14379 => x"e40884b8",
         14380 => x"e40ca73d",
         14381 => x"0d04b817",
         14382 => x"5d981908",
         14383 => x"56805ab4",
         14384 => x"1708762e",
         14385 => x"82b93883",
         14386 => x"17337a59",
         14387 => x"55747a2e",
         14388 => x"09810680",
         14389 => x"dd388154",
         14390 => x"7553b817",
         14391 => x"52811733",
         14392 => x"51fef1ee",
         14393 => x"3f84b8e4",
         14394 => x"08802e85",
         14395 => x"38ff5681",
         14396 => x"5875b418",
         14397 => x"0c775677",
         14398 => x"ab389c19",
         14399 => x"0858e578",
         14400 => x"34810b83",
         14401 => x"18349019",
         14402 => x"087c27fe",
         14403 => x"ec388052",
         14404 => x"7851ff8b",
         14405 => x"de3f84b8",
         14406 => x"e4085684",
         14407 => x"b8e40880",
         14408 => x"2eff9638",
         14409 => x"75842e09",
         14410 => x"8106fecd",
         14411 => x"388256fe",
         14412 => x"c8398154",
         14413 => x"b4170853",
         14414 => x"7c528117",
         14415 => x"3351fef2",
         14416 => x"903f8158",
         14417 => x"84b8e408",
         14418 => x"7a2e0981",
         14419 => x"06ffa638",
         14420 => x"84b8e408",
         14421 => x"831834b4",
         14422 => x"1708a818",
         14423 => x"083184b8",
         14424 => x"e4085955",
         14425 => x"74a01808",
         14426 => x"27feeb38",
         14427 => x"82173355",
         14428 => x"74822e09",
         14429 => x"8106fede",
         14430 => x"388154b4",
         14431 => x"1708a018",
         14432 => x"0805537c",
         14433 => x"52811733",
         14434 => x"51fef1c5",
         14435 => x"3f7958fe",
         14436 => x"c5397955",
         14437 => x"79782780",
         14438 => x"e1387452",
         14439 => x"7851fef6",
         14440 => x"e43f84b8",
         14441 => x"e4085a84",
         14442 => x"b8e40880",
         14443 => x"2e80cb38",
         14444 => x"84b8e408",
         14445 => x"812efde6",
         14446 => x"3884b8e4",
         14447 => x"08ff2e80",
         14448 => x"cb388053",
         14449 => x"74527651",
         14450 => x"fefd9b3f",
         14451 => x"84b8e408",
         14452 => x"b3389c17",
         14453 => x"08fe1194",
         14454 => x"1908585c",
         14455 => x"58757b27",
         14456 => x"ffb03881",
         14457 => x"1694180c",
         14458 => x"84173381",
         14459 => x"075c7b84",
         14460 => x"18347955",
         14461 => x"777a26ff",
         14462 => x"a1388056",
         14463 => x"fda23979",
         14464 => x"56fdf739",
         14465 => x"84b8e408",
         14466 => x"56fd9539",
         14467 => x"8156fd90",
         14468 => x"39e33d0d",
         14469 => x"82539f3d",
         14470 => x"ffbc0552",
         14471 => x"a03d51ff",
         14472 => x"b2c03f84",
         14473 => x"b8e40856",
         14474 => x"84b8e408",
         14475 => x"802e8a38",
         14476 => x"7584b8e4",
         14477 => x"0c9f3d0d",
         14478 => x"047d436f",
         14479 => x"52933d70",
         14480 => x"525affa6",
         14481 => x"bf3f84b8",
         14482 => x"e4085684",
         14483 => x"b8e4088b",
         14484 => x"38880b84",
         14485 => x"b8e40c9f",
         14486 => x"3d0d0484",
         14487 => x"b8e40884",
         14488 => x"2e098106",
         14489 => x"cb380280",
         14490 => x"f3053370",
         14491 => x"852a8106",
         14492 => x"56588656",
         14493 => x"74ffb938",
         14494 => x"7d5f7452",
         14495 => x"8f3d7052",
         14496 => x"5dff83c0",
         14497 => x"3f84b8e4",
         14498 => x"0875575c",
         14499 => x"84b8e408",
         14500 => x"83388756",
         14501 => x"84b8e408",
         14502 => x"812e80f9",
         14503 => x"3884b8e4",
         14504 => x"08ff2e81",
         14505 => x"cb387581",
         14506 => x"c9387d84",
         14507 => x"b8e40883",
         14508 => x"12335d5a",
         14509 => x"577a80e2",
         14510 => x"38fe199c",
         14511 => x"1808fe05",
         14512 => x"5a56805b",
         14513 => x"7579278d",
         14514 => x"388a1722",
         14515 => x"767129b0",
         14516 => x"1908055c",
         14517 => x"587ab418",
         14518 => x"0cb81759",
         14519 => x"84807957",
         14520 => x"55807670",
         14521 => x"81055834",
         14522 => x"ff155574",
         14523 => x"f4387458",
         14524 => x"8a172255",
         14525 => x"77752781",
         14526 => x"f9388154",
         14527 => x"771b5378",
         14528 => x"52811733",
         14529 => x"51feeec9",
         14530 => x"3f84b8e4",
         14531 => x"0881df38",
         14532 => x"811858dc",
         14533 => x"398256ff",
         14534 => x"84398154",
         14535 => x"b4170853",
         14536 => x"b8177053",
         14537 => x"81183352",
         14538 => x"58feeea5",
         14539 => x"3f815684",
         14540 => x"b8e408be",
         14541 => x"3884b8e4",
         14542 => x"08831834",
         14543 => x"b41708a8",
         14544 => x"18083155",
         14545 => x"74a01808",
         14546 => x"27feee38",
         14547 => x"8217335b",
         14548 => x"7a822e09",
         14549 => x"8106fee1",
         14550 => x"387554b4",
         14551 => x"1708a018",
         14552 => x"08055377",
         14553 => x"52811733",
         14554 => x"51feede5",
         14555 => x"3ffeca39",
         14556 => x"81567b7d",
         14557 => x"08585581",
         14558 => x"7c27fdb4",
         14559 => x"387b9c18",
         14560 => x"0827fdac",
         14561 => x"3874527c",
         14562 => x"51fef2f9",
         14563 => x"3f84b8e4",
         14564 => x"085a84b8",
         14565 => x"e408802e",
         14566 => x"fd963884",
         14567 => x"b8e40881",
         14568 => x"2efd8d38",
         14569 => x"84b8e408",
         14570 => x"ff2efd84",
         14571 => x"38805374",
         14572 => x"527651fe",
         14573 => x"f9b03f84",
         14574 => x"b8e408fc",
         14575 => x"f3389c17",
         14576 => x"08fe1194",
         14577 => x"19085a5c",
         14578 => x"59777b27",
         14579 => x"90388118",
         14580 => x"94180c84",
         14581 => x"17338107",
         14582 => x"5c7b8418",
         14583 => x"34795578",
         14584 => x"7a26ffa1",
         14585 => x"387584b8",
         14586 => x"e40c9f3d",
         14587 => x"0d048a17",
         14588 => x"22557483",
         14589 => x"ffff0657",
         14590 => x"81567678",
         14591 => x"2e098106",
         14592 => x"fef0388b",
         14593 => x"0bb81f56",
         14594 => x"56a07570",
         14595 => x"81055734",
         14596 => x"ff165675",
         14597 => x"f4387d57",
         14598 => x"ae0bb818",
         14599 => x"347d5890",
         14600 => x"0b80c319",
         14601 => x"347d5975",
         14602 => x"80ce1a34",
         14603 => x"7580cf1a",
         14604 => x"34a10b80",
         14605 => x"d01a3480",
         14606 => x"cc0b80d1",
         14607 => x"1a347d7c",
         14608 => x"83ffff06",
         14609 => x"59567780",
         14610 => x"d2173477",
         14611 => x"882a5b7a",
         14612 => x"80d31734",
         14613 => x"75335574",
         14614 => x"832e81cc",
         14615 => x"387d59a0",
         14616 => x"0b80d81a",
         14617 => x"b81b5758",
         14618 => x"56747081",
         14619 => x"05563377",
         14620 => x"70810559",
         14621 => x"34ff1656",
         14622 => x"75ef387d",
         14623 => x"56ae0b80",
         14624 => x"d9173464",
         14625 => x"7e7183ff",
         14626 => x"ff065b57",
         14627 => x"577880f2",
         14628 => x"17347888",
         14629 => x"2a5b7a80",
         14630 => x"f3173475",
         14631 => x"33557483",
         14632 => x"2e80f038",
         14633 => x"7d5b810b",
         14634 => x"831c3479",
         14635 => x"51ff9296",
         14636 => x"3f84b8e4",
         14637 => x"085684b8",
         14638 => x"e408fdb6",
         14639 => x"38695684",
         14640 => x"b8e40896",
         14641 => x"173484b8",
         14642 => x"e4089717",
         14643 => x"34a10b98",
         14644 => x"173480cc",
         14645 => x"0b991734",
         14646 => x"7d6a585d",
         14647 => x"779a1834",
         14648 => x"77882a59",
         14649 => x"789b1834",
         14650 => x"7c335a79",
         14651 => x"832e80d9",
         14652 => x"38695590",
         14653 => x"0b8b1634",
         14654 => x"7d57810b",
         14655 => x"8318347d",
         14656 => x"51feed80",
         14657 => x"3f84b8e4",
         14658 => x"08567584",
         14659 => x"b8e40c9f",
         14660 => x"3d0d0476",
         14661 => x"902a5574",
         14662 => x"80ec1734",
         14663 => x"74882a57",
         14664 => x"7680ed17",
         14665 => x"34fefd39",
         14666 => x"7b902a5b",
         14667 => x"7a80cc17",
         14668 => x"347a882a",
         14669 => x"557480cd",
         14670 => x"17347d59",
         14671 => x"a00b80d8",
         14672 => x"1ab81b57",
         14673 => x"5856fea1",
         14674 => x"397b902a",
         14675 => x"58779418",
         14676 => x"3477882a",
         14677 => x"5c7b9518",
         14678 => x"34695590",
         14679 => x"0b8b1634",
         14680 => x"7d57810b",
         14681 => x"8318347d",
         14682 => x"51feec98",
         14683 => x"3f84b8e4",
         14684 => x"0856ff96",
         14685 => x"39d13d0d",
         14686 => x"b33db43d",
         14687 => x"0870595b",
         14688 => x"5f79802e",
         14689 => x"9b387970",
         14690 => x"81055b33",
         14691 => x"709f2656",
         14692 => x"5675ba2e",
         14693 => x"81b83874",
         14694 => x"ed3875ba",
         14695 => x"2e81af38",
         14696 => x"8253b13d",
         14697 => x"fefc0552",
         14698 => x"b23d51ff",
         14699 => x"abb43f84",
         14700 => x"b8e40856",
         14701 => x"84b8e408",
         14702 => x"802e8a38",
         14703 => x"7584b8e4",
         14704 => x"0cb13d0d",
         14705 => x"047fa63d",
         14706 => x"0cb23d08",
         14707 => x"52a53d70",
         14708 => x"5259ff9f",
         14709 => x"af3f84b8",
         14710 => x"e4085684",
         14711 => x"b8e408dc",
         14712 => x"380281bb",
         14713 => x"053381a0",
         14714 => x"065d8656",
         14715 => x"7cce38a0",
         14716 => x"0b923dae",
         14717 => x"3d085858",
         14718 => x"55757081",
         14719 => x"05573377",
         14720 => x"70810559",
         14721 => x"34ff1555",
         14722 => x"74ef3899",
         14723 => x"3d58b078",
         14724 => x"7a585855",
         14725 => x"75708105",
         14726 => x"57337770",
         14727 => x"81055934",
         14728 => x"ff155574",
         14729 => x"ef38b33d",
         14730 => x"08527751",
         14731 => x"ff9ed53f",
         14732 => x"84b8e408",
         14733 => x"5684b8e4",
         14734 => x"0885d838",
         14735 => x"6aa83d08",
         14736 => x"2e81cb38",
         14737 => x"880b84b8",
         14738 => x"e40cb13d",
         14739 => x"0d047633",
         14740 => x"d0117081",
         14741 => x"ff065757",
         14742 => x"58748926",
         14743 => x"91388217",
         14744 => x"7881ff06",
         14745 => x"d0055d59",
         14746 => x"787a2e80",
         14747 => x"fa38807f",
         14748 => x"0883e4d4",
         14749 => x"7008725d",
         14750 => x"5e5f5f5c",
         14751 => x"7a708105",
         14752 => x"5c337970",
         14753 => x"81055b33",
         14754 => x"ff9f125a",
         14755 => x"58567799",
         14756 => x"268938e0",
         14757 => x"167081ff",
         14758 => x"065755ff",
         14759 => x"9f175877",
         14760 => x"99268938",
         14761 => x"e0177081",
         14762 => x"ff065855",
         14763 => x"7530709f",
         14764 => x"2a595575",
         14765 => x"772e0981",
         14766 => x"06853877",
         14767 => x"ffbe3878",
         14768 => x"7a327030",
         14769 => x"7072079f",
         14770 => x"2a7a075d",
         14771 => x"58557a80",
         14772 => x"2e953881",
         14773 => x"1c841e5e",
         14774 => x"5c7b8324",
         14775 => x"fdc2387c",
         14776 => x"087e5a5b",
         14777 => x"ff96397b",
         14778 => x"8324fdb4",
         14779 => x"38797f0c",
         14780 => x"8253b13d",
         14781 => x"fefc0552",
         14782 => x"b23d51ff",
         14783 => x"a8e43f84",
         14784 => x"b8e40856",
         14785 => x"84b8e408",
         14786 => x"fdb238fd",
         14787 => x"b8396caa",
         14788 => x"3d082e09",
         14789 => x"8106feac",
         14790 => x"387751ff",
         14791 => x"8da83f84",
         14792 => x"b8e40856",
         14793 => x"84b8e408",
         14794 => x"fd92386f",
         14795 => x"58930b8d",
         14796 => x"19028805",
         14797 => x"80cd0558",
         14798 => x"565a7570",
         14799 => x"81055733",
         14800 => x"75708105",
         14801 => x"5734ff1a",
         14802 => x"5a79ef38",
         14803 => x"0280cb05",
         14804 => x"338b1934",
         14805 => x"8b183370",
         14806 => x"842a8106",
         14807 => x"40567e89",
         14808 => x"3875a007",
         14809 => x"57768b19",
         14810 => x"347f5d81",
         14811 => x"0b831e34",
         14812 => x"8b183370",
         14813 => x"842a8106",
         14814 => x"575c7580",
         14815 => x"2e81c538",
         14816 => x"a73d086b",
         14817 => x"2e81bd38",
         14818 => x"7f9b1933",
         14819 => x"9a1a3371",
         14820 => x"882b0772",
         14821 => x"3341585c",
         14822 => x"577d832e",
         14823 => x"82e038fe",
         14824 => x"169c1808",
         14825 => x"fe055e56",
         14826 => x"757d2782",
         14827 => x"c7388a17",
         14828 => x"22767129",
         14829 => x"b0190805",
         14830 => x"575e7580",
         14831 => x"2e82b538",
         14832 => x"757a5d58",
         14833 => x"b4170876",
         14834 => x"2eaa3883",
         14835 => x"17335f7e",
         14836 => x"83bc3881",
         14837 => x"547553b8",
         14838 => x"17528117",
         14839 => x"3351fee3",
         14840 => x"f13f84b8",
         14841 => x"e408802e",
         14842 => x"8538ff58",
         14843 => x"815c77b4",
         14844 => x"180c7f57",
         14845 => x"7b80d818",
         14846 => x"56567bfb",
         14847 => x"bf388115",
         14848 => x"335a79ae",
         14849 => x"2e098106",
         14850 => x"bb386a70",
         14851 => x"83ffff06",
         14852 => x"5d567b80",
         14853 => x"f218347b",
         14854 => x"882a5877",
         14855 => x"80f31834",
         14856 => x"76335b7a",
         14857 => x"832e0981",
         14858 => x"06933875",
         14859 => x"902a5e7d",
         14860 => x"80ec1834",
         14861 => x"7d882a56",
         14862 => x"7580ed18",
         14863 => x"347f5781",
         14864 => x"0b831834",
         14865 => x"7808aa3d",
         14866 => x"08b23d08",
         14867 => x"575c5674",
         14868 => x"ff2e9538",
         14869 => x"74527851",
         14870 => x"fefba23f",
         14871 => x"84b8e408",
         14872 => x"5584b8e4",
         14873 => x"0880f538",
         14874 => x"b8165c98",
         14875 => x"19085780",
         14876 => x"5ab41608",
         14877 => x"772eb438",
         14878 => x"8316337a",
         14879 => x"595f7e7a",
         14880 => x"2e098106",
         14881 => x"81a83881",
         14882 => x"547653b8",
         14883 => x"16528116",
         14884 => x"3351fee2",
         14885 => x"bd3f84b8",
         14886 => x"e408802e",
         14887 => x"8538ff57",
         14888 => x"815876b4",
         14889 => x"170c7755",
         14890 => x"77aa389c",
         14891 => x"19085ae5",
         14892 => x"7a34810b",
         14893 => x"83173490",
         14894 => x"19087b27",
         14895 => x"a5388052",
         14896 => x"7851fefc",
         14897 => x"ae3f84b8",
         14898 => x"e4085584",
         14899 => x"b8e40880",
         14900 => x"2eff9838",
         14901 => x"82567484",
         14902 => x"2ef9e138",
         14903 => x"745674f9",
         14904 => x"db387f51",
         14905 => x"fee59d3f",
         14906 => x"84b8e408",
         14907 => x"84b8e40c",
         14908 => x"b13d0d04",
         14909 => x"820b84b8",
         14910 => x"e40cb13d",
         14911 => x"0d049518",
         14912 => x"33941933",
         14913 => x"71982b71",
         14914 => x"902b0778",
         14915 => x"0758565c",
         14916 => x"fd8d3984",
         14917 => x"b8e40884",
         14918 => x"2efbfe38",
         14919 => x"84b8e408",
         14920 => x"802efea0",
         14921 => x"387584b8",
         14922 => x"e40cb13d",
         14923 => x"0d048154",
         14924 => x"b4160853",
         14925 => x"7b528116",
         14926 => x"3351fee2",
         14927 => x"943f8158",
         14928 => x"84b8e408",
         14929 => x"7a2e0981",
         14930 => x"06fedb38",
         14931 => x"84b8e408",
         14932 => x"831734b4",
         14933 => x"1608a817",
         14934 => x"083184b8",
         14935 => x"e4085955",
         14936 => x"74a01708",
         14937 => x"27fea038",
         14938 => x"8216335d",
         14939 => x"7c822e09",
         14940 => x"8106fe93",
         14941 => x"388154b4",
         14942 => x"1608a017",
         14943 => x"0805537b",
         14944 => x"52811633",
         14945 => x"51fee1c9",
         14946 => x"3f7958fd",
         14947 => x"fa398154",
         14948 => x"b4170853",
         14949 => x"b8177053",
         14950 => x"81183352",
         14951 => x"5bfee1b1",
         14952 => x"3f815c84",
         14953 => x"b8e408fc",
         14954 => x"c93884b8",
         14955 => x"e4088318",
         14956 => x"34b41708",
         14957 => x"a8180831",
         14958 => x"84b8e408",
         14959 => x"5d5574a0",
         14960 => x"180827fc",
         14961 => x"8e388217",
         14962 => x"335d7c82",
         14963 => x"2e098106",
         14964 => x"fc813881",
         14965 => x"54b41708",
         14966 => x"a0180805",
         14967 => x"537a5281",
         14968 => x"173351fe",
         14969 => x"e0eb3f79",
         14970 => x"5cfbe839",
         14971 => x"ec3d0d02",
         14972 => x"80df0533",
         14973 => x"02840580",
         14974 => x"e3053356",
         14975 => x"57825396",
         14976 => x"3dcc0552",
         14977 => x"973d51ff",
         14978 => x"a2d83f84",
         14979 => x"b8e40856",
         14980 => x"84b8e408",
         14981 => x"802e8a38",
         14982 => x"7584b8e4",
         14983 => x"0c963d0d",
         14984 => x"04785a66",
         14985 => x"52963dd0",
         14986 => x"0551ff96",
         14987 => x"d73f84b8",
         14988 => x"e4085684",
         14989 => x"b8e408e0",
         14990 => x"380280cf",
         14991 => x"053381a0",
         14992 => x"06548656",
         14993 => x"73d23874",
         14994 => x"a7066171",
         14995 => x"098b1233",
         14996 => x"71067a74",
         14997 => x"06075156",
         14998 => x"5755738b",
         14999 => x"17347855",
         15000 => x"810b8316",
         15001 => x"347851fe",
         15002 => x"e29a3f84",
         15003 => x"b8e40884",
         15004 => x"b8e40c96",
         15005 => x"3d0d04ec",
         15006 => x"3d0d6757",
         15007 => x"8253963d",
         15008 => x"cc055297",
         15009 => x"3d51ffa1",
         15010 => x"d93f84b8",
         15011 => x"e4085584",
         15012 => x"b8e40880",
         15013 => x"2e8a3874",
         15014 => x"84b8e40c",
         15015 => x"963d0d04",
         15016 => x"785a6652",
         15017 => x"963dd005",
         15018 => x"51ff95d8",
         15019 => x"3f84b8e4",
         15020 => x"085584b8",
         15021 => x"e408e038",
         15022 => x"0280cf05",
         15023 => x"3381a006",
         15024 => x"56865575",
         15025 => x"d2386084",
         15026 => x"18228619",
         15027 => x"2271902b",
         15028 => x"07595956",
         15029 => x"76961734",
         15030 => x"76882a55",
         15031 => x"74971734",
         15032 => x"76902a58",
         15033 => x"77981734",
         15034 => x"76982a54",
         15035 => x"73991734",
         15036 => x"7857810b",
         15037 => x"83183478",
         15038 => x"51fee188",
         15039 => x"3f84b8e4",
         15040 => x"0884b8e4",
         15041 => x"0c963d0d",
         15042 => x"04e83d0d",
         15043 => x"6b6d5d5b",
         15044 => x"80539a3d",
         15045 => x"cc05529b",
         15046 => x"3d51ffa0",
         15047 => x"c53f84b8",
         15048 => x"e40884b8",
         15049 => x"e4083070",
         15050 => x"84b8e408",
         15051 => x"07802551",
         15052 => x"56577a80",
         15053 => x"2e8b3881",
         15054 => x"7076065a",
         15055 => x"567881a4",
         15056 => x"38763070",
         15057 => x"78078025",
         15058 => x"565b7b80",
         15059 => x"2e818c38",
         15060 => x"81707606",
         15061 => x"5a587880",
         15062 => x"2e818038",
         15063 => x"7ca41108",
         15064 => x"5856805a",
         15065 => x"b4160877",
         15066 => x"2e82f638",
         15067 => x"8316337a",
         15068 => x"5a55747a",
         15069 => x"2e098106",
         15070 => x"81983881",
         15071 => x"547653b8",
         15072 => x"16528116",
         15073 => x"3351fedc",
         15074 => x"c93f84b8",
         15075 => x"e408802e",
         15076 => x"8538ff57",
         15077 => x"815976b4",
         15078 => x"170c7857",
         15079 => x"78bd387c",
         15080 => x"70335658",
         15081 => x"80c35674",
         15082 => x"832e8b38",
         15083 => x"80e45674",
         15084 => x"842e8338",
         15085 => x"a7567518",
         15086 => x"b8058311",
         15087 => x"33821233",
         15088 => x"71902b71",
         15089 => x"882b0781",
         15090 => x"14337072",
         15091 => x"07882b75",
         15092 => x"33710762",
         15093 => x"0c5f5d5e",
         15094 => x"57595676",
         15095 => x"84b8e40c",
         15096 => x"9a3d0d04",
         15097 => x"7c5e8040",
         15098 => x"80528e3d",
         15099 => x"705255fe",
         15100 => x"f48b3f84",
         15101 => x"b8e40857",
         15102 => x"84b8e408",
         15103 => x"802e818d",
         15104 => x"3876842e",
         15105 => x"098106fe",
         15106 => x"b838807b",
         15107 => x"348057fe",
         15108 => x"b0397754",
         15109 => x"b4160853",
         15110 => x"b8167053",
         15111 => x"81173352",
         15112 => x"5bfedcad",
         15113 => x"3f775984",
         15114 => x"b8e4087a",
         15115 => x"2e098106",
         15116 => x"fee83884",
         15117 => x"b8e40883",
         15118 => x"1734b416",
         15119 => x"08a81708",
         15120 => x"3184b8e4",
         15121 => x"085a5574",
         15122 => x"a0170827",
         15123 => x"fead3882",
         15124 => x"16335574",
         15125 => x"822e0981",
         15126 => x"06fea038",
         15127 => x"7754b416",
         15128 => x"08a01708",
         15129 => x"05537a52",
         15130 => x"81163351",
         15131 => x"fedbe23f",
         15132 => x"79598154",
         15133 => x"7653b816",
         15134 => x"52811633",
         15135 => x"51fedad2",
         15136 => x"3f84b8e4",
         15137 => x"08802efe",
         15138 => x"8d38fe86",
         15139 => x"39755274",
         15140 => x"51fef8bb",
         15141 => x"3f84b8e4",
         15142 => x"085784b8",
         15143 => x"e408fee1",
         15144 => x"3884b8e4",
         15145 => x"0884b8e4",
         15146 => x"08665c59",
         15147 => x"59791881",
         15148 => x"197c1b57",
         15149 => x"59567533",
         15150 => x"75348119",
         15151 => x"598a7827",
         15152 => x"ec388b70",
         15153 => x"1c575880",
         15154 => x"76347780",
         15155 => x"2efcf238",
         15156 => x"ff187b11",
         15157 => x"70335c57",
         15158 => x"5879a02e",
         15159 => x"ea38fce1",
         15160 => x"397957fd",
         15161 => x"ba39e13d",
         15162 => x"0d8253a1",
         15163 => x"3dffb405",
         15164 => x"52a23d51",
         15165 => x"ff9ceb3f",
         15166 => x"84b8e408",
         15167 => x"5684b8e4",
         15168 => x"0882a638",
         15169 => x"8f3d5d8b",
         15170 => x"7d5755a0",
         15171 => x"76708105",
         15172 => x"5834ff15",
         15173 => x"5574f438",
         15174 => x"74a33d08",
         15175 => x"70337081",
         15176 => x"ff065b58",
         15177 => x"585a9f78",
         15178 => x"2781b738",
         15179 => x"a23d903d",
         15180 => x"5c5c7581",
         15181 => x"ff068118",
         15182 => x"57557481",
         15183 => x"f538757c",
         15184 => x"0c7483ff",
         15185 => x"ff2681ff",
         15186 => x"387451a1",
         15187 => x"953f83b5",
         15188 => x"5284b8e4",
         15189 => x"08519fdc",
         15190 => x"3f84b8e4",
         15191 => x"0883ffff",
         15192 => x"06577680",
         15193 => x"2e81e038",
         15194 => x"83e5f40b",
         15195 => x"83e5f433",
         15196 => x"7081ff06",
         15197 => x"5b565878",
         15198 => x"802e81d6",
         15199 => x"38745678",
         15200 => x"772e9938",
         15201 => x"81187033",
         15202 => x"7081ff06",
         15203 => x"57575874",
         15204 => x"802e8938",
         15205 => x"74772e09",
         15206 => x"8106e938",
         15207 => x"7581ff06",
         15208 => x"597881a3",
         15209 => x"3881ff77",
         15210 => x"2781f838",
         15211 => x"79892681",
         15212 => x"963881ff",
         15213 => x"77278f38",
         15214 => x"76882a55",
         15215 => x"747b7081",
         15216 => x"055d3481",
         15217 => x"1a5a767b",
         15218 => x"7081055d",
         15219 => x"34811aa3",
         15220 => x"3d087033",
         15221 => x"7081ff06",
         15222 => x"5b58585a",
         15223 => x"779f26fe",
         15224 => x"d1388f3d",
         15225 => x"33578656",
         15226 => x"7681e52e",
         15227 => x"bc387980",
         15228 => x"2e993802",
         15229 => x"b7055679",
         15230 => x"1670335c",
         15231 => x"5c7aa02e",
         15232 => x"09810687",
         15233 => x"38ff1a5a",
         15234 => x"79ed387d",
         15235 => x"45804780",
         15236 => x"52953d70",
         15237 => x"5256feef",
         15238 => x"e43f84b8",
         15239 => x"e4085584",
         15240 => x"b8e40880",
         15241 => x"2eb43874",
         15242 => x"567584b8",
         15243 => x"e40ca13d",
         15244 => x"0d0483b5",
         15245 => x"5274519e",
         15246 => x"e73f84b8",
         15247 => x"e40883ff",
         15248 => x"ff065574",
         15249 => x"fdf83886",
         15250 => x"567584b8",
         15251 => x"e40ca13d",
         15252 => x"0d0483e5",
         15253 => x"f43356fe",
         15254 => x"c3398152",
         15255 => x"7551fef4",
         15256 => x"ee3f84b8",
         15257 => x"e4085584",
         15258 => x"b8e40880",
         15259 => x"c1387980",
         15260 => x"2e82c438",
         15261 => x"8b6c7e59",
         15262 => x"57557670",
         15263 => x"81055833",
         15264 => x"76708105",
         15265 => x"5834ff15",
         15266 => x"5574ef38",
         15267 => x"7d5d810b",
         15268 => x"831e347d",
         15269 => x"51fed9ec",
         15270 => x"3f84b8e4",
         15271 => x"08557456",
         15272 => x"ff87398a",
         15273 => x"7a27fe8a",
         15274 => x"388656ff",
         15275 => x"9c3984b8",
         15276 => x"e408842e",
         15277 => x"098106fe",
         15278 => x"ee388055",
         15279 => x"79752efe",
         15280 => x"e6387508",
         15281 => x"75537652",
         15282 => x"58feeeb1",
         15283 => x"3f84b8e4",
         15284 => x"085784b8",
         15285 => x"e408752e",
         15286 => x"09810681",
         15287 => x"843884b8",
         15288 => x"e408b819",
         15289 => x"5c5a9816",
         15290 => x"08578059",
         15291 => x"b4180877",
         15292 => x"2eb23883",
         15293 => x"18335574",
         15294 => x"792e0981",
         15295 => x"0681d738",
         15296 => x"81547653",
         15297 => x"b8185281",
         15298 => x"183351fe",
         15299 => x"d5c43f84",
         15300 => x"b8e40880",
         15301 => x"2e8538ff",
         15302 => x"57815976",
         15303 => x"b4190c78",
         15304 => x"5778be38",
         15305 => x"789c1708",
         15306 => x"7033575a",
         15307 => x"577481e5",
         15308 => x"2e819e38",
         15309 => x"74307080",
         15310 => x"25780756",
         15311 => x"5c74802e",
         15312 => x"81d73881",
         15313 => x"1a5a7981",
         15314 => x"2ea53881",
         15315 => x"527551fe",
         15316 => x"efa13f84",
         15317 => x"b8e40857",
         15318 => x"84b8e408",
         15319 => x"802eff86",
         15320 => x"38875576",
         15321 => x"842efdbf",
         15322 => x"38765576",
         15323 => x"fdb938a0",
         15324 => x"6c575580",
         15325 => x"76708105",
         15326 => x"5834ff15",
         15327 => x"5574f438",
         15328 => x"6b56880b",
         15329 => x"8b17348b",
         15330 => x"6c7e5957",
         15331 => x"55767081",
         15332 => x"05583376",
         15333 => x"70810558",
         15334 => x"34ff1555",
         15335 => x"74802efd",
         15336 => x"eb387670",
         15337 => x"81055833",
         15338 => x"76708105",
         15339 => x"5834ff15",
         15340 => x"5574da38",
         15341 => x"fdd6396b",
         15342 => x"5ae57a34",
         15343 => x"7d5d810b",
         15344 => x"831e347d",
         15345 => x"51fed7bc",
         15346 => x"3f84b8e4",
         15347 => x"0855fdce",
         15348 => x"398157fe",
         15349 => x"df398154",
         15350 => x"b4180853",
         15351 => x"7a528118",
         15352 => x"3351fed4",
         15353 => x"ec3f84b8",
         15354 => x"e408792e",
         15355 => x"09810680",
         15356 => x"c33884b8",
         15357 => x"e4088319",
         15358 => x"34b41808",
         15359 => x"a8190831",
         15360 => x"5c7ba019",
         15361 => x"08278a38",
         15362 => x"82183355",
         15363 => x"74822eb1",
         15364 => x"3884b8e4",
         15365 => x"0859fde8",
         15366 => x"39745a81",
         15367 => x"527551fe",
         15368 => x"edd13f84",
         15369 => x"b8e40857",
         15370 => x"84b8e408",
         15371 => x"802efdb6",
         15372 => x"38feae39",
         15373 => x"81705859",
         15374 => x"78802efd",
         15375 => x"e738fea1",
         15376 => x"398154b4",
         15377 => x"1808a019",
         15378 => x"0805537a",
         15379 => x"52811833",
         15380 => x"51fed3fd",
         15381 => x"3ffda939",
         15382 => x"f23d0d60",
         15383 => x"62028805",
         15384 => x"80cb0533",
         15385 => x"5e5b5789",
         15386 => x"5676802e",
         15387 => x"9f387608",
         15388 => x"5574802e",
         15389 => x"97387433",
         15390 => x"5473802e",
         15391 => x"8f388615",
         15392 => x"22841822",
         15393 => x"59597878",
         15394 => x"2e81c238",
         15395 => x"8054735f",
         15396 => x"7581a538",
         15397 => x"91173356",
         15398 => x"75819d38",
         15399 => x"79802e81",
         15400 => x"a2388c17",
         15401 => x"08819c38",
         15402 => x"90173370",
         15403 => x"812a8106",
         15404 => x"565d7480",
         15405 => x"2e818c38",
         15406 => x"7e8a1122",
         15407 => x"70892b70",
         15408 => x"557c5457",
         15409 => x"5c59fd87",
         15410 => x"dc3fff15",
         15411 => x"7a067030",
         15412 => x"7072079f",
         15413 => x"2a84b8e4",
         15414 => x"0805901c",
         15415 => x"08794253",
         15416 => x"5f555881",
         15417 => x"78278838",
         15418 => x"9c190878",
         15419 => x"26833882",
         15420 => x"58777856",
         15421 => x"5b805974",
         15422 => x"527651fe",
         15423 => x"d8873f81",
         15424 => x"157f5555",
         15425 => x"9c140875",
         15426 => x"26833882",
         15427 => x"5584b8e4",
         15428 => x"08812e81",
         15429 => x"dc3884b8",
         15430 => x"e408ff2e",
         15431 => x"81d83884",
         15432 => x"b8e40881",
         15433 => x"c5388119",
         15434 => x"59787d2e",
         15435 => x"bb387478",
         15436 => x"2e098106",
         15437 => x"c2388756",
         15438 => x"75547384",
         15439 => x"b8e40c90",
         15440 => x"3d0d0487",
         15441 => x"0b84b8e4",
         15442 => x"0c903d0d",
         15443 => x"04811533",
         15444 => x"51fed0ac",
         15445 => x"3f84b8e4",
         15446 => x"08810654",
         15447 => x"73fead38",
         15448 => x"73770855",
         15449 => x"56fea739",
         15450 => x"7b802e81",
         15451 => x"8e387a7d",
         15452 => x"56587c80",
         15453 => x"2eab3881",
         15454 => x"18547481",
         15455 => x"2e80e638",
         15456 => x"73537752",
         15457 => x"7e51fedd",
         15458 => x"dd3f84b8",
         15459 => x"e4085684",
         15460 => x"b8e408ff",
         15461 => x"a3387781",
         15462 => x"19ff1757",
         15463 => x"595e74d7",
         15464 => x"387e7e90",
         15465 => x"120c557b",
         15466 => x"802eff8c",
         15467 => x"387a8818",
         15468 => x"0c798c18",
         15469 => x"0c901733",
         15470 => x"80c0075c",
         15471 => x"7b901834",
         15472 => x"9c1508fe",
         15473 => x"05941608",
         15474 => x"585a767a",
         15475 => x"26fee938",
         15476 => x"767d3194",
         15477 => x"160c8415",
         15478 => x"3381075d",
         15479 => x"7c841634",
         15480 => x"7554fed6",
         15481 => x"39ff54ff",
         15482 => x"9739745b",
         15483 => x"8059febe",
         15484 => x"398254fe",
         15485 => x"c5398154",
         15486 => x"fec039ff",
         15487 => x"1b5effa1",
         15488 => x"3984b8f0",
         15489 => x"08e33d0d",
         15490 => x"a33d08a5",
         15491 => x"3d080288",
         15492 => x"05818705",
         15493 => x"3344425f",
         15494 => x"ff0ba23d",
         15495 => x"08705f5b",
         15496 => x"4079802e",
         15497 => x"858a3879",
         15498 => x"7081055b",
         15499 => x"33709f26",
         15500 => x"565675ba",
         15501 => x"2e859b38",
         15502 => x"74ed3875",
         15503 => x"ba2e8592",
         15504 => x"3884d0c0",
         15505 => x"33568076",
         15506 => x"2484e538",
         15507 => x"75101084",
         15508 => x"d0ac0570",
         15509 => x"08565a74",
         15510 => x"802e8438",
         15511 => x"80753475",
         15512 => x"1684b8d8",
         15513 => x"113384b8",
         15514 => x"d9123340",
         15515 => x"5b5d8152",
         15516 => x"7951fece",
         15517 => x"a93f84b8",
         15518 => x"e40881ff",
         15519 => x"06708106",
         15520 => x"5d568357",
         15521 => x"7b84ab38",
         15522 => x"75822a81",
         15523 => x"06408a57",
         15524 => x"7f849f38",
         15525 => x"9f3dfc05",
         15526 => x"53835279",
         15527 => x"51fed0b0",
         15528 => x"3f84b8e4",
         15529 => x"08849838",
         15530 => x"6d557480",
         15531 => x"2e849038",
         15532 => x"74828080",
         15533 => x"26848838",
         15534 => x"ff157506",
         15535 => x"557483ff",
         15536 => x"387e802e",
         15537 => x"88388480",
         15538 => x"7f2683f8",
         15539 => x"387e8180",
         15540 => x"0a2683f0",
         15541 => x"38ff1f7f",
         15542 => x"06557483",
         15543 => x"e7387e89",
         15544 => x"2aa63d08",
         15545 => x"892a7089",
         15546 => x"2b77594c",
         15547 => x"475b6080",
         15548 => x"2e85ab38",
         15549 => x"65307080",
         15550 => x"25770756",
         15551 => x"5f915774",
         15552 => x"83b0387d",
         15553 => x"802e84df",
         15554 => x"38815474",
         15555 => x"53605279",
         15556 => x"51fecdbe",
         15557 => x"3f815784",
         15558 => x"b8e40883",
         15559 => x"95386083",
         15560 => x"ff053361",
         15561 => x"83fe0533",
         15562 => x"71882b07",
         15563 => x"59568e57",
         15564 => x"7782d4d5",
         15565 => x"2e098106",
         15566 => x"82f8387d",
         15567 => x"90296105",
         15568 => x"83b21133",
         15569 => x"44586280",
         15570 => x"2e82e738",
         15571 => x"83b61883",
         15572 => x"11338212",
         15573 => x"3371902b",
         15574 => x"71882b07",
         15575 => x"81143370",
         15576 => x"7207882b",
         15577 => x"75337107",
         15578 => x"83ba1f83",
         15579 => x"11338212",
         15580 => x"3371902b",
         15581 => x"71882b07",
         15582 => x"81143370",
         15583 => x"7207882b",
         15584 => x"75337107",
         15585 => x"5ca23d0c",
         15586 => x"42a33d0c",
         15587 => x"a33d0c44",
         15588 => x"4e544559",
         15589 => x"4f415a4b",
         15590 => x"784d8e57",
         15591 => x"80ff7927",
         15592 => x"82903893",
         15593 => x"577a8180",
         15594 => x"26828738",
         15595 => x"61812a70",
         15596 => x"81064549",
         15597 => x"63802e83",
         15598 => x"f9386187",
         15599 => x"06456482",
         15600 => x"2e893861",
         15601 => x"81064766",
         15602 => x"83f43883",
         15603 => x"6e70304a",
         15604 => x"46437a58",
         15605 => x"62832e8a",
         15606 => x"c2387aae",
         15607 => x"38788c2a",
         15608 => x"57810b83",
         15609 => x"e6882256",
         15610 => x"5874802e",
         15611 => x"9d387477",
         15612 => x"26983883",
         15613 => x"e6885677",
         15614 => x"10821770",
         15615 => x"22575758",
         15616 => x"74802e86",
         15617 => x"38767527",
         15618 => x"ee387752",
         15619 => x"7851fd81",
         15620 => x"943f84b8",
         15621 => x"e4081084",
         15622 => x"055584b8",
         15623 => x"e4089ff5",
         15624 => x"26963881",
         15625 => x"0b84b8e4",
         15626 => x"081084b8",
         15627 => x"e4080571",
         15628 => x"11722a83",
         15629 => x"05574c43",
         15630 => x"83ff1589",
         15631 => x"2a5d815c",
         15632 => x"a0477b1f",
         15633 => x"7d116805",
         15634 => x"6611ff05",
         15635 => x"706b0672",
         15636 => x"31584e57",
         15637 => x"4462832e",
         15638 => x"89b83874",
         15639 => x"1d5d7790",
         15640 => x"29167060",
         15641 => x"31565774",
         15642 => x"792682f2",
         15643 => x"38787c31",
         15644 => x"7d317853",
         15645 => x"70683152",
         15646 => x"56fd80a9",
         15647 => x"3f84b8e4",
         15648 => x"08406283",
         15649 => x"2e89f638",
         15650 => x"62822e09",
         15651 => x"810682dd",
         15652 => x"3883fff5",
         15653 => x"0b84b8e4",
         15654 => x"082782ac",
         15655 => x"387a89f9",
         15656 => x"38771855",
         15657 => x"7480c026",
         15658 => x"89ef3874",
         15659 => x"5bfea339",
         15660 => x"8b577684",
         15661 => x"b8e40c9f",
         15662 => x"3d0d84b8",
         15663 => x"f00c0481",
         15664 => x"4efbfe39",
         15665 => x"930b84b8",
         15666 => x"e40c9f3d",
         15667 => x"0d84b8f0",
         15668 => x"0c047c33",
         15669 => x"d0117081",
         15670 => x"ff065757",
         15671 => x"57748926",
         15672 => x"9138821d",
         15673 => x"7781ff06",
         15674 => x"d0055d58",
         15675 => x"777a2e81",
         15676 => x"b238800b",
         15677 => x"83e4d45f",
         15678 => x"5c7d087d",
         15679 => x"575b7a70",
         15680 => x"81055c33",
         15681 => x"76708105",
         15682 => x"5833ff9f",
         15683 => x"12455957",
         15684 => x"62992689",
         15685 => x"38e01770",
         15686 => x"81ff0658",
         15687 => x"44ff9f18",
         15688 => x"45649926",
         15689 => x"8938e018",
         15690 => x"7081ff06",
         15691 => x"59467630",
         15692 => x"709f2a5a",
         15693 => x"4776782e",
         15694 => x"09810685",
         15695 => x"3878ffbe",
         15696 => x"38757a32",
         15697 => x"70307072",
         15698 => x"079f2a7b",
         15699 => x"075d4a4a",
         15700 => x"7a802e80",
         15701 => x"ce38811c",
         15702 => x"841f5f5c",
         15703 => x"837c25ff",
         15704 => x"98387f56",
         15705 => x"f9e0399f",
         15706 => x"3df80553",
         15707 => x"81527951",
         15708 => x"fecadd3f",
         15709 => x"815784b8",
         15710 => x"e408feb6",
         15711 => x"3861832a",
         15712 => x"770684b8",
         15713 => x"e4084056",
         15714 => x"758338bf",
         15715 => x"5f6c558e",
         15716 => x"577e7526",
         15717 => x"fe9c3874",
         15718 => x"7f3159fb",
         15719 => x"fb398156",
         15720 => x"fad2397b",
         15721 => x"8324ffba",
         15722 => x"387b7aa3",
         15723 => x"3d0c56f9",
         15724 => x"95396181",
         15725 => x"06489357",
         15726 => x"67802efd",
         15727 => x"f538826e",
         15728 => x"70304a46",
         15729 => x"43fc8b39",
         15730 => x"84b8e408",
         15731 => x"9ff5269d",
         15732 => x"387a8b38",
         15733 => x"77185b81",
         15734 => x"807b27fb",
         15735 => x"f5388e57",
         15736 => x"7684b8e4",
         15737 => x"0c9f3d0d",
         15738 => x"84b8f00c",
         15739 => x"04805562",
         15740 => x"812e8699",
         15741 => x"389ff560",
         15742 => x"278b3874",
         15743 => x"81065b8e",
         15744 => x"577afdae",
         15745 => x"38848061",
         15746 => x"57558076",
         15747 => x"70810558",
         15748 => x"34ff1555",
         15749 => x"74f4388b",
         15750 => x"6183e4a0",
         15751 => x"59575576",
         15752 => x"70810558",
         15753 => x"33767081",
         15754 => x"055834ff",
         15755 => x"155574ef",
         15756 => x"38608b05",
         15757 => x"45746534",
         15758 => x"82618c05",
         15759 => x"3477618d",
         15760 => x"05347b83",
         15761 => x"ffff064b",
         15762 => x"6a618e05",
         15763 => x"346a882a",
         15764 => x"5c7b618f",
         15765 => x"05348161",
         15766 => x"90053462",
         15767 => x"83327030",
         15768 => x"5a488061",
         15769 => x"91053478",
         15770 => x"9e2a8206",
         15771 => x"49686192",
         15772 => x"05346c56",
         15773 => x"7583ffff",
         15774 => x"2686ad38",
         15775 => x"7583ffff",
         15776 => x"06557461",
         15777 => x"93053474",
         15778 => x"882a4c6b",
         15779 => x"61940534",
         15780 => x"f8619505",
         15781 => x"34bf6198",
         15782 => x"05348061",
         15783 => x"990534ff",
         15784 => x"619a0534",
         15785 => x"80619b05",
         15786 => x"347e619c",
         15787 => x"05347e88",
         15788 => x"2a486761",
         15789 => x"9d05347e",
         15790 => x"902a4c6b",
         15791 => x"619e0534",
         15792 => x"7e982a84",
         15793 => x"b8f00c84",
         15794 => x"b8f00861",
         15795 => x"9f053462",
         15796 => x"832e85f7",
         15797 => x"388061a7",
         15798 => x"05348061",
         15799 => x"a80534a1",
         15800 => x"61a90534",
         15801 => x"80cc61aa",
         15802 => x"05347c83",
         15803 => x"ffff0655",
         15804 => x"74619605",
         15805 => x"3474882a",
         15806 => x"4b6a6197",
         15807 => x"0534ff80",
         15808 => x"61a40534",
         15809 => x"a961a605",
         15810 => x"349361ab",
         15811 => x"0583e4ac",
         15812 => x"59575576",
         15813 => x"70810558",
         15814 => x"33767081",
         15815 => x"055834ff",
         15816 => x"155574ef",
         15817 => x"386083fe",
         15818 => x"054980d5",
         15819 => x"69346083",
         15820 => x"ff054bff",
         15821 => x"aa6b3481",
         15822 => x"547e5360",
         15823 => x"527951fe",
         15824 => x"c68f3f81",
         15825 => x"5784b8e4",
         15826 => x"08fae738",
         15827 => x"60175c62",
         15828 => x"832e879c",
         15829 => x"38696157",
         15830 => x"55807670",
         15831 => x"81055834",
         15832 => x"ff155574",
         15833 => x"f4386375",
         15834 => x"415b6283",
         15835 => x"2e86c038",
         15836 => x"87fffff8",
         15837 => x"5762812e",
         15838 => x"8338f857",
         15839 => x"76613476",
         15840 => x"882a7c45",
         15841 => x"55746470",
         15842 => x"81054634",
         15843 => x"76902a59",
         15844 => x"78647081",
         15845 => x"05463476",
         15846 => x"982a5675",
         15847 => x"64347c57",
         15848 => x"65597666",
         15849 => x"26833876",
         15850 => x"5978547a",
         15851 => x"53605279",
         15852 => x"51fec59d",
         15853 => x"3f84b8e4",
         15854 => x"0885e638",
         15855 => x"84806157",
         15856 => x"55807670",
         15857 => x"81055834",
         15858 => x"ff155574",
         15859 => x"f438781b",
         15860 => x"777a3158",
         15861 => x"5b76c938",
         15862 => x"7f810540",
         15863 => x"7f802eff",
         15864 => x"89387756",
         15865 => x"62832e83",
         15866 => x"38665665",
         15867 => x"55756626",
         15868 => x"83387555",
         15869 => x"74547a53",
         15870 => x"60527951",
         15871 => x"fec4d23f",
         15872 => x"84b8e408",
         15873 => x"859b3874",
         15874 => x"1b767631",
         15875 => x"575b75db",
         15876 => x"388c5862",
         15877 => x"832e9338",
         15878 => x"86586c83",
         15879 => x"ffff268a",
         15880 => x"38845862",
         15881 => x"822e8338",
         15882 => x"81587d84",
         15883 => x"c1386183",
         15884 => x"2a81065e",
         15885 => x"7d81b338",
         15886 => x"84806156",
         15887 => x"59807570",
         15888 => x"81055734",
         15889 => x"ff195978",
         15890 => x"f43880d5",
         15891 => x"6934ffaa",
         15892 => x"6b346083",
         15893 => x"be054778",
         15894 => x"67348167",
         15895 => x"81053481",
         15896 => x"67820534",
         15897 => x"78678305",
         15898 => x"34776784",
         15899 => x"05346c43",
         15900 => x"80fdc152",
         15901 => x"621f51fc",
         15902 => x"f8ab3ffe",
         15903 => x"67850534",
         15904 => x"84b8e408",
         15905 => x"822abf07",
         15906 => x"57766786",
         15907 => x"053484b8",
         15908 => x"e4086787",
         15909 => x"05347e61",
         15910 => x"83c60534",
         15911 => x"676183c7",
         15912 => x"05346b61",
         15913 => x"83c80534",
         15914 => x"84b8f008",
         15915 => x"6183c905",
         15916 => x"34626183",
         15917 => x"ca053462",
         15918 => x"882a4564",
         15919 => x"6183cb05",
         15920 => x"3462902a",
         15921 => x"58776183",
         15922 => x"cc053462",
         15923 => x"982a5f7e",
         15924 => x"6183cd05",
         15925 => x"34815478",
         15926 => x"53605279",
         15927 => x"51fec2f1",
         15928 => x"3f815784",
         15929 => x"b8e408f7",
         15930 => x"c9388053",
         15931 => x"80527951",
         15932 => x"fec3dd3f",
         15933 => x"815784b8",
         15934 => x"e408f7b6",
         15935 => x"3884b8e4",
         15936 => x"0884b8e4",
         15937 => x"0c9f3d0d",
         15938 => x"84b8f00c",
         15939 => x"046255f9",
         15940 => x"e439741c",
         15941 => x"6416455c",
         15942 => x"f6c4397a",
         15943 => x"ae387891",
         15944 => x"2a57810b",
         15945 => x"83e69822",
         15946 => x"56587480",
         15947 => x"2e9d3874",
         15948 => x"77269838",
         15949 => x"83e69856",
         15950 => x"77108217",
         15951 => x"70225757",
         15952 => x"5874802e",
         15953 => x"86387675",
         15954 => x"27ee3877",
         15955 => x"527851fc",
         15956 => x"f6d33f84",
         15957 => x"b8e40810",
         15958 => x"10848705",
         15959 => x"70892a5e",
         15960 => x"5ca05c80",
         15961 => x"0b84b8e4",
         15962 => x"08fc808a",
         15963 => x"055847fd",
         15964 => x"fff00a77",
         15965 => x"27f5cb38",
         15966 => x"8e57f8e4",
         15967 => x"3984b8e4",
         15968 => x"0883fff5",
         15969 => x"26f8e638",
         15970 => x"7af8d338",
         15971 => x"77812a5b",
         15972 => x"7af4bf38",
         15973 => x"8e57f8c8",
         15974 => x"39688106",
         15975 => x"4463802e",
         15976 => x"f8af3883",
         15977 => x"43f4ab39",
         15978 => x"7561a005",
         15979 => x"3475882a",
         15980 => x"496861a1",
         15981 => x"05347590",
         15982 => x"2a5b7a61",
         15983 => x"a2053475",
         15984 => x"982a5776",
         15985 => x"61a30534",
         15986 => x"f9c63980",
         15987 => x"6180c305",
         15988 => x"34806180",
         15989 => x"c40534a1",
         15990 => x"6180c505",
         15991 => x"3480cc61",
         15992 => x"80c60534",
         15993 => x"7c61a405",
         15994 => x"347c882a",
         15995 => x"5c7b61a5",
         15996 => x"05347c90",
         15997 => x"2a597861",
         15998 => x"a605347c",
         15999 => x"982a5675",
         16000 => x"61a70534",
         16001 => x"8261ac05",
         16002 => x"348061ad",
         16003 => x"05348061",
         16004 => x"ae053480",
         16005 => x"61af0534",
         16006 => x"8161b005",
         16007 => x"348061b1",
         16008 => x"05348661",
         16009 => x"b2053480",
         16010 => x"61b30534",
         16011 => x"ff806180",
         16012 => x"c00534a9",
         16013 => x"6180c205",
         16014 => x"34936180",
         16015 => x"c70583e4",
         16016 => x"c0595755",
         16017 => x"76708105",
         16018 => x"58337670",
         16019 => x"81055834",
         16020 => x"ff155574",
         16021 => x"802ef9cd",
         16022 => x"38767081",
         16023 => x"05583376",
         16024 => x"70810558",
         16025 => x"34ff1555",
         16026 => x"74da38f9",
         16027 => x"b8398154",
         16028 => x"80536052",
         16029 => x"7951febe",
         16030 => x"d93f8157",
         16031 => x"84b8e408",
         16032 => x"f4b0387d",
         16033 => x"90296105",
         16034 => x"42776283",
         16035 => x"b2053476",
         16036 => x"5484b8e4",
         16037 => x"08536052",
         16038 => x"7951febf",
         16039 => x"b43ffcc3",
         16040 => x"39810b84",
         16041 => x"b8e40c9f",
         16042 => x"3d0d84b8",
         16043 => x"f00c04f8",
         16044 => x"61347b4a",
         16045 => x"ff6a7081",
         16046 => x"054c34ff",
         16047 => x"6a708105",
         16048 => x"4c34ff6a",
         16049 => x"34ff6184",
         16050 => x"0534ff61",
         16051 => x"850534ff",
         16052 => x"61860534",
         16053 => x"ff618705",
         16054 => x"34ff6188",
         16055 => x"0534ff61",
         16056 => x"890534ff",
         16057 => x"618a0534",
         16058 => x"8f65347c",
         16059 => x"57f9b139",
         16060 => x"7654861f",
         16061 => x"53605279",
         16062 => x"51febed5",
         16063 => x"3f848061",
         16064 => x"56578075",
         16065 => x"70810557",
         16066 => x"34ff1757",
         16067 => x"76f43860",
         16068 => x"5c80d27c",
         16069 => x"7081055e",
         16070 => x"347b5580",
         16071 => x"d2757081",
         16072 => x"05573480",
         16073 => x"e1757081",
         16074 => x"05573480",
         16075 => x"c1753480",
         16076 => x"f26183e4",
         16077 => x"053480f2",
         16078 => x"6183e505",
         16079 => x"3480c161",
         16080 => x"83e60534",
         16081 => x"80e16183",
         16082 => x"e705347f",
         16083 => x"ff055b7a",
         16084 => x"6183e805",
         16085 => x"347a882a",
         16086 => x"59786183",
         16087 => x"e905347a",
         16088 => x"902a5675",
         16089 => x"6183ea05",
         16090 => x"347a982a",
         16091 => x"407f6183",
         16092 => x"eb053482",
         16093 => x"6183ec05",
         16094 => x"34766183",
         16095 => x"ed053476",
         16096 => x"6183ee05",
         16097 => x"34766183",
         16098 => x"ef053480",
         16099 => x"d56934ff",
         16100 => x"aa6b3481",
         16101 => x"54871f53",
         16102 => x"60527951",
         16103 => x"febdb23f",
         16104 => x"8154811f",
         16105 => x"53605279",
         16106 => x"51febda5",
         16107 => x"3f696157",
         16108 => x"55f7a639",
         16109 => x"f43d0d7e",
         16110 => x"615b5b80",
         16111 => x"7b61ff05",
         16112 => x"5a575776",
         16113 => x"7825b838",
         16114 => x"8d3d598e",
         16115 => x"3df80554",
         16116 => x"81537852",
         16117 => x"7951ff9a",
         16118 => x"b43f7b81",
         16119 => x"2e098106",
         16120 => x"9e388d3d",
         16121 => x"3355748d",
         16122 => x"2e903874",
         16123 => x"76708105",
         16124 => x"58348117",
         16125 => x"57748a2e",
         16126 => x"86387777",
         16127 => x"24cd3880",
         16128 => x"76347a55",
         16129 => x"76833876",
         16130 => x"557484b8",
         16131 => x"e40c8e3d",
         16132 => x"0d04f73d",
         16133 => x"0d7b0284",
         16134 => x"05b30533",
         16135 => x"5957778a",
         16136 => x"2e80d538",
         16137 => x"84170856",
         16138 => x"8076249e",
         16139 => x"38881708",
         16140 => x"77178c05",
         16141 => x"56597775",
         16142 => x"34811655",
         16143 => x"74bb248e",
         16144 => x"38748418",
         16145 => x"0c811988",
         16146 => x"180c8b3d",
         16147 => x"0d048b3d",
         16148 => x"fc055474",
         16149 => x"538c1752",
         16150 => x"760851ff",
         16151 => x"9ed13f74",
         16152 => x"7a327030",
         16153 => x"7072079f",
         16154 => x"2a703084",
         16155 => x"1b0c811c",
         16156 => x"881b0c5a",
         16157 => x"5656d339",
         16158 => x"8d527651",
         16159 => x"ff943fff",
         16160 => x"a339e33d",
         16161 => x"0d0280ff",
         16162 => x"05338d3d",
         16163 => x"585880cc",
         16164 => x"77575580",
         16165 => x"76708105",
         16166 => x"5834ff15",
         16167 => x"5574f438",
         16168 => x"a13d0877",
         16169 => x"0c778a2e",
         16170 => x"80f7387c",
         16171 => x"56807624",
         16172 => x"80c0387d",
         16173 => x"77178c05",
         16174 => x"56597775",
         16175 => x"34811655",
         16176 => x"74bb24b8",
         16177 => x"38748418",
         16178 => x"0c811988",
         16179 => x"180c7c55",
         16180 => x"8075249e",
         16181 => x"389f3dff",
         16182 => x"ac115575",
         16183 => x"54c00552",
         16184 => x"760851ff",
         16185 => x"9dc93f84",
         16186 => x"b8e40886",
         16187 => x"387c7a2e",
         16188 => x"ba38ff0b",
         16189 => x"84b8e40c",
         16190 => x"9f3d0d04",
         16191 => x"9f3dffb0",
         16192 => x"11557554",
         16193 => x"c0055276",
         16194 => x"0851ff9d",
         16195 => x"a23f747b",
         16196 => x"32703070",
         16197 => x"72079f2a",
         16198 => x"7030525a",
         16199 => x"5656ffa5",
         16200 => x"398d5276",
         16201 => x"51fdeb3f",
         16202 => x"ff81397d",
         16203 => x"84b8e40c",
         16204 => x"9f3d0d04",
         16205 => x"fd3d0d75",
         16206 => x"0284059a",
         16207 => x"05225253",
         16208 => x"80527280",
         16209 => x"ff269038",
         16210 => x"7283ffff",
         16211 => x"06527184",
         16212 => x"b8e40c85",
         16213 => x"3d0d0483",
         16214 => x"ffff7327",
         16215 => x"547083b5",
         16216 => x"2e098106",
         16217 => x"e9387380",
         16218 => x"2ee43883",
         16219 => x"e6a82251",
         16220 => x"72712e9c",
         16221 => x"38811270",
         16222 => x"83ffff06",
         16223 => x"53547180",
         16224 => x"ff268d38",
         16225 => x"711083e6",
         16226 => x"a8057022",
         16227 => x"5151e139",
         16228 => x"81801270",
         16229 => x"81ff0684",
         16230 => x"b8e40c53",
         16231 => x"853d0d04",
         16232 => x"fe3d0d02",
         16233 => x"92052202",
         16234 => x"84059605",
         16235 => x"22535180",
         16236 => x"537080ff",
         16237 => x"268c3870",
         16238 => x"537284b8",
         16239 => x"e40c843d",
         16240 => x"0d047183",
         16241 => x"b52e0981",
         16242 => x"06ef3870",
         16243 => x"81ff26e9",
         16244 => x"38701083",
         16245 => x"e4a80570",
         16246 => x"2284b8e4",
         16247 => x"0c51843d",
         16248 => x"0d04fb3d",
         16249 => x"0d775170",
         16250 => x"83ffff26",
         16251 => x"80e13870",
         16252 => x"83ffff06",
         16253 => x"83e8a856",
         16254 => x"56759fff",
         16255 => x"2680d938",
         16256 => x"74708205",
         16257 => x"56227571",
         16258 => x"30708025",
         16259 => x"737a2607",
         16260 => x"54565353",
         16261 => x"70b73871",
         16262 => x"70820553",
         16263 => x"22727188",
         16264 => x"2a545681",
         16265 => x"ff067014",
         16266 => x"52547076",
         16267 => x"24b13871",
         16268 => x"cf387310",
         16269 => x"15707082",
         16270 => x"05522254",
         16271 => x"73307080",
         16272 => x"25757926",
         16273 => x"07535552",
         16274 => x"70802ecb",
         16275 => x"38755170",
         16276 => x"84b8e40c",
         16277 => x"873d0d04",
         16278 => x"83ec9c55",
         16279 => x"ffa23971",
         16280 => x"8826ea38",
         16281 => x"71101083",
         16282 => x"c9d00554",
         16283 => x"730804c7",
         16284 => x"a0167083",
         16285 => x"ffff0657",
         16286 => x"517551d3",
         16287 => x"39ffb016",
         16288 => x"7083ffff",
         16289 => x"065751f1",
         16290 => x"39881670",
         16291 => x"83ffff06",
         16292 => x"5751e639",
         16293 => x"e6167083",
         16294 => x"ffff0657",
         16295 => x"51db39d0",
         16296 => x"167083ff",
         16297 => x"ff065751",
         16298 => x"d039e016",
         16299 => x"7083ffff",
         16300 => x"065751c5",
         16301 => x"39f01670",
         16302 => x"83ffff06",
         16303 => x"5751ffb9",
         16304 => x"39757331",
         16305 => x"81067671",
         16306 => x"317083ff",
         16307 => x"ff065852",
         16308 => x"55ffa639",
         16309 => x"75733110",
         16310 => x"75057022",
         16311 => x"5252feef",
         16312 => x"39000000",
         16313 => x"00ffffff",
         16314 => x"ff00ffff",
         16315 => x"ffff00ff",
         16316 => x"ffffff00",
         16317 => x"0000198b",
         16318 => x"00001980",
         16319 => x"00001975",
         16320 => x"0000196a",
         16321 => x"0000195f",
         16322 => x"00001954",
         16323 => x"00001949",
         16324 => x"0000193e",
         16325 => x"00001933",
         16326 => x"00001928",
         16327 => x"0000191d",
         16328 => x"00001912",
         16329 => x"00001907",
         16330 => x"000018fc",
         16331 => x"000018f1",
         16332 => x"000018e6",
         16333 => x"000018db",
         16334 => x"000018d0",
         16335 => x"000018c5",
         16336 => x"000018ba",
         16337 => x"00001ebf",
         16338 => x"00001f59",
         16339 => x"00001f59",
         16340 => x"00001f59",
         16341 => x"00001f59",
         16342 => x"00001f59",
         16343 => x"00001f59",
         16344 => x"00001f59",
         16345 => x"00001f59",
         16346 => x"00001f59",
         16347 => x"00001f59",
         16348 => x"00001f59",
         16349 => x"00001f59",
         16350 => x"00001f59",
         16351 => x"00001f59",
         16352 => x"00001f59",
         16353 => x"00001f59",
         16354 => x"00001f59",
         16355 => x"00001f59",
         16356 => x"00001f59",
         16357 => x"00001f59",
         16358 => x"00001f59",
         16359 => x"00001f59",
         16360 => x"00001f59",
         16361 => x"00001f59",
         16362 => x"00001f59",
         16363 => x"00001f59",
         16364 => x"00001f59",
         16365 => x"00001f59",
         16366 => x"00001f59",
         16367 => x"00001f59",
         16368 => x"00001f59",
         16369 => x"00001f59",
         16370 => x"00001f59",
         16371 => x"00001f59",
         16372 => x"00001f59",
         16373 => x"00001f59",
         16374 => x"00001f59",
         16375 => x"00001f59",
         16376 => x"00001f59",
         16377 => x"00001f59",
         16378 => x"00001f59",
         16379 => x"00001f59",
         16380 => x"00002471",
         16381 => x"00001f59",
         16382 => x"00001f59",
         16383 => x"00001f59",
         16384 => x"00001f59",
         16385 => x"00001f59",
         16386 => x"00001f59",
         16387 => x"00001f59",
         16388 => x"00001f59",
         16389 => x"00001f59",
         16390 => x"00001f59",
         16391 => x"00001f59",
         16392 => x"00001f59",
         16393 => x"00001f59",
         16394 => x"00001f59",
         16395 => x"00001f59",
         16396 => x"00001f59",
         16397 => x"00002407",
         16398 => x"00002306",
         16399 => x"00001f59",
         16400 => x"0000228a",
         16401 => x"000024a8",
         16402 => x"00002367",
         16403 => x"0000222c",
         16404 => x"000021ce",
         16405 => x"00001f59",
         16406 => x"00001f59",
         16407 => x"00001f59",
         16408 => x"00001f59",
         16409 => x"00001f59",
         16410 => x"00001f59",
         16411 => x"00001f59",
         16412 => x"00001f59",
         16413 => x"00001f59",
         16414 => x"00001f59",
         16415 => x"00001f59",
         16416 => x"00001f59",
         16417 => x"00001f59",
         16418 => x"00001f59",
         16419 => x"00001f59",
         16420 => x"00001f59",
         16421 => x"00001f59",
         16422 => x"00001f59",
         16423 => x"00001f59",
         16424 => x"00001f59",
         16425 => x"00001f59",
         16426 => x"00001f59",
         16427 => x"00001f59",
         16428 => x"00001f59",
         16429 => x"00001f59",
         16430 => x"00001f59",
         16431 => x"00001f59",
         16432 => x"00001f59",
         16433 => x"00001f59",
         16434 => x"00001f59",
         16435 => x"00001f59",
         16436 => x"00001f59",
         16437 => x"00001f59",
         16438 => x"00001f59",
         16439 => x"00001f59",
         16440 => x"00001f59",
         16441 => x"00001f59",
         16442 => x"00001f59",
         16443 => x"00001f59",
         16444 => x"00001f59",
         16445 => x"00001f59",
         16446 => x"00001f59",
         16447 => x"00001f59",
         16448 => x"00001f59",
         16449 => x"00001f59",
         16450 => x"00001f59",
         16451 => x"00001f59",
         16452 => x"00001f59",
         16453 => x"00001f59",
         16454 => x"00001f59",
         16455 => x"00001f59",
         16456 => x"00001f59",
         16457 => x"000021ab",
         16458 => x"00002170",
         16459 => x"00001f59",
         16460 => x"00001f59",
         16461 => x"00001f59",
         16462 => x"00001f59",
         16463 => x"00001f59",
         16464 => x"00001f59",
         16465 => x"00001f59",
         16466 => x"00001f59",
         16467 => x"00002163",
         16468 => x"00002158",
         16469 => x"00001f59",
         16470 => x"00002141",
         16471 => x"00001f59",
         16472 => x"00002151",
         16473 => x"00002147",
         16474 => x"0000213a",
         16475 => x"00003212",
         16476 => x"0000322a",
         16477 => x"00003236",
         16478 => x"00003242",
         16479 => x"0000324e",
         16480 => x"0000321e",
         16481 => x"00003b86",
         16482 => x"00003a74",
         16483 => x"000038f0",
         16484 => x"0000363e",
         16485 => x"00003a10",
         16486 => x"000034cd",
         16487 => x"0000378a",
         16488 => x"00003663",
         16489 => x"000039ba",
         16490 => x"00003692",
         16491 => x"00003701",
         16492 => x"00003919",
         16493 => x"000034cd",
         16494 => x"000038f0",
         16495 => x"000037fa",
         16496 => x"0000378a",
         16497 => x"000034cd",
         16498 => x"000034cd",
         16499 => x"00003701",
         16500 => x"00003692",
         16501 => x"00003663",
         16502 => x"0000363e",
         16503 => x"0000466b",
         16504 => x"00004684",
         16505 => x"000046a9",
         16506 => x"000046ca",
         16507 => x"0000462b",
         16508 => x"000046ef",
         16509 => x"00004644",
         16510 => x"00004794",
         16511 => x"00004751",
         16512 => x"00004751",
         16513 => x"00004751",
         16514 => x"00004751",
         16515 => x"00004751",
         16516 => x"00004751",
         16517 => x"0000472a",
         16518 => x"00004751",
         16519 => x"00004751",
         16520 => x"00004751",
         16521 => x"00004751",
         16522 => x"00004751",
         16523 => x"00004751",
         16524 => x"00004751",
         16525 => x"00004751",
         16526 => x"00004751",
         16527 => x"00004751",
         16528 => x"00004751",
         16529 => x"00004751",
         16530 => x"00004751",
         16531 => x"00004751",
         16532 => x"00004751",
         16533 => x"00004751",
         16534 => x"00004751",
         16535 => x"00004751",
         16536 => x"00004751",
         16537 => x"00004751",
         16538 => x"00004751",
         16539 => x"00004751",
         16540 => x"00004869",
         16541 => x"00004857",
         16542 => x"00004844",
         16543 => x"00004831",
         16544 => x"0000475b",
         16545 => x"0000481f",
         16546 => x"0000480c",
         16547 => x"00004774",
         16548 => x"00004751",
         16549 => x"00004774",
         16550 => x"000047fc",
         16551 => x"00004879",
         16552 => x"000047a5",
         16553 => x"00004783",
         16554 => x"000047ea",
         16555 => x"000047d8",
         16556 => x"000047c6",
         16557 => x"000047b7",
         16558 => x"00004751",
         16559 => x"0000475b",
         16560 => x"000053f7",
         16561 => x"00005566",
         16562 => x"00005538",
         16563 => x"0000548f",
         16564 => x"0000546c",
         16565 => x"0000544b",
         16566 => x"00005421",
         16567 => x"000055f1",
         16568 => x"00005278",
         16569 => x"000055cb",
         16570 => x"000057ba",
         16571 => x"00005278",
         16572 => x"00005278",
         16573 => x"00005278",
         16574 => x"00005278",
         16575 => x"00005278",
         16576 => x"00005278",
         16577 => x"00005594",
         16578 => x"000057a2",
         16579 => x"00005659",
         16580 => x"00005278",
         16581 => x"00005278",
         16582 => x"00005278",
         16583 => x"00005278",
         16584 => x"00005278",
         16585 => x"00005278",
         16586 => x"00005278",
         16587 => x"00005278",
         16588 => x"00005278",
         16589 => x"00005278",
         16590 => x"00005278",
         16591 => x"00005278",
         16592 => x"00005278",
         16593 => x"00005278",
         16594 => x"00005278",
         16595 => x"00005278",
         16596 => x"00005278",
         16597 => x"00005278",
         16598 => x"00005278",
         16599 => x"00005516",
         16600 => x"00005278",
         16601 => x"00005278",
         16602 => x"00005278",
         16603 => x"000054b9",
         16604 => x"000053c8",
         16605 => x"0000536a",
         16606 => x"00005278",
         16607 => x"00005278",
         16608 => x"00005278",
         16609 => x"00005278",
         16610 => x"0000534f",
         16611 => x"00005278",
         16612 => x"00005332",
         16613 => x"0000599b",
         16614 => x"00005910",
         16615 => x"00005910",
         16616 => x"00005910",
         16617 => x"00005910",
         16618 => x"00005910",
         16619 => x"00005910",
         16620 => x"000058eb",
         16621 => x"00005910",
         16622 => x"00005910",
         16623 => x"00005910",
         16624 => x"00005910",
         16625 => x"00005910",
         16626 => x"00005910",
         16627 => x"00005910",
         16628 => x"00005910",
         16629 => x"00005910",
         16630 => x"00005910",
         16631 => x"00005910",
         16632 => x"00005910",
         16633 => x"00005910",
         16634 => x"00005910",
         16635 => x"00005910",
         16636 => x"00005910",
         16637 => x"00005910",
         16638 => x"00005910",
         16639 => x"00005910",
         16640 => x"00005910",
         16641 => x"00005910",
         16642 => x"00005910",
         16643 => x"000059ad",
         16644 => x"000059f5",
         16645 => x"000059e2",
         16646 => x"000059cf",
         16647 => x"000059bd",
         16648 => x"00005a80",
         16649 => x"00005a6d",
         16650 => x"00005a5d",
         16651 => x"00005910",
         16652 => x"00005a4d",
         16653 => x"00005a3d",
         16654 => x"00005a2b",
         16655 => x"00005a19",
         16656 => x"00005a07",
         16657 => x"00005978",
         16658 => x"00005967",
         16659 => x"00005956",
         16660 => x"0000593f",
         16661 => x"00005910",
         16662 => x"00005989",
         16663 => x"0000636a",
         16664 => x"000061c6",
         16665 => x"000061c6",
         16666 => x"000061c6",
         16667 => x"000061c6",
         16668 => x"000061c6",
         16669 => x"000061c6",
         16670 => x"000061c6",
         16671 => x"000061c6",
         16672 => x"000061c6",
         16673 => x"000061c6",
         16674 => x"000061c6",
         16675 => x"000061c6",
         16676 => x"000061c6",
         16677 => x"00005ee8",
         16678 => x"000061c6",
         16679 => x"000061c6",
         16680 => x"000061c6",
         16681 => x"000061c6",
         16682 => x"000061c6",
         16683 => x"000061c6",
         16684 => x"000063b4",
         16685 => x"000061c6",
         16686 => x"000061c6",
         16687 => x"0000633f",
         16688 => x"000061c6",
         16689 => x"00006356",
         16690 => x"00005ec7",
         16691 => x"00006328",
         16692 => x"0000ded4",
         16693 => x"0000dec1",
         16694 => x"0000deb5",
         16695 => x"0000deaa",
         16696 => x"0000de9f",
         16697 => x"0000de94",
         16698 => x"0000de89",
         16699 => x"0000de7d",
         16700 => x"0000de6f",
         16701 => x"00000e01",
         16702 => x"00000bfd",
         16703 => x"00000bfd",
         16704 => x"00000f49",
         16705 => x"00000bfd",
         16706 => x"00000bfd",
         16707 => x"00000bfd",
         16708 => x"00000bfd",
         16709 => x"00000bfd",
         16710 => x"00000bfd",
         16711 => x"00000bfd",
         16712 => x"00000dfd",
         16713 => x"00000bfd",
         16714 => x"00000f7f",
         16715 => x"00000f0d",
         16716 => x"00000bfd",
         16717 => x"00000bfd",
         16718 => x"00000bfd",
         16719 => x"00000bfd",
         16720 => x"00000bfd",
         16721 => x"00000bfd",
         16722 => x"00000bfd",
         16723 => x"00000bfd",
         16724 => x"00000bfd",
         16725 => x"00000bfd",
         16726 => x"00000bfd",
         16727 => x"00000bfd",
         16728 => x"00000bfd",
         16729 => x"00000bfd",
         16730 => x"00000bfd",
         16731 => x"00000bfd",
         16732 => x"00000bfd",
         16733 => x"00000bfd",
         16734 => x"00000bfd",
         16735 => x"00000bfd",
         16736 => x"00000bfd",
         16737 => x"00000bfd",
         16738 => x"00000bfd",
         16739 => x"00000bfd",
         16740 => x"00000bfd",
         16741 => x"00000bfd",
         16742 => x"00000bfd",
         16743 => x"00000bfd",
         16744 => x"00000bfd",
         16745 => x"00000bfd",
         16746 => x"00000bfd",
         16747 => x"00000bfd",
         16748 => x"00000bfd",
         16749 => x"00000bfd",
         16750 => x"00000bfd",
         16751 => x"00000bfd",
         16752 => x"00000f1d",
         16753 => x"00000bfd",
         16754 => x"00000bfd",
         16755 => x"00000bfd",
         16756 => x"00000bfd",
         16757 => x"00000e17",
         16758 => x"00000bfd",
         16759 => x"00000bfd",
         16760 => x"00000bfd",
         16761 => x"00000bfd",
         16762 => x"00000bfd",
         16763 => x"00000bfd",
         16764 => x"00000bfd",
         16765 => x"00000bfd",
         16766 => x"00000bfd",
         16767 => x"00000bfd",
         16768 => x"00000e2b",
         16769 => x"00000ee1",
         16770 => x"00000eb8",
         16771 => x"00000eb8",
         16772 => x"00000eb8",
         16773 => x"00000bfd",
         16774 => x"00000ee1",
         16775 => x"00000bfd",
         16776 => x"00000bfd",
         16777 => x"00000eff",
         16778 => x"00000bfd",
         16779 => x"00000bfd",
         16780 => x"00000c16",
         16781 => x"00000e0f",
         16782 => x"00000bfd",
         16783 => x"00000bfd",
         16784 => x"00000f58",
         16785 => x"00000bfd",
         16786 => x"00000c18",
         16787 => x"00000bfd",
         16788 => x"00000bfd",
         16789 => x"00000e17",
         16790 => x"64696e69",
         16791 => x"74000000",
         16792 => x"64696f63",
         16793 => x"746c0000",
         16794 => x"66696e69",
         16795 => x"74000000",
         16796 => x"666c6f61",
         16797 => x"64000000",
         16798 => x"66657865",
         16799 => x"63000000",
         16800 => x"6d636c65",
         16801 => x"61720000",
         16802 => x"6d636f70",
         16803 => x"79000000",
         16804 => x"6d646966",
         16805 => x"66000000",
         16806 => x"6d64756d",
         16807 => x"70000000",
         16808 => x"6d656200",
         16809 => x"6d656800",
         16810 => x"6d657700",
         16811 => x"68696400",
         16812 => x"68696500",
         16813 => x"68666400",
         16814 => x"68666500",
         16815 => x"63616c6c",
         16816 => x"00000000",
         16817 => x"6a6d7000",
         16818 => x"72657374",
         16819 => x"61727400",
         16820 => x"72657365",
         16821 => x"74000000",
         16822 => x"696e666f",
         16823 => x"00000000",
         16824 => x"74657374",
         16825 => x"00000000",
         16826 => x"636c7300",
         16827 => x"7a383000",
         16828 => x"74626173",
         16829 => x"69630000",
         16830 => x"6d626173",
         16831 => x"69630000",
         16832 => x"6b696c6f",
         16833 => x"00000000",
         16834 => x"65640000",
         16835 => x"556e6b6e",
         16836 => x"6f776e20",
         16837 => x"6572726f",
         16838 => x"722e0000",
         16839 => x"50617261",
         16840 => x"6d657465",
         16841 => x"72732069",
         16842 => x"6e636f72",
         16843 => x"72656374",
         16844 => x"2e000000",
         16845 => x"546f6f20",
         16846 => x"6d616e79",
         16847 => x"206f7065",
         16848 => x"6e206669",
         16849 => x"6c65732e",
         16850 => x"00000000",
         16851 => x"496e7375",
         16852 => x"66666963",
         16853 => x"69656e74",
         16854 => x"206d656d",
         16855 => x"6f72792e",
         16856 => x"00000000",
         16857 => x"46696c65",
         16858 => x"20697320",
         16859 => x"6c6f636b",
         16860 => x"65642e00",
         16861 => x"54696d65",
         16862 => x"6f75742c",
         16863 => x"206f7065",
         16864 => x"72617469",
         16865 => x"6f6e2063",
         16866 => x"616e6365",
         16867 => x"6c6c6564",
         16868 => x"2e000000",
         16869 => x"466f726d",
         16870 => x"61742061",
         16871 => x"626f7274",
         16872 => x"65642e00",
         16873 => x"4e6f2063",
         16874 => x"6f6d7061",
         16875 => x"7469626c",
         16876 => x"65206669",
         16877 => x"6c657379",
         16878 => x"7374656d",
         16879 => x"20666f75",
         16880 => x"6e64206f",
         16881 => x"6e206469",
         16882 => x"736b2e00",
         16883 => x"4469736b",
         16884 => x"206e6f74",
         16885 => x"20656e61",
         16886 => x"626c6564",
         16887 => x"2e000000",
         16888 => x"44726976",
         16889 => x"65206e75",
         16890 => x"6d626572",
         16891 => x"20697320",
         16892 => x"696e7661",
         16893 => x"6c69642e",
         16894 => x"00000000",
         16895 => x"53442069",
         16896 => x"73207772",
         16897 => x"69746520",
         16898 => x"70726f74",
         16899 => x"65637465",
         16900 => x"642e0000",
         16901 => x"46696c65",
         16902 => x"2068616e",
         16903 => x"646c6520",
         16904 => x"696e7661",
         16905 => x"6c69642e",
         16906 => x"00000000",
         16907 => x"46696c65",
         16908 => x"20616c72",
         16909 => x"65616479",
         16910 => x"20657869",
         16911 => x"7374732e",
         16912 => x"00000000",
         16913 => x"41636365",
         16914 => x"73732064",
         16915 => x"656e6965",
         16916 => x"642e0000",
         16917 => x"496e7661",
         16918 => x"6c696420",
         16919 => x"66696c65",
         16920 => x"6e616d65",
         16921 => x"2e000000",
         16922 => x"4e6f2070",
         16923 => x"61746820",
         16924 => x"666f756e",
         16925 => x"642e0000",
         16926 => x"4e6f2066",
         16927 => x"696c6520",
         16928 => x"666f756e",
         16929 => x"642e0000",
         16930 => x"4469736b",
         16931 => x"206e6f74",
         16932 => x"20726561",
         16933 => x"64792e00",
         16934 => x"496e7465",
         16935 => x"726e616c",
         16936 => x"20657272",
         16937 => x"6f722e00",
         16938 => x"4469736b",
         16939 => x"20457272",
         16940 => x"6f720000",
         16941 => x"53756363",
         16942 => x"6573732e",
         16943 => x"00000000",
         16944 => x"0a256c75",
         16945 => x"20627974",
         16946 => x"65732025",
         16947 => x"73206174",
         16948 => x"20256c75",
         16949 => x"20627974",
         16950 => x"65732f73",
         16951 => x"65632e0a",
         16952 => x"00000000",
         16953 => x"72656164",
         16954 => x"00000000",
         16955 => x"2530386c",
         16956 => x"58000000",
         16957 => x"3a202000",
         16958 => x"25303258",
         16959 => x"00000000",
         16960 => x"207c0000",
         16961 => x"7c000000",
         16962 => x"20200000",
         16963 => x"25303458",
         16964 => x"00000000",
         16965 => x"20202020",
         16966 => x"20202020",
         16967 => x"00000000",
         16968 => x"7a4f5300",
         16969 => x"2a2a2025",
         16970 => x"73202800",
         16971 => x"31312f30",
         16972 => x"332f3230",
         16973 => x"32310000",
         16974 => x"76312e31",
         16975 => x"6b000000",
         16976 => x"205a5055",
         16977 => x"2c207265",
         16978 => x"76202530",
         16979 => x"32782920",
         16980 => x"25732025",
         16981 => x"73202a2a",
         16982 => x"0a0a0000",
         16983 => x"5a505520",
         16984 => x"496e7465",
         16985 => x"72727570",
         16986 => x"74204861",
         16987 => x"6e646c65",
         16988 => x"72000000",
         16989 => x"55415254",
         16990 => x"31205458",
         16991 => x"20696e74",
         16992 => x"65727275",
         16993 => x"70740000",
         16994 => x"55415254",
         16995 => x"31205258",
         16996 => x"20696e74",
         16997 => x"65727275",
         16998 => x"70740000",
         16999 => x"55415254",
         17000 => x"30205458",
         17001 => x"20696e74",
         17002 => x"65727275",
         17003 => x"70740000",
         17004 => x"55415254",
         17005 => x"30205258",
         17006 => x"20696e74",
         17007 => x"65727275",
         17008 => x"70740000",
         17009 => x"494f4354",
         17010 => x"4c205752",
         17011 => x"20696e74",
         17012 => x"65727275",
         17013 => x"70740000",
         17014 => x"494f4354",
         17015 => x"4c205244",
         17016 => x"20696e74",
         17017 => x"65727275",
         17018 => x"70740000",
         17019 => x"50533220",
         17020 => x"696e7465",
         17021 => x"72727570",
         17022 => x"74000000",
         17023 => x"54696d65",
         17024 => x"7220696e",
         17025 => x"74657272",
         17026 => x"75707400",
         17027 => x"53657474",
         17028 => x"696e6720",
         17029 => x"75702074",
         17030 => x"696d6572",
         17031 => x"2e2e2e00",
         17032 => x"456e6162",
         17033 => x"6c696e67",
         17034 => x"2074696d",
         17035 => x"65722e2e",
         17036 => x"2e000000",
         17037 => x"6175746f",
         17038 => x"65786563",
         17039 => x"2e626174",
         17040 => x"00000000",
         17041 => x"7a4f535f",
         17042 => x"7a70752e",
         17043 => x"68737400",
         17044 => x"4661696c",
         17045 => x"65642074",
         17046 => x"6f20696e",
         17047 => x"69746961",
         17048 => x"6c697365",
         17049 => x"20736420",
         17050 => x"63617264",
         17051 => x"20302c20",
         17052 => x"706c6561",
         17053 => x"73652069",
         17054 => x"6e697420",
         17055 => x"6d616e75",
         17056 => x"616c6c79",
         17057 => x"2e000000",
         17058 => x"2a200000",
         17059 => x"25643a5c",
         17060 => x"25730000",
         17061 => x"303a0000",
         17062 => x"42616420",
         17063 => x"636f6d6d",
         17064 => x"616e642e",
         17065 => x"00000000",
         17066 => x"5a505500",
         17067 => x"62696e00",
         17068 => x"25643a5c",
         17069 => x"25735c25",
         17070 => x"732e2573",
         17071 => x"00000000",
         17072 => x"436f6c64",
         17073 => x"20726562",
         17074 => x"6f6f7469",
         17075 => x"6e672e2e",
         17076 => x"2e000000",
         17077 => x"52657374",
         17078 => x"61727469",
         17079 => x"6e672061",
         17080 => x"70706c69",
         17081 => x"63617469",
         17082 => x"6f6e2e2e",
         17083 => x"2e000000",
         17084 => x"43616c6c",
         17085 => x"696e6720",
         17086 => x"636f6465",
         17087 => x"20402025",
         17088 => x"30386c78",
         17089 => x"202e2e2e",
         17090 => x"0a000000",
         17091 => x"43616c6c",
         17092 => x"20726574",
         17093 => x"75726e65",
         17094 => x"6420636f",
         17095 => x"64652028",
         17096 => x"2564292e",
         17097 => x"0a000000",
         17098 => x"45786563",
         17099 => x"7574696e",
         17100 => x"6720636f",
         17101 => x"64652040",
         17102 => x"20253038",
         17103 => x"6c78202e",
         17104 => x"2e2e0a00",
         17105 => x"2530386c",
         17106 => x"58202530",
         17107 => x"386c582d",
         17108 => x"00000000",
         17109 => x"2530386c",
         17110 => x"58202530",
         17111 => x"34582d00",
         17112 => x"436f6d70",
         17113 => x"6172696e",
         17114 => x"672e2e2e",
         17115 => x"00000000",
         17116 => x"2530386c",
         17117 => x"78282530",
         17118 => x"3878292d",
         17119 => x"3e253038",
         17120 => x"6c782825",
         17121 => x"30387829",
         17122 => x"0a000000",
         17123 => x"436f7079",
         17124 => x"696e672e",
         17125 => x"2e2e0000",
         17126 => x"2530386c",
         17127 => x"58202530",
         17128 => x"32582d00",
         17129 => x"436c6561",
         17130 => x"72696e67",
         17131 => x"2e2e2e2e",
         17132 => x"00000000",
         17133 => x"44756d70",
         17134 => x"204d656d",
         17135 => x"6f727900",
         17136 => x"0a436f6d",
         17137 => x"706c6574",
         17138 => x"652e0000",
         17139 => x"25643a5c",
         17140 => x"25735c25",
         17141 => x"73000000",
         17142 => x"4d656d6f",
         17143 => x"72792065",
         17144 => x"78686175",
         17145 => x"73746564",
         17146 => x"2c206361",
         17147 => x"6e6e6f74",
         17148 => x"2070726f",
         17149 => x"63657373",
         17150 => x"20636f6d",
         17151 => x"6d616e64",
         17152 => x"2e000000",
         17153 => x"3f3f3f00",
         17154 => x"25642f25",
         17155 => x"642f2564",
         17156 => x"2025643a",
         17157 => x"25643a25",
         17158 => x"642e2564",
         17159 => x"25640a00",
         17160 => x"536f4320",
         17161 => x"436f6e66",
         17162 => x"69677572",
         17163 => x"6174696f",
         17164 => x"6e000000",
         17165 => x"3a0a4465",
         17166 => x"76696365",
         17167 => x"7320696d",
         17168 => x"706c656d",
         17169 => x"656e7465",
         17170 => x"643a0000",
         17171 => x"41646472",
         17172 => x"65737365",
         17173 => x"733a0000",
         17174 => x"20202020",
         17175 => x"43505520",
         17176 => x"52657365",
         17177 => x"74205665",
         17178 => x"63746f72",
         17179 => x"20416464",
         17180 => x"72657373",
         17181 => x"203d2025",
         17182 => x"3038580a",
         17183 => x"00000000",
         17184 => x"20202020",
         17185 => x"43505520",
         17186 => x"4d656d6f",
         17187 => x"72792053",
         17188 => x"74617274",
         17189 => x"20416464",
         17190 => x"72657373",
         17191 => x"203d2025",
         17192 => x"3038580a",
         17193 => x"00000000",
         17194 => x"20202020",
         17195 => x"53746163",
         17196 => x"6b205374",
         17197 => x"61727420",
         17198 => x"41646472",
         17199 => x"65737320",
         17200 => x"20202020",
         17201 => x"203d2025",
         17202 => x"3038580a",
         17203 => x"00000000",
         17204 => x"4d697363",
         17205 => x"3a000000",
         17206 => x"20202020",
         17207 => x"5a505520",
         17208 => x"49642020",
         17209 => x"20202020",
         17210 => x"20202020",
         17211 => x"20202020",
         17212 => x"20202020",
         17213 => x"203d2025",
         17214 => x"3034580a",
         17215 => x"00000000",
         17216 => x"20202020",
         17217 => x"53797374",
         17218 => x"656d2043",
         17219 => x"6c6f636b",
         17220 => x"20467265",
         17221 => x"71202020",
         17222 => x"20202020",
         17223 => x"203d2025",
         17224 => x"642e2530",
         17225 => x"34644d48",
         17226 => x"7a0a0000",
         17227 => x"20202020",
         17228 => x"57697368",
         17229 => x"626f6e65",
         17230 => x"20534452",
         17231 => x"414d2043",
         17232 => x"6c6f636b",
         17233 => x"20467265",
         17234 => x"713d2025",
         17235 => x"642e2530",
         17236 => x"34644d48",
         17237 => x"7a0a0000",
         17238 => x"20202020",
         17239 => x"53445241",
         17240 => x"4d20436c",
         17241 => x"6f636b20",
         17242 => x"46726571",
         17243 => x"20202020",
         17244 => x"20202020",
         17245 => x"203d2025",
         17246 => x"642e2530",
         17247 => x"34644d48",
         17248 => x"7a0a0000",
         17249 => x"20202020",
         17250 => x"53504900",
         17251 => x"20202020",
         17252 => x"50533200",
         17253 => x"20202020",
         17254 => x"494f4354",
         17255 => x"4c000000",
         17256 => x"20202020",
         17257 => x"57422049",
         17258 => x"32430000",
         17259 => x"20202020",
         17260 => x"57495348",
         17261 => x"424f4e45",
         17262 => x"20425553",
         17263 => x"00000000",
         17264 => x"20202020",
         17265 => x"494e5452",
         17266 => x"20435452",
         17267 => x"4c202843",
         17268 => x"68616e6e",
         17269 => x"656c733d",
         17270 => x"25303264",
         17271 => x"292e0a00",
         17272 => x"20202020",
         17273 => x"54494d45",
         17274 => x"52312020",
         17275 => x"20202854",
         17276 => x"696d6572",
         17277 => x"7320203d",
         17278 => x"25303264",
         17279 => x"292e0a00",
         17280 => x"20202020",
         17281 => x"53442043",
         17282 => x"41524420",
         17283 => x"20202844",
         17284 => x"65766963",
         17285 => x"6573203d",
         17286 => x"25303264",
         17287 => x"292e0a00",
         17288 => x"20202020",
         17289 => x"52414d20",
         17290 => x"20202020",
         17291 => x"20202825",
         17292 => x"3038583a",
         17293 => x"25303858",
         17294 => x"292e0a00",
         17295 => x"20202020",
         17296 => x"4252414d",
         17297 => x"20202020",
         17298 => x"20202825",
         17299 => x"3038583a",
         17300 => x"25303858",
         17301 => x"292e0a00",
         17302 => x"20202020",
         17303 => x"494e534e",
         17304 => x"20425241",
         17305 => x"4d202825",
         17306 => x"3038583a",
         17307 => x"25303858",
         17308 => x"292e0a00",
         17309 => x"20202020",
         17310 => x"53445241",
         17311 => x"4d202020",
         17312 => x"20202825",
         17313 => x"3038583a",
         17314 => x"25303858",
         17315 => x"292e0a00",
         17316 => x"20202020",
         17317 => x"57422053",
         17318 => x"4452414d",
         17319 => x"20202825",
         17320 => x"3038583a",
         17321 => x"25303858",
         17322 => x"292e0a00",
         17323 => x"20286672",
         17324 => x"6f6d2053",
         17325 => x"6f432063",
         17326 => x"6f6e6669",
         17327 => x"67290000",
         17328 => x"556e6b6e",
         17329 => x"6f776e00",
         17330 => x"45564f6d",
         17331 => x"00000000",
         17332 => x"536d616c",
         17333 => x"6c000000",
         17334 => x"4d656469",
         17335 => x"756d0000",
         17336 => x"466c6578",
         17337 => x"00000000",
         17338 => x"45564f00",
         17339 => x"0000f048",
         17340 => x"01000000",
         17341 => x"00000002",
         17342 => x"0000f044",
         17343 => x"01000000",
         17344 => x"00000003",
         17345 => x"0000f040",
         17346 => x"01000000",
         17347 => x"00000004",
         17348 => x"0000f03c",
         17349 => x"01000000",
         17350 => x"00000005",
         17351 => x"0000f038",
         17352 => x"01000000",
         17353 => x"00000006",
         17354 => x"0000f034",
         17355 => x"01000000",
         17356 => x"00000007",
         17357 => x"0000f030",
         17358 => x"01000000",
         17359 => x"00000001",
         17360 => x"0000f02c",
         17361 => x"01000000",
         17362 => x"00000008",
         17363 => x"0000f028",
         17364 => x"01000000",
         17365 => x"0000000b",
         17366 => x"0000f024",
         17367 => x"01000000",
         17368 => x"00000009",
         17369 => x"0000f020",
         17370 => x"01000000",
         17371 => x"0000000a",
         17372 => x"0000f01c",
         17373 => x"04000000",
         17374 => x"0000000d",
         17375 => x"0000f018",
         17376 => x"04000000",
         17377 => x"0000000c",
         17378 => x"0000f014",
         17379 => x"04000000",
         17380 => x"0000000e",
         17381 => x"0000f010",
         17382 => x"03000000",
         17383 => x"0000000f",
         17384 => x"0000f00c",
         17385 => x"04000000",
         17386 => x"0000000f",
         17387 => x"0000f008",
         17388 => x"04000000",
         17389 => x"00000010",
         17390 => x"0000f004",
         17391 => x"04000000",
         17392 => x"00000011",
         17393 => x"0000f000",
         17394 => x"03000000",
         17395 => x"00000012",
         17396 => x"0000effc",
         17397 => x"03000000",
         17398 => x"00000013",
         17399 => x"0000eff8",
         17400 => x"03000000",
         17401 => x"00000014",
         17402 => x"0000eff4",
         17403 => x"03000000",
         17404 => x"00000015",
         17405 => x"1b5b4400",
         17406 => x"1b5b4300",
         17407 => x"1b5b4200",
         17408 => x"1b5b4100",
         17409 => x"1b5b367e",
         17410 => x"1b5b357e",
         17411 => x"1b5b347e",
         17412 => x"1b304600",
         17413 => x"1b5b337e",
         17414 => x"1b5b327e",
         17415 => x"1b5b317e",
         17416 => x"10000000",
         17417 => x"0e000000",
         17418 => x"0d000000",
         17419 => x"0b000000",
         17420 => x"08000000",
         17421 => x"06000000",
         17422 => x"05000000",
         17423 => x"04000000",
         17424 => x"03000000",
         17425 => x"02000000",
         17426 => x"01000000",
         17427 => x"43616e6e",
         17428 => x"6f74206f",
         17429 => x"70656e2f",
         17430 => x"63726561",
         17431 => x"74652068",
         17432 => x"6973746f",
         17433 => x"72792066",
         17434 => x"696c652c",
         17435 => x"20646973",
         17436 => x"61626c69",
         17437 => x"6e672e00",
         17438 => x"68697374",
         17439 => x"6f727900",
         17440 => x"68697374",
         17441 => x"00000000",
         17442 => x"21000000",
         17443 => x"2530366c",
         17444 => x"75202025",
         17445 => x"730a0000",
         17446 => x"4661696c",
         17447 => x"65642074",
         17448 => x"6f207265",
         17449 => x"73657420",
         17450 => x"74686520",
         17451 => x"68697374",
         17452 => x"6f727920",
         17453 => x"66696c65",
         17454 => x"20746f20",
         17455 => x"454f462e",
         17456 => x"00000000",
         17457 => x"3e25730a",
         17458 => x"00000000",
         17459 => x"1b5b317e",
         17460 => x"00000000",
         17461 => x"1b5b4100",
         17462 => x"1b5b4200",
         17463 => x"1b5b4300",
         17464 => x"1b5b4400",
         17465 => x"1b5b3130",
         17466 => x"7e000000",
         17467 => x"1b5b3131",
         17468 => x"7e000000",
         17469 => x"1b5b3132",
         17470 => x"7e000000",
         17471 => x"1b5b3133",
         17472 => x"7e000000",
         17473 => x"1b5b3134",
         17474 => x"7e000000",
         17475 => x"1b5b3135",
         17476 => x"7e000000",
         17477 => x"1b5b3137",
         17478 => x"7e000000",
         17479 => x"1b5b3138",
         17480 => x"7e000000",
         17481 => x"1b5b3139",
         17482 => x"7e000000",
         17483 => x"1b5b3230",
         17484 => x"7e000000",
         17485 => x"1b5b327e",
         17486 => x"00000000",
         17487 => x"1b5b337e",
         17488 => x"00000000",
         17489 => x"1b5b4600",
         17490 => x"1b5b357e",
         17491 => x"00000000",
         17492 => x"1b5b367e",
         17493 => x"00000000",
         17494 => x"583a2564",
         17495 => x"2c25642c",
         17496 => x"25642c25",
         17497 => x"642c2564",
         17498 => x"2c25643a",
         17499 => x"25303278",
         17500 => x"00000000",
         17501 => x"443a2564",
         17502 => x"2d25642d",
         17503 => x"25643a25",
         17504 => x"633a2564",
         17505 => x"2c25642c",
         17506 => x"25643a00",
         17507 => x"25642c00",
         17508 => x"4b3a2564",
         17509 => x"3a000000",
         17510 => x"25303278",
         17511 => x"2c000000",
         17512 => x"25635b25",
         17513 => x"643b2564",
         17514 => x"52000000",
         17515 => x"5265706f",
         17516 => x"72742043",
         17517 => x"7572736f",
         17518 => x"723a0000",
         17519 => x"55703a25",
         17520 => x"30327820",
         17521 => x"25303278",
         17522 => x"00000000",
         17523 => x"44773a25",
         17524 => x"30327820",
         17525 => x"25303278",
         17526 => x"00000000",
         17527 => x"48643a25",
         17528 => x"30327820",
         17529 => x"00000000",
         17530 => x"4e6f2074",
         17531 => x"65737420",
         17532 => x"64656669",
         17533 => x"6e65642e",
         17534 => x"00000000",
         17535 => x"53440000",
         17536 => x"222a3a3c",
         17537 => x"3e3f7c7f",
         17538 => x"00000000",
         17539 => x"2b2c3b3d",
         17540 => x"5b5d0000",
         17541 => x"46415400",
         17542 => x"46415433",
         17543 => x"32000000",
         17544 => x"ebfe904d",
         17545 => x"53444f53",
         17546 => x"352e3000",
         17547 => x"4e4f204e",
         17548 => x"414d4520",
         17549 => x"20202046",
         17550 => x"41542020",
         17551 => x"20202000",
         17552 => x"4e4f204e",
         17553 => x"414d4520",
         17554 => x"20202046",
         17555 => x"41543332",
         17556 => x"20202000",
         17557 => x"0000f1fc",
         17558 => x"00000000",
         17559 => x"00000000",
         17560 => x"00000000",
         17561 => x"01030507",
         17562 => x"090e1012",
         17563 => x"1416181c",
         17564 => x"1e000000",
         17565 => x"809a4541",
         17566 => x"8e418f80",
         17567 => x"45454549",
         17568 => x"49498e8f",
         17569 => x"9092924f",
         17570 => x"994f5555",
         17571 => x"59999a9b",
         17572 => x"9c9d9e9f",
         17573 => x"41494f55",
         17574 => x"a5a5a6a7",
         17575 => x"a8a9aaab",
         17576 => x"acadaeaf",
         17577 => x"b0b1b2b3",
         17578 => x"b4b5b6b7",
         17579 => x"b8b9babb",
         17580 => x"bcbdbebf",
         17581 => x"c0c1c2c3",
         17582 => x"c4c5c6c7",
         17583 => x"c8c9cacb",
         17584 => x"cccdcecf",
         17585 => x"d0d1d2d3",
         17586 => x"d4d5d6d7",
         17587 => x"d8d9dadb",
         17588 => x"dcdddedf",
         17589 => x"e0e1e2e3",
         17590 => x"e4e5e6e7",
         17591 => x"e8e9eaeb",
         17592 => x"ecedeeef",
         17593 => x"f0f1f2f3",
         17594 => x"f4f5f6f7",
         17595 => x"f8f9fafb",
         17596 => x"fcfdfeff",
         17597 => x"2b2e2c3b",
         17598 => x"3d5b5d2f",
         17599 => x"5c222a3a",
         17600 => x"3c3e3f7c",
         17601 => x"7f000000",
         17602 => x"00010004",
         17603 => x"00100040",
         17604 => x"01000200",
         17605 => x"00000000",
         17606 => x"00010002",
         17607 => x"00040008",
         17608 => x"00100020",
         17609 => x"00000000",
         17610 => x"00c700fc",
         17611 => x"00e900e2",
         17612 => x"00e400e0",
         17613 => x"00e500e7",
         17614 => x"00ea00eb",
         17615 => x"00e800ef",
         17616 => x"00ee00ec",
         17617 => x"00c400c5",
         17618 => x"00c900e6",
         17619 => x"00c600f4",
         17620 => x"00f600f2",
         17621 => x"00fb00f9",
         17622 => x"00ff00d6",
         17623 => x"00dc00a2",
         17624 => x"00a300a5",
         17625 => x"20a70192",
         17626 => x"00e100ed",
         17627 => x"00f300fa",
         17628 => x"00f100d1",
         17629 => x"00aa00ba",
         17630 => x"00bf2310",
         17631 => x"00ac00bd",
         17632 => x"00bc00a1",
         17633 => x"00ab00bb",
         17634 => x"25912592",
         17635 => x"25932502",
         17636 => x"25242561",
         17637 => x"25622556",
         17638 => x"25552563",
         17639 => x"25512557",
         17640 => x"255d255c",
         17641 => x"255b2510",
         17642 => x"25142534",
         17643 => x"252c251c",
         17644 => x"2500253c",
         17645 => x"255e255f",
         17646 => x"255a2554",
         17647 => x"25692566",
         17648 => x"25602550",
         17649 => x"256c2567",
         17650 => x"25682564",
         17651 => x"25652559",
         17652 => x"25582552",
         17653 => x"2553256b",
         17654 => x"256a2518",
         17655 => x"250c2588",
         17656 => x"2584258c",
         17657 => x"25902580",
         17658 => x"03b100df",
         17659 => x"039303c0",
         17660 => x"03a303c3",
         17661 => x"00b503c4",
         17662 => x"03a60398",
         17663 => x"03a903b4",
         17664 => x"221e03c6",
         17665 => x"03b52229",
         17666 => x"226100b1",
         17667 => x"22652264",
         17668 => x"23202321",
         17669 => x"00f72248",
         17670 => x"00b02219",
         17671 => x"00b7221a",
         17672 => x"207f00b2",
         17673 => x"25a000a0",
         17674 => x"0061031a",
         17675 => x"00e00317",
         17676 => x"00f80307",
         17677 => x"00ff0001",
         17678 => x"01780100",
         17679 => x"01300132",
         17680 => x"01060139",
         17681 => x"0110014a",
         17682 => x"012e0179",
         17683 => x"01060180",
         17684 => x"004d0243",
         17685 => x"01810182",
         17686 => x"01820184",
         17687 => x"01840186",
         17688 => x"01870187",
         17689 => x"0189018a",
         17690 => x"018b018b",
         17691 => x"018d018e",
         17692 => x"018f0190",
         17693 => x"01910191",
         17694 => x"01930194",
         17695 => x"01f60196",
         17696 => x"01970198",
         17697 => x"0198023d",
         17698 => x"019b019c",
         17699 => x"019d0220",
         17700 => x"019f01a0",
         17701 => x"01a001a2",
         17702 => x"01a201a4",
         17703 => x"01a401a6",
         17704 => x"01a701a7",
         17705 => x"01a901aa",
         17706 => x"01ab01ac",
         17707 => x"01ac01ae",
         17708 => x"01af01af",
         17709 => x"01b101b2",
         17710 => x"01b301b3",
         17711 => x"01b501b5",
         17712 => x"01b701b8",
         17713 => x"01b801ba",
         17714 => x"01bb01bc",
         17715 => x"01bc01be",
         17716 => x"01f701c0",
         17717 => x"01c101c2",
         17718 => x"01c301c4",
         17719 => x"01c501c4",
         17720 => x"01c701c8",
         17721 => x"01c701ca",
         17722 => x"01cb01ca",
         17723 => x"01cd0110",
         17724 => x"01dd0001",
         17725 => x"018e01de",
         17726 => x"011201f3",
         17727 => x"000301f1",
         17728 => x"01f401f4",
         17729 => x"01f80128",
         17730 => x"02220112",
         17731 => x"023a0009",
         17732 => x"2c65023b",
         17733 => x"023b023d",
         17734 => x"2c66023f",
         17735 => x"02400241",
         17736 => x"02410246",
         17737 => x"010a0253",
         17738 => x"00400181",
         17739 => x"01860255",
         17740 => x"0189018a",
         17741 => x"0258018f",
         17742 => x"025a0190",
         17743 => x"025c025d",
         17744 => x"025e025f",
         17745 => x"01930261",
         17746 => x"02620194",
         17747 => x"02640265",
         17748 => x"02660267",
         17749 => x"01970196",
         17750 => x"026a2c62",
         17751 => x"026c026d",
         17752 => x"026e019c",
         17753 => x"02700271",
         17754 => x"019d0273",
         17755 => x"0274019f",
         17756 => x"02760277",
         17757 => x"02780279",
         17758 => x"027a027b",
         17759 => x"027c2c64",
         17760 => x"027e027f",
         17761 => x"01a60281",
         17762 => x"028201a9",
         17763 => x"02840285",
         17764 => x"02860287",
         17765 => x"01ae0244",
         17766 => x"01b101b2",
         17767 => x"0245028d",
         17768 => x"028e028f",
         17769 => x"02900291",
         17770 => x"01b7037b",
         17771 => x"000303fd",
         17772 => x"03fe03ff",
         17773 => x"03ac0004",
         17774 => x"03860388",
         17775 => x"0389038a",
         17776 => x"03b10311",
         17777 => x"03c20002",
         17778 => x"03a303a3",
         17779 => x"03c40308",
         17780 => x"03cc0003",
         17781 => x"038c038e",
         17782 => x"038f03d8",
         17783 => x"011803f2",
         17784 => x"000a03f9",
         17785 => x"03f303f4",
         17786 => x"03f503f6",
         17787 => x"03f703f7",
         17788 => x"03f903fa",
         17789 => x"03fa0430",
         17790 => x"03200450",
         17791 => x"07100460",
         17792 => x"0122048a",
         17793 => x"013604c1",
         17794 => x"010e04cf",
         17795 => x"000104c0",
         17796 => x"04d00144",
         17797 => x"05610426",
         17798 => x"00000000",
         17799 => x"1d7d0001",
         17800 => x"2c631e00",
         17801 => x"01961ea0",
         17802 => x"015a1f00",
         17803 => x"06081f10",
         17804 => x"06061f20",
         17805 => x"06081f30",
         17806 => x"06081f40",
         17807 => x"06061f51",
         17808 => x"00071f59",
         17809 => x"1f521f5b",
         17810 => x"1f541f5d",
         17811 => x"1f561f5f",
         17812 => x"1f600608",
         17813 => x"1f70000e",
         17814 => x"1fba1fbb",
         17815 => x"1fc81fc9",
         17816 => x"1fca1fcb",
         17817 => x"1fda1fdb",
         17818 => x"1ff81ff9",
         17819 => x"1fea1feb",
         17820 => x"1ffa1ffb",
         17821 => x"1f800608",
         17822 => x"1f900608",
         17823 => x"1fa00608",
         17824 => x"1fb00004",
         17825 => x"1fb81fb9",
         17826 => x"1fb21fbc",
         17827 => x"1fcc0001",
         17828 => x"1fc31fd0",
         17829 => x"06021fe0",
         17830 => x"06021fe5",
         17831 => x"00011fec",
         17832 => x"1ff30001",
         17833 => x"1ffc214e",
         17834 => x"00012132",
         17835 => x"21700210",
         17836 => x"21840001",
         17837 => x"218324d0",
         17838 => x"051a2c30",
         17839 => x"042f2c60",
         17840 => x"01022c67",
         17841 => x"01062c75",
         17842 => x"01022c80",
         17843 => x"01642d00",
         17844 => x"0826ff41",
         17845 => x"031a0000",
         17846 => x"00000000",
         17847 => x"0000e658",
         17848 => x"01020100",
         17849 => x"00000000",
         17850 => x"00000000",
         17851 => x"0000e660",
         17852 => x"01040100",
         17853 => x"00000000",
         17854 => x"00000000",
         17855 => x"0000e668",
         17856 => x"01140300",
         17857 => x"00000000",
         17858 => x"00000000",
         17859 => x"0000e670",
         17860 => x"012b0300",
         17861 => x"00000000",
         17862 => x"00000000",
         17863 => x"0000e678",
         17864 => x"01300300",
         17865 => x"00000000",
         17866 => x"00000000",
         17867 => x"0000e680",
         17868 => x"013c0400",
         17869 => x"00000000",
         17870 => x"00000000",
         17871 => x"0000e688",
         17872 => x"013d0400",
         17873 => x"00000000",
         17874 => x"00000000",
         17875 => x"0000e690",
         17876 => x"013f0400",
         17877 => x"00000000",
         17878 => x"00000000",
         17879 => x"0000e698",
         17880 => x"01400400",
         17881 => x"00000000",
         17882 => x"00000000",
         17883 => x"0000e6a0",
         17884 => x"01410400",
         17885 => x"00000000",
         17886 => x"00000000",
         17887 => x"0000e6a4",
         17888 => x"01420400",
         17889 => x"00000000",
         17890 => x"00000000",
         17891 => x"0000e6a8",
         17892 => x"01430400",
         17893 => x"00000000",
         17894 => x"00000000",
         17895 => x"0000e6ac",
         17896 => x"01500500",
         17897 => x"00000000",
         17898 => x"00000000",
         17899 => x"0000e6b0",
         17900 => x"01510500",
         17901 => x"00000000",
         17902 => x"00000000",
         17903 => x"0000e6b4",
         17904 => x"01540500",
         17905 => x"00000000",
         17906 => x"00000000",
         17907 => x"0000e6b8",
         17908 => x"01550500",
         17909 => x"00000000",
         17910 => x"00000000",
         17911 => x"0000e6bc",
         17912 => x"01790700",
         17913 => x"00000000",
         17914 => x"00000000",
         17915 => x"0000e6c4",
         17916 => x"01780700",
         17917 => x"00000000",
         17918 => x"00000000",
         17919 => x"0000e6c8",
         17920 => x"01820800",
         17921 => x"00000000",
         17922 => x"00000000",
         17923 => x"0000e6d0",
         17924 => x"01830800",
         17925 => x"00000000",
         17926 => x"00000000",
         17927 => x"0000e6d8",
         17928 => x"01850800",
         17929 => x"00000000",
         17930 => x"00000000",
         17931 => x"0000e6e0",
         17932 => x"01870800",
         17933 => x"00000000",
         17934 => x"00000000",
         17935 => x"0000e6e8",
         17936 => x"01880800",
         17937 => x"00000000",
         17938 => x"00000000",
         17939 => x"0000e6ec",
         17940 => x"01890800",
         17941 => x"00000000",
         17942 => x"00000000",
         17943 => x"0000e6f0",
         17944 => x"018c0900",
         17945 => x"00000000",
         17946 => x"00000000",
         17947 => x"0000e6f8",
         17948 => x"018d0900",
         17949 => x"00000000",
         17950 => x"00000000",
         17951 => x"0000e700",
         17952 => x"018e0900",
         17953 => x"00000000",
         17954 => x"00000000",
         17955 => x"0000e708",
         17956 => x"018f0900",
         17957 => x"00000000",
         17958 => x"00000000",
         17959 => x"00000000",
         17960 => x"00000000",
         17961 => x"00007fff",
         17962 => x"00000000",
         17963 => x"00007fff",
         17964 => x"00010000",
         17965 => x"00007fff",
         17966 => x"00010000",
         17967 => x"00810000",
         17968 => x"01000000",
         17969 => x"017fffff",
         17970 => x"00000000",
         17971 => x"00000000",
         17972 => x"00007800",
         17973 => x"00000000",
         17974 => x"05f5e100",
         17975 => x"05f5e100",
         17976 => x"05f5e100",
         17977 => x"00000000",
         17978 => x"01010101",
         17979 => x"01010101",
         17980 => x"01011001",
         17981 => x"01000000",
         17982 => x"00000000",
         17983 => x"00000000",
         17984 => x"00000000",
         17985 => x"00000000",
         17986 => x"00000000",
         17987 => x"00000000",
         17988 => x"00000000",
         17989 => x"00000000",
         17990 => x"00000000",
         17991 => x"00000000",
         17992 => x"00000000",
         17993 => x"00000000",
         17994 => x"00000000",
         17995 => x"00000000",
         17996 => x"00000000",
         17997 => x"00000000",
         17998 => x"00000000",
         17999 => x"00000000",
         18000 => x"00000000",
         18001 => x"00000000",
         18002 => x"00000000",
         18003 => x"00000000",
         18004 => x"00000000",
         18005 => x"00000000",
         18006 => x"0000f078",
         18007 => x"01000000",
         18008 => x"0000f080",
         18009 => x"01000000",
         18010 => x"0000f088",
         18011 => x"02000000",
         18012 => x"0001fd80",
         18013 => x"1bfc5ffd",
         18014 => x"f03b3a0d",
         18015 => x"797a405b",
         18016 => x"5df0f0f0",
         18017 => x"71727374",
         18018 => x"75767778",
         18019 => x"696a6b6c",
         18020 => x"6d6e6f70",
         18021 => x"61626364",
         18022 => x"65666768",
         18023 => x"31323334",
         18024 => x"35363738",
         18025 => x"5cf32d20",
         18026 => x"30392c2e",
         18027 => x"f67ff3f4",
         18028 => x"f1f23f2f",
         18029 => x"08f0f0f0",
         18030 => x"f0f0f0f0",
         18031 => x"80818283",
         18032 => x"84f0f0f0",
         18033 => x"1bfc58fd",
         18034 => x"f03a3b0d",
         18035 => x"595a405b",
         18036 => x"5df0f0f0",
         18037 => x"51525354",
         18038 => x"55565758",
         18039 => x"494a4b4c",
         18040 => x"4d4e4f50",
         18041 => x"41424344",
         18042 => x"45464748",
         18043 => x"31323334",
         18044 => x"35363738",
         18045 => x"5cf32d20",
         18046 => x"30392c2e",
         18047 => x"f67ff3f4",
         18048 => x"f1f23f2f",
         18049 => x"08f0f0f0",
         18050 => x"f0f0f0f0",
         18051 => x"80818283",
         18052 => x"84f0f0f0",
         18053 => x"1bfc58fd",
         18054 => x"f02b2a0d",
         18055 => x"595a607b",
         18056 => x"7df0f0f0",
         18057 => x"51525354",
         18058 => x"55565758",
         18059 => x"494a4b4c",
         18060 => x"4d4e4f50",
         18061 => x"41424344",
         18062 => x"45464748",
         18063 => x"21222324",
         18064 => x"25262728",
         18065 => x"7c7e3d20",
         18066 => x"20293c3e",
         18067 => x"f7e2e0e1",
         18068 => x"f9f83f2f",
         18069 => x"fbf0f0f0",
         18070 => x"f0f0f0f0",
         18071 => x"85868788",
         18072 => x"89f0f0f0",
         18073 => x"1bfe1efa",
         18074 => x"f0f0f0f0",
         18075 => x"191a001b",
         18076 => x"1df0f0f0",
         18077 => x"11121314",
         18078 => x"15161718",
         18079 => x"090a0b0c",
         18080 => x"0d0e0f10",
         18081 => x"01020304",
         18082 => x"05060708",
         18083 => x"f0f0f0f0",
         18084 => x"f0f0f0f0",
         18085 => x"f01ef0f0",
         18086 => x"f01ff0f0",
         18087 => x"f0f0f0f0",
         18088 => x"f0f0f01c",
         18089 => x"f0f0f0f0",
         18090 => x"f0f0f0f0",
         18091 => x"80818283",
         18092 => x"84f0f0f0",
         18093 => x"bff0cfc9",
         18094 => x"f0b54dcd",
         18095 => x"3577d7b3",
         18096 => x"b7f0f0f0",
         18097 => x"7c704131",
         18098 => x"39a678dd",
         18099 => x"3d5d6c56",
         18100 => x"1d33d5b1",
         18101 => x"466ed948",
         18102 => x"74434c73",
         18103 => x"3f367e3b",
         18104 => x"7a1e5fa2",
         18105 => x"d39fd100",
         18106 => x"9da3d0b9",
         18107 => x"c6c5c2c1",
         18108 => x"c3c4bbbe",
         18109 => x"f0f0f0f0",
         18110 => x"f0f0f0f0",
         18111 => x"80818283",
         18112 => x"84f0f0f0",
         18113 => x"00000000",
         18114 => x"00000000",
         18115 => x"00000000",
         18116 => x"00000000",
         18117 => x"00000000",
         18118 => x"00000000",
         18119 => x"00000000",
         18120 => x"00000000",
         18121 => x"00000000",
         18122 => x"00000000",
         18123 => x"00000000",
         18124 => x"00000000",
         18125 => x"00000000",
         18126 => x"00000000",
         18127 => x"00000000",
         18128 => x"00000000",
         18129 => x"00000000",
         18130 => x"00000000",
         18131 => x"00000000",
         18132 => x"00000000",
         18133 => x"00000000",
         18134 => x"00000000",
         18135 => x"00000000",
         18136 => x"00000000",
         18137 => x"00000000",
         18138 => x"00010000",
         18139 => x"00000000",
         18140 => x"f8000000",
         18141 => x"0000f0cc",
         18142 => x"f3000000",
         18143 => x"0000f0d4",
         18144 => x"f4000000",
         18145 => x"0000f0d8",
         18146 => x"f1000000",
         18147 => x"0000f0dc",
         18148 => x"f2000000",
         18149 => x"0000f0e0",
         18150 => x"80000000",
         18151 => x"0000f0e4",
         18152 => x"81000000",
         18153 => x"0000f0ec",
         18154 => x"82000000",
         18155 => x"0000f0f4",
         18156 => x"83000000",
         18157 => x"0000f0fc",
         18158 => x"84000000",
         18159 => x"0000f104",
         18160 => x"85000000",
         18161 => x"0000f10c",
         18162 => x"86000000",
         18163 => x"0000f114",
         18164 => x"87000000",
         18165 => x"0000f11c",
         18166 => x"88000000",
         18167 => x"0000f124",
         18168 => x"89000000",
         18169 => x"0000f12c",
         18170 => x"f6000000",
         18171 => x"0000f134",
         18172 => x"7f000000",
         18173 => x"0000f13c",
         18174 => x"f9000000",
         18175 => x"0000f144",
         18176 => x"e0000000",
         18177 => x"0000f148",
         18178 => x"e1000000",
         18179 => x"0000f150",
         18180 => x"71000000",
         18181 => x"00000000",
         18182 => x"00000000",
         18183 => x"00000000",
         18184 => x"00000000",
         18185 => x"00000000",
         18186 => x"00000000",
         18187 => x"00000000",
         18188 => x"00000000",
         18189 => x"00000000",
         18190 => x"00000000",
         18191 => x"00000000",
         18192 => x"00000000",
         18193 => x"00000000",
         18194 => x"00000000",
         18195 => x"00000000",
         18196 => x"00000000",
         18197 => x"00000000",
         18198 => x"00000000",
         18199 => x"00000000",
         18200 => x"00000000",
         18201 => x"00000000",
         18202 => x"00000000",
         18203 => x"00000000",
         18204 => x"00000000",
         18205 => x"00000000",
         18206 => x"00000000",
         18207 => x"00000000",
         18208 => x"00000000",
         18209 => x"00000000",
         18210 => x"00000000",
         18211 => x"00000000",
         18212 => x"00000000",
         18213 => x"00000000",
         18214 => x"00000000",
         18215 => x"00000000",
         18216 => x"00000000",
         18217 => x"00000000",
         18218 => x"00000000",
         18219 => x"00000000",
         18220 => x"00000000",
         18221 => x"00000000",
         18222 => x"00000000",
         18223 => x"00000000",
         18224 => x"00000000",
         18225 => x"00000000",
         18226 => x"00000000",
         18227 => x"00000000",
         18228 => x"00000000",
         18229 => x"00000000",
         18230 => x"00000000",
         18231 => x"00000000",
         18232 => x"00000000",
         18233 => x"00000000",
         18234 => x"00000000",
         18235 => x"00000000",
         18236 => x"00000000",
         18237 => x"00000000",
         18238 => x"00000000",
         18239 => x"00000000",
         18240 => x"00000000",
         18241 => x"00000000",
         18242 => x"00000000",
         18243 => x"00000000",
         18244 => x"00000000",
         18245 => x"00000000",
         18246 => x"00000000",
         18247 => x"00000000",
         18248 => x"00000000",
         18249 => x"00000000",
         18250 => x"00000000",
         18251 => x"00000000",
         18252 => x"00000000",
         18253 => x"00000000",
         18254 => x"00000000",
         18255 => x"00000000",
         18256 => x"00000000",
         18257 => x"00000000",
         18258 => x"00000000",
         18259 => x"00000000",
         18260 => x"00000000",
         18261 => x"00000000",
         18262 => x"00000000",
         18263 => x"00000000",
         18264 => x"00000000",
         18265 => x"00000000",
         18266 => x"00000000",
         18267 => x"00000000",
         18268 => x"00000000",
         18269 => x"00000000",
         18270 => x"00000000",
         18271 => x"00000000",
         18272 => x"00000000",
         18273 => x"00000000",
         18274 => x"00000000",
         18275 => x"00000000",
         18276 => x"00000000",
         18277 => x"00000000",
         18278 => x"00000000",
         18279 => x"00000000",
         18280 => x"00000000",
         18281 => x"00000000",
         18282 => x"00000000",
         18283 => x"00000000",
         18284 => x"00000000",
         18285 => x"00000000",
         18286 => x"00000000",
         18287 => x"00000000",
         18288 => x"00000000",
         18289 => x"00000000",
         18290 => x"00000000",
         18291 => x"00000000",
         18292 => x"00000000",
         18293 => x"00000000",
         18294 => x"00000000",
         18295 => x"00000000",
         18296 => x"00000000",
         18297 => x"00000000",
         18298 => x"00000000",
         18299 => x"00000000",
         18300 => x"00000000",
         18301 => x"00000000",
         18302 => x"00000000",
         18303 => x"00000000",
         18304 => x"00000000",
         18305 => x"00000000",
         18306 => x"00000000",
         18307 => x"00000000",
         18308 => x"00000000",
         18309 => x"00000000",
         18310 => x"00000000",
         18311 => x"00000000",
         18312 => x"00000000",
         18313 => x"00000000",
         18314 => x"00000000",
         18315 => x"00000000",
         18316 => x"00000000",
         18317 => x"00000000",
         18318 => x"00000000",
         18319 => x"00000000",
         18320 => x"00000000",
         18321 => x"00000000",
         18322 => x"00000000",
         18323 => x"00000000",
         18324 => x"00000000",
         18325 => x"00000000",
         18326 => x"00000000",
         18327 => x"00000000",
         18328 => x"00000000",
         18329 => x"00000000",
         18330 => x"00000000",
         18331 => x"00000000",
         18332 => x"00000000",
         18333 => x"00000000",
         18334 => x"00000000",
         18335 => x"00000000",
         18336 => x"00000000",
         18337 => x"00000000",
         18338 => x"00000000",
         18339 => x"00000000",
         18340 => x"00000000",
         18341 => x"00000000",
         18342 => x"00000000",
         18343 => x"00000000",
         18344 => x"00000000",
         18345 => x"00000000",
         18346 => x"00000000",
         18347 => x"00000000",
         18348 => x"00000000",
         18349 => x"00000000",
         18350 => x"00000000",
         18351 => x"00000000",
         18352 => x"00000000",
         18353 => x"00000000",
         18354 => x"00000000",
         18355 => x"00000000",
         18356 => x"00000000",
         18357 => x"00000000",
         18358 => x"00000000",
         18359 => x"00000000",
         18360 => x"00000000",
         18361 => x"00000000",
         18362 => x"00000000",
         18363 => x"00000000",
         18364 => x"00000000",
         18365 => x"00000000",
         18366 => x"00000000",
         18367 => x"00000000",
         18368 => x"00000000",
         18369 => x"00000000",
         18370 => x"00000000",
         18371 => x"00000000",
         18372 => x"00000000",
         18373 => x"00000000",
         18374 => x"00000000",
         18375 => x"00000000",
         18376 => x"00000000",
         18377 => x"00000000",
         18378 => x"00000000",
         18379 => x"00000000",
         18380 => x"00000000",
         18381 => x"00000000",
         18382 => x"00000000",
         18383 => x"00000000",
         18384 => x"00000000",
         18385 => x"00000000",
         18386 => x"00000000",
         18387 => x"00000000",
         18388 => x"00000000",
         18389 => x"00000000",
         18390 => x"00000000",
         18391 => x"00000000",
         18392 => x"00000000",
         18393 => x"00000000",
         18394 => x"00000000",
         18395 => x"00000000",
         18396 => x"00000000",
         18397 => x"00000000",
         18398 => x"00000000",
         18399 => x"00000000",
         18400 => x"00000000",
         18401 => x"00000000",
         18402 => x"00000000",
         18403 => x"00000000",
         18404 => x"00000000",
         18405 => x"00000000",
         18406 => x"00000000",
         18407 => x"00000000",
         18408 => x"00000000",
         18409 => x"00000000",
         18410 => x"00000000",
         18411 => x"00000000",
         18412 => x"00000000",
         18413 => x"00000000",
         18414 => x"00000000",
         18415 => x"00000000",
         18416 => x"00000000",
         18417 => x"00000000",
         18418 => x"00000000",
         18419 => x"00000000",
         18420 => x"00000000",
         18421 => x"00000000",
         18422 => x"00000000",
         18423 => x"00000000",
         18424 => x"00000000",
         18425 => x"00000000",
         18426 => x"00000000",
         18427 => x"00000000",
         18428 => x"00000000",
         18429 => x"00000000",
         18430 => x"00000000",
         18431 => x"00000000",
         18432 => x"00000000",
         18433 => x"00000000",
         18434 => x"00000000",
         18435 => x"00000000",
         18436 => x"00000000",
         18437 => x"00000000",
         18438 => x"00000000",
         18439 => x"00000000",
         18440 => x"00000000",
         18441 => x"00000000",
         18442 => x"00000000",
         18443 => x"00000000",
         18444 => x"00000000",
         18445 => x"00000000",
         18446 => x"00000000",
         18447 => x"00000000",
         18448 => x"00000000",
         18449 => x"00000000",
         18450 => x"00000000",
         18451 => x"00000000",
         18452 => x"00000000",
         18453 => x"00000000",
         18454 => x"00000000",
         18455 => x"00000000",
         18456 => x"00000000",
         18457 => x"00000000",
         18458 => x"00000000",
         18459 => x"00000000",
         18460 => x"00000000",
         18461 => x"00000000",
         18462 => x"00000000",
         18463 => x"00000000",
         18464 => x"00000000",
         18465 => x"00000000",
         18466 => x"00000000",
         18467 => x"00000000",
         18468 => x"00000000",
         18469 => x"00000000",
         18470 => x"00000000",
         18471 => x"00000000",
         18472 => x"00000000",
         18473 => x"00000000",
         18474 => x"00000000",
         18475 => x"00000000",
         18476 => x"00000000",
         18477 => x"00000000",
         18478 => x"00000000",
         18479 => x"00000000",
         18480 => x"00000000",
         18481 => x"00000000",
         18482 => x"00000000",
         18483 => x"00000000",
         18484 => x"00000000",
         18485 => x"00000000",
         18486 => x"00000000",
         18487 => x"00000000",
         18488 => x"00000000",
         18489 => x"00000000",
         18490 => x"00000000",
         18491 => x"00000000",
         18492 => x"00000000",
         18493 => x"00000000",
         18494 => x"00000000",
         18495 => x"00000000",
         18496 => x"00000000",
         18497 => x"00000000",
         18498 => x"00000000",
         18499 => x"00000000",
         18500 => x"00000000",
         18501 => x"00000000",
         18502 => x"00000000",
         18503 => x"00000000",
         18504 => x"00000000",
         18505 => x"00000000",
         18506 => x"00000000",
         18507 => x"00000000",
         18508 => x"00000000",
         18509 => x"00000000",
         18510 => x"00000000",
         18511 => x"00000000",
         18512 => x"00000000",
         18513 => x"00000000",
         18514 => x"00000000",
         18515 => x"00000000",
         18516 => x"00000000",
         18517 => x"00000000",
         18518 => x"00000000",
         18519 => x"00000000",
         18520 => x"00000000",
         18521 => x"00000000",
         18522 => x"00000000",
         18523 => x"00000000",
         18524 => x"00000000",
         18525 => x"00000000",
         18526 => x"00000000",
         18527 => x"00000000",
         18528 => x"00000000",
         18529 => x"00000000",
         18530 => x"00000000",
         18531 => x"00000000",
         18532 => x"00000000",
         18533 => x"00000000",
         18534 => x"00000000",
         18535 => x"00000000",
         18536 => x"00000000",
         18537 => x"00000000",
         18538 => x"00000000",
         18539 => x"00000000",
         18540 => x"00000000",
         18541 => x"00000000",
         18542 => x"00000000",
         18543 => x"00000000",
         18544 => x"00000000",
         18545 => x"00000000",
         18546 => x"00000000",
         18547 => x"00000000",
         18548 => x"00000000",
         18549 => x"00000000",
         18550 => x"00000000",
         18551 => x"00000000",
         18552 => x"00000000",
         18553 => x"00000000",
         18554 => x"00000000",
         18555 => x"00000000",
         18556 => x"00000000",
         18557 => x"00000000",
         18558 => x"00000000",
         18559 => x"00000000",
         18560 => x"00000000",
         18561 => x"00000000",
         18562 => x"00000000",
         18563 => x"00000000",
         18564 => x"00000000",
         18565 => x"00000000",
         18566 => x"00000000",
         18567 => x"00000000",
         18568 => x"00000000",
         18569 => x"00000000",
         18570 => x"00000000",
         18571 => x"00000000",
         18572 => x"00000000",
         18573 => x"00000000",
         18574 => x"00000000",
         18575 => x"00000000",
         18576 => x"00000000",
         18577 => x"00000000",
         18578 => x"00000000",
         18579 => x"00000000",
         18580 => x"00000000",
         18581 => x"00000000",
         18582 => x"00000000",
         18583 => x"00000000",
         18584 => x"00000000",
         18585 => x"00000000",
         18586 => x"00000000",
         18587 => x"00000000",
         18588 => x"00000000",
         18589 => x"00000000",
         18590 => x"00000000",
         18591 => x"00000000",
         18592 => x"00000000",
         18593 => x"00000000",
         18594 => x"00000000",
         18595 => x"00000000",
         18596 => x"00000000",
         18597 => x"00000000",
         18598 => x"00000000",
         18599 => x"00000000",
         18600 => x"00000000",
         18601 => x"00000000",
         18602 => x"00000000",
         18603 => x"00000000",
         18604 => x"00000000",
         18605 => x"00000000",
         18606 => x"00000000",
         18607 => x"00000000",
         18608 => x"00000000",
         18609 => x"00000000",
         18610 => x"00000000",
         18611 => x"00000000",
         18612 => x"00000000",
         18613 => x"00000000",
         18614 => x"00000000",
         18615 => x"00000000",
         18616 => x"00000000",
         18617 => x"00000000",
         18618 => x"00000000",
         18619 => x"00000000",
         18620 => x"00000000",
         18621 => x"00000000",
         18622 => x"00000000",
         18623 => x"00000000",
         18624 => x"00000000",
         18625 => x"00000000",
         18626 => x"00000000",
         18627 => x"00000000",
         18628 => x"00000000",
         18629 => x"00000000",
         18630 => x"00000000",
         18631 => x"00000000",
         18632 => x"00000000",
         18633 => x"00000000",
         18634 => x"00000000",
         18635 => x"00000000",
         18636 => x"00000000",
         18637 => x"00000000",
         18638 => x"00000000",
         18639 => x"00000000",
         18640 => x"00000000",
         18641 => x"00000000",
         18642 => x"00000000",
         18643 => x"00000000",
         18644 => x"00000000",
         18645 => x"00000000",
         18646 => x"00000000",
         18647 => x"00000000",
         18648 => x"00000000",
         18649 => x"00000000",
         18650 => x"00000000",
         18651 => x"00000000",
         18652 => x"00000000",
         18653 => x"00000000",
         18654 => x"00000000",
         18655 => x"00000000",
         18656 => x"00000000",
         18657 => x"00000000",
         18658 => x"00000000",
         18659 => x"00000000",
         18660 => x"00000000",
         18661 => x"00000000",
         18662 => x"00000000",
         18663 => x"00000000",
         18664 => x"00000000",
         18665 => x"00000000",
         18666 => x"00000000",
         18667 => x"00000000",
         18668 => x"00000000",
         18669 => x"00000000",
         18670 => x"00000000",
         18671 => x"00000000",
         18672 => x"00000000",
         18673 => x"00000000",
         18674 => x"00000000",
         18675 => x"00000000",
         18676 => x"00000000",
         18677 => x"00000000",
         18678 => x"00000000",
         18679 => x"00000000",
         18680 => x"00000000",
         18681 => x"00000000",
         18682 => x"00000000",
         18683 => x"00000000",
         18684 => x"00000000",
         18685 => x"00000000",
         18686 => x"00000000",
         18687 => x"00000000",
         18688 => x"00000000",
         18689 => x"00000000",
         18690 => x"00000000",
         18691 => x"00000000",
         18692 => x"00000000",
         18693 => x"00000000",
         18694 => x"00000000",
         18695 => x"00000000",
         18696 => x"00000000",
         18697 => x"00000000",
         18698 => x"00000000",
         18699 => x"00000000",
         18700 => x"00000000",
         18701 => x"00000000",
         18702 => x"00000000",
         18703 => x"00000000",
         18704 => x"00000000",
         18705 => x"00000000",
         18706 => x"00000000",
         18707 => x"00000000",
         18708 => x"00000000",
         18709 => x"00000000",
         18710 => x"00000000",
         18711 => x"00000000",
         18712 => x"00000000",
         18713 => x"00000000",
         18714 => x"00000000",
         18715 => x"00000000",
         18716 => x"00000000",
         18717 => x"00000000",
         18718 => x"00000000",
         18719 => x"00000000",
         18720 => x"00000000",
         18721 => x"00000000",
         18722 => x"00000000",
         18723 => x"00000000",
         18724 => x"00000000",
         18725 => x"00000000",
         18726 => x"00000000",
         18727 => x"00000000",
         18728 => x"00000000",
         18729 => x"00000000",
         18730 => x"00000000",
         18731 => x"00000000",
         18732 => x"00000000",
         18733 => x"00000000",
         18734 => x"00000000",
         18735 => x"00000000",
         18736 => x"00000000",
         18737 => x"00000000",
         18738 => x"00000000",
         18739 => x"00000000",
         18740 => x"00000000",
         18741 => x"00000000",
         18742 => x"00000000",
         18743 => x"00000000",
         18744 => x"00000000",
         18745 => x"00000000",
         18746 => x"00000000",
         18747 => x"00000000",
         18748 => x"00000000",
         18749 => x"00000000",
         18750 => x"00000000",
         18751 => x"00000000",
         18752 => x"00000000",
         18753 => x"00000000",
         18754 => x"00000000",
         18755 => x"00000000",
         18756 => x"00000000",
         18757 => x"00000000",
         18758 => x"00000000",
         18759 => x"00000000",
         18760 => x"00000000",
         18761 => x"00000000",
         18762 => x"00000000",
         18763 => x"00000000",
         18764 => x"00000000",
         18765 => x"00000000",
         18766 => x"00000000",
         18767 => x"00000000",
         18768 => x"00000000",
         18769 => x"00000000",
         18770 => x"00000000",
         18771 => x"00000000",
         18772 => x"00000000",
         18773 => x"00000000",
         18774 => x"00000000",
         18775 => x"00000000",
         18776 => x"00000000",
         18777 => x"00000000",
         18778 => x"00000000",
         18779 => x"00000000",
         18780 => x"00000000",
         18781 => x"00000000",
         18782 => x"00000000",
         18783 => x"00000000",
         18784 => x"00000000",
         18785 => x"00000000",
         18786 => x"00000000",
         18787 => x"00000000",
         18788 => x"00000000",
         18789 => x"00000000",
         18790 => x"00000000",
         18791 => x"00000000",
         18792 => x"00000000",
         18793 => x"00000000",
         18794 => x"00000000",
         18795 => x"00000000",
         18796 => x"00000000",
         18797 => x"00000000",
         18798 => x"00000000",
         18799 => x"00000000",
         18800 => x"00000000",
         18801 => x"00000000",
         18802 => x"00000000",
         18803 => x"00000000",
         18804 => x"00000000",
         18805 => x"00000000",
         18806 => x"00000000",
         18807 => x"00000000",
         18808 => x"00000000",
         18809 => x"00000000",
         18810 => x"00000000",
         18811 => x"00000000",
         18812 => x"00000000",
         18813 => x"00000000",
         18814 => x"00000000",
         18815 => x"00000000",
         18816 => x"00000000",
         18817 => x"00000000",
         18818 => x"00000000",
         18819 => x"00000000",
         18820 => x"00000000",
         18821 => x"00000000",
         18822 => x"00000000",
         18823 => x"00000000",
         18824 => x"00000000",
         18825 => x"00000000",
         18826 => x"00000000",
         18827 => x"00000000",
         18828 => x"00000000",
         18829 => x"00000000",
         18830 => x"00000000",
         18831 => x"00000000",
         18832 => x"00000000",
         18833 => x"00000000",
         18834 => x"00000000",
         18835 => x"00000000",
         18836 => x"00000000",
         18837 => x"00000000",
         18838 => x"00000000",
         18839 => x"00000000",
         18840 => x"00000000",
         18841 => x"00000000",
         18842 => x"00000000",
         18843 => x"00000000",
         18844 => x"00000000",
         18845 => x"00000000",
         18846 => x"00000000",
         18847 => x"00000000",
         18848 => x"00000000",
         18849 => x"00000000",
         18850 => x"00000000",
         18851 => x"00000000",
         18852 => x"00000000",
         18853 => x"00000000",
         18854 => x"00000000",
         18855 => x"00000000",
         18856 => x"00000000",
         18857 => x"00000000",
         18858 => x"00000000",
         18859 => x"00000000",
         18860 => x"00000000",
         18861 => x"00000000",
         18862 => x"00000000",
         18863 => x"00000000",
         18864 => x"00000000",
         18865 => x"00000000",
         18866 => x"00000000",
         18867 => x"00000000",
         18868 => x"00000000",
         18869 => x"00000000",
         18870 => x"00000000",
         18871 => x"00000000",
         18872 => x"00000000",
         18873 => x"00000000",
         18874 => x"00000000",
         18875 => x"00000000",
         18876 => x"00000000",
         18877 => x"00000000",
         18878 => x"00000000",
         18879 => x"00000000",
         18880 => x"00000000",
         18881 => x"00000000",
         18882 => x"00000000",
         18883 => x"00000000",
         18884 => x"00000000",
         18885 => x"00000000",
         18886 => x"00000000",
         18887 => x"00000000",
         18888 => x"00000000",
         18889 => x"00000000",
         18890 => x"00000000",
         18891 => x"00000000",
         18892 => x"00000000",
         18893 => x"00000000",
         18894 => x"00000000",
         18895 => x"00000000",
         18896 => x"00000000",
         18897 => x"00000000",
         18898 => x"00000000",
         18899 => x"00000000",
         18900 => x"00000000",
         18901 => x"00000000",
         18902 => x"00000000",
         18903 => x"00000000",
         18904 => x"00000000",
         18905 => x"00000000",
         18906 => x"00000000",
         18907 => x"00000000",
         18908 => x"00000000",
         18909 => x"00000000",
         18910 => x"00000000",
         18911 => x"00000000",
         18912 => x"00000000",
         18913 => x"00000000",
         18914 => x"00000000",
         18915 => x"00000000",
         18916 => x"00000000",
         18917 => x"00000000",
         18918 => x"00000000",
         18919 => x"00000000",
         18920 => x"00000000",
         18921 => x"00000000",
         18922 => x"00000000",
         18923 => x"00000000",
         18924 => x"00000000",
         18925 => x"00000000",
         18926 => x"00000000",
         18927 => x"00000000",
         18928 => x"00000000",
         18929 => x"00000000",
         18930 => x"00000000",
         18931 => x"00000000",
         18932 => x"00000000",
         18933 => x"00000000",
         18934 => x"00000000",
         18935 => x"00000000",
         18936 => x"00000000",
         18937 => x"00000000",
         18938 => x"00000000",
         18939 => x"00000000",
         18940 => x"00000000",
         18941 => x"00000000",
         18942 => x"00000000",
         18943 => x"00000000",
         18944 => x"00000000",
         18945 => x"00000000",
         18946 => x"00000000",
         18947 => x"00000000",
         18948 => x"00000000",
         18949 => x"00000000",
         18950 => x"00000000",
         18951 => x"00000000",
         18952 => x"00000000",
         18953 => x"00000000",
         18954 => x"00000000",
         18955 => x"00000000",
         18956 => x"00000000",
         18957 => x"00000000",
         18958 => x"00000000",
         18959 => x"00000000",
         18960 => x"00000000",
         18961 => x"00000000",
         18962 => x"00000000",
         18963 => x"00000000",
         18964 => x"00000000",
         18965 => x"00000000",
         18966 => x"00000000",
         18967 => x"00000000",
         18968 => x"00000000",
         18969 => x"00000000",
         18970 => x"00000000",
         18971 => x"00000000",
         18972 => x"00000000",
         18973 => x"00000000",
         18974 => x"00000000",
         18975 => x"00000000",
         18976 => x"00000000",
         18977 => x"00000000",
         18978 => x"00000000",
         18979 => x"00000000",
         18980 => x"00000000",
         18981 => x"00000000",
         18982 => x"00000000",
         18983 => x"00000000",
         18984 => x"00000000",
         18985 => x"00000000",
         18986 => x"00000000",
         18987 => x"00000000",
         18988 => x"00000000",
         18989 => x"00000000",
         18990 => x"00000000",
         18991 => x"00000000",
         18992 => x"00000000",
         18993 => x"00000000",
         18994 => x"00000000",
         18995 => x"00000000",
         18996 => x"00000000",
         18997 => x"00000000",
         18998 => x"00000000",
         18999 => x"00000000",
         19000 => x"00000000",
         19001 => x"00000000",
         19002 => x"00000000",
         19003 => x"00000000",
         19004 => x"00000000",
         19005 => x"00000000",
         19006 => x"00000000",
         19007 => x"00000000",
         19008 => x"00000000",
         19009 => x"00000000",
         19010 => x"00000000",
         19011 => x"00000000",
         19012 => x"00000000",
         19013 => x"00000000",
         19014 => x"00000000",
         19015 => x"00000000",
         19016 => x"00000000",
         19017 => x"00000000",
         19018 => x"00000000",
         19019 => x"00000000",
         19020 => x"00000000",
         19021 => x"00000000",
         19022 => x"00000000",
         19023 => x"00000000",
         19024 => x"00000000",
         19025 => x"00000000",
         19026 => x"00000000",
         19027 => x"00000000",
         19028 => x"00000000",
         19029 => x"00000000",
         19030 => x"00000000",
         19031 => x"00000000",
         19032 => x"00000000",
         19033 => x"00000000",
         19034 => x"00000000",
         19035 => x"00000000",
         19036 => x"00000000",
         19037 => x"00000000",
         19038 => x"00000000",
         19039 => x"00000000",
         19040 => x"00000000",
         19041 => x"00000000",
         19042 => x"00000000",
         19043 => x"00000000",
         19044 => x"00000000",
         19045 => x"00000000",
         19046 => x"00000000",
         19047 => x"00000000",
         19048 => x"00000000",
         19049 => x"00000000",
         19050 => x"00000000",
         19051 => x"00000000",
         19052 => x"00000000",
         19053 => x"00000000",
         19054 => x"00000000",
         19055 => x"00000000",
         19056 => x"00000000",
         19057 => x"00000000",
         19058 => x"00000000",
         19059 => x"00000000",
         19060 => x"00000000",
         19061 => x"00000000",
         19062 => x"00000000",
         19063 => x"00000000",
         19064 => x"00000000",
         19065 => x"00000000",
         19066 => x"00000000",
         19067 => x"00000000",
         19068 => x"00000000",
         19069 => x"00000000",
         19070 => x"00000000",
         19071 => x"00000000",
         19072 => x"00000000",
         19073 => x"00000000",
         19074 => x"00000000",
         19075 => x"00000000",
         19076 => x"00000000",
         19077 => x"00000000",
         19078 => x"00000000",
         19079 => x"00000000",
         19080 => x"00000000",
         19081 => x"00000000",
         19082 => x"00000000",
         19083 => x"00000000",
         19084 => x"00000000",
         19085 => x"00000000",
         19086 => x"00000000",
         19087 => x"00000000",
         19088 => x"00000000",
         19089 => x"00000000",
         19090 => x"00000000",
         19091 => x"00000000",
         19092 => x"00000000",
         19093 => x"00000000",
         19094 => x"00000000",
         19095 => x"00000000",
         19096 => x"00000000",
         19097 => x"00000000",
         19098 => x"00000000",
         19099 => x"00000000",
         19100 => x"00000000",
         19101 => x"00000000",
         19102 => x"00000000",
         19103 => x"00000000",
         19104 => x"00000000",
         19105 => x"00000000",
         19106 => x"00000000",
         19107 => x"00000000",
         19108 => x"00000000",
         19109 => x"00000000",
         19110 => x"00000000",
         19111 => x"00000000",
         19112 => x"00000000",
         19113 => x"00000000",
         19114 => x"00000000",
         19115 => x"00000000",
         19116 => x"00000000",
         19117 => x"00000000",
         19118 => x"00000000",
         19119 => x"00000000",
         19120 => x"00000000",
         19121 => x"00000000",
         19122 => x"00000000",
         19123 => x"00000000",
         19124 => x"00000000",
         19125 => x"00000000",
         19126 => x"00000000",
         19127 => x"00000000",
         19128 => x"00000000",
         19129 => x"00000000",
         19130 => x"00000000",
         19131 => x"00000000",
         19132 => x"00000000",
         19133 => x"00000000",
         19134 => x"00000000",
         19135 => x"00000000",
         19136 => x"00000000",
         19137 => x"00000000",
         19138 => x"00000000",
         19139 => x"00000000",
         19140 => x"00000000",
         19141 => x"00000000",
         19142 => x"00000000",
         19143 => x"00000000",
         19144 => x"00000000",
         19145 => x"00000000",
         19146 => x"00000000",
         19147 => x"00000000",
         19148 => x"00000000",
         19149 => x"00000000",
         19150 => x"00000000",
         19151 => x"00000000",
         19152 => x"00000000",
         19153 => x"00000000",
         19154 => x"00000000",
         19155 => x"00000000",
         19156 => x"00000000",
         19157 => x"00000000",
         19158 => x"00000000",
         19159 => x"00000000",
         19160 => x"00000000",
         19161 => x"00000000",
         19162 => x"00000000",
         19163 => x"00000000",
         19164 => x"00000000",
         19165 => x"00000000",
         19166 => x"00000000",
         19167 => x"00000000",
         19168 => x"00000000",
         19169 => x"00000000",
         19170 => x"00000000",
         19171 => x"00000000",
         19172 => x"00000000",
         19173 => x"00000000",
         19174 => x"00000000",
         19175 => x"00000000",
         19176 => x"00000000",
         19177 => x"00000000",
         19178 => x"00000000",
         19179 => x"00000000",
         19180 => x"00000000",
         19181 => x"00000000",
         19182 => x"00000000",
         19183 => x"00000000",
         19184 => x"00000000",
         19185 => x"00000000",
         19186 => x"00000000",
         19187 => x"00000000",
         19188 => x"00000000",
         19189 => x"00000000",
         19190 => x"00000000",
         19191 => x"00000000",
         19192 => x"00000000",
         19193 => x"00000000",
         19194 => x"00000000",
         19195 => x"00000000",
         19196 => x"00000000",
         19197 => x"00000000",
         19198 => x"00000000",
         19199 => x"00000000",
         19200 => x"00000000",
         19201 => x"00000000",
         19202 => x"00000000",
         19203 => x"00000000",
         19204 => x"00000000",
         19205 => x"00000000",
         19206 => x"00000000",
         19207 => x"00000000",
         19208 => x"00000000",
         19209 => x"00000000",
         19210 => x"00000000",
         19211 => x"00000000",
         19212 => x"00000000",
         19213 => x"00000000",
         19214 => x"00000000",
         19215 => x"00000000",
         19216 => x"00000000",
         19217 => x"00000000",
         19218 => x"00000000",
         19219 => x"00000000",
         19220 => x"00000000",
         19221 => x"00000000",
         19222 => x"00000000",
         19223 => x"00000000",
         19224 => x"00000000",
         19225 => x"00000000",
         19226 => x"00000000",
         19227 => x"00000000",
         19228 => x"00000000",
         19229 => x"00000000",
         19230 => x"00000000",
         19231 => x"00000000",
         19232 => x"00000000",
         19233 => x"00000000",
         19234 => x"00000000",
         19235 => x"00000000",
         19236 => x"00000000",
         19237 => x"00000000",
         19238 => x"00000000",
         19239 => x"00000000",
         19240 => x"00000000",
         19241 => x"00000000",
         19242 => x"00000000",
         19243 => x"00000000",
         19244 => x"00000000",
         19245 => x"00000000",
         19246 => x"00000000",
         19247 => x"00000000",
         19248 => x"00000000",
         19249 => x"00000000",
         19250 => x"00000000",
         19251 => x"00000000",
         19252 => x"00000000",
         19253 => x"00000000",
         19254 => x"00000000",
         19255 => x"00000000",
         19256 => x"00000000",
         19257 => x"00000000",
         19258 => x"00000000",
         19259 => x"00000000",
         19260 => x"00000000",
         19261 => x"00000000",
         19262 => x"00000000",
         19263 => x"00000000",
         19264 => x"00000000",
         19265 => x"00000000",
         19266 => x"00000000",
         19267 => x"00000000",
         19268 => x"00000000",
         19269 => x"00000000",
         19270 => x"00000000",
         19271 => x"00000000",
         19272 => x"00000000",
         19273 => x"00000000",
         19274 => x"00000000",
         19275 => x"00000000",
         19276 => x"00000000",
         19277 => x"00000000",
         19278 => x"00000000",
         19279 => x"00000000",
         19280 => x"00000000",
         19281 => x"00000000",
         19282 => x"00000000",
         19283 => x"00000000",
         19284 => x"00000000",
         19285 => x"00000000",
         19286 => x"00000000",
         19287 => x"00000000",
         19288 => x"00000000",
         19289 => x"00000000",
         19290 => x"00000000",
         19291 => x"00000000",
         19292 => x"00000000",
         19293 => x"00000000",
         19294 => x"00000000",
         19295 => x"00000000",
         19296 => x"00000000",
         19297 => x"00000000",
         19298 => x"00000000",
         19299 => x"00000000",
         19300 => x"00000000",
         19301 => x"00000000",
         19302 => x"00000000",
         19303 => x"00000000",
         19304 => x"00000000",
         19305 => x"00000000",
         19306 => x"00000000",
         19307 => x"00000000",
         19308 => x"00000000",
         19309 => x"00000000",
         19310 => x"00000000",
         19311 => x"00000000",
         19312 => x"00000000",
         19313 => x"00000000",
         19314 => x"00000000",
         19315 => x"00000000",
         19316 => x"00000000",
         19317 => x"00000000",
         19318 => x"00000000",
         19319 => x"00000000",
         19320 => x"00000000",
         19321 => x"00000000",
         19322 => x"00000000",
         19323 => x"00000000",
         19324 => x"00000000",
         19325 => x"00000000",
         19326 => x"00000000",
         19327 => x"00000000",
         19328 => x"00000000",
         19329 => x"00000000",
         19330 => x"00000000",
         19331 => x"00000000",
         19332 => x"00000000",
         19333 => x"00000000",
         19334 => x"00000000",
         19335 => x"00000000",
         19336 => x"00000000",
         19337 => x"00000000",
         19338 => x"00000000",
         19339 => x"00000000",
         19340 => x"00000000",
         19341 => x"00000000",
         19342 => x"00000000",
         19343 => x"00000000",
         19344 => x"00000000",
         19345 => x"00000000",
         19346 => x"00000000",
         19347 => x"00000000",
         19348 => x"00000000",
         19349 => x"00000000",
         19350 => x"00000000",
         19351 => x"00000000",
         19352 => x"00000000",
         19353 => x"00000000",
         19354 => x"00000000",
         19355 => x"00000000",
         19356 => x"00000000",
         19357 => x"00000000",
         19358 => x"00000000",
         19359 => x"00000000",
         19360 => x"00000000",
         19361 => x"00000000",
         19362 => x"00000000",
         19363 => x"00000000",
         19364 => x"00000000",
         19365 => x"00000000",
         19366 => x"00000000",
         19367 => x"00000000",
         19368 => x"00000000",
         19369 => x"00000000",
         19370 => x"00000000",
         19371 => x"00000000",
         19372 => x"00000000",
         19373 => x"00000000",
         19374 => x"00000000",
         19375 => x"00000000",
         19376 => x"00000000",
         19377 => x"00000000",
         19378 => x"00000000",
         19379 => x"00000000",
         19380 => x"00000000",
         19381 => x"00000000",
         19382 => x"00000000",
         19383 => x"00000000",
         19384 => x"00000000",
         19385 => x"00000000",
         19386 => x"00000000",
         19387 => x"00000000",
         19388 => x"00000000",
         19389 => x"00000000",
         19390 => x"00000000",
         19391 => x"00000000",
         19392 => x"00000000",
         19393 => x"00000000",
         19394 => x"00000000",
         19395 => x"00000000",
         19396 => x"00000000",
         19397 => x"00000000",
         19398 => x"00000000",
         19399 => x"00000000",
         19400 => x"00000000",
         19401 => x"00000000",
         19402 => x"00000000",
         19403 => x"00000000",
         19404 => x"00000000",
         19405 => x"00000000",
         19406 => x"00000000",
         19407 => x"00000000",
         19408 => x"00000000",
         19409 => x"00000000",
         19410 => x"00000000",
         19411 => x"00000000",
         19412 => x"00000000",
         19413 => x"00000000",
         19414 => x"00000000",
         19415 => x"00000000",
         19416 => x"00000000",
         19417 => x"00000000",
         19418 => x"00000000",
         19419 => x"00000000",
         19420 => x"00000000",
         19421 => x"00000000",
         19422 => x"00000000",
         19423 => x"00000000",
         19424 => x"00000000",
         19425 => x"00000000",
         19426 => x"00000000",
         19427 => x"00000000",
         19428 => x"00000000",
         19429 => x"00000000",
         19430 => x"00000000",
         19431 => x"00000000",
         19432 => x"00000000",
         19433 => x"00000000",
         19434 => x"00000000",
         19435 => x"00000000",
         19436 => x"00000000",
         19437 => x"00000000",
         19438 => x"00000000",
         19439 => x"00000000",
         19440 => x"00000000",
         19441 => x"00000000",
         19442 => x"00000000",
         19443 => x"00000000",
         19444 => x"00000000",
         19445 => x"00000000",
         19446 => x"00000000",
         19447 => x"00000000",
         19448 => x"00000000",
         19449 => x"00000000",
         19450 => x"00000000",
         19451 => x"00000000",
         19452 => x"00000000",
         19453 => x"00000000",
         19454 => x"00000000",
         19455 => x"00000000",
         19456 => x"00000000",
         19457 => x"00000000",
         19458 => x"00000000",
         19459 => x"00000000",
         19460 => x"00000000",
         19461 => x"00000000",
         19462 => x"00000000",
         19463 => x"00000000",
         19464 => x"00000000",
         19465 => x"00000000",
         19466 => x"00000000",
         19467 => x"00000000",
         19468 => x"00000000",
         19469 => x"00000000",
         19470 => x"00000000",
         19471 => x"00000000",
         19472 => x"00000000",
         19473 => x"00000000",
         19474 => x"00000000",
         19475 => x"00000000",
         19476 => x"00000000",
         19477 => x"00000000",
         19478 => x"00000000",
         19479 => x"00000000",
         19480 => x"00000000",
         19481 => x"00000000",
         19482 => x"00000000",
         19483 => x"00000000",
         19484 => x"00000000",
         19485 => x"00000000",
         19486 => x"00000000",
         19487 => x"00000000",
         19488 => x"00000000",
         19489 => x"00000000",
         19490 => x"00000000",
         19491 => x"00000000",
         19492 => x"00000000",
         19493 => x"00000000",
         19494 => x"00000000",
         19495 => x"00000000",
         19496 => x"00000000",
         19497 => x"00000000",
         19498 => x"00000000",
         19499 => x"00000000",
         19500 => x"00000000",
         19501 => x"00000000",
         19502 => x"00000000",
         19503 => x"00000000",
         19504 => x"00000000",
         19505 => x"00000000",
         19506 => x"00000000",
         19507 => x"00000000",
         19508 => x"00000000",
         19509 => x"00000000",
         19510 => x"00000000",
         19511 => x"00000000",
         19512 => x"00000000",
         19513 => x"00000000",
         19514 => x"00000000",
         19515 => x"00000000",
         19516 => x"00000000",
         19517 => x"00000000",
         19518 => x"00000000",
         19519 => x"00000000",
         19520 => x"00000000",
         19521 => x"00000000",
         19522 => x"00000000",
         19523 => x"00000000",
         19524 => x"00000000",
         19525 => x"00000000",
         19526 => x"00000000",
         19527 => x"00000000",
         19528 => x"00000000",
         19529 => x"00000000",
         19530 => x"00000000",
         19531 => x"00000000",
         19532 => x"00000000",
         19533 => x"00000000",
         19534 => x"00000000",
         19535 => x"00000000",
         19536 => x"00000000",
         19537 => x"00000000",
         19538 => x"00000000",
         19539 => x"00000000",
         19540 => x"00000000",
         19541 => x"00000000",
         19542 => x"00000000",
         19543 => x"00000000",
         19544 => x"00000000",
         19545 => x"00000000",
         19546 => x"00000000",
         19547 => x"00000000",
         19548 => x"00000000",
         19549 => x"00000000",
         19550 => x"00000000",
         19551 => x"00000000",
         19552 => x"00000000",
         19553 => x"00000000",
         19554 => x"00000000",
         19555 => x"00000000",
         19556 => x"00000000",
         19557 => x"00000000",
         19558 => x"00000000",
         19559 => x"00000000",
         19560 => x"00000000",
         19561 => x"00000000",
         19562 => x"00000000",
         19563 => x"00000000",
         19564 => x"00000000",
         19565 => x"00000000",
         19566 => x"00000000",
         19567 => x"00000000",
         19568 => x"00000000",
         19569 => x"00000000",
         19570 => x"00000000",
         19571 => x"00000000",
         19572 => x"00000000",
         19573 => x"00000000",
         19574 => x"00000000",
         19575 => x"00000000",
         19576 => x"00000000",
         19577 => x"00000000",
         19578 => x"00000000",
         19579 => x"00000000",
         19580 => x"00000000",
         19581 => x"00000000",
         19582 => x"00000000",
         19583 => x"00000000",
         19584 => x"00000000",
         19585 => x"00000000",
         19586 => x"00000000",
         19587 => x"00000000",
         19588 => x"00000000",
         19589 => x"00000000",
         19590 => x"00000000",
         19591 => x"00000000",
         19592 => x"00000000",
         19593 => x"00000000",
         19594 => x"00000000",
         19595 => x"00000000",
         19596 => x"00000000",
         19597 => x"00000000",
         19598 => x"00000000",
         19599 => x"00000000",
         19600 => x"00000000",
         19601 => x"00000000",
         19602 => x"00000000",
         19603 => x"00000000",
         19604 => x"00000000",
         19605 => x"00000000",
         19606 => x"00000000",
         19607 => x"00000000",
         19608 => x"00000000",
         19609 => x"00000000",
         19610 => x"00000000",
         19611 => x"00000000",
         19612 => x"00000000",
         19613 => x"00000000",
         19614 => x"00000000",
         19615 => x"00000000",
         19616 => x"00000000",
         19617 => x"00000000",
         19618 => x"00000000",
         19619 => x"00000000",
         19620 => x"00000000",
         19621 => x"00000000",
         19622 => x"00000000",
         19623 => x"00000000",
         19624 => x"00000000",
         19625 => x"00000000",
         19626 => x"00000000",
         19627 => x"00000000",
         19628 => x"00000000",
         19629 => x"00000000",
         19630 => x"00000000",
         19631 => x"00000000",
         19632 => x"00000000",
         19633 => x"00000000",
         19634 => x"00000000",
         19635 => x"00000000",
         19636 => x"00000000",
         19637 => x"00000000",
         19638 => x"00000000",
         19639 => x"00000000",
         19640 => x"00000000",
         19641 => x"00000000",
         19642 => x"00000000",
         19643 => x"00000000",
         19644 => x"00000000",
         19645 => x"00000000",
         19646 => x"00000000",
         19647 => x"00000000",
         19648 => x"00000000",
         19649 => x"00000000",
         19650 => x"00000000",
         19651 => x"00000000",
         19652 => x"00000000",
         19653 => x"00000000",
         19654 => x"00000000",
         19655 => x"00000000",
         19656 => x"00000000",
         19657 => x"00000000",
         19658 => x"00000000",
         19659 => x"00000000",
         19660 => x"00000000",
         19661 => x"00000000",
         19662 => x"00000000",
         19663 => x"00000000",
         19664 => x"00000000",
         19665 => x"00000000",
         19666 => x"00000000",
         19667 => x"00000000",
         19668 => x"00000000",
         19669 => x"00000000",
         19670 => x"00000000",
         19671 => x"00000000",
         19672 => x"00000000",
         19673 => x"00000000",
         19674 => x"00000000",
         19675 => x"00000000",
         19676 => x"00000000",
         19677 => x"00000000",
         19678 => x"00000000",
         19679 => x"00000000",
         19680 => x"00000000",
         19681 => x"00000000",
         19682 => x"00000000",
         19683 => x"00000000",
         19684 => x"00000000",
         19685 => x"00000000",
         19686 => x"00000000",
         19687 => x"00000000",
         19688 => x"00000000",
         19689 => x"00000000",
         19690 => x"00000000",
         19691 => x"00000000",
         19692 => x"00000000",
         19693 => x"00000000",
         19694 => x"00000000",
         19695 => x"00000000",
         19696 => x"00000000",
         19697 => x"00000000",
         19698 => x"00000000",
         19699 => x"00000000",
         19700 => x"00000000",
         19701 => x"00000000",
         19702 => x"00000000",
         19703 => x"00000000",
         19704 => x"00000000",
         19705 => x"00000000",
         19706 => x"00000000",
         19707 => x"00000000",
         19708 => x"00000000",
         19709 => x"00000000",
         19710 => x"00000000",
         19711 => x"00000000",
         19712 => x"00000000",
         19713 => x"00000000",
         19714 => x"00000000",
         19715 => x"00000000",
         19716 => x"00000000",
         19717 => x"00000000",
         19718 => x"00000000",
         19719 => x"00000000",
         19720 => x"00000000",
         19721 => x"00000000",
         19722 => x"00000000",
         19723 => x"00000000",
         19724 => x"00000000",
         19725 => x"00000000",
         19726 => x"00000000",
         19727 => x"00000000",
         19728 => x"00000000",
         19729 => x"00000000",
         19730 => x"00000000",
         19731 => x"00000000",
         19732 => x"00000000",
         19733 => x"00000000",
         19734 => x"00000000",
         19735 => x"00000000",
         19736 => x"00000000",
         19737 => x"00000000",
         19738 => x"00000000",
         19739 => x"00000000",
         19740 => x"00000000",
         19741 => x"00000000",
         19742 => x"00000000",
         19743 => x"00000000",
         19744 => x"00000000",
         19745 => x"00000000",
         19746 => x"00000000",
         19747 => x"00000000",
         19748 => x"00000000",
         19749 => x"00000000",
         19750 => x"00000000",
         19751 => x"00000000",
         19752 => x"00000000",
         19753 => x"00000000",
         19754 => x"00000000",
         19755 => x"00000000",
         19756 => x"00000000",
         19757 => x"00000000",
         19758 => x"00000000",
         19759 => x"00000000",
         19760 => x"00000000",
         19761 => x"00000000",
         19762 => x"00000000",
         19763 => x"00000000",
         19764 => x"00000000",
         19765 => x"00000000",
         19766 => x"00000000",
         19767 => x"00000000",
         19768 => x"00000000",
         19769 => x"00000000",
         19770 => x"00000000",
         19771 => x"00000000",
         19772 => x"00000000",
         19773 => x"00000000",
         19774 => x"00000000",
         19775 => x"00000000",
         19776 => x"00000000",
         19777 => x"00000000",
         19778 => x"00000000",
         19779 => x"00000000",
         19780 => x"00000000",
         19781 => x"00000000",
         19782 => x"00000000",
         19783 => x"00000000",
         19784 => x"00000000",
         19785 => x"00000000",
         19786 => x"00000000",
         19787 => x"00000000",
         19788 => x"00000000",
         19789 => x"00000000",
         19790 => x"00000000",
         19791 => x"00000000",
         19792 => x"00000000",
         19793 => x"00000000",
         19794 => x"00000000",
         19795 => x"00000000",
         19796 => x"00000000",
         19797 => x"00000000",
         19798 => x"00000000",
         19799 => x"00000000",
         19800 => x"00000000",
         19801 => x"00000000",
         19802 => x"00000000",
         19803 => x"00000000",
         19804 => x"00000000",
         19805 => x"00000000",
         19806 => x"00000000",
         19807 => x"00000000",
         19808 => x"00000000",
         19809 => x"00000000",
         19810 => x"00000000",
         19811 => x"00000000",
         19812 => x"00000000",
         19813 => x"00000000",
         19814 => x"00000000",
         19815 => x"00000000",
         19816 => x"00000000",
         19817 => x"00000000",
         19818 => x"00000000",
         19819 => x"00000000",
         19820 => x"00000000",
         19821 => x"00000000",
         19822 => x"00000000",
         19823 => x"00000000",
         19824 => x"00000000",
         19825 => x"00000000",
         19826 => x"00000000",
         19827 => x"00000000",
         19828 => x"00000000",
         19829 => x"00000000",
         19830 => x"00000000",
         19831 => x"00000000",
         19832 => x"00000000",
         19833 => x"00000000",
         19834 => x"00000000",
         19835 => x"00000000",
         19836 => x"00000000",
         19837 => x"00000000",
         19838 => x"00000000",
         19839 => x"00000000",
         19840 => x"00000000",
         19841 => x"00000000",
         19842 => x"00000000",
         19843 => x"00000000",
         19844 => x"00000000",
         19845 => x"00000000",
         19846 => x"00000000",
         19847 => x"00000000",
         19848 => x"00000000",
         19849 => x"00000000",
         19850 => x"00000000",
         19851 => x"00000000",
         19852 => x"00000000",
         19853 => x"00000000",
         19854 => x"00000000",
         19855 => x"00000000",
         19856 => x"00000000",
         19857 => x"00000000",
         19858 => x"00000000",
         19859 => x"00000000",
         19860 => x"00000000",
         19861 => x"00000000",
         19862 => x"00000000",
         19863 => x"00000000",
         19864 => x"00000000",
         19865 => x"00000000",
         19866 => x"00000000",
         19867 => x"00000000",
         19868 => x"00000000",
         19869 => x"00000000",
         19870 => x"00000000",
         19871 => x"00000000",
         19872 => x"00000000",
         19873 => x"00000000",
         19874 => x"00000000",
         19875 => x"00000000",
         19876 => x"00000000",
         19877 => x"00000000",
         19878 => x"00000000",
         19879 => x"00000000",
         19880 => x"00000000",
         19881 => x"00000000",
         19882 => x"00000000",
         19883 => x"00000000",
         19884 => x"00000000",
         19885 => x"00000000",
         19886 => x"00000000",
         19887 => x"00000000",
         19888 => x"00000000",
         19889 => x"00000000",
         19890 => x"00000000",
         19891 => x"00000000",
         19892 => x"00000000",
         19893 => x"00000000",
         19894 => x"00000000",
         19895 => x"00000000",
         19896 => x"00000000",
         19897 => x"00000000",
         19898 => x"00000000",
         19899 => x"00000000",
         19900 => x"00000000",
         19901 => x"00000000",
         19902 => x"00000000",
         19903 => x"00000000",
         19904 => x"00000000",
         19905 => x"00000000",
         19906 => x"00000000",
         19907 => x"00000000",
         19908 => x"00000000",
         19909 => x"00000000",
         19910 => x"00000000",
         19911 => x"00000000",
         19912 => x"00000000",
         19913 => x"00000000",
         19914 => x"00000000",
         19915 => x"00000000",
         19916 => x"00000000",
         19917 => x"00000000",
         19918 => x"00000000",
         19919 => x"00000000",
         19920 => x"00000000",
         19921 => x"00000000",
         19922 => x"00000000",
         19923 => x"00000000",
         19924 => x"00000000",
         19925 => x"00000000",
         19926 => x"00000000",
         19927 => x"00000000",
         19928 => x"00000000",
         19929 => x"00000000",
         19930 => x"00000000",
         19931 => x"00000000",
         19932 => x"00000000",
         19933 => x"00000000",
         19934 => x"00000000",
         19935 => x"00000000",
         19936 => x"00000000",
         19937 => x"00000000",
         19938 => x"00000000",
         19939 => x"00000000",
         19940 => x"00000000",
         19941 => x"00000000",
         19942 => x"00000000",
         19943 => x"00000000",
         19944 => x"00000000",
         19945 => x"00000000",
         19946 => x"00000000",
         19947 => x"00000000",
         19948 => x"00000000",
         19949 => x"00000000",
         19950 => x"00000000",
         19951 => x"00000000",
         19952 => x"00000000",
         19953 => x"00000000",
         19954 => x"00000000",
         19955 => x"00000000",
         19956 => x"00000000",
         19957 => x"00000000",
         19958 => x"00000000",
         19959 => x"00000000",
         19960 => x"00000000",
         19961 => x"00000000",
         19962 => x"00000000",
         19963 => x"00000000",
         19964 => x"00000000",
         19965 => x"00000000",
         19966 => x"00000000",
         19967 => x"00000000",
         19968 => x"00000000",
         19969 => x"00000000",
         19970 => x"00000000",
         19971 => x"00000000",
         19972 => x"00000000",
         19973 => x"00000000",
         19974 => x"00000000",
         19975 => x"00000000",
         19976 => x"00000000",
         19977 => x"00000000",
         19978 => x"00000000",
         19979 => x"00000000",
         19980 => x"00000000",
         19981 => x"00000000",
         19982 => x"00000000",
         19983 => x"00000000",
         19984 => x"00000000",
         19985 => x"00000000",
         19986 => x"00000000",
         19987 => x"00000000",
         19988 => x"00000000",
         19989 => x"00000000",
         19990 => x"00000000",
         19991 => x"00000000",
         19992 => x"00000000",
         19993 => x"00000000",
         19994 => x"00000000",
         19995 => x"00000000",
         19996 => x"00000000",
         19997 => x"00000000",
         19998 => x"00000000",
         19999 => x"00000000",
         20000 => x"00000000",
         20001 => x"00000000",
         20002 => x"00000000",
         20003 => x"00000000",
         20004 => x"00000000",
         20005 => x"00000000",
         20006 => x"00000000",
         20007 => x"00000000",
         20008 => x"00000000",
         20009 => x"00000000",
         20010 => x"00000000",
         20011 => x"00000000",
         20012 => x"00000000",
         20013 => x"00000000",
         20014 => x"00000000",
         20015 => x"00000000",
         20016 => x"00000000",
         20017 => x"00000000",
         20018 => x"00000000",
         20019 => x"00000000",
         20020 => x"00000000",
         20021 => x"00000000",
         20022 => x"00000000",
         20023 => x"00000000",
         20024 => x"00000000",
         20025 => x"00000000",
         20026 => x"00000000",
         20027 => x"00000000",
         20028 => x"00000000",
         20029 => x"00000000",
         20030 => x"00000000",
         20031 => x"00000000",
         20032 => x"00000000",
         20033 => x"00000000",
         20034 => x"00000000",
         20035 => x"00000000",
         20036 => x"00000000",
         20037 => x"00000000",
         20038 => x"00000000",
         20039 => x"00000000",
         20040 => x"00000000",
         20041 => x"00000000",
         20042 => x"00000000",
         20043 => x"00000000",
         20044 => x"00000000",
         20045 => x"00000000",
         20046 => x"00000000",
         20047 => x"00000000",
         20048 => x"00000000",
         20049 => x"00000000",
         20050 => x"00000000",
         20051 => x"00000000",
         20052 => x"00000000",
         20053 => x"00000000",
         20054 => x"00000000",
         20055 => x"00000000",
         20056 => x"00000000",
         20057 => x"00000000",
         20058 => x"00000000",
         20059 => x"00000000",
         20060 => x"00000000",
         20061 => x"00000000",
         20062 => x"00000000",
         20063 => x"00000000",
         20064 => x"00000000",
         20065 => x"00000000",
         20066 => x"00000000",
         20067 => x"00000000",
         20068 => x"00000000",
         20069 => x"00000000",
         20070 => x"00000000",
         20071 => x"00000000",
         20072 => x"00000000",
         20073 => x"00000000",
         20074 => x"00000000",
         20075 => x"00000000",
         20076 => x"00000000",
         20077 => x"00000000",
         20078 => x"00000000",
         20079 => x"00000000",
         20080 => x"00000000",
         20081 => x"00000000",
         20082 => x"00000000",
         20083 => x"00000000",
         20084 => x"00000000",
         20085 => x"00000000",
         20086 => x"00000000",
         20087 => x"00000000",
         20088 => x"00000000",
         20089 => x"00000000",
         20090 => x"00000000",
         20091 => x"00000000",
         20092 => x"00000000",
         20093 => x"00000000",
         20094 => x"00000000",
         20095 => x"00000000",
         20096 => x"00000000",
         20097 => x"00000000",
         20098 => x"00000000",
         20099 => x"00000000",
         20100 => x"00000000",
         20101 => x"00000000",
         20102 => x"00000000",
         20103 => x"00000000",
         20104 => x"00000000",
         20105 => x"00000000",
         20106 => x"00000000",
         20107 => x"00000000",
         20108 => x"00000000",
         20109 => x"00000000",
         20110 => x"00000000",
         20111 => x"00000000",
         20112 => x"00000000",
         20113 => x"00000000",
         20114 => x"00000000",
         20115 => x"00000000",
         20116 => x"00000000",
         20117 => x"00000000",
         20118 => x"00000000",
         20119 => x"00000000",
         20120 => x"00000000",
         20121 => x"00000000",
         20122 => x"00000000",
         20123 => x"00000000",
         20124 => x"00000000",
         20125 => x"00000000",
         20126 => x"00000000",
         20127 => x"00000000",
         20128 => x"00000000",
         20129 => x"00000000",
         20130 => x"00000000",
         20131 => x"00000000",
         20132 => x"00000000",
         20133 => x"00000000",
         20134 => x"00000000",
         20135 => x"00000000",
         20136 => x"00000000",
         20137 => x"00000000",
         20138 => x"00000000",
         20139 => x"00000000",
         20140 => x"00000000",
         20141 => x"00000000",
         20142 => x"00000000",
         20143 => x"00000000",
         20144 => x"00000000",
         20145 => x"00000000",
         20146 => x"00000000",
         20147 => x"00000000",
         20148 => x"00000000",
         20149 => x"00000000",
         20150 => x"00000000",
         20151 => x"00000000",
         20152 => x"00000000",
         20153 => x"00000000",
         20154 => x"00000000",
         20155 => x"00000000",
         20156 => x"00000000",
         20157 => x"00000000",
         20158 => x"00000000",
         20159 => x"00000000",
         20160 => x"00000000",
         20161 => x"00000000",
         20162 => x"00000000",
         20163 => x"00000000",
         20164 => x"00000000",
         20165 => x"00000000",
         20166 => x"00000000",
         20167 => x"00000000",
         20168 => x"00000000",
         20169 => x"00000000",
         20170 => x"00000000",
         20171 => x"00000000",
         20172 => x"00000000",
         20173 => x"00000000",
         20174 => x"00000000",
         20175 => x"00000000",
         20176 => x"00000000",
         20177 => x"00000000",
         20178 => x"00000000",
         20179 => x"00000000",
         20180 => x"00000000",
         20181 => x"00003219",
         20182 => x"50000100",
         20183 => x"00000000",
         20184 => x"cce0f2f3",
         20185 => x"cecff6f7",
         20186 => x"f8f9fafb",
         20187 => x"fcfdfeff",
         20188 => x"e1c1c2c3",
         20189 => x"c4c5c6e2",
         20190 => x"e3e4e5e6",
         20191 => x"ebeeeff4",
         20192 => x"00616263",
         20193 => x"64656667",
         20194 => x"68696b6a",
         20195 => x"2f2a2e2d",
         20196 => x"20212223",
         20197 => x"24252627",
         20198 => x"28294f2c",
         20199 => x"512b5749",
         20200 => x"55010203",
         20201 => x"04050607",
         20202 => x"08090a0b",
         20203 => x"0c0d0e0f",
         20204 => x"10111213",
         20205 => x"14151617",
         20206 => x"18191a52",
         20207 => x"5954be3c",
         20208 => x"c7818283",
         20209 => x"84858687",
         20210 => x"88898a8b",
         20211 => x"8c8d8e8f",
         20212 => x"90919293",
         20213 => x"94959697",
         20214 => x"98999abc",
         20215 => x"8040a5c0",
         20216 => x"00000000",
         20217 => x"00000000",
         20218 => x"00000000",
         20219 => x"00000000",
         20220 => x"00000000",
         20221 => x"00000000",
         20222 => x"00000000",
         20223 => x"00000000",
         20224 => x"00000000",
         20225 => x"00000000",
         20226 => x"00000000",
         20227 => x"00000000",
         20228 => x"00000000",
         20229 => x"00000000",
         20230 => x"00000000",
         20231 => x"00000000",
         20232 => x"00000000",
         20233 => x"00000000",
         20234 => x"00000000",
         20235 => x"00000000",
         20236 => x"00000000",
         20237 => x"00000000",
         20238 => x"00000000",
         20239 => x"00000000",
         20240 => x"00000000",
         20241 => x"00000000",
         20242 => x"00000000",
         20243 => x"00000000",
         20244 => x"00000000",
         20245 => x"00000000",
         20246 => x"00020003",
         20247 => x"00040101",
         20248 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

