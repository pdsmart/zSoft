-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b83ff",
          2049 => x"f80d0b0b",
          2050 => x"0b93b704",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b93",
          2121 => x"9b040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b92fe",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b8294",
          2210 => x"b0738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"93830400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b80cf",
          2219 => x"942d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b80d1",
          2227 => x"802d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"95040b0b",
          2317 => x"0b8ca404",
          2318 => x"0b0b0b8c",
          2319 => x"b3040b0b",
          2320 => x"0b8cc204",
          2321 => x"0b0b0b8c",
          2322 => x"d1040b0b",
          2323 => x"0b8ce004",
          2324 => x"0b0b0b8c",
          2325 => x"ef040b0b",
          2326 => x"0b8cfe04",
          2327 => x"0b0b0b8d",
          2328 => x"8d040b0b",
          2329 => x"0b8d9c04",
          2330 => x"0b0b0b8d",
          2331 => x"ab040b0b",
          2332 => x"0b8dbb04",
          2333 => x"0b0b0b8d",
          2334 => x"cb040b0b",
          2335 => x"0b8ddb04",
          2336 => x"0b0b0b8d",
          2337 => x"eb040b0b",
          2338 => x"0b8dfb04",
          2339 => x"0b0b0b8e",
          2340 => x"8b040b0b",
          2341 => x"0b8e9b04",
          2342 => x"0b0b0b8e",
          2343 => x"ab040b0b",
          2344 => x"0b8ebb04",
          2345 => x"0b0b0b8e",
          2346 => x"cb040b0b",
          2347 => x"0b8edb04",
          2348 => x"0b0b0b8e",
          2349 => x"eb040b0b",
          2350 => x"0b8efb04",
          2351 => x"0b0b0b8f",
          2352 => x"8b040b0b",
          2353 => x"0b8f9b04",
          2354 => x"0b0b0b8f",
          2355 => x"ab040b0b",
          2356 => x"0b8fbb04",
          2357 => x"0b0b0b8f",
          2358 => x"cb040b0b",
          2359 => x"0b8fdb04",
          2360 => x"0b0b0b8f",
          2361 => x"eb040b0b",
          2362 => x"0b8ffb04",
          2363 => x"0b0b0b90",
          2364 => x"8b040b0b",
          2365 => x"0b909b04",
          2366 => x"0b0b0b90",
          2367 => x"ab040b0b",
          2368 => x"0b90bb04",
          2369 => x"0b0b0b90",
          2370 => x"cb040b0b",
          2371 => x"0b90db04",
          2372 => x"0b0b0b90",
          2373 => x"eb040b0b",
          2374 => x"0b90fb04",
          2375 => x"0b0b0b91",
          2376 => x"8b040b0b",
          2377 => x"0b919b04",
          2378 => x"0b0b0b91",
          2379 => x"ab040b0b",
          2380 => x"0b91bb04",
          2381 => x"0b0b0b91",
          2382 => x"cb040b0b",
          2383 => x"0b91db04",
          2384 => x"0b0b0b91",
          2385 => x"eb040b0b",
          2386 => x"0b91fb04",
          2387 => x"0b0b0b92",
          2388 => x"8b040b0b",
          2389 => x"0b929b04",
          2390 => x"0b0b0b92",
          2391 => x"ab040b0b",
          2392 => x"0b92bb04",
          2393 => x"0b0b0b92",
          2394 => x"cb04ffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0482b5b4",
          2434 => x"0c80f4c6",
          2435 => x"2d82b5b4",
          2436 => x"0882d090",
          2437 => x"0482b5b4",
          2438 => x"0cbed22d",
          2439 => x"82b5b408",
          2440 => x"82d09004",
          2441 => x"82b5b40c",
          2442 => x"bb832d82",
          2443 => x"b5b40882",
          2444 => x"d0900482",
          2445 => x"b5b40cb4",
          2446 => x"fc2d82b5",
          2447 => x"b40882d0",
          2448 => x"900482b5",
          2449 => x"b40c94ab",
          2450 => x"2d82b5b4",
          2451 => x"0882d090",
          2452 => x"0482b5b4",
          2453 => x"0cbce22d",
          2454 => x"82b5b408",
          2455 => x"82d09004",
          2456 => x"82b5b40c",
          2457 => x"b5b22d82",
          2458 => x"b5b40882",
          2459 => x"d0900482",
          2460 => x"b5b40caf",
          2461 => x"ab2d82b5",
          2462 => x"b40882d0",
          2463 => x"900482b5",
          2464 => x"b40c93d6",
          2465 => x"2d82b5b4",
          2466 => x"0882d090",
          2467 => x"0482b5b4",
          2468 => x"0c96be2d",
          2469 => x"82b5b408",
          2470 => x"82d09004",
          2471 => x"82b5b40c",
          2472 => x"97cb2d82",
          2473 => x"b5b40882",
          2474 => x"d0900482",
          2475 => x"b5b40c80",
          2476 => x"f7f02d82",
          2477 => x"b5b40882",
          2478 => x"d0900482",
          2479 => x"b5b40c80",
          2480 => x"f8ce2d82",
          2481 => x"b5b40882",
          2482 => x"d0900482",
          2483 => x"b5b40c80",
          2484 => x"f08a2d82",
          2485 => x"b5b40882",
          2486 => x"d0900482",
          2487 => x"b5b40c80",
          2488 => x"f2822d82",
          2489 => x"b5b40882",
          2490 => x"d0900482",
          2491 => x"b5b40c80",
          2492 => x"f3b52d82",
          2493 => x"b5b40882",
          2494 => x"d0900482",
          2495 => x"b5b40c81",
          2496 => x"d7912d82",
          2497 => x"b5b40882",
          2498 => x"d0900482",
          2499 => x"b5b40c81",
          2500 => x"e4822d82",
          2501 => x"b5b40882",
          2502 => x"d0900482",
          2503 => x"b5b40c81",
          2504 => x"dbf62d82",
          2505 => x"b5b40882",
          2506 => x"d0900482",
          2507 => x"b5b40c81",
          2508 => x"def32d82",
          2509 => x"b5b40882",
          2510 => x"d0900482",
          2511 => x"b5b40c81",
          2512 => x"e9912d82",
          2513 => x"b5b40882",
          2514 => x"d0900482",
          2515 => x"b5b40c81",
          2516 => x"f1f12d82",
          2517 => x"b5b40882",
          2518 => x"d0900482",
          2519 => x"b5b40c81",
          2520 => x"e2e42d82",
          2521 => x"b5b40882",
          2522 => x"d0900482",
          2523 => x"b5b40c81",
          2524 => x"ecb02d82",
          2525 => x"b5b40882",
          2526 => x"d0900482",
          2527 => x"b5b40c81",
          2528 => x"edcf2d82",
          2529 => x"b5b40882",
          2530 => x"d0900482",
          2531 => x"b5b40c81",
          2532 => x"edee2d82",
          2533 => x"b5b40882",
          2534 => x"d0900482",
          2535 => x"b5b40c81",
          2536 => x"f5d82d82",
          2537 => x"b5b40882",
          2538 => x"d0900482",
          2539 => x"b5b40c81",
          2540 => x"f3be2d82",
          2541 => x"b5b40882",
          2542 => x"d0900482",
          2543 => x"b5b40c81",
          2544 => x"f8ac2d82",
          2545 => x"b5b40882",
          2546 => x"d0900482",
          2547 => x"b5b40c81",
          2548 => x"eef22d82",
          2549 => x"b5b40882",
          2550 => x"d0900482",
          2551 => x"b5b40c81",
          2552 => x"fbac2d82",
          2553 => x"b5b40882",
          2554 => x"d0900482",
          2555 => x"b5b40c81",
          2556 => x"fcad2d82",
          2557 => x"b5b40882",
          2558 => x"d0900482",
          2559 => x"b5b40c81",
          2560 => x"e4e22d82",
          2561 => x"b5b40882",
          2562 => x"d0900482",
          2563 => x"b5b40c81",
          2564 => x"e4bb2d82",
          2565 => x"b5b40882",
          2566 => x"d0900482",
          2567 => x"b5b40c81",
          2568 => x"e5e62d82",
          2569 => x"b5b40882",
          2570 => x"d0900482",
          2571 => x"b5b40c81",
          2572 => x"efc92d82",
          2573 => x"b5b40882",
          2574 => x"d0900482",
          2575 => x"b5b40c81",
          2576 => x"fd9e2d82",
          2577 => x"b5b40882",
          2578 => x"d0900482",
          2579 => x"b5b40c81",
          2580 => x"ffa82d82",
          2581 => x"b5b40882",
          2582 => x"d0900482",
          2583 => x"b5b40c82",
          2584 => x"82ea2d82",
          2585 => x"b5b40882",
          2586 => x"d0900482",
          2587 => x"b5b40c81",
          2588 => x"d6b02d82",
          2589 => x"b5b40882",
          2590 => x"d0900482",
          2591 => x"b5b40c82",
          2592 => x"85d62d82",
          2593 => x"b5b40882",
          2594 => x"d0900482",
          2595 => x"b5b40c82",
          2596 => x"948b2d82",
          2597 => x"b5b40882",
          2598 => x"d0900482",
          2599 => x"b5b40c82",
          2600 => x"91f72d82",
          2601 => x"b5b40882",
          2602 => x"d0900482",
          2603 => x"b5b40c81",
          2604 => x"a7eb2d82",
          2605 => x"b5b40882",
          2606 => x"d0900482",
          2607 => x"b5b40c81",
          2608 => x"a9d52d82",
          2609 => x"b5b40882",
          2610 => x"d0900482",
          2611 => x"b5b40c81",
          2612 => x"abb92d82",
          2613 => x"b5b40882",
          2614 => x"d0900482",
          2615 => x"b5b40c80",
          2616 => x"f0b32d82",
          2617 => x"b5b40882",
          2618 => x"d0900482",
          2619 => x"b5b40c80",
          2620 => x"f1d72d82",
          2621 => x"b5b40882",
          2622 => x"d0900482",
          2623 => x"b5b40c80",
          2624 => x"f5bb2d82",
          2625 => x"b5b40882",
          2626 => x"d0900482",
          2627 => x"b5b40c80",
          2628 => x"d6962d82",
          2629 => x"b5b40882",
          2630 => x"d0900482",
          2631 => x"b5b40c81",
          2632 => x"a1ff2d82",
          2633 => x"b5b40882",
          2634 => x"d0900482",
          2635 => x"b5b40c81",
          2636 => x"a2a72d82",
          2637 => x"b5b40882",
          2638 => x"d0900482",
          2639 => x"b5b40c81",
          2640 => x"a69f2d82",
          2641 => x"b5b40882",
          2642 => x"d0900482",
          2643 => x"b5b40c81",
          2644 => x"9ee92d82",
          2645 => x"b5b40882",
          2646 => x"d090043c",
          2647 => x"04000010",
          2648 => x"10101010",
          2649 => x"10101010",
          2650 => x"10101010",
          2651 => x"10101010",
          2652 => x"10101010",
          2653 => x"10101010",
          2654 => x"10101010",
          2655 => x"10105351",
          2656 => x"04000073",
          2657 => x"81ff0673",
          2658 => x"83060981",
          2659 => x"05830510",
          2660 => x"10102b07",
          2661 => x"72fc060c",
          2662 => x"51510472",
          2663 => x"72807281",
          2664 => x"06ff0509",
          2665 => x"72060571",
          2666 => x"1052720a",
          2667 => x"100a5372",
          2668 => x"ed385151",
          2669 => x"53510482",
          2670 => x"b5a87082",
          2671 => x"cd84278e",
          2672 => x"38807170",
          2673 => x"8405530c",
          2674 => x"0b0b0b93",
          2675 => x"ba048c81",
          2676 => x"5180eecb",
          2677 => x"040082b5",
          2678 => x"b4080282",
          2679 => x"b5b40cfb",
          2680 => x"3d0d82b5",
          2681 => x"b4088c05",
          2682 => x"7082b5b4",
          2683 => x"08fc050c",
          2684 => x"82b5b408",
          2685 => x"fc050854",
          2686 => x"82b5b408",
          2687 => x"88050853",
          2688 => x"82ccfc08",
          2689 => x"5254849a",
          2690 => x"3f82b5a8",
          2691 => x"087082b5",
          2692 => x"b408f805",
          2693 => x"0c82b5b4",
          2694 => x"08f80508",
          2695 => x"7082b5a8",
          2696 => x"0c515487",
          2697 => x"3d0d82b5",
          2698 => x"b40c0482",
          2699 => x"b5b40802",
          2700 => x"82b5b40c",
          2701 => x"fb3d0d82",
          2702 => x"b5b40890",
          2703 => x"05088511",
          2704 => x"33708132",
          2705 => x"70810651",
          2706 => x"51515271",
          2707 => x"8f38800b",
          2708 => x"82b5b408",
          2709 => x"8c050825",
          2710 => x"83388d39",
          2711 => x"800b82b5",
          2712 => x"b408f405",
          2713 => x"0c81c439",
          2714 => x"82b5b408",
          2715 => x"8c0508ff",
          2716 => x"0582b5b4",
          2717 => x"088c050c",
          2718 => x"800b82b5",
          2719 => x"b408f805",
          2720 => x"0c82b5b4",
          2721 => x"08880508",
          2722 => x"82b5b408",
          2723 => x"fc050c82",
          2724 => x"b5b408f8",
          2725 => x"05088a2e",
          2726 => x"80f63880",
          2727 => x"0b82b5b4",
          2728 => x"088c0508",
          2729 => x"2580e938",
          2730 => x"82b5b408",
          2731 => x"90050851",
          2732 => x"abb23f82",
          2733 => x"b5a80870",
          2734 => x"82b5b408",
          2735 => x"f8050c52",
          2736 => x"82b5b408",
          2737 => x"f80508ff",
          2738 => x"2e098106",
          2739 => x"8d38800b",
          2740 => x"82b5b408",
          2741 => x"f4050c80",
          2742 => x"d23982b5",
          2743 => x"b408fc05",
          2744 => x"0882b5b4",
          2745 => x"08f80508",
          2746 => x"53537173",
          2747 => x"3482b5b4",
          2748 => x"088c0508",
          2749 => x"ff0582b5",
          2750 => x"b4088c05",
          2751 => x"0c82b5b4",
          2752 => x"08fc0508",
          2753 => x"810582b5",
          2754 => x"b408fc05",
          2755 => x"0cff8039",
          2756 => x"82b5b408",
          2757 => x"fc050852",
          2758 => x"80723482",
          2759 => x"b5b40888",
          2760 => x"05087082",
          2761 => x"b5b408f4",
          2762 => x"050c5282",
          2763 => x"b5b408f4",
          2764 => x"050882b5",
          2765 => x"a80c873d",
          2766 => x"0d82b5b4",
          2767 => x"0c0482b5",
          2768 => x"b4080282",
          2769 => x"b5b40cf4",
          2770 => x"3d0d860b",
          2771 => x"82b5b408",
          2772 => x"e5053482",
          2773 => x"b5b40888",
          2774 => x"050882b5",
          2775 => x"b408e005",
          2776 => x"0cfe0a0b",
          2777 => x"82b5b408",
          2778 => x"e8050c82",
          2779 => x"b5b40890",
          2780 => x"057082b5",
          2781 => x"b408fc05",
          2782 => x"0c82b5b4",
          2783 => x"08fc0508",
          2784 => x"5482b5b4",
          2785 => x"088c0508",
          2786 => x"5382b5b4",
          2787 => x"08e00570",
          2788 => x"53515481",
          2789 => x"8d3f82b5",
          2790 => x"a8087082",
          2791 => x"b5b408dc",
          2792 => x"050c82b5",
          2793 => x"b408ec05",
          2794 => x"0882b5b4",
          2795 => x"08880508",
          2796 => x"05515480",
          2797 => x"743482b5",
          2798 => x"b408dc05",
          2799 => x"087082b5",
          2800 => x"a80c548e",
          2801 => x"3d0d82b5",
          2802 => x"b40c0482",
          2803 => x"b5b40802",
          2804 => x"82b5b40c",
          2805 => x"fb3d0d82",
          2806 => x"b5b40890",
          2807 => x"057082b5",
          2808 => x"b408fc05",
          2809 => x"0c82b5b4",
          2810 => x"08fc0508",
          2811 => x"5482b5b4",
          2812 => x"088c0508",
          2813 => x"5382b5b4",
          2814 => x"08880508",
          2815 => x"5254a33f",
          2816 => x"82b5a808",
          2817 => x"7082b5b4",
          2818 => x"08f8050c",
          2819 => x"82b5b408",
          2820 => x"f8050870",
          2821 => x"82b5a80c",
          2822 => x"5154873d",
          2823 => x"0d82b5b4",
          2824 => x"0c0482b5",
          2825 => x"b4080282",
          2826 => x"b5b40ced",
          2827 => x"3d0d800b",
          2828 => x"82b5b408",
          2829 => x"e4052382",
          2830 => x"b5b40888",
          2831 => x"05085380",
          2832 => x"0b8c140c",
          2833 => x"82b5b408",
          2834 => x"88050885",
          2835 => x"11337081",
          2836 => x"2a708132",
          2837 => x"70810651",
          2838 => x"51515153",
          2839 => x"72802e8d",
          2840 => x"38ff0b82",
          2841 => x"b5b408e0",
          2842 => x"050c96ac",
          2843 => x"3982b5b4",
          2844 => x"088c0508",
          2845 => x"53723353",
          2846 => x"7282b5b4",
          2847 => x"08f80534",
          2848 => x"7281ff06",
          2849 => x"5372802e",
          2850 => x"95fa3882",
          2851 => x"b5b4088c",
          2852 => x"05088105",
          2853 => x"82b5b408",
          2854 => x"8c050c82",
          2855 => x"b5b408e4",
          2856 => x"05227081",
          2857 => x"06515372",
          2858 => x"802e958b",
          2859 => x"3882b5b4",
          2860 => x"08f80533",
          2861 => x"53af7327",
          2862 => x"81fc3882",
          2863 => x"b5b408f8",
          2864 => x"05335372",
          2865 => x"b92681ee",
          2866 => x"3882b5b4",
          2867 => x"08f80533",
          2868 => x"5372b02e",
          2869 => x"09810680",
          2870 => x"c53882b5",
          2871 => x"b408e805",
          2872 => x"3370982b",
          2873 => x"70982c51",
          2874 => x"515372b2",
          2875 => x"3882b5b4",
          2876 => x"08e40522",
          2877 => x"70832a70",
          2878 => x"81327081",
          2879 => x"06515151",
          2880 => x"5372802e",
          2881 => x"993882b5",
          2882 => x"b408e405",
          2883 => x"22708280",
          2884 => x"07515372",
          2885 => x"82b5b408",
          2886 => x"e40523fe",
          2887 => x"d03982b5",
          2888 => x"b408e805",
          2889 => x"3370982b",
          2890 => x"70982c70",
          2891 => x"70832b72",
          2892 => x"11731151",
          2893 => x"51515351",
          2894 => x"55537282",
          2895 => x"b5b408e8",
          2896 => x"053482b5",
          2897 => x"b408e805",
          2898 => x"335482b5",
          2899 => x"b408f805",
          2900 => x"337015d0",
          2901 => x"11515153",
          2902 => x"7282b5b4",
          2903 => x"08e80534",
          2904 => x"82b5b408",
          2905 => x"e8053370",
          2906 => x"982b7098",
          2907 => x"2c515153",
          2908 => x"7280258b",
          2909 => x"3880ff0b",
          2910 => x"82b5b408",
          2911 => x"e8053482",
          2912 => x"b5b408e4",
          2913 => x"05227083",
          2914 => x"2a708106",
          2915 => x"51515372",
          2916 => x"fddb3882",
          2917 => x"b5b408e8",
          2918 => x"05337088",
          2919 => x"2b70902b",
          2920 => x"70902c70",
          2921 => x"882c5151",
          2922 => x"51515372",
          2923 => x"82b5b408",
          2924 => x"ec0523fd",
          2925 => x"b83982b5",
          2926 => x"b408e405",
          2927 => x"2270832a",
          2928 => x"70810651",
          2929 => x"51537280",
          2930 => x"2e9d3882",
          2931 => x"b5b408e8",
          2932 => x"05337098",
          2933 => x"2b70982c",
          2934 => x"51515372",
          2935 => x"8a38810b",
          2936 => x"82b5b408",
          2937 => x"e8053482",
          2938 => x"b5b408f8",
          2939 => x"0533e011",
          2940 => x"82b5b408",
          2941 => x"c4050c53",
          2942 => x"82b5b408",
          2943 => x"c4050880",
          2944 => x"d8269294",
          2945 => x"3882b5b4",
          2946 => x"08c40508",
          2947 => x"70822b82",
          2948 => x"95fc1170",
          2949 => x"08515151",
          2950 => x"53720482",
          2951 => x"b5b408e4",
          2952 => x"05227090",
          2953 => x"07515372",
          2954 => x"82b5b408",
          2955 => x"e4052382",
          2956 => x"b5b408e4",
          2957 => x"052270a0",
          2958 => x"07515372",
          2959 => x"82b5b408",
          2960 => x"e40523fc",
          2961 => x"a83982b5",
          2962 => x"b408e405",
          2963 => x"22708180",
          2964 => x"07515372",
          2965 => x"82b5b408",
          2966 => x"e40523fc",
          2967 => x"903982b5",
          2968 => x"b408e405",
          2969 => x"227080c0",
          2970 => x"07515372",
          2971 => x"82b5b408",
          2972 => x"e40523fb",
          2973 => x"f83982b5",
          2974 => x"b408e405",
          2975 => x"22708807",
          2976 => x"51537282",
          2977 => x"b5b408e4",
          2978 => x"0523800b",
          2979 => x"82b5b408",
          2980 => x"e80534fb",
          2981 => x"d83982b5",
          2982 => x"b408e405",
          2983 => x"22708407",
          2984 => x"51537282",
          2985 => x"b5b408e4",
          2986 => x"0523fbc1",
          2987 => x"39bf0b82",
          2988 => x"b5b408fc",
          2989 => x"053482b5",
          2990 => x"b408ec05",
          2991 => x"22ff1151",
          2992 => x"537282b5",
          2993 => x"b408ec05",
          2994 => x"2380e30b",
          2995 => x"82b5b408",
          2996 => x"f805348d",
          2997 => x"a83982b5",
          2998 => x"b4089005",
          2999 => x"0882b5b4",
          3000 => x"08900508",
          3001 => x"840582b5",
          3002 => x"b4089005",
          3003 => x"0c700851",
          3004 => x"537282b5",
          3005 => x"b408fc05",
          3006 => x"3482b5b4",
          3007 => x"08ec0522",
          3008 => x"ff115153",
          3009 => x"7282b5b4",
          3010 => x"08ec0523",
          3011 => x"8cef3982",
          3012 => x"b5b40890",
          3013 => x"050882b5",
          3014 => x"b4089005",
          3015 => x"08840582",
          3016 => x"b5b40890",
          3017 => x"050c7008",
          3018 => x"82b5b408",
          3019 => x"fc050c82",
          3020 => x"b5b408e4",
          3021 => x"05227083",
          3022 => x"2a708106",
          3023 => x"51515153",
          3024 => x"72802eab",
          3025 => x"3882b5b4",
          3026 => x"08e80533",
          3027 => x"70982b53",
          3028 => x"72982c53",
          3029 => x"82b5b408",
          3030 => x"fc050852",
          3031 => x"53adfa3f",
          3032 => x"82b5a808",
          3033 => x"537282b5",
          3034 => x"b408f405",
          3035 => x"23993982",
          3036 => x"b5b408fc",
          3037 => x"050851a8",
          3038 => x"ac3f82b5",
          3039 => x"a8085372",
          3040 => x"82b5b408",
          3041 => x"f4052382",
          3042 => x"b5b408ec",
          3043 => x"05225382",
          3044 => x"b5b408f4",
          3045 => x"05227371",
          3046 => x"31545472",
          3047 => x"82b5b408",
          3048 => x"ec05238b",
          3049 => x"d83982b5",
          3050 => x"b4089005",
          3051 => x"0882b5b4",
          3052 => x"08900508",
          3053 => x"840582b5",
          3054 => x"b4089005",
          3055 => x"0c700882",
          3056 => x"b5b408fc",
          3057 => x"050c82b5",
          3058 => x"b408e405",
          3059 => x"2270832a",
          3060 => x"70810651",
          3061 => x"51515372",
          3062 => x"802eab38",
          3063 => x"82b5b408",
          3064 => x"e8053370",
          3065 => x"982b5372",
          3066 => x"982c5382",
          3067 => x"b5b408fc",
          3068 => x"05085253",
          3069 => x"ace33f82",
          3070 => x"b5a80853",
          3071 => x"7282b5b4",
          3072 => x"08f40523",
          3073 => x"993982b5",
          3074 => x"b408fc05",
          3075 => x"0851a795",
          3076 => x"3f82b5a8",
          3077 => x"08537282",
          3078 => x"b5b408f4",
          3079 => x"052382b5",
          3080 => x"b408ec05",
          3081 => x"225382b5",
          3082 => x"b408f405",
          3083 => x"22737131",
          3084 => x"54547282",
          3085 => x"b5b408ec",
          3086 => x"05238ac1",
          3087 => x"3982b5b4",
          3088 => x"08e40522",
          3089 => x"70822a70",
          3090 => x"81065151",
          3091 => x"5372802e",
          3092 => x"a43882b5",
          3093 => x"b4089005",
          3094 => x"0882b5b4",
          3095 => x"08900508",
          3096 => x"840582b5",
          3097 => x"b4089005",
          3098 => x"0c700882",
          3099 => x"b5b408dc",
          3100 => x"050c53a2",
          3101 => x"3982b5b4",
          3102 => x"08900508",
          3103 => x"82b5b408",
          3104 => x"90050884",
          3105 => x"0582b5b4",
          3106 => x"0890050c",
          3107 => x"700882b5",
          3108 => x"b408dc05",
          3109 => x"0c5382b5",
          3110 => x"b408dc05",
          3111 => x"0882b5b4",
          3112 => x"08fc050c",
          3113 => x"82b5b408",
          3114 => x"fc050880",
          3115 => x"25a43882",
          3116 => x"b5b408e4",
          3117 => x"05227082",
          3118 => x"07515372",
          3119 => x"82b5b408",
          3120 => x"e4052382",
          3121 => x"b5b408fc",
          3122 => x"05083082",
          3123 => x"b5b408fc",
          3124 => x"050c82b5",
          3125 => x"b408e405",
          3126 => x"2270ffbf",
          3127 => x"06515372",
          3128 => x"82b5b408",
          3129 => x"e4052381",
          3130 => x"af39880b",
          3131 => x"82b5b408",
          3132 => x"f40523a9",
          3133 => x"3982b5b4",
          3134 => x"08e40522",
          3135 => x"7080c007",
          3136 => x"51537282",
          3137 => x"b5b408e4",
          3138 => x"052380f8",
          3139 => x"0b82b5b4",
          3140 => x"08f80534",
          3141 => x"900b82b5",
          3142 => x"b408f405",
          3143 => x"2382b5b4",
          3144 => x"08e40522",
          3145 => x"70822a70",
          3146 => x"81065151",
          3147 => x"5372802e",
          3148 => x"a43882b5",
          3149 => x"b4089005",
          3150 => x"0882b5b4",
          3151 => x"08900508",
          3152 => x"840582b5",
          3153 => x"b4089005",
          3154 => x"0c700882",
          3155 => x"b5b408d8",
          3156 => x"050c53a2",
          3157 => x"3982b5b4",
          3158 => x"08900508",
          3159 => x"82b5b408",
          3160 => x"90050884",
          3161 => x"0582b5b4",
          3162 => x"0890050c",
          3163 => x"700882b5",
          3164 => x"b408d805",
          3165 => x"0c5382b5",
          3166 => x"b408d805",
          3167 => x"0882b5b4",
          3168 => x"08fc050c",
          3169 => x"82b5b408",
          3170 => x"e4052270",
          3171 => x"cf065153",
          3172 => x"7282b5b4",
          3173 => x"08e40523",
          3174 => x"82b5b80b",
          3175 => x"82b5b408",
          3176 => x"f0050c82",
          3177 => x"b5b408f0",
          3178 => x"050882b5",
          3179 => x"b408f405",
          3180 => x"2282b5b4",
          3181 => x"08fc0508",
          3182 => x"71557054",
          3183 => x"565455af",
          3184 => x"953f82b5",
          3185 => x"a8085372",
          3186 => x"753482b5",
          3187 => x"b408f005",
          3188 => x"0882b5b4",
          3189 => x"08d4050c",
          3190 => x"82b5b408",
          3191 => x"f0050870",
          3192 => x"33515389",
          3193 => x"7327a438",
          3194 => x"82b5b408",
          3195 => x"f0050853",
          3196 => x"72335482",
          3197 => x"b5b408f8",
          3198 => x"05337015",
          3199 => x"df115151",
          3200 => x"537282b5",
          3201 => x"b408d005",
          3202 => x"34973982",
          3203 => x"b5b408f0",
          3204 => x"05085372",
          3205 => x"33b01151",
          3206 => x"537282b5",
          3207 => x"b408d005",
          3208 => x"3482b5b4",
          3209 => x"08d40508",
          3210 => x"5382b5b4",
          3211 => x"08d00533",
          3212 => x"733482b5",
          3213 => x"b408f005",
          3214 => x"08810582",
          3215 => x"b5b408f0",
          3216 => x"050c82b5",
          3217 => x"b408f405",
          3218 => x"22705382",
          3219 => x"b5b408fc",
          3220 => x"05085253",
          3221 => x"adcd3f82",
          3222 => x"b5a80870",
          3223 => x"82b5b408",
          3224 => x"fc050c53",
          3225 => x"82b5b408",
          3226 => x"fc050880",
          3227 => x"2e8438fe",
          3228 => x"b23982b5",
          3229 => x"b408f005",
          3230 => x"0882b5b8",
          3231 => x"54557254",
          3232 => x"74707531",
          3233 => x"51537282",
          3234 => x"b5b408fc",
          3235 => x"053482b5",
          3236 => x"b408e405",
          3237 => x"2270b206",
          3238 => x"51537280",
          3239 => x"2e943882",
          3240 => x"b5b408ec",
          3241 => x"0522ff11",
          3242 => x"51537282",
          3243 => x"b5b408ec",
          3244 => x"052382b5",
          3245 => x"b408e405",
          3246 => x"2270862a",
          3247 => x"70810651",
          3248 => x"51537280",
          3249 => x"2e80e738",
          3250 => x"82b5b408",
          3251 => x"ec052270",
          3252 => x"902b82b5",
          3253 => x"b408cc05",
          3254 => x"0c82b5b4",
          3255 => x"08cc0508",
          3256 => x"902c82b5",
          3257 => x"b408cc05",
          3258 => x"0c82b5b4",
          3259 => x"08f40522",
          3260 => x"51537290",
          3261 => x"2e098106",
          3262 => x"953882b5",
          3263 => x"b408cc05",
          3264 => x"08fe0553",
          3265 => x"7282b5b4",
          3266 => x"08c80523",
          3267 => x"933982b5",
          3268 => x"b408cc05",
          3269 => x"08ff0553",
          3270 => x"7282b5b4",
          3271 => x"08c80523",
          3272 => x"82b5b408",
          3273 => x"c8052282",
          3274 => x"b5b408ec",
          3275 => x"052382b5",
          3276 => x"b408e405",
          3277 => x"2270832a",
          3278 => x"70810651",
          3279 => x"51537280",
          3280 => x"2e80d038",
          3281 => x"82b5b408",
          3282 => x"e8053370",
          3283 => x"982b7098",
          3284 => x"2c82b5b4",
          3285 => x"08fc0533",
          3286 => x"57515153",
          3287 => x"72742497",
          3288 => x"3882b5b4",
          3289 => x"08e40522",
          3290 => x"70f70651",
          3291 => x"537282b5",
          3292 => x"b408e405",
          3293 => x"239d3982",
          3294 => x"b5b408e8",
          3295 => x"05335382",
          3296 => x"b5b408fc",
          3297 => x"05337371",
          3298 => x"31545472",
          3299 => x"82b5b408",
          3300 => x"e8053482",
          3301 => x"b5b408e4",
          3302 => x"05227083",
          3303 => x"2a708106",
          3304 => x"51515372",
          3305 => x"802eb138",
          3306 => x"82b5b408",
          3307 => x"e8053370",
          3308 => x"882b7090",
          3309 => x"2b70902c",
          3310 => x"70882c51",
          3311 => x"51515153",
          3312 => x"725482b5",
          3313 => x"b408ec05",
          3314 => x"22707531",
          3315 => x"51537282",
          3316 => x"b5b408ec",
          3317 => x"0523af39",
          3318 => x"82b5b408",
          3319 => x"fc053370",
          3320 => x"882b7090",
          3321 => x"2b70902c",
          3322 => x"70882c51",
          3323 => x"51515153",
          3324 => x"725482b5",
          3325 => x"b408ec05",
          3326 => x"22707531",
          3327 => x"51537282",
          3328 => x"b5b408ec",
          3329 => x"052382b5",
          3330 => x"b408e405",
          3331 => x"22708380",
          3332 => x"06515372",
          3333 => x"b03882b5",
          3334 => x"b408ec05",
          3335 => x"22ff1154",
          3336 => x"547282b5",
          3337 => x"b408ec05",
          3338 => x"2373902b",
          3339 => x"70902c51",
          3340 => x"53807325",
          3341 => x"903882b5",
          3342 => x"b4088805",
          3343 => x"0852a051",
          3344 => x"96903fd2",
          3345 => x"3982b5b4",
          3346 => x"08e40522",
          3347 => x"70812a70",
          3348 => x"81065151",
          3349 => x"5372802e",
          3350 => x"913882b5",
          3351 => x"b4088805",
          3352 => x"0852ad51",
          3353 => x"95ec3f80",
          3354 => x"c73982b5",
          3355 => x"b408e405",
          3356 => x"2270842a",
          3357 => x"70810651",
          3358 => x"51537280",
          3359 => x"2e903882",
          3360 => x"b5b40888",
          3361 => x"050852ab",
          3362 => x"5195c73f",
          3363 => x"a33982b5",
          3364 => x"b408e405",
          3365 => x"2270852a",
          3366 => x"70810651",
          3367 => x"51537280",
          3368 => x"2e8e3882",
          3369 => x"b5b40888",
          3370 => x"050852a0",
          3371 => x"5195a33f",
          3372 => x"82b5b408",
          3373 => x"e4052270",
          3374 => x"862a7081",
          3375 => x"06515153",
          3376 => x"72802eb1",
          3377 => x"3882b5b4",
          3378 => x"08880508",
          3379 => x"52b05195",
          3380 => x"813f82b5",
          3381 => x"b408f405",
          3382 => x"22537290",
          3383 => x"2e098106",
          3384 => x"943882b5",
          3385 => x"b4088805",
          3386 => x"085282b5",
          3387 => x"b408f805",
          3388 => x"335194de",
          3389 => x"3f82b5b4",
          3390 => x"08e40522",
          3391 => x"70882a70",
          3392 => x"81065151",
          3393 => x"5372802e",
          3394 => x"b03882b5",
          3395 => x"b408ec05",
          3396 => x"22ff1154",
          3397 => x"547282b5",
          3398 => x"b408ec05",
          3399 => x"2373902b",
          3400 => x"70902c51",
          3401 => x"53807325",
          3402 => x"903882b5",
          3403 => x"b4088805",
          3404 => x"0852b051",
          3405 => x"949c3fd2",
          3406 => x"3982b5b4",
          3407 => x"08e40522",
          3408 => x"70832a70",
          3409 => x"81065151",
          3410 => x"5372802e",
          3411 => x"b03882b5",
          3412 => x"b408e805",
          3413 => x"33ff1154",
          3414 => x"547282b5",
          3415 => x"b408e805",
          3416 => x"3473982b",
          3417 => x"70982c51",
          3418 => x"53807325",
          3419 => x"903882b5",
          3420 => x"b4088805",
          3421 => x"0852b051",
          3422 => x"93d83fd2",
          3423 => x"3982b5b4",
          3424 => x"08e40522",
          3425 => x"70872a70",
          3426 => x"81065151",
          3427 => x"5372b038",
          3428 => x"82b5b408",
          3429 => x"ec0522ff",
          3430 => x"11545472",
          3431 => x"82b5b408",
          3432 => x"ec052373",
          3433 => x"902b7090",
          3434 => x"2c515380",
          3435 => x"73259038",
          3436 => x"82b5b408",
          3437 => x"88050852",
          3438 => x"a0519396",
          3439 => x"3fd23982",
          3440 => x"b5b408f8",
          3441 => x"05335372",
          3442 => x"80e32e09",
          3443 => x"81069738",
          3444 => x"82b5b408",
          3445 => x"88050852",
          3446 => x"82b5b408",
          3447 => x"fc053351",
          3448 => x"92f03f81",
          3449 => x"ee3982b5",
          3450 => x"b408f805",
          3451 => x"33537280",
          3452 => x"f32e0981",
          3453 => x"0680cb38",
          3454 => x"82b5b408",
          3455 => x"f40522ff",
          3456 => x"11515372",
          3457 => x"82b5b408",
          3458 => x"f4052372",
          3459 => x"83ffff06",
          3460 => x"537283ff",
          3461 => x"ff2e81bb",
          3462 => x"3882b5b4",
          3463 => x"08880508",
          3464 => x"5282b5b4",
          3465 => x"08fc0508",
          3466 => x"70335282",
          3467 => x"b5b408fc",
          3468 => x"05088105",
          3469 => x"82b5b408",
          3470 => x"fc050c53",
          3471 => x"92943fff",
          3472 => x"b73982b5",
          3473 => x"b408f805",
          3474 => x"33537280",
          3475 => x"d32e0981",
          3476 => x"0680cb38",
          3477 => x"82b5b408",
          3478 => x"f40522ff",
          3479 => x"11515372",
          3480 => x"82b5b408",
          3481 => x"f4052372",
          3482 => x"83ffff06",
          3483 => x"537283ff",
          3484 => x"ff2e80df",
          3485 => x"3882b5b4",
          3486 => x"08880508",
          3487 => x"5282b5b4",
          3488 => x"08fc0508",
          3489 => x"70335253",
          3490 => x"91c83f82",
          3491 => x"b5b408fc",
          3492 => x"05088105",
          3493 => x"82b5b408",
          3494 => x"fc050cff",
          3495 => x"b73982b5",
          3496 => x"b408f005",
          3497 => x"0882b5b8",
          3498 => x"2ea93882",
          3499 => x"b5b40888",
          3500 => x"05085282",
          3501 => x"b5b408f0",
          3502 => x"0508ff05",
          3503 => x"82b5b408",
          3504 => x"f0050c82",
          3505 => x"b5b408f0",
          3506 => x"05087033",
          3507 => x"52539182",
          3508 => x"3fcc3982",
          3509 => x"b5b408e4",
          3510 => x"05227087",
          3511 => x"2a708106",
          3512 => x"51515372",
          3513 => x"802e80c3",
          3514 => x"3882b5b4",
          3515 => x"08ec0522",
          3516 => x"ff115454",
          3517 => x"7282b5b4",
          3518 => x"08ec0523",
          3519 => x"73902b70",
          3520 => x"902c5153",
          3521 => x"807325a3",
          3522 => x"3882b5b4",
          3523 => x"08880508",
          3524 => x"52a05190",
          3525 => x"bd3fd239",
          3526 => x"82b5b408",
          3527 => x"88050852",
          3528 => x"82b5b408",
          3529 => x"f8053351",
          3530 => x"90a83f80",
          3531 => x"0b82b5b4",
          3532 => x"08e40523",
          3533 => x"eab73982",
          3534 => x"b5b408f8",
          3535 => x"05335372",
          3536 => x"a52e0981",
          3537 => x"06a83881",
          3538 => x"0b82b5b4",
          3539 => x"08e40523",
          3540 => x"800b82b5",
          3541 => x"b408ec05",
          3542 => x"23800b82",
          3543 => x"b5b408e8",
          3544 => x"05348a0b",
          3545 => x"82b5b408",
          3546 => x"f40523ea",
          3547 => x"803982b5",
          3548 => x"b4088805",
          3549 => x"085282b5",
          3550 => x"b408f805",
          3551 => x"33518fd2",
          3552 => x"3fe9ea39",
          3553 => x"82b5b408",
          3554 => x"8805088c",
          3555 => x"11087082",
          3556 => x"b5b408e0",
          3557 => x"050c5153",
          3558 => x"82b5b408",
          3559 => x"e0050882",
          3560 => x"b5a80c95",
          3561 => x"3d0d82b5",
          3562 => x"b40c0482",
          3563 => x"b5b40802",
          3564 => x"82b5b40c",
          3565 => x"f73d0d80",
          3566 => x"0b82b5b4",
          3567 => x"08f00534",
          3568 => x"82b5b408",
          3569 => x"8c050853",
          3570 => x"80730c82",
          3571 => x"b5b40888",
          3572 => x"05087008",
          3573 => x"51537233",
          3574 => x"537282b5",
          3575 => x"b408f805",
          3576 => x"347281ff",
          3577 => x"065372a0",
          3578 => x"2e098106",
          3579 => x"913882b5",
          3580 => x"b4088805",
          3581 => x"08700881",
          3582 => x"05710c53",
          3583 => x"ce3982b5",
          3584 => x"b408f805",
          3585 => x"335372ad",
          3586 => x"2e098106",
          3587 => x"a438810b",
          3588 => x"82b5b408",
          3589 => x"f0053482",
          3590 => x"b5b40888",
          3591 => x"05087008",
          3592 => x"8105710c",
          3593 => x"70085153",
          3594 => x"723382b5",
          3595 => x"b408f805",
          3596 => x"3482b5b4",
          3597 => x"08f80533",
          3598 => x"5372b02e",
          3599 => x"09810681",
          3600 => x"dc3882b5",
          3601 => x"b4088805",
          3602 => x"08700881",
          3603 => x"05710c70",
          3604 => x"08515372",
          3605 => x"3382b5b4",
          3606 => x"08f80534",
          3607 => x"82b5b408",
          3608 => x"f8053382",
          3609 => x"b5b408e8",
          3610 => x"050c82b5",
          3611 => x"b408e805",
          3612 => x"0880e22e",
          3613 => x"b63882b5",
          3614 => x"b408e805",
          3615 => x"0880f82e",
          3616 => x"843880cd",
          3617 => x"39900b82",
          3618 => x"b5b408f4",
          3619 => x"053482b5",
          3620 => x"b4088805",
          3621 => x"08700881",
          3622 => x"05710c70",
          3623 => x"08515372",
          3624 => x"3382b5b4",
          3625 => x"08f80534",
          3626 => x"81a43982",
          3627 => x"0b82b5b4",
          3628 => x"08f40534",
          3629 => x"82b5b408",
          3630 => x"88050870",
          3631 => x"08810571",
          3632 => x"0c700851",
          3633 => x"53723382",
          3634 => x"b5b408f8",
          3635 => x"053480fe",
          3636 => x"3982b5b4",
          3637 => x"08f80533",
          3638 => x"5372a026",
          3639 => x"8d38810b",
          3640 => x"82b5b408",
          3641 => x"ec050c83",
          3642 => x"803982b5",
          3643 => x"b408f805",
          3644 => x"3353af73",
          3645 => x"27903882",
          3646 => x"b5b408f8",
          3647 => x"05335372",
          3648 => x"b9268338",
          3649 => x"8d39800b",
          3650 => x"82b5b408",
          3651 => x"ec050c82",
          3652 => x"d839880b",
          3653 => x"82b5b408",
          3654 => x"f40534b2",
          3655 => x"3982b5b4",
          3656 => x"08f80533",
          3657 => x"53af7327",
          3658 => x"903882b5",
          3659 => x"b408f805",
          3660 => x"335372b9",
          3661 => x"2683388d",
          3662 => x"39800b82",
          3663 => x"b5b408ec",
          3664 => x"050c82a5",
          3665 => x"398a0b82",
          3666 => x"b5b408f4",
          3667 => x"0534800b",
          3668 => x"82b5b408",
          3669 => x"fc050c82",
          3670 => x"b5b408f8",
          3671 => x"053353a0",
          3672 => x"732781cf",
          3673 => x"3882b5b4",
          3674 => x"08f80533",
          3675 => x"5380e073",
          3676 => x"27943882",
          3677 => x"b5b408f8",
          3678 => x"0533e011",
          3679 => x"51537282",
          3680 => x"b5b408f8",
          3681 => x"053482b5",
          3682 => x"b408f805",
          3683 => x"33d01151",
          3684 => x"537282b5",
          3685 => x"b408f805",
          3686 => x"3482b5b4",
          3687 => x"08f80533",
          3688 => x"53907327",
          3689 => x"ad3882b5",
          3690 => x"b408f805",
          3691 => x"33f91151",
          3692 => x"537282b5",
          3693 => x"b408f805",
          3694 => x"3482b5b4",
          3695 => x"08f80533",
          3696 => x"53728926",
          3697 => x"8d38800b",
          3698 => x"82b5b408",
          3699 => x"ec050c81",
          3700 => x"983982b5",
          3701 => x"b408f805",
          3702 => x"3382b5b4",
          3703 => x"08f40533",
          3704 => x"54547274",
          3705 => x"268d3880",
          3706 => x"0b82b5b4",
          3707 => x"08ec050c",
          3708 => x"80f73982",
          3709 => x"b5b408f4",
          3710 => x"05337082",
          3711 => x"b5b408fc",
          3712 => x"05082982",
          3713 => x"b5b408f8",
          3714 => x"05337012",
          3715 => x"82b5b408",
          3716 => x"fc050c82",
          3717 => x"b5b40888",
          3718 => x"05087008",
          3719 => x"8105710c",
          3720 => x"70085151",
          3721 => x"52555372",
          3722 => x"3382b5b4",
          3723 => x"08f80534",
          3724 => x"fea53982",
          3725 => x"b5b408f0",
          3726 => x"05335372",
          3727 => x"802e9038",
          3728 => x"82b5b408",
          3729 => x"fc050830",
          3730 => x"82b5b408",
          3731 => x"fc050c82",
          3732 => x"b5b4088c",
          3733 => x"050882b5",
          3734 => x"b408fc05",
          3735 => x"08710c53",
          3736 => x"810b82b5",
          3737 => x"b408ec05",
          3738 => x"0c82b5b4",
          3739 => x"08ec0508",
          3740 => x"82b5a80c",
          3741 => x"8b3d0d82",
          3742 => x"b5b40c04",
          3743 => x"82b5b408",
          3744 => x"0282b5b4",
          3745 => x"0cfd3d0d",
          3746 => x"82ccf808",
          3747 => x"5382b5b4",
          3748 => x"088c0508",
          3749 => x"5282b5b4",
          3750 => x"08880508",
          3751 => x"51df8c3f",
          3752 => x"82b5a808",
          3753 => x"7082b5a8",
          3754 => x"0c54853d",
          3755 => x"0d82b5b4",
          3756 => x"0c0482b5",
          3757 => x"b4080282",
          3758 => x"b5b40cf7",
          3759 => x"3d0d800b",
          3760 => x"82b5b408",
          3761 => x"f0053482",
          3762 => x"b5b4088c",
          3763 => x"05085380",
          3764 => x"730c82b5",
          3765 => x"b4088805",
          3766 => x"08700851",
          3767 => x"53723353",
          3768 => x"7282b5b4",
          3769 => x"08f80534",
          3770 => x"7281ff06",
          3771 => x"5372a02e",
          3772 => x"09810691",
          3773 => x"3882b5b4",
          3774 => x"08880508",
          3775 => x"70088105",
          3776 => x"710c53ce",
          3777 => x"3982b5b4",
          3778 => x"08f80533",
          3779 => x"5372ad2e",
          3780 => x"098106a4",
          3781 => x"38810b82",
          3782 => x"b5b408f0",
          3783 => x"053482b5",
          3784 => x"b4088805",
          3785 => x"08700881",
          3786 => x"05710c70",
          3787 => x"08515372",
          3788 => x"3382b5b4",
          3789 => x"08f80534",
          3790 => x"82b5b408",
          3791 => x"f8053353",
          3792 => x"72b02e09",
          3793 => x"810681dc",
          3794 => x"3882b5b4",
          3795 => x"08880508",
          3796 => x"70088105",
          3797 => x"710c7008",
          3798 => x"51537233",
          3799 => x"82b5b408",
          3800 => x"f8053482",
          3801 => x"b5b408f8",
          3802 => x"053382b5",
          3803 => x"b408e805",
          3804 => x"0c82b5b4",
          3805 => x"08e80508",
          3806 => x"80e22eb6",
          3807 => x"3882b5b4",
          3808 => x"08e80508",
          3809 => x"80f82e84",
          3810 => x"3880cd39",
          3811 => x"900b82b5",
          3812 => x"b408f405",
          3813 => x"3482b5b4",
          3814 => x"08880508",
          3815 => x"70088105",
          3816 => x"710c7008",
          3817 => x"51537233",
          3818 => x"82b5b408",
          3819 => x"f8053481",
          3820 => x"a439820b",
          3821 => x"82b5b408",
          3822 => x"f4053482",
          3823 => x"b5b40888",
          3824 => x"05087008",
          3825 => x"8105710c",
          3826 => x"70085153",
          3827 => x"723382b5",
          3828 => x"b408f805",
          3829 => x"3480fe39",
          3830 => x"82b5b408",
          3831 => x"f8053353",
          3832 => x"72a0268d",
          3833 => x"38810b82",
          3834 => x"b5b408ec",
          3835 => x"050c8380",
          3836 => x"3982b5b4",
          3837 => x"08f80533",
          3838 => x"53af7327",
          3839 => x"903882b5",
          3840 => x"b408f805",
          3841 => x"335372b9",
          3842 => x"2683388d",
          3843 => x"39800b82",
          3844 => x"b5b408ec",
          3845 => x"050c82d8",
          3846 => x"39880b82",
          3847 => x"b5b408f4",
          3848 => x"0534b239",
          3849 => x"82b5b408",
          3850 => x"f8053353",
          3851 => x"af732790",
          3852 => x"3882b5b4",
          3853 => x"08f80533",
          3854 => x"5372b926",
          3855 => x"83388d39",
          3856 => x"800b82b5",
          3857 => x"b408ec05",
          3858 => x"0c82a539",
          3859 => x"8a0b82b5",
          3860 => x"b408f405",
          3861 => x"34800b82",
          3862 => x"b5b408fc",
          3863 => x"050c82b5",
          3864 => x"b408f805",
          3865 => x"3353a073",
          3866 => x"2781cf38",
          3867 => x"82b5b408",
          3868 => x"f8053353",
          3869 => x"80e07327",
          3870 => x"943882b5",
          3871 => x"b408f805",
          3872 => x"33e01151",
          3873 => x"537282b5",
          3874 => x"b408f805",
          3875 => x"3482b5b4",
          3876 => x"08f80533",
          3877 => x"d0115153",
          3878 => x"7282b5b4",
          3879 => x"08f80534",
          3880 => x"82b5b408",
          3881 => x"f8053353",
          3882 => x"907327ad",
          3883 => x"3882b5b4",
          3884 => x"08f80533",
          3885 => x"f9115153",
          3886 => x"7282b5b4",
          3887 => x"08f80534",
          3888 => x"82b5b408",
          3889 => x"f8053353",
          3890 => x"7289268d",
          3891 => x"38800b82",
          3892 => x"b5b408ec",
          3893 => x"050c8198",
          3894 => x"3982b5b4",
          3895 => x"08f80533",
          3896 => x"82b5b408",
          3897 => x"f4053354",
          3898 => x"54727426",
          3899 => x"8d38800b",
          3900 => x"82b5b408",
          3901 => x"ec050c80",
          3902 => x"f73982b5",
          3903 => x"b408f405",
          3904 => x"337082b5",
          3905 => x"b408fc05",
          3906 => x"082982b5",
          3907 => x"b408f805",
          3908 => x"33701282",
          3909 => x"b5b408fc",
          3910 => x"050c82b5",
          3911 => x"b4088805",
          3912 => x"08700881",
          3913 => x"05710c70",
          3914 => x"08515152",
          3915 => x"55537233",
          3916 => x"82b5b408",
          3917 => x"f80534fe",
          3918 => x"a53982b5",
          3919 => x"b408f005",
          3920 => x"33537280",
          3921 => x"2e903882",
          3922 => x"b5b408fc",
          3923 => x"05083082",
          3924 => x"b5b408fc",
          3925 => x"050c82b5",
          3926 => x"b4088c05",
          3927 => x"0882b5b4",
          3928 => x"08fc0508",
          3929 => x"710c5381",
          3930 => x"0b82b5b4",
          3931 => x"08ec050c",
          3932 => x"82b5b408",
          3933 => x"ec050882",
          3934 => x"b5a80c8b",
          3935 => x"3d0d82b5",
          3936 => x"b40c0482",
          3937 => x"b5b40802",
          3938 => x"82b5b40c",
          3939 => x"fb3d0d80",
          3940 => x"0b82b5b4",
          3941 => x"08f8050c",
          3942 => x"82ccfc08",
          3943 => x"85113370",
          3944 => x"812a7081",
          3945 => x"32708106",
          3946 => x"51515151",
          3947 => x"5372802e",
          3948 => x"8d38ff0b",
          3949 => x"82b5b408",
          3950 => x"f4050c81",
          3951 => x"923982b5",
          3952 => x"b4088805",
          3953 => x"08537233",
          3954 => x"82b5b408",
          3955 => x"88050881",
          3956 => x"0582b5b4",
          3957 => x"0888050c",
          3958 => x"537282b5",
          3959 => x"b408fc05",
          3960 => x"347281ff",
          3961 => x"06537280",
          3962 => x"2eb03882",
          3963 => x"ccfc0882",
          3964 => x"ccfc0853",
          3965 => x"82b5b408",
          3966 => x"fc053352",
          3967 => x"90110851",
          3968 => x"53722d82",
          3969 => x"b5a80853",
          3970 => x"72802eff",
          3971 => x"b138ff0b",
          3972 => x"82b5b408",
          3973 => x"f8050cff",
          3974 => x"a53982cc",
          3975 => x"fc0882cc",
          3976 => x"fc085353",
          3977 => x"8a519013",
          3978 => x"0853722d",
          3979 => x"82b5a808",
          3980 => x"5372802e",
          3981 => x"8a38ff0b",
          3982 => x"82b5b408",
          3983 => x"f8050c82",
          3984 => x"b5b408f8",
          3985 => x"05087082",
          3986 => x"b5b408f4",
          3987 => x"050c5382",
          3988 => x"b5b408f4",
          3989 => x"050882b5",
          3990 => x"a80c873d",
          3991 => x"0d82b5b4",
          3992 => x"0c0482b5",
          3993 => x"b4080282",
          3994 => x"b5b40cfb",
          3995 => x"3d0d800b",
          3996 => x"82b5b408",
          3997 => x"f8050c82",
          3998 => x"b5b4088c",
          3999 => x"05088511",
          4000 => x"3370812a",
          4001 => x"70813270",
          4002 => x"81065151",
          4003 => x"51515372",
          4004 => x"802e8d38",
          4005 => x"ff0b82b5",
          4006 => x"b408f405",
          4007 => x"0c80f339",
          4008 => x"82b5b408",
          4009 => x"88050853",
          4010 => x"723382b5",
          4011 => x"b4088805",
          4012 => x"08810582",
          4013 => x"b5b40888",
          4014 => x"050c5372",
          4015 => x"82b5b408",
          4016 => x"fc053472",
          4017 => x"81ff0653",
          4018 => x"72802eb6",
          4019 => x"3882b5b4",
          4020 => x"088c0508",
          4021 => x"82b5b408",
          4022 => x"8c050853",
          4023 => x"82b5b408",
          4024 => x"fc053352",
          4025 => x"90110851",
          4026 => x"53722d82",
          4027 => x"b5a80853",
          4028 => x"72802eff",
          4029 => x"ab38ff0b",
          4030 => x"82b5b408",
          4031 => x"f8050cff",
          4032 => x"9f3982b5",
          4033 => x"b408f805",
          4034 => x"087082b5",
          4035 => x"b408f405",
          4036 => x"0c5382b5",
          4037 => x"b408f405",
          4038 => x"0882b5a8",
          4039 => x"0c873d0d",
          4040 => x"82b5b40c",
          4041 => x"0482b5b4",
          4042 => x"080282b5",
          4043 => x"b40cfe3d",
          4044 => x"0d82ccfc",
          4045 => x"085282b5",
          4046 => x"b4088805",
          4047 => x"0851933f",
          4048 => x"82b5a808",
          4049 => x"7082b5a8",
          4050 => x"0c53843d",
          4051 => x"0d82b5b4",
          4052 => x"0c0482b5",
          4053 => x"b4080282",
          4054 => x"b5b40cfb",
          4055 => x"3d0d82b5",
          4056 => x"b4088c05",
          4057 => x"08851133",
          4058 => x"70812a70",
          4059 => x"81327081",
          4060 => x"06515151",
          4061 => x"51537280",
          4062 => x"2e8d38ff",
          4063 => x"0b82b5b4",
          4064 => x"08fc050c",
          4065 => x"81cb3982",
          4066 => x"b5b4088c",
          4067 => x"05088511",
          4068 => x"3370822a",
          4069 => x"70810651",
          4070 => x"51515372",
          4071 => x"802e80db",
          4072 => x"3882b5b4",
          4073 => x"088c0508",
          4074 => x"82b5b408",
          4075 => x"8c050854",
          4076 => x"548c1408",
          4077 => x"88140825",
          4078 => x"9f3882b5",
          4079 => x"b4088c05",
          4080 => x"08700870",
          4081 => x"82b5b408",
          4082 => x"88050852",
          4083 => x"57545472",
          4084 => x"75347308",
          4085 => x"8105740c",
          4086 => x"82b5b408",
          4087 => x"8c05088c",
          4088 => x"11088105",
          4089 => x"8c120c82",
          4090 => x"b5b40888",
          4091 => x"05087082",
          4092 => x"b5b408fc",
          4093 => x"050c5153",
          4094 => x"80d73982",
          4095 => x"b5b4088c",
          4096 => x"050882b5",
          4097 => x"b4088c05",
          4098 => x"085382b5",
          4099 => x"b4088805",
          4100 => x"087081ff",
          4101 => x"06539012",
          4102 => x"08515454",
          4103 => x"722d82b5",
          4104 => x"a8085372",
          4105 => x"a33882b5",
          4106 => x"b4088c05",
          4107 => x"088c1108",
          4108 => x"81058c12",
          4109 => x"0c82b5b4",
          4110 => x"08880508",
          4111 => x"7082b5b4",
          4112 => x"08fc050c",
          4113 => x"51538a39",
          4114 => x"ff0b82b5",
          4115 => x"b408fc05",
          4116 => x"0c82b5b4",
          4117 => x"08fc0508",
          4118 => x"82b5a80c",
          4119 => x"873d0d82",
          4120 => x"b5b40c04",
          4121 => x"82b5b408",
          4122 => x"0282b5b4",
          4123 => x"0cf93d0d",
          4124 => x"82b5b408",
          4125 => x"88050885",
          4126 => x"11337081",
          4127 => x"32708106",
          4128 => x"51515152",
          4129 => x"71802e8d",
          4130 => x"38ff0b82",
          4131 => x"b5b408f8",
          4132 => x"050c8394",
          4133 => x"3982b5b4",
          4134 => x"08880508",
          4135 => x"85113370",
          4136 => x"862a7081",
          4137 => x"06515151",
          4138 => x"5271802e",
          4139 => x"80c53882",
          4140 => x"b5b40888",
          4141 => x"050882b5",
          4142 => x"b4088805",
          4143 => x"08535385",
          4144 => x"123370ff",
          4145 => x"bf065152",
          4146 => x"71851434",
          4147 => x"82b5b408",
          4148 => x"8805088c",
          4149 => x"11088105",
          4150 => x"8c120c82",
          4151 => x"b5b40888",
          4152 => x"05088411",
          4153 => x"337082b5",
          4154 => x"b408f805",
          4155 => x"0c515152",
          4156 => x"82b63982",
          4157 => x"b5b40888",
          4158 => x"05088511",
          4159 => x"3370822a",
          4160 => x"70810651",
          4161 => x"51515271",
          4162 => x"802e80d7",
          4163 => x"3882b5b4",
          4164 => x"08880508",
          4165 => x"70087033",
          4166 => x"82b5b408",
          4167 => x"fc050c51",
          4168 => x"5282b5b4",
          4169 => x"08fc0508",
          4170 => x"a93882b5",
          4171 => x"b4088805",
          4172 => x"0882b5b4",
          4173 => x"08880508",
          4174 => x"53538512",
          4175 => x"3370a007",
          4176 => x"51527185",
          4177 => x"1434ff0b",
          4178 => x"82b5b408",
          4179 => x"f8050c81",
          4180 => x"d73982b5",
          4181 => x"b4088805",
          4182 => x"08700881",
          4183 => x"05710c52",
          4184 => x"81a13982",
          4185 => x"b5b40888",
          4186 => x"050882b5",
          4187 => x"b4088805",
          4188 => x"08529411",
          4189 => x"08515271",
          4190 => x"2d82b5a8",
          4191 => x"087082b5",
          4192 => x"b408fc05",
          4193 => x"0c5282b5",
          4194 => x"b408fc05",
          4195 => x"08802580",
          4196 => x"f23882b5",
          4197 => x"b4088805",
          4198 => x"0882b5b4",
          4199 => x"08f4050c",
          4200 => x"82b5b408",
          4201 => x"88050885",
          4202 => x"113382b5",
          4203 => x"b408f005",
          4204 => x"0c5282b5",
          4205 => x"b408fc05",
          4206 => x"08ff2e09",
          4207 => x"81069538",
          4208 => x"82b5b408",
          4209 => x"f0050890",
          4210 => x"07527182",
          4211 => x"b5b408ec",
          4212 => x"05349339",
          4213 => x"82b5b408",
          4214 => x"f00508a0",
          4215 => x"07527182",
          4216 => x"b5b408ec",
          4217 => x"053482b5",
          4218 => x"b408f405",
          4219 => x"085282b5",
          4220 => x"b408ec05",
          4221 => x"33851334",
          4222 => x"ff0b82b5",
          4223 => x"b408f805",
          4224 => x"0ca63982",
          4225 => x"b5b40888",
          4226 => x"05088c11",
          4227 => x"0881058c",
          4228 => x"120c82b5",
          4229 => x"b408fc05",
          4230 => x"087081ff",
          4231 => x"067082b5",
          4232 => x"b408f805",
          4233 => x"0c515152",
          4234 => x"82b5b408",
          4235 => x"f8050882",
          4236 => x"b5a80c89",
          4237 => x"3d0d82b5",
          4238 => x"b40c0482",
          4239 => x"b5b40802",
          4240 => x"82b5b40c",
          4241 => x"fd3d0d82",
          4242 => x"b5b40888",
          4243 => x"050882b5",
          4244 => x"b408fc05",
          4245 => x"0c82b5b4",
          4246 => x"088c0508",
          4247 => x"82b5b408",
          4248 => x"f8050c82",
          4249 => x"b5b40890",
          4250 => x"0508802e",
          4251 => x"82a23882",
          4252 => x"b5b408f8",
          4253 => x"050882b5",
          4254 => x"b408fc05",
          4255 => x"082681ac",
          4256 => x"3882b5b4",
          4257 => x"08f80508",
          4258 => x"82b5b408",
          4259 => x"90050805",
          4260 => x"5182b5b4",
          4261 => x"08fc0508",
          4262 => x"71278190",
          4263 => x"3882b5b4",
          4264 => x"08fc0508",
          4265 => x"82b5b408",
          4266 => x"90050805",
          4267 => x"82b5b408",
          4268 => x"fc050c82",
          4269 => x"b5b408f8",
          4270 => x"050882b5",
          4271 => x"b4089005",
          4272 => x"080582b5",
          4273 => x"b408f805",
          4274 => x"0c82b5b4",
          4275 => x"08900508",
          4276 => x"810582b5",
          4277 => x"b4089005",
          4278 => x"0c82b5b4",
          4279 => x"08900508",
          4280 => x"ff0582b5",
          4281 => x"b4089005",
          4282 => x"0c82b5b4",
          4283 => x"08900508",
          4284 => x"802e819c",
          4285 => x"3882b5b4",
          4286 => x"08fc0508",
          4287 => x"ff0582b5",
          4288 => x"b408fc05",
          4289 => x"0c82b5b4",
          4290 => x"08f80508",
          4291 => x"ff0582b5",
          4292 => x"b408f805",
          4293 => x"0c82b5b4",
          4294 => x"08fc0508",
          4295 => x"82b5b408",
          4296 => x"f8050853",
          4297 => x"51713371",
          4298 => x"34ffae39",
          4299 => x"82b5b408",
          4300 => x"90050881",
          4301 => x"0582b5b4",
          4302 => x"0890050c",
          4303 => x"82b5b408",
          4304 => x"900508ff",
          4305 => x"0582b5b4",
          4306 => x"0890050c",
          4307 => x"82b5b408",
          4308 => x"90050880",
          4309 => x"2eba3882",
          4310 => x"b5b408f8",
          4311 => x"05085170",
          4312 => x"3382b5b4",
          4313 => x"08f80508",
          4314 => x"810582b5",
          4315 => x"b408f805",
          4316 => x"0c82b5b4",
          4317 => x"08fc0508",
          4318 => x"52527171",
          4319 => x"3482b5b4",
          4320 => x"08fc0508",
          4321 => x"810582b5",
          4322 => x"b408fc05",
          4323 => x"0cffad39",
          4324 => x"82b5b408",
          4325 => x"88050870",
          4326 => x"82b5a80c",
          4327 => x"51853d0d",
          4328 => x"82b5b40c",
          4329 => x"0482b5b4",
          4330 => x"080282b5",
          4331 => x"b40cfe3d",
          4332 => x"0d82b5b4",
          4333 => x"08880508",
          4334 => x"82b5b408",
          4335 => x"fc050c82",
          4336 => x"b5b408fc",
          4337 => x"05085271",
          4338 => x"3382b5b4",
          4339 => x"08fc0508",
          4340 => x"810582b5",
          4341 => x"b408fc05",
          4342 => x"0c7081ff",
          4343 => x"06515170",
          4344 => x"802e8338",
          4345 => x"da3982b5",
          4346 => x"b408fc05",
          4347 => x"08ff0582",
          4348 => x"b5b408fc",
          4349 => x"050c82b5",
          4350 => x"b408fc05",
          4351 => x"0882b5b4",
          4352 => x"08880508",
          4353 => x"317082b5",
          4354 => x"a80c5184",
          4355 => x"3d0d82b5",
          4356 => x"b40c0482",
          4357 => x"b5b40802",
          4358 => x"82b5b40c",
          4359 => x"fe3d0d82",
          4360 => x"b5b40888",
          4361 => x"050882b5",
          4362 => x"b408fc05",
          4363 => x"0c82b5b4",
          4364 => x"088c0508",
          4365 => x"52713382",
          4366 => x"b5b4088c",
          4367 => x"05088105",
          4368 => x"82b5b408",
          4369 => x"8c050c82",
          4370 => x"b5b408fc",
          4371 => x"05085351",
          4372 => x"70723482",
          4373 => x"b5b408fc",
          4374 => x"05088105",
          4375 => x"82b5b408",
          4376 => x"fc050c70",
          4377 => x"81ff0651",
          4378 => x"70802e84",
          4379 => x"38ffbe39",
          4380 => x"82b5b408",
          4381 => x"88050870",
          4382 => x"82b5a80c",
          4383 => x"51843d0d",
          4384 => x"82b5b40c",
          4385 => x"0482b5b4",
          4386 => x"080282b5",
          4387 => x"b40cfd3d",
          4388 => x"0d82b5b4",
          4389 => x"08880508",
          4390 => x"82b5b408",
          4391 => x"fc050c82",
          4392 => x"b5b4088c",
          4393 => x"050882b5",
          4394 => x"b408f805",
          4395 => x"0c82b5b4",
          4396 => x"08900508",
          4397 => x"802e80e5",
          4398 => x"3882b5b4",
          4399 => x"08900508",
          4400 => x"810582b5",
          4401 => x"b4089005",
          4402 => x"0c82b5b4",
          4403 => x"08900508",
          4404 => x"ff0582b5",
          4405 => x"b4089005",
          4406 => x"0c82b5b4",
          4407 => x"08900508",
          4408 => x"802eba38",
          4409 => x"82b5b408",
          4410 => x"f8050851",
          4411 => x"703382b5",
          4412 => x"b408f805",
          4413 => x"08810582",
          4414 => x"b5b408f8",
          4415 => x"050c82b5",
          4416 => x"b408fc05",
          4417 => x"08525271",
          4418 => x"713482b5",
          4419 => x"b408fc05",
          4420 => x"08810582",
          4421 => x"b5b408fc",
          4422 => x"050cffad",
          4423 => x"3982b5b4",
          4424 => x"08880508",
          4425 => x"7082b5a8",
          4426 => x"0c51853d",
          4427 => x"0d82b5b4",
          4428 => x"0c0482b5",
          4429 => x"b4080282",
          4430 => x"b5b40cfd",
          4431 => x"3d0d82b5",
          4432 => x"b4089005",
          4433 => x"08802e81",
          4434 => x"f43882b5",
          4435 => x"b4088c05",
          4436 => x"08527133",
          4437 => x"82b5b408",
          4438 => x"8c050881",
          4439 => x"0582b5b4",
          4440 => x"088c050c",
          4441 => x"82b5b408",
          4442 => x"88050870",
          4443 => x"337281ff",
          4444 => x"06535454",
          4445 => x"5171712e",
          4446 => x"843880ce",
          4447 => x"3982b5b4",
          4448 => x"08880508",
          4449 => x"52713382",
          4450 => x"b5b40888",
          4451 => x"05088105",
          4452 => x"82b5b408",
          4453 => x"88050c70",
          4454 => x"81ff0651",
          4455 => x"51708d38",
          4456 => x"800b82b5",
          4457 => x"b408fc05",
          4458 => x"0c819b39",
          4459 => x"82b5b408",
          4460 => x"900508ff",
          4461 => x"0582b5b4",
          4462 => x"0890050c",
          4463 => x"82b5b408",
          4464 => x"90050880",
          4465 => x"2e8438ff",
          4466 => x"813982b5",
          4467 => x"b4089005",
          4468 => x"08802e80",
          4469 => x"e83882b5",
          4470 => x"b4088805",
          4471 => x"08703352",
          4472 => x"53708d38",
          4473 => x"ff0b82b5",
          4474 => x"b408fc05",
          4475 => x"0c80d739",
          4476 => x"82b5b408",
          4477 => x"8c0508ff",
          4478 => x"0582b5b4",
          4479 => x"088c050c",
          4480 => x"82b5b408",
          4481 => x"8c050870",
          4482 => x"33525270",
          4483 => x"8c38810b",
          4484 => x"82b5b408",
          4485 => x"fc050cae",
          4486 => x"3982b5b4",
          4487 => x"08880508",
          4488 => x"703382b5",
          4489 => x"b4088c05",
          4490 => x"08703372",
          4491 => x"71317082",
          4492 => x"b5b408fc",
          4493 => x"050c5355",
          4494 => x"5252538a",
          4495 => x"39800b82",
          4496 => x"b5b408fc",
          4497 => x"050c82b5",
          4498 => x"b408fc05",
          4499 => x"0882b5a8",
          4500 => x"0c853d0d",
          4501 => x"82b5b40c",
          4502 => x"0482b5b4",
          4503 => x"080282b5",
          4504 => x"b40cfd3d",
          4505 => x"0d82b5b4",
          4506 => x"08880508",
          4507 => x"82b5b408",
          4508 => x"f8050c82",
          4509 => x"b5b4088c",
          4510 => x"05088d38",
          4511 => x"800b82b5",
          4512 => x"b408fc05",
          4513 => x"0c80ec39",
          4514 => x"82b5b408",
          4515 => x"f8050852",
          4516 => x"713382b5",
          4517 => x"b408f805",
          4518 => x"08810582",
          4519 => x"b5b408f8",
          4520 => x"050c7081",
          4521 => x"ff065151",
          4522 => x"70802e9f",
          4523 => x"3882b5b4",
          4524 => x"088c0508",
          4525 => x"ff0582b5",
          4526 => x"b4088c05",
          4527 => x"0c82b5b4",
          4528 => x"088c0508",
          4529 => x"ff2e8438",
          4530 => x"ffbe3982",
          4531 => x"b5b408f8",
          4532 => x"0508ff05",
          4533 => x"82b5b408",
          4534 => x"f8050c82",
          4535 => x"b5b408f8",
          4536 => x"050882b5",
          4537 => x"b4088805",
          4538 => x"08317082",
          4539 => x"b5b408fc",
          4540 => x"050c5182",
          4541 => x"b5b408fc",
          4542 => x"050882b5",
          4543 => x"a80c853d",
          4544 => x"0d82b5b4",
          4545 => x"0c0482b5",
          4546 => x"b4080282",
          4547 => x"b5b40cfe",
          4548 => x"3d0d82b5",
          4549 => x"b4088805",
          4550 => x"0882b5b4",
          4551 => x"08fc050c",
          4552 => x"82b5b408",
          4553 => x"90050880",
          4554 => x"2e80d438",
          4555 => x"82b5b408",
          4556 => x"90050881",
          4557 => x"0582b5b4",
          4558 => x"0890050c",
          4559 => x"82b5b408",
          4560 => x"900508ff",
          4561 => x"0582b5b4",
          4562 => x"0890050c",
          4563 => x"82b5b408",
          4564 => x"90050880",
          4565 => x"2ea93882",
          4566 => x"b5b4088c",
          4567 => x"05085170",
          4568 => x"82b5b408",
          4569 => x"fc050852",
          4570 => x"52717134",
          4571 => x"82b5b408",
          4572 => x"fc050881",
          4573 => x"0582b5b4",
          4574 => x"08fc050c",
          4575 => x"ffbe3982",
          4576 => x"b5b40888",
          4577 => x"05087082",
          4578 => x"b5a80c51",
          4579 => x"843d0d82",
          4580 => x"b5b40c04",
          4581 => x"82b5b408",
          4582 => x"0282b5b4",
          4583 => x"0cf93d0d",
          4584 => x"800b82b5",
          4585 => x"b408fc05",
          4586 => x"0c82b5b4",
          4587 => x"08880508",
          4588 => x"8025b938",
          4589 => x"82b5b408",
          4590 => x"88050830",
          4591 => x"82b5b408",
          4592 => x"88050c80",
          4593 => x"0b82b5b4",
          4594 => x"08f4050c",
          4595 => x"82b5b408",
          4596 => x"fc05088a",
          4597 => x"38810b82",
          4598 => x"b5b408f4",
          4599 => x"050c82b5",
          4600 => x"b408f405",
          4601 => x"0882b5b4",
          4602 => x"08fc050c",
          4603 => x"82b5b408",
          4604 => x"8c050880",
          4605 => x"25b93882",
          4606 => x"b5b4088c",
          4607 => x"05083082",
          4608 => x"b5b4088c",
          4609 => x"050c800b",
          4610 => x"82b5b408",
          4611 => x"f0050c82",
          4612 => x"b5b408fc",
          4613 => x"05088a38",
          4614 => x"810b82b5",
          4615 => x"b408f005",
          4616 => x"0c82b5b4",
          4617 => x"08f00508",
          4618 => x"82b5b408",
          4619 => x"fc050c80",
          4620 => x"5382b5b4",
          4621 => x"088c0508",
          4622 => x"5282b5b4",
          4623 => x"08880508",
          4624 => x"5182c53f",
          4625 => x"82b5a808",
          4626 => x"7082b5b4",
          4627 => x"08f8050c",
          4628 => x"5482b5b4",
          4629 => x"08fc0508",
          4630 => x"802e9038",
          4631 => x"82b5b408",
          4632 => x"f8050830",
          4633 => x"82b5b408",
          4634 => x"f8050c82",
          4635 => x"b5b408f8",
          4636 => x"05087082",
          4637 => x"b5a80c54",
          4638 => x"893d0d82",
          4639 => x"b5b40c04",
          4640 => x"82b5b408",
          4641 => x"0282b5b4",
          4642 => x"0cfb3d0d",
          4643 => x"800b82b5",
          4644 => x"b408fc05",
          4645 => x"0c82b5b4",
          4646 => x"08880508",
          4647 => x"80259938",
          4648 => x"82b5b408",
          4649 => x"88050830",
          4650 => x"82b5b408",
          4651 => x"88050c81",
          4652 => x"0b82b5b4",
          4653 => x"08fc050c",
          4654 => x"82b5b408",
          4655 => x"8c050880",
          4656 => x"25903882",
          4657 => x"b5b4088c",
          4658 => x"05083082",
          4659 => x"b5b4088c",
          4660 => x"050c8153",
          4661 => x"82b5b408",
          4662 => x"8c050852",
          4663 => x"82b5b408",
          4664 => x"88050851",
          4665 => x"81a23f82",
          4666 => x"b5a80870",
          4667 => x"82b5b408",
          4668 => x"f8050c54",
          4669 => x"82b5b408",
          4670 => x"fc050880",
          4671 => x"2e903882",
          4672 => x"b5b408f8",
          4673 => x"05083082",
          4674 => x"b5b408f8",
          4675 => x"050c82b5",
          4676 => x"b408f805",
          4677 => x"087082b5",
          4678 => x"a80c5487",
          4679 => x"3d0d82b5",
          4680 => x"b40c0482",
          4681 => x"b5b40802",
          4682 => x"82b5b40c",
          4683 => x"fd3d0d80",
          4684 => x"5382b5b4",
          4685 => x"088c0508",
          4686 => x"5282b5b4",
          4687 => x"08880508",
          4688 => x"5180c53f",
          4689 => x"82b5a808",
          4690 => x"7082b5a8",
          4691 => x"0c54853d",
          4692 => x"0d82b5b4",
          4693 => x"0c0482b5",
          4694 => x"b4080282",
          4695 => x"b5b40cfd",
          4696 => x"3d0d8153",
          4697 => x"82b5b408",
          4698 => x"8c050852",
          4699 => x"82b5b408",
          4700 => x"88050851",
          4701 => x"933f82b5",
          4702 => x"a8087082",
          4703 => x"b5a80c54",
          4704 => x"853d0d82",
          4705 => x"b5b40c04",
          4706 => x"82b5b408",
          4707 => x"0282b5b4",
          4708 => x"0cfd3d0d",
          4709 => x"810b82b5",
          4710 => x"b408fc05",
          4711 => x"0c800b82",
          4712 => x"b5b408f8",
          4713 => x"050c82b5",
          4714 => x"b4088c05",
          4715 => x"0882b5b4",
          4716 => x"08880508",
          4717 => x"27b93882",
          4718 => x"b5b408fc",
          4719 => x"0508802e",
          4720 => x"ae38800b",
          4721 => x"82b5b408",
          4722 => x"8c050824",
          4723 => x"a23882b5",
          4724 => x"b4088c05",
          4725 => x"081082b5",
          4726 => x"b4088c05",
          4727 => x"0c82b5b4",
          4728 => x"08fc0508",
          4729 => x"1082b5b4",
          4730 => x"08fc050c",
          4731 => x"ffb83982",
          4732 => x"b5b408fc",
          4733 => x"0508802e",
          4734 => x"80e13882",
          4735 => x"b5b4088c",
          4736 => x"050882b5",
          4737 => x"b4088805",
          4738 => x"0826ad38",
          4739 => x"82b5b408",
          4740 => x"88050882",
          4741 => x"b5b4088c",
          4742 => x"05083182",
          4743 => x"b5b40888",
          4744 => x"050c82b5",
          4745 => x"b408f805",
          4746 => x"0882b5b4",
          4747 => x"08fc0508",
          4748 => x"0782b5b4",
          4749 => x"08f8050c",
          4750 => x"82b5b408",
          4751 => x"fc050881",
          4752 => x"2a82b5b4",
          4753 => x"08fc050c",
          4754 => x"82b5b408",
          4755 => x"8c050881",
          4756 => x"2a82b5b4",
          4757 => x"088c050c",
          4758 => x"ff953982",
          4759 => x"b5b40890",
          4760 => x"0508802e",
          4761 => x"933882b5",
          4762 => x"b4088805",
          4763 => x"087082b5",
          4764 => x"b408f405",
          4765 => x"0c519139",
          4766 => x"82b5b408",
          4767 => x"f8050870",
          4768 => x"82b5b408",
          4769 => x"f4050c51",
          4770 => x"82b5b408",
          4771 => x"f4050882",
          4772 => x"b5a80c85",
          4773 => x"3d0d82b5",
          4774 => x"b40c04f9",
          4775 => x"3d0d7970",
          4776 => x"08705656",
          4777 => x"5874802e",
          4778 => x"80e33895",
          4779 => x"39750851",
          4780 => x"f1f33f82",
          4781 => x"b5a80815",
          4782 => x"780c8516",
          4783 => x"335480cd",
          4784 => x"39743354",
          4785 => x"73a02e09",
          4786 => x"81068638",
          4787 => x"811555f1",
          4788 => x"39805776",
          4789 => x"902982b0",
          4790 => x"a8057008",
          4791 => x"5256f1c5",
          4792 => x"3f82b5a8",
          4793 => x"08537452",
          4794 => x"750851f4",
          4795 => x"c53f82b5",
          4796 => x"a8088b38",
          4797 => x"84163354",
          4798 => x"73812eff",
          4799 => x"b0388117",
          4800 => x"7081ff06",
          4801 => x"58549977",
          4802 => x"27c938ff",
          4803 => x"547382b5",
          4804 => x"a80c893d",
          4805 => x"0d04ff3d",
          4806 => x"0d735271",
          4807 => x"9326818e",
          4808 => x"38718429",
          4809 => x"8294c005",
          4810 => x"52710804",
          4811 => x"829a8c51",
          4812 => x"81803982",
          4813 => x"9a985180",
          4814 => x"f939829a",
          4815 => x"ac5180f2",
          4816 => x"39829ac0",
          4817 => x"5180eb39",
          4818 => x"829ad051",
          4819 => x"80e43982",
          4820 => x"9ae05180",
          4821 => x"dd39829a",
          4822 => x"f45180d6",
          4823 => x"39829b84",
          4824 => x"5180cf39",
          4825 => x"829b9c51",
          4826 => x"80c83982",
          4827 => x"9bb45180",
          4828 => x"c139829b",
          4829 => x"cc51bb39",
          4830 => x"829be851",
          4831 => x"b539829b",
          4832 => x"fc51af39",
          4833 => x"829ca851",
          4834 => x"a939829c",
          4835 => x"bc51a339",
          4836 => x"829cdc51",
          4837 => x"9d39829c",
          4838 => x"f0519739",
          4839 => x"829d8851",
          4840 => x"9139829d",
          4841 => x"a0518b39",
          4842 => x"829db851",
          4843 => x"8539829d",
          4844 => x"c451e3cf",
          4845 => x"3f833d0d",
          4846 => x"04fb3d0d",
          4847 => x"77795656",
          4848 => x"7487e726",
          4849 => x"8a387452",
          4850 => x"7587e829",
          4851 => x"51903987",
          4852 => x"e8527451",
          4853 => x"facd3f82",
          4854 => x"b5a80852",
          4855 => x"7551fac3",
          4856 => x"3f82b5a8",
          4857 => x"08547953",
          4858 => x"7552829d",
          4859 => x"d451ffbb",
          4860 => x"e53f873d",
          4861 => x"0d04ec3d",
          4862 => x"0d660284",
          4863 => x"0580e305",
          4864 => x"335b5780",
          4865 => x"68783070",
          4866 => x"7a077325",
          4867 => x"51575959",
          4868 => x"78567787",
          4869 => x"ff268338",
          4870 => x"81567476",
          4871 => x"077081ff",
          4872 => x"06515593",
          4873 => x"56748182",
          4874 => x"38815376",
          4875 => x"528c3d70",
          4876 => x"525680fe",
          4877 => x"dc3f82b5",
          4878 => x"a8085782",
          4879 => x"b5a808b9",
          4880 => x"3882b5a8",
          4881 => x"0887c098",
          4882 => x"880c82b5",
          4883 => x"a8085996",
          4884 => x"3dd40554",
          4885 => x"84805377",
          4886 => x"52755181",
          4887 => x"83983f82",
          4888 => x"b5a80857",
          4889 => x"82b5a808",
          4890 => x"90387a55",
          4891 => x"74802e89",
          4892 => x"38741975",
          4893 => x"195959d7",
          4894 => x"39963dd8",
          4895 => x"0551818b",
          4896 => x"813f7630",
          4897 => x"70780780",
          4898 => x"257b3070",
          4899 => x"9f2a7206",
          4900 => x"51575156",
          4901 => x"74802e90",
          4902 => x"38829df8",
          4903 => x"5387c098",
          4904 => x"88085278",
          4905 => x"51fe923f",
          4906 => x"76567582",
          4907 => x"b5a80c96",
          4908 => x"3d0d04f8",
          4909 => x"3d0d7c02",
          4910 => x"8405b705",
          4911 => x"335859ff",
          4912 => x"5880537b",
          4913 => x"527a51fe",
          4914 => x"ad3f82b5",
          4915 => x"a808a638",
          4916 => x"76802e88",
          4917 => x"3876812e",
          4918 => x"9a389a39",
          4919 => x"62566155",
          4920 => x"605482b5",
          4921 => x"a8537f52",
          4922 => x"7e51782d",
          4923 => x"82b5a808",
          4924 => x"58833978",
          4925 => x"047782b5",
          4926 => x"a80c8a3d",
          4927 => x"0d04f33d",
          4928 => x"0d7f6163",
          4929 => x"028c0580",
          4930 => x"cf053373",
          4931 => x"73156841",
          4932 => x"5f5c5c5e",
          4933 => x"5e5e7a52",
          4934 => x"829e8051",
          4935 => x"ffb9b73f",
          4936 => x"829e8851",
          4937 => x"e0dd3f80",
          4938 => x"55747927",
          4939 => x"80fd387b",
          4940 => x"902e8938",
          4941 => x"7ba02ea6",
          4942 => x"3880c439",
          4943 => x"74185372",
          4944 => x"7a278e38",
          4945 => x"72225282",
          4946 => x"9e8c51ff",
          4947 => x"b9883f88",
          4948 => x"39829e98",
          4949 => x"51e0ac3f",
          4950 => x"82155580",
          4951 => x"c1397418",
          4952 => x"53727a27",
          4953 => x"8e387208",
          4954 => x"52829e80",
          4955 => x"51ffb8e6",
          4956 => x"3f883982",
          4957 => x"9e9451e0",
          4958 => x"8a3f8415",
          4959 => x"55a03974",
          4960 => x"1853727a",
          4961 => x"278e3872",
          4962 => x"3352829e",
          4963 => x"a051ffb8",
          4964 => x"c53f8839",
          4965 => x"829ea851",
          4966 => x"dfe93f81",
          4967 => x"155582cc",
          4968 => x"fc0852a0",
          4969 => x"51e3ab3f",
          4970 => x"feff3982",
          4971 => x"9eac51df",
          4972 => x"d23f8055",
          4973 => x"74792780",
          4974 => x"c6387418",
          4975 => x"70335553",
          4976 => x"8056727a",
          4977 => x"27833881",
          4978 => x"5680539f",
          4979 => x"74278338",
          4980 => x"81537573",
          4981 => x"067081ff",
          4982 => x"06515372",
          4983 => x"802e9038",
          4984 => x"7380fe26",
          4985 => x"8a3882cc",
          4986 => x"fc085273",
          4987 => x"51883982",
          4988 => x"ccfc0852",
          4989 => x"a051e2da",
          4990 => x"3f811555",
          4991 => x"ffb63982",
          4992 => x"9eb051de",
          4993 => x"fe3f7818",
          4994 => x"791c5c58",
          4995 => x"9cc03f82",
          4996 => x"b5a80898",
          4997 => x"2b70982c",
          4998 => x"515776a0",
          4999 => x"2e098106",
          5000 => x"aa389caa",
          5001 => x"3f82b5a8",
          5002 => x"08982b70",
          5003 => x"982c70a0",
          5004 => x"32703072",
          5005 => x"9b327030",
          5006 => x"70720773",
          5007 => x"75070651",
          5008 => x"58585957",
          5009 => x"51578073",
          5010 => x"24d83876",
          5011 => x"9b2e0981",
          5012 => x"06853880",
          5013 => x"538c397c",
          5014 => x"1e537278",
          5015 => x"26fdb738",
          5016 => x"ff537282",
          5017 => x"b5a80c8f",
          5018 => x"3d0d04fc",
          5019 => x"3d0d029b",
          5020 => x"0533829e",
          5021 => x"b453829e",
          5022 => x"b85255ff",
          5023 => x"b6d83f82",
          5024 => x"b4802251",
          5025 => x"a59b3f82",
          5026 => x"9ec45482",
          5027 => x"9ed05382",
          5028 => x"b4813352",
          5029 => x"829ed851",
          5030 => x"ffb6bb3f",
          5031 => x"74802e84",
          5032 => x"38a0cd3f",
          5033 => x"863d0d04",
          5034 => x"fe3d0d87",
          5035 => x"c0968008",
          5036 => x"53a5b73f",
          5037 => x"81519883",
          5038 => x"3f829ef4",
          5039 => x"5199983f",
          5040 => x"805197f7",
          5041 => x"3f72812a",
          5042 => x"70810651",
          5043 => x"5271802e",
          5044 => x"92388151",
          5045 => x"97e53f82",
          5046 => x"9f8c5198",
          5047 => x"fa3f8051",
          5048 => x"97d93f72",
          5049 => x"822a7081",
          5050 => x"06515271",
          5051 => x"802e9238",
          5052 => x"815197c7",
          5053 => x"3f829fa0",
          5054 => x"5198dc3f",
          5055 => x"805197bb",
          5056 => x"3f72832a",
          5057 => x"70810651",
          5058 => x"5271802e",
          5059 => x"92388151",
          5060 => x"97a93f82",
          5061 => x"9fb05198",
          5062 => x"be3f8051",
          5063 => x"979d3f72",
          5064 => x"842a7081",
          5065 => x"06515271",
          5066 => x"802e9238",
          5067 => x"8151978b",
          5068 => x"3f829fc4",
          5069 => x"5198a03f",
          5070 => x"805196ff",
          5071 => x"3f72852a",
          5072 => x"70810651",
          5073 => x"5271802e",
          5074 => x"92388151",
          5075 => x"96ed3f82",
          5076 => x"9fd85198",
          5077 => x"823f8051",
          5078 => x"96e13f72",
          5079 => x"862a7081",
          5080 => x"06515271",
          5081 => x"802e9238",
          5082 => x"815196cf",
          5083 => x"3f829fec",
          5084 => x"5197e43f",
          5085 => x"805196c3",
          5086 => x"3f72872a",
          5087 => x"70810651",
          5088 => x"5271802e",
          5089 => x"92388151",
          5090 => x"96b13f82",
          5091 => x"a0805197",
          5092 => x"c63f8051",
          5093 => x"96a53f72",
          5094 => x"882a7081",
          5095 => x"06515271",
          5096 => x"802e9238",
          5097 => x"81519693",
          5098 => x"3f82a094",
          5099 => x"5197a83f",
          5100 => x"80519687",
          5101 => x"3fa3bb3f",
          5102 => x"843d0d04",
          5103 => x"fb3d0d77",
          5104 => x"028405a3",
          5105 => x"05337055",
          5106 => x"56568052",
          5107 => x"7551eeb6",
          5108 => x"3f0b0b82",
          5109 => x"b0a43354",
          5110 => x"73a93881",
          5111 => x"5382a0d4",
          5112 => x"5282cca8",
          5113 => x"5180f7a9",
          5114 => x"3f82b5a8",
          5115 => x"08307082",
          5116 => x"b5a80807",
          5117 => x"80258271",
          5118 => x"31515154",
          5119 => x"730b0b82",
          5120 => x"b0a4340b",
          5121 => x"0b82b0a4",
          5122 => x"33547381",
          5123 => x"2e098106",
          5124 => x"af3882cc",
          5125 => x"a8537452",
          5126 => x"755181b1",
          5127 => x"da3f82b5",
          5128 => x"a808802e",
          5129 => x"8b3882b5",
          5130 => x"a80851da",
          5131 => x"d63f9139",
          5132 => x"82cca851",
          5133 => x"8183cb3f",
          5134 => x"820b0b0b",
          5135 => x"82b0a434",
          5136 => x"0b0b82b0",
          5137 => x"a4335473",
          5138 => x"822e0981",
          5139 => x"068c3882",
          5140 => x"a0e45374",
          5141 => x"527551a9",
          5142 => x"a23f800b",
          5143 => x"82b5a80c",
          5144 => x"873d0d04",
          5145 => x"cd3d0d80",
          5146 => x"707182cc",
          5147 => x"a40c405e",
          5148 => x"81527d51",
          5149 => x"80c5f53f",
          5150 => x"82b5a808",
          5151 => x"81ff065a",
          5152 => x"797e2e09",
          5153 => x"8106a338",
          5154 => x"973d5a83",
          5155 => x"5382a0ec",
          5156 => x"527951e7",
          5157 => x"f03f7d53",
          5158 => x"795282b6",
          5159 => x"d45180f5",
          5160 => x"8f3f82b5",
          5161 => x"a8087e2e",
          5162 => x"883882a0",
          5163 => x"f0518d95",
          5164 => x"39817040",
          5165 => x"5e82a1a8",
          5166 => x"51d9c83f",
          5167 => x"973d7047",
          5168 => x"5b80f852",
          5169 => x"7a51fdf4",
          5170 => x"3fb53dff",
          5171 => x"840551f3",
          5172 => x"ca3f82b5",
          5173 => x"a808902b",
          5174 => x"70902c51",
          5175 => x"5a7980c2",
          5176 => x"2e879938",
          5177 => x"7980c224",
          5178 => x"b23879bd",
          5179 => x"2e81d138",
          5180 => x"79bd2490",
          5181 => x"3879802e",
          5182 => x"ffbb3879",
          5183 => x"bc2e80da",
          5184 => x"388ac039",
          5185 => x"7980c02e",
          5186 => x"83953879",
          5187 => x"80c02485",
          5188 => x"c93879bf",
          5189 => x"2e828a38",
          5190 => x"8aa93979",
          5191 => x"80f92e89",
          5192 => x"c5387980",
          5193 => x"f9249238",
          5194 => x"7980c32e",
          5195 => x"87fa3879",
          5196 => x"80f82e89",
          5197 => x"8d388a8b",
          5198 => x"39798183",
          5199 => x"2e89f238",
          5200 => x"79818324",
          5201 => x"8b387981",
          5202 => x"822e89d7",
          5203 => x"3889f439",
          5204 => x"7981852e",
          5205 => x"89e73889",
          5206 => x"ea39b53d",
          5207 => x"ff801153",
          5208 => x"ff840551",
          5209 => x"d2cc3f82",
          5210 => x"b5a80880",
          5211 => x"2efec638",
          5212 => x"b53dfefc",
          5213 => x"1153ff84",
          5214 => x"0551d2b6",
          5215 => x"3f82b5a8",
          5216 => x"08802efe",
          5217 => x"b038b53d",
          5218 => x"fef81153",
          5219 => x"ff840551",
          5220 => x"d2a03f82",
          5221 => x"b5a80886",
          5222 => x"3882b5a8",
          5223 => x"084382a1",
          5224 => x"ac51d7df",
          5225 => x"3f64645d",
          5226 => x"5b7a7c27",
          5227 => x"81ea3862",
          5228 => x"5a797b70",
          5229 => x"84055d0c",
          5230 => x"7b7b26f5",
          5231 => x"3881d939",
          5232 => x"b53dff80",
          5233 => x"1153ff84",
          5234 => x"0551d1e6",
          5235 => x"3f82b5a8",
          5236 => x"08802efd",
          5237 => x"e038b53d",
          5238 => x"fefc1153",
          5239 => x"ff840551",
          5240 => x"d1d03f82",
          5241 => x"b5a80880",
          5242 => x"2efdca38",
          5243 => x"b53dfef8",
          5244 => x"1153ff84",
          5245 => x"0551d1ba",
          5246 => x"3f82b5a8",
          5247 => x"08802efd",
          5248 => x"b43882a1",
          5249 => x"bc51d6fb",
          5250 => x"3f645b7a",
          5251 => x"64278188",
          5252 => x"38625a7a",
          5253 => x"7081055c",
          5254 => x"337a3462",
          5255 => x"810543eb",
          5256 => x"39b53dff",
          5257 => x"801153ff",
          5258 => x"840551d1",
          5259 => x"853f82b5",
          5260 => x"a808802e",
          5261 => x"fcff38b5",
          5262 => x"3dfefc11",
          5263 => x"53ff8405",
          5264 => x"51d0ef3f",
          5265 => x"82b5a808",
          5266 => x"802efce9",
          5267 => x"38b53dfe",
          5268 => x"f81153ff",
          5269 => x"840551d0",
          5270 => x"d93f82b5",
          5271 => x"a808802e",
          5272 => x"fcd33882",
          5273 => x"a1c851d6",
          5274 => x"9a3f645b",
          5275 => x"7a6427a8",
          5276 => x"38627033",
          5277 => x"7c335f5b",
          5278 => x"5c797d2e",
          5279 => x"92387955",
          5280 => x"7b547a33",
          5281 => x"537a5282",
          5282 => x"a1d851ff",
          5283 => x"aec83f81",
          5284 => x"1b638105",
          5285 => x"445bd539",
          5286 => x"82a1f051",
          5287 => x"89a739b5",
          5288 => x"3dff8011",
          5289 => x"53ff8405",
          5290 => x"51d0873f",
          5291 => x"82b5a808",
          5292 => x"80df3882",
          5293 => x"b494335a",
          5294 => x"79802e89",
          5295 => x"3882b3cc",
          5296 => x"084580cd",
          5297 => x"3982b495",
          5298 => x"335a7980",
          5299 => x"2e883882",
          5300 => x"b3d40845",
          5301 => x"bc3982b4",
          5302 => x"96335a79",
          5303 => x"802e8838",
          5304 => x"82b3dc08",
          5305 => x"45ab3982",
          5306 => x"b497335a",
          5307 => x"79802e88",
          5308 => x"3882b3e4",
          5309 => x"08459a39",
          5310 => x"82b49233",
          5311 => x"5a79802e",
          5312 => x"883882b3",
          5313 => x"ec084589",
          5314 => x"3982b3fc",
          5315 => x"08fc8005",
          5316 => x"45b53dfe",
          5317 => x"fc1153ff",
          5318 => x"840551cf",
          5319 => x"953f82b5",
          5320 => x"a80880de",
          5321 => x"3882b494",
          5322 => x"335a7980",
          5323 => x"2e893882",
          5324 => x"b3d00844",
          5325 => x"80cc3982",
          5326 => x"b495335a",
          5327 => x"79802e88",
          5328 => x"3882b3d8",
          5329 => x"0844bb39",
          5330 => x"82b49633",
          5331 => x"5a79802e",
          5332 => x"883882b3",
          5333 => x"e00844aa",
          5334 => x"3982b497",
          5335 => x"335a7980",
          5336 => x"2e883882",
          5337 => x"b3e80844",
          5338 => x"993982b4",
          5339 => x"92335a79",
          5340 => x"802e8838",
          5341 => x"82b3f008",
          5342 => x"44883982",
          5343 => x"b3fc0888",
          5344 => x"0544b53d",
          5345 => x"fef81153",
          5346 => x"ff840551",
          5347 => x"cea43f82",
          5348 => x"b5a80880",
          5349 => x"2ea73880",
          5350 => x"635d5d7b",
          5351 => x"882e8338",
          5352 => x"815d7b90",
          5353 => x"32703070",
          5354 => x"72079f2a",
          5355 => x"70600651",
          5356 => x"515b5b79",
          5357 => x"802e8838",
          5358 => x"7ba02e83",
          5359 => x"38884382",
          5360 => x"a1f451d3",
          5361 => x"be3fa055",
          5362 => x"64546253",
          5363 => x"63526451",
          5364 => x"f2ac3f82",
          5365 => x"a2845186",
          5366 => x"ec39b53d",
          5367 => x"ff801153",
          5368 => x"ff840551",
          5369 => x"cdcc3f82",
          5370 => x"b5a80880",
          5371 => x"2ef9c638",
          5372 => x"b53dfefc",
          5373 => x"1153ff84",
          5374 => x"0551cdb6",
          5375 => x"3f82b5a8",
          5376 => x"08802ea4",
          5377 => x"38645a02",
          5378 => x"80cf0533",
          5379 => x"7a346481",
          5380 => x"0545b53d",
          5381 => x"fefc1153",
          5382 => x"ff840551",
          5383 => x"cd943f82",
          5384 => x"b5a808e1",
          5385 => x"38f98e39",
          5386 => x"64703354",
          5387 => x"5282a290",
          5388 => x"51ffaba2",
          5389 => x"3f80f852",
          5390 => x"7a51ccc0",
          5391 => x"3f7a467a",
          5392 => x"335a79ae",
          5393 => x"2ef8ee38",
          5394 => x"9f7a279f",
          5395 => x"38b53dfe",
          5396 => x"fc1153ff",
          5397 => x"840551cc",
          5398 => x"d93f82b5",
          5399 => x"a808802e",
          5400 => x"9138645a",
          5401 => x"0280cf05",
          5402 => x"337a3464",
          5403 => x"810545ff",
          5404 => x"b73982a2",
          5405 => x"9c51d28b",
          5406 => x"3fffad39",
          5407 => x"b53dfef4",
          5408 => x"1153ff84",
          5409 => x"0551c6a3",
          5410 => x"3f82b5a8",
          5411 => x"08802ef8",
          5412 => x"a438b53d",
          5413 => x"fef01153",
          5414 => x"ff840551",
          5415 => x"c68d3f82",
          5416 => x"b5a80880",
          5417 => x"2ea63861",
          5418 => x"5a0280c2",
          5419 => x"05227a70",
          5420 => x"82055c23",
          5421 => x"7942b53d",
          5422 => x"fef01153",
          5423 => x"ff840551",
          5424 => x"c5e93f82",
          5425 => x"b5a808df",
          5426 => x"38f7ea39",
          5427 => x"61702254",
          5428 => x"5282a2a4",
          5429 => x"51ffa9fe",
          5430 => x"3f80f852",
          5431 => x"7a51cb9c",
          5432 => x"3f7a467a",
          5433 => x"335a79ae",
          5434 => x"2ef7ca38",
          5435 => x"799f2687",
          5436 => x"38618205",
          5437 => x"42d639b5",
          5438 => x"3dfef011",
          5439 => x"53ff8405",
          5440 => x"51c5a83f",
          5441 => x"82b5a808",
          5442 => x"802e9338",
          5443 => x"615a0280",
          5444 => x"c205227a",
          5445 => x"7082055c",
          5446 => x"237942ff",
          5447 => x"af3982a2",
          5448 => x"9c51d0df",
          5449 => x"3fffa539",
          5450 => x"b53dfef4",
          5451 => x"1153ff84",
          5452 => x"0551c4f7",
          5453 => x"3f82b5a8",
          5454 => x"08802ef6",
          5455 => x"f838b53d",
          5456 => x"fef01153",
          5457 => x"ff840551",
          5458 => x"c4e13f82",
          5459 => x"b5a80880",
          5460 => x"2ea03861",
          5461 => x"61710c5a",
          5462 => x"61840542",
          5463 => x"b53dfef0",
          5464 => x"1153ff84",
          5465 => x"0551c4c3",
          5466 => x"3f82b5a8",
          5467 => x"08e538f6",
          5468 => x"c4396170",
          5469 => x"08545282",
          5470 => x"a2b051ff",
          5471 => x"a8d83f80",
          5472 => x"f8527a51",
          5473 => x"c9f63f7a",
          5474 => x"467a335a",
          5475 => x"79ae2ef6",
          5476 => x"a4389f7a",
          5477 => x"279b38b5",
          5478 => x"3dfef011",
          5479 => x"53ff8405",
          5480 => x"51c4883f",
          5481 => x"82b5a808",
          5482 => x"802e8d38",
          5483 => x"6161710c",
          5484 => x"5a618405",
          5485 => x"42ffbb39",
          5486 => x"82a29c51",
          5487 => x"cfc53fff",
          5488 => x"b139b53d",
          5489 => x"ff801153",
          5490 => x"ff840551",
          5491 => x"c9e43f82",
          5492 => x"b5a80880",
          5493 => x"2ef5de38",
          5494 => x"645282a2",
          5495 => x"bc51ffa7",
          5496 => x"f53f645a",
          5497 => x"7904b53d",
          5498 => x"ff801153",
          5499 => x"ff840551",
          5500 => x"c9c03f82",
          5501 => x"b5a80880",
          5502 => x"2ef5ba38",
          5503 => x"645282a2",
          5504 => x"d851ffa7",
          5505 => x"d13f645a",
          5506 => x"792d82b5",
          5507 => x"a808802e",
          5508 => x"f5a33882",
          5509 => x"b5a80852",
          5510 => x"82a2f451",
          5511 => x"ffa7b73f",
          5512 => x"f5933982",
          5513 => x"a39051ce",
          5514 => x"da3fffa7",
          5515 => x"8a3ff585",
          5516 => x"3982a3ac",
          5517 => x"51cecc3f",
          5518 => x"805affa8",
          5519 => x"3991b13f",
          5520 => x"f4f3397a",
          5521 => x"467a335a",
          5522 => x"79802ef4",
          5523 => x"e8387e7e",
          5524 => x"065a7980",
          5525 => x"2e81d638",
          5526 => x"b53dff84",
          5527 => x"055183d3",
          5528 => x"3f82b5a8",
          5529 => x"085d815c",
          5530 => x"7b822eb2",
          5531 => x"387b8224",
          5532 => x"89387b81",
          5533 => x"2e8c3880",
          5534 => x"cd397b83",
          5535 => x"2eb03880",
          5536 => x"c53982a3",
          5537 => x"c0567c55",
          5538 => x"82a3c454",
          5539 => x"805382a3",
          5540 => x"c852b53d",
          5541 => x"ffb00551",
          5542 => x"ffa9a33f",
          5543 => x"bb3982a3",
          5544 => x"e852b53d",
          5545 => x"ffb00551",
          5546 => x"ffa9933f",
          5547 => x"ab397c55",
          5548 => x"82a3c454",
          5549 => x"805382a3",
          5550 => x"d852b53d",
          5551 => x"ffb00551",
          5552 => x"ffa8fb3f",
          5553 => x"93397c54",
          5554 => x"805382a3",
          5555 => x"e452b53d",
          5556 => x"ffb00551",
          5557 => x"ffa8e73f",
          5558 => x"82ccf859",
          5559 => x"82b3cc58",
          5560 => x"82b5d857",
          5561 => x"80566555",
          5562 => x"805482d0",
          5563 => x"805382d0",
          5564 => x"8052b53d",
          5565 => x"ffb00551",
          5566 => x"ebb93f82",
          5567 => x"b5a80882",
          5568 => x"b5a80809",
          5569 => x"70307072",
          5570 => x"07802551",
          5571 => x"5c5c4080",
          5572 => x"5b7b8326",
          5573 => x"8338815b",
          5574 => x"797b065a",
          5575 => x"79802e8d",
          5576 => x"38811c70",
          5577 => x"81ff065d",
          5578 => x"5a7bfebc",
          5579 => x"387e8132",
          5580 => x"7e813207",
          5581 => x"5a798a38",
          5582 => x"7fff2e09",
          5583 => x"8106f2f5",
          5584 => x"3882a3ec",
          5585 => x"51ccbc3f",
          5586 => x"f2eb39f5",
          5587 => x"3d0d800b",
          5588 => x"82b5d834",
          5589 => x"87c0948c",
          5590 => x"70085455",
          5591 => x"87848052",
          5592 => x"7251e3bf",
          5593 => x"3f82b5a8",
          5594 => x"08902b75",
          5595 => x"08555387",
          5596 => x"84805273",
          5597 => x"51e3ac3f",
          5598 => x"7282b5a8",
          5599 => x"0807750c",
          5600 => x"87c0949c",
          5601 => x"70085455",
          5602 => x"87848052",
          5603 => x"7251e393",
          5604 => x"3f82b5a8",
          5605 => x"08902b75",
          5606 => x"08555387",
          5607 => x"84805273",
          5608 => x"51e3803f",
          5609 => x"7282b5a8",
          5610 => x"0807750c",
          5611 => x"8c80830b",
          5612 => x"87c09484",
          5613 => x"0c8c8083",
          5614 => x"0b87c094",
          5615 => x"940c82a3",
          5616 => x"fc51cbbf",
          5617 => x"3f80f5d3",
          5618 => x"5a80f8bf",
          5619 => x"5b830284",
          5620 => x"05990534",
          5621 => x"805c8d3d",
          5622 => x"e40582cc",
          5623 => x"fc0c89c4",
          5624 => x"3f93873f",
          5625 => x"82a49051",
          5626 => x"cb993f82",
          5627 => x"a4a451cb",
          5628 => x"923f82a4",
          5629 => x"b051cb8b",
          5630 => x"3f80dda8",
          5631 => x"5192e63f",
          5632 => x"8151ece7",
          5633 => x"3ff0dd3f",
          5634 => x"8004fe3d",
          5635 => x"0d805283",
          5636 => x"5371882b",
          5637 => x"5287d93f",
          5638 => x"82b5a808",
          5639 => x"81ff0672",
          5640 => x"07ff1454",
          5641 => x"52728025",
          5642 => x"e8387182",
          5643 => x"b5a80c84",
          5644 => x"3d0d04fc",
          5645 => x"3d0d7670",
          5646 => x"08545580",
          5647 => x"73525472",
          5648 => x"742e818a",
          5649 => x"38723351",
          5650 => x"70a02e09",
          5651 => x"81068638",
          5652 => x"811353f1",
          5653 => x"39723351",
          5654 => x"70a22e09",
          5655 => x"81068638",
          5656 => x"81135381",
          5657 => x"54725273",
          5658 => x"812e0981",
          5659 => x"069f3884",
          5660 => x"39811252",
          5661 => x"80723352",
          5662 => x"5470a22e",
          5663 => x"83388154",
          5664 => x"70802e9d",
          5665 => x"3873ea38",
          5666 => x"98398112",
          5667 => x"52807233",
          5668 => x"525470a0",
          5669 => x"2e833881",
          5670 => x"5470802e",
          5671 => x"843873ea",
          5672 => x"38807233",
          5673 => x"525470a0",
          5674 => x"2e098106",
          5675 => x"83388154",
          5676 => x"70a23270",
          5677 => x"30708025",
          5678 => x"76075151",
          5679 => x"5170802e",
          5680 => x"88388072",
          5681 => x"70810554",
          5682 => x"3471750c",
          5683 => x"72517082",
          5684 => x"b5a80c86",
          5685 => x"3d0d04fc",
          5686 => x"3d0d7653",
          5687 => x"7208802e",
          5688 => x"9238863d",
          5689 => x"fc055272",
          5690 => x"51ffbdbf",
          5691 => x"3f82b5a8",
          5692 => x"08853880",
          5693 => x"53833974",
          5694 => x"537282b5",
          5695 => x"a80c863d",
          5696 => x"0d04fc3d",
          5697 => x"0d768211",
          5698 => x"33ff0552",
          5699 => x"53815270",
          5700 => x"8b268198",
          5701 => x"38831333",
          5702 => x"ff055182",
          5703 => x"52709e26",
          5704 => x"818a3884",
          5705 => x"13335183",
          5706 => x"52709726",
          5707 => x"80fe3885",
          5708 => x"13335184",
          5709 => x"5270bb26",
          5710 => x"80f23886",
          5711 => x"13335185",
          5712 => x"5270bb26",
          5713 => x"80e63888",
          5714 => x"13225586",
          5715 => x"527487e7",
          5716 => x"2680d938",
          5717 => x"8a132254",
          5718 => x"87527387",
          5719 => x"e72680cc",
          5720 => x"38810b87",
          5721 => x"c0989c0c",
          5722 => x"722287c0",
          5723 => x"98bc0c82",
          5724 => x"133387c0",
          5725 => x"98b80c83",
          5726 => x"133387c0",
          5727 => x"98b40c84",
          5728 => x"133387c0",
          5729 => x"98b00c85",
          5730 => x"133387c0",
          5731 => x"98ac0c86",
          5732 => x"133387c0",
          5733 => x"98a80c74",
          5734 => x"87c098a4",
          5735 => x"0c7387c0",
          5736 => x"98a00c80",
          5737 => x"0b87c098",
          5738 => x"9c0c8052",
          5739 => x"7182b5a8",
          5740 => x"0c863d0d",
          5741 => x"04f33d0d",
          5742 => x"7f5b87c0",
          5743 => x"989c5d81",
          5744 => x"7d0c87c0",
          5745 => x"98bc085e",
          5746 => x"7d7b2387",
          5747 => x"c098b808",
          5748 => x"5a79821c",
          5749 => x"3487c098",
          5750 => x"b4085a79",
          5751 => x"831c3487",
          5752 => x"c098b008",
          5753 => x"5a79841c",
          5754 => x"3487c098",
          5755 => x"ac085a79",
          5756 => x"851c3487",
          5757 => x"c098a808",
          5758 => x"5a79861c",
          5759 => x"3487c098",
          5760 => x"a4085c7b",
          5761 => x"881c2387",
          5762 => x"c098a008",
          5763 => x"5a798a1c",
          5764 => x"23807d0c",
          5765 => x"7983ffff",
          5766 => x"06597b83",
          5767 => x"ffff0658",
          5768 => x"861b3357",
          5769 => x"851b3356",
          5770 => x"841b3355",
          5771 => x"831b3354",
          5772 => x"821b3353",
          5773 => x"7d83ffff",
          5774 => x"065282a4",
          5775 => x"c851ff9f",
          5776 => x"953f8f3d",
          5777 => x"0d04fb3d",
          5778 => x"0d029f05",
          5779 => x"3382b3c8",
          5780 => x"337081ff",
          5781 => x"06585555",
          5782 => x"87c09484",
          5783 => x"5175802e",
          5784 => x"863887c0",
          5785 => x"94945170",
          5786 => x"0870962a",
          5787 => x"70810653",
          5788 => x"54527080",
          5789 => x"2e8c3871",
          5790 => x"912a7081",
          5791 => x"06515170",
          5792 => x"d7387281",
          5793 => x"32708106",
          5794 => x"51517080",
          5795 => x"2e8d3871",
          5796 => x"932a7081",
          5797 => x"06515170",
          5798 => x"ffbe3873",
          5799 => x"81ff0651",
          5800 => x"87c09480",
          5801 => x"5270802e",
          5802 => x"863887c0",
          5803 => x"94905274",
          5804 => x"720c7482",
          5805 => x"b5a80c87",
          5806 => x"3d0d04ff",
          5807 => x"3d0d028f",
          5808 => x"05337030",
          5809 => x"709f2a51",
          5810 => x"52527082",
          5811 => x"b3c83483",
          5812 => x"3d0d04f9",
          5813 => x"3d0d02a7",
          5814 => x"05335877",
          5815 => x"8a2e0981",
          5816 => x"0687387a",
          5817 => x"528d51eb",
          5818 => x"3f82b3c8",
          5819 => x"337081ff",
          5820 => x"06585687",
          5821 => x"c0948453",
          5822 => x"76802e86",
          5823 => x"3887c094",
          5824 => x"94537208",
          5825 => x"70962a70",
          5826 => x"81065556",
          5827 => x"5472802e",
          5828 => x"8c387391",
          5829 => x"2a708106",
          5830 => x"515372d7",
          5831 => x"38748132",
          5832 => x"70810651",
          5833 => x"5372802e",
          5834 => x"8d387393",
          5835 => x"2a708106",
          5836 => x"515372ff",
          5837 => x"be387581",
          5838 => x"ff065387",
          5839 => x"c0948054",
          5840 => x"72802e86",
          5841 => x"3887c094",
          5842 => x"90547774",
          5843 => x"0c800b82",
          5844 => x"b5a80c89",
          5845 => x"3d0d04f9",
          5846 => x"3d0d7954",
          5847 => x"80743370",
          5848 => x"81ff0653",
          5849 => x"53577077",
          5850 => x"2e80fc38",
          5851 => x"7181ff06",
          5852 => x"811582b3",
          5853 => x"c8337081",
          5854 => x"ff065957",
          5855 => x"555887c0",
          5856 => x"94845175",
          5857 => x"802e8638",
          5858 => x"87c09494",
          5859 => x"51700870",
          5860 => x"962a7081",
          5861 => x"06535452",
          5862 => x"70802e8c",
          5863 => x"3871912a",
          5864 => x"70810651",
          5865 => x"5170d738",
          5866 => x"72813270",
          5867 => x"81065151",
          5868 => x"70802e8d",
          5869 => x"3871932a",
          5870 => x"70810651",
          5871 => x"5170ffbe",
          5872 => x"387481ff",
          5873 => x"065187c0",
          5874 => x"94805270",
          5875 => x"802e8638",
          5876 => x"87c09490",
          5877 => x"5277720c",
          5878 => x"81177433",
          5879 => x"7081ff06",
          5880 => x"53535770",
          5881 => x"ff863876",
          5882 => x"82b5a80c",
          5883 => x"893d0d04",
          5884 => x"fe3d0d82",
          5885 => x"b3c83370",
          5886 => x"81ff0654",
          5887 => x"5287c094",
          5888 => x"84517280",
          5889 => x"2e863887",
          5890 => x"c0949451",
          5891 => x"70087082",
          5892 => x"2a708106",
          5893 => x"51515170",
          5894 => x"802ee238",
          5895 => x"7181ff06",
          5896 => x"5187c094",
          5897 => x"80527080",
          5898 => x"2e863887",
          5899 => x"c0949052",
          5900 => x"71087081",
          5901 => x"ff0682b5",
          5902 => x"a80c5184",
          5903 => x"3d0d04ff",
          5904 => x"af3f82b5",
          5905 => x"a80881ff",
          5906 => x"0682b5a8",
          5907 => x"0c04fe3d",
          5908 => x"0d82b3c8",
          5909 => x"337081ff",
          5910 => x"06525387",
          5911 => x"c0948452",
          5912 => x"70802e86",
          5913 => x"3887c094",
          5914 => x"94527108",
          5915 => x"70822a70",
          5916 => x"81065151",
          5917 => x"51ff5270",
          5918 => x"802ea038",
          5919 => x"7281ff06",
          5920 => x"5187c094",
          5921 => x"80527080",
          5922 => x"2e863887",
          5923 => x"c0949052",
          5924 => x"71087098",
          5925 => x"2b70982c",
          5926 => x"51535171",
          5927 => x"82b5a80c",
          5928 => x"843d0d04",
          5929 => x"ff3d0d87",
          5930 => x"c09e8008",
          5931 => x"709c2a8a",
          5932 => x"06515170",
          5933 => x"802e84b4",
          5934 => x"3887c09e",
          5935 => x"a40882b3",
          5936 => x"cc0c87c0",
          5937 => x"9ea80882",
          5938 => x"b3d00c87",
          5939 => x"c09e9408",
          5940 => x"82b3d40c",
          5941 => x"87c09e98",
          5942 => x"0882b3d8",
          5943 => x"0c87c09e",
          5944 => x"9c0882b3",
          5945 => x"dc0c87c0",
          5946 => x"9ea00882",
          5947 => x"b3e00c87",
          5948 => x"c09eac08",
          5949 => x"82b3e40c",
          5950 => x"87c09eb0",
          5951 => x"0882b3e8",
          5952 => x"0c87c09e",
          5953 => x"b40882b3",
          5954 => x"ec0c87c0",
          5955 => x"9eb80882",
          5956 => x"b3f00c87",
          5957 => x"c09ebc08",
          5958 => x"82b3f40c",
          5959 => x"87c09ec0",
          5960 => x"0882b3f8",
          5961 => x"0c87c09e",
          5962 => x"c40882b3",
          5963 => x"fc0c87c0",
          5964 => x"9e800851",
          5965 => x"7082b480",
          5966 => x"2387c09e",
          5967 => x"840882b4",
          5968 => x"840c87c0",
          5969 => x"9e880882",
          5970 => x"b4880c87",
          5971 => x"c09e8c08",
          5972 => x"82b48c0c",
          5973 => x"810b82b4",
          5974 => x"9034800b",
          5975 => x"87c09e90",
          5976 => x"08708480",
          5977 => x"0a065152",
          5978 => x"5270802e",
          5979 => x"83388152",
          5980 => x"7182b491",
          5981 => x"34800b87",
          5982 => x"c09e9008",
          5983 => x"7088800a",
          5984 => x"06515252",
          5985 => x"70802e83",
          5986 => x"38815271",
          5987 => x"82b49234",
          5988 => x"800b87c0",
          5989 => x"9e900870",
          5990 => x"90800a06",
          5991 => x"51525270",
          5992 => x"802e8338",
          5993 => x"81527182",
          5994 => x"b4933480",
          5995 => x"0b87c09e",
          5996 => x"90087088",
          5997 => x"80800651",
          5998 => x"52527080",
          5999 => x"2e833881",
          6000 => x"527182b4",
          6001 => x"9434800b",
          6002 => x"87c09e90",
          6003 => x"0870a080",
          6004 => x"80065152",
          6005 => x"5270802e",
          6006 => x"83388152",
          6007 => x"7182b495",
          6008 => x"34800b87",
          6009 => x"c09e9008",
          6010 => x"70908080",
          6011 => x"06515252",
          6012 => x"70802e83",
          6013 => x"38815271",
          6014 => x"82b49634",
          6015 => x"800b87c0",
          6016 => x"9e900870",
          6017 => x"84808006",
          6018 => x"51525270",
          6019 => x"802e8338",
          6020 => x"81527182",
          6021 => x"b4973480",
          6022 => x"0b87c09e",
          6023 => x"90087082",
          6024 => x"80800651",
          6025 => x"52527080",
          6026 => x"2e833881",
          6027 => x"527182b4",
          6028 => x"9834800b",
          6029 => x"87c09e90",
          6030 => x"08708180",
          6031 => x"80065152",
          6032 => x"5270802e",
          6033 => x"83388152",
          6034 => x"7182b499",
          6035 => x"34800b87",
          6036 => x"c09e9008",
          6037 => x"7080c080",
          6038 => x"06515252",
          6039 => x"70802e83",
          6040 => x"38815271",
          6041 => x"82b49a34",
          6042 => x"800b87c0",
          6043 => x"9e900870",
          6044 => x"a0800651",
          6045 => x"52527080",
          6046 => x"2e833881",
          6047 => x"527182b4",
          6048 => x"9b3487c0",
          6049 => x"9e900870",
          6050 => x"98800670",
          6051 => x"8a2a5151",
          6052 => x"517082b4",
          6053 => x"9c34800b",
          6054 => x"87c09e90",
          6055 => x"08708480",
          6056 => x"06515252",
          6057 => x"70802e83",
          6058 => x"38815271",
          6059 => x"82b49d34",
          6060 => x"87c09e90",
          6061 => x"087083f0",
          6062 => x"0670842a",
          6063 => x"51515170",
          6064 => x"82b49e34",
          6065 => x"800b87c0",
          6066 => x"9e900870",
          6067 => x"88065152",
          6068 => x"5270802e",
          6069 => x"83388152",
          6070 => x"7182b49f",
          6071 => x"3487c09e",
          6072 => x"90087087",
          6073 => x"06515170",
          6074 => x"82b4a034",
          6075 => x"833d0d04",
          6076 => x"fb3d0d82",
          6077 => x"a4e051ff",
          6078 => x"bd893f82",
          6079 => x"b4903354",
          6080 => x"73802e89",
          6081 => x"3882a4f4",
          6082 => x"51ffbcf7",
          6083 => x"3f82a588",
          6084 => x"51ffbcef",
          6085 => x"3f82b492",
          6086 => x"33547380",
          6087 => x"2e943882",
          6088 => x"b3ec0882",
          6089 => x"b3f00811",
          6090 => x"545282a5",
          6091 => x"a051ff95",
          6092 => x"a53f82b4",
          6093 => x"97335473",
          6094 => x"802e9438",
          6095 => x"82b3e408",
          6096 => x"82b3e808",
          6097 => x"11545282",
          6098 => x"a5bc51ff",
          6099 => x"95883f82",
          6100 => x"b4943354",
          6101 => x"73802e94",
          6102 => x"3882b3cc",
          6103 => x"0882b3d0",
          6104 => x"08115452",
          6105 => x"82a5d851",
          6106 => x"ff94eb3f",
          6107 => x"82b49533",
          6108 => x"5473802e",
          6109 => x"943882b3",
          6110 => x"d40882b3",
          6111 => x"d8081154",
          6112 => x"5282a5f4",
          6113 => x"51ff94ce",
          6114 => x"3f82b496",
          6115 => x"33547380",
          6116 => x"2e943882",
          6117 => x"b3dc0882",
          6118 => x"b3e00811",
          6119 => x"545282a6",
          6120 => x"9051ff94",
          6121 => x"b13f82b4",
          6122 => x"9b335473",
          6123 => x"802e8e38",
          6124 => x"82b49c33",
          6125 => x"5282a6ac",
          6126 => x"51ff949a",
          6127 => x"3f82b49f",
          6128 => x"33547380",
          6129 => x"2e8e3882",
          6130 => x"b4a03352",
          6131 => x"82a6cc51",
          6132 => x"ff94833f",
          6133 => x"82b49d33",
          6134 => x"5473802e",
          6135 => x"8e3882b4",
          6136 => x"9e335282",
          6137 => x"a6ec51ff",
          6138 => x"93ec3f82",
          6139 => x"b4913354",
          6140 => x"73802e89",
          6141 => x"3882a78c",
          6142 => x"51ffbb87",
          6143 => x"3f82b493",
          6144 => x"33547380",
          6145 => x"2e893882",
          6146 => x"a7a051ff",
          6147 => x"baf53f82",
          6148 => x"b4983354",
          6149 => x"73802e89",
          6150 => x"3882a7ac",
          6151 => x"51ffbae3",
          6152 => x"3f82b499",
          6153 => x"33547380",
          6154 => x"2e893882",
          6155 => x"a7b851ff",
          6156 => x"bad13f82",
          6157 => x"b49a3354",
          6158 => x"73802e89",
          6159 => x"3882a7c4",
          6160 => x"51ffbabf",
          6161 => x"3f82a7d0",
          6162 => x"51ffbab7",
          6163 => x"3f82b3f4",
          6164 => x"085282a7",
          6165 => x"dc51ff92",
          6166 => x"fd3f82b3",
          6167 => x"f8085282",
          6168 => x"a88451ff",
          6169 => x"92f03f82",
          6170 => x"b3fc0852",
          6171 => x"82a8ac51",
          6172 => x"ff92e33f",
          6173 => x"82a8d451",
          6174 => x"ffba883f",
          6175 => x"82b48022",
          6176 => x"5282a8dc",
          6177 => x"51ff92ce",
          6178 => x"3f82b484",
          6179 => x"0856bd84",
          6180 => x"c0527551",
          6181 => x"d18d3f82",
          6182 => x"b5a808bd",
          6183 => x"84c02976",
          6184 => x"71315454",
          6185 => x"82b5a808",
          6186 => x"5282a984",
          6187 => x"51ff92a6",
          6188 => x"3f82b497",
          6189 => x"33547380",
          6190 => x"2ea93882",
          6191 => x"b4880856",
          6192 => x"bd84c052",
          6193 => x"7551d0db",
          6194 => x"3f82b5a8",
          6195 => x"08bd84c0",
          6196 => x"29767131",
          6197 => x"545482b5",
          6198 => x"a8085282",
          6199 => x"a9b051ff",
          6200 => x"91f43f82",
          6201 => x"b4923354",
          6202 => x"73802ea9",
          6203 => x"3882b48c",
          6204 => x"0856bd84",
          6205 => x"c0527551",
          6206 => x"d0a93f82",
          6207 => x"b5a808bd",
          6208 => x"84c02976",
          6209 => x"71315454",
          6210 => x"82b5a808",
          6211 => x"5282a9dc",
          6212 => x"51ff91c2",
          6213 => x"3f82a1f0",
          6214 => x"51ffb8e7",
          6215 => x"3f873d0d",
          6216 => x"04fe3d0d",
          6217 => x"02920533",
          6218 => x"ff055271",
          6219 => x"8426aa38",
          6220 => x"71842982",
          6221 => x"95900552",
          6222 => x"71080482",
          6223 => x"aa88519d",
          6224 => x"3982aa90",
          6225 => x"51973982",
          6226 => x"aa985191",
          6227 => x"3982aaa0",
          6228 => x"518b3982",
          6229 => x"aaa45185",
          6230 => x"3982aaac",
          6231 => x"51ffb8a3",
          6232 => x"3f843d0d",
          6233 => x"04718880",
          6234 => x"0c04800b",
          6235 => x"87c09684",
          6236 => x"0c0482b4",
          6237 => x"a40887c0",
          6238 => x"96840c04",
          6239 => x"fd3d0d76",
          6240 => x"982b7098",
          6241 => x"2c79982b",
          6242 => x"70982c72",
          6243 => x"10137082",
          6244 => x"2b515351",
          6245 => x"54515180",
          6246 => x"0b82aab8",
          6247 => x"12335553",
          6248 => x"7174259c",
          6249 => x"3882aab4",
          6250 => x"11081202",
          6251 => x"84059705",
          6252 => x"33713352",
          6253 => x"52527072",
          6254 => x"2e098106",
          6255 => x"83388153",
          6256 => x"7282b5a8",
          6257 => x"0c853d0d",
          6258 => x"04fc3d0d",
          6259 => x"78028405",
          6260 => x"9f053371",
          6261 => x"33545553",
          6262 => x"71802ea2",
          6263 => x"388851ff",
          6264 => x"bac33fa0",
          6265 => x"51ffbabd",
          6266 => x"3f8851ff",
          6267 => x"bab73f72",
          6268 => x"33ff0552",
          6269 => x"71733471",
          6270 => x"81ff0652",
          6271 => x"db397651",
          6272 => x"ffb7803f",
          6273 => x"73733486",
          6274 => x"3d0d04f6",
          6275 => x"3d0d7c02",
          6276 => x"8405b705",
          6277 => x"33028805",
          6278 => x"bb053382",
          6279 => x"b5803370",
          6280 => x"842982b4",
          6281 => x"a8057008",
          6282 => x"5159595a",
          6283 => x"58597480",
          6284 => x"2e863874",
          6285 => x"519ab23f",
          6286 => x"82b58033",
          6287 => x"70842982",
          6288 => x"b4a80581",
          6289 => x"19705458",
          6290 => x"565a9db3",
          6291 => x"3f82b5a8",
          6292 => x"08750c82",
          6293 => x"b5803370",
          6294 => x"842982b4",
          6295 => x"a8057008",
          6296 => x"51565a74",
          6297 => x"802ea638",
          6298 => x"75537852",
          6299 => x"7451c495",
          6300 => x"3f82b580",
          6301 => x"33810555",
          6302 => x"7482b580",
          6303 => x"347481ff",
          6304 => x"06559375",
          6305 => x"27873880",
          6306 => x"0b82b580",
          6307 => x"3477802e",
          6308 => x"b63882b4",
          6309 => x"fc085675",
          6310 => x"802eac38",
          6311 => x"82b4f833",
          6312 => x"5574a438",
          6313 => x"8c3dfc05",
          6314 => x"54765378",
          6315 => x"52755180",
          6316 => x"d9c13f82",
          6317 => x"b4fc0852",
          6318 => x"8a51818e",
          6319 => x"ce3f82b4",
          6320 => x"fc085180",
          6321 => x"dd9e3f8c",
          6322 => x"3d0d04fd",
          6323 => x"3d0d82b4",
          6324 => x"a8539354",
          6325 => x"72085271",
          6326 => x"802e8938",
          6327 => x"71519989",
          6328 => x"3f80730c",
          6329 => x"ff148414",
          6330 => x"54547380",
          6331 => x"25e63880",
          6332 => x"0b82b580",
          6333 => x"3482b4fc",
          6334 => x"08527180",
          6335 => x"2e953871",
          6336 => x"5180ddfe",
          6337 => x"3f82b4fc",
          6338 => x"085198dd",
          6339 => x"3f800b82",
          6340 => x"b4fc0c85",
          6341 => x"3d0d04dc",
          6342 => x"3d0d8157",
          6343 => x"805282b4",
          6344 => x"fc085180",
          6345 => x"e2eb3f82",
          6346 => x"b5a80880",
          6347 => x"d23882b4",
          6348 => x"fc085380",
          6349 => x"f852883d",
          6350 => x"70525681",
          6351 => x"8bb93f82",
          6352 => x"b5a80880",
          6353 => x"2eb93875",
          6354 => x"51c0da3f",
          6355 => x"82b5a808",
          6356 => x"55800b82",
          6357 => x"b5a80825",
          6358 => x"9d3882b5",
          6359 => x"a808ff05",
          6360 => x"70175555",
          6361 => x"80743475",
          6362 => x"53765281",
          6363 => x"1782ada8",
          6364 => x"5257ff8c",
          6365 => x"e13f74ff",
          6366 => x"2e098106",
          6367 => x"ffb038a6",
          6368 => x"3d0d04d9",
          6369 => x"3d0daa3d",
          6370 => x"08ad3d08",
          6371 => x"5a5a8170",
          6372 => x"58588052",
          6373 => x"82b4fc08",
          6374 => x"5180e1f5",
          6375 => x"3f82b5a8",
          6376 => x"08819538",
          6377 => x"ff0b82b4",
          6378 => x"fc085455",
          6379 => x"80f8528b",
          6380 => x"3d705256",
          6381 => x"818ac03f",
          6382 => x"82b5a808",
          6383 => x"802ea538",
          6384 => x"7551ffbf",
          6385 => x"e03f82b5",
          6386 => x"a8088118",
          6387 => x"5855800b",
          6388 => x"82b5a808",
          6389 => x"258e3882",
          6390 => x"b5a808ff",
          6391 => x"05701755",
          6392 => x"55807434",
          6393 => x"74097030",
          6394 => x"7072079f",
          6395 => x"2a515555",
          6396 => x"78772e85",
          6397 => x"3873ffac",
          6398 => x"3882b4fc",
          6399 => x"088c1108",
          6400 => x"535180e1",
          6401 => x"8c3f82b5",
          6402 => x"a808802e",
          6403 => x"893882ad",
          6404 => x"b451ffb2",
          6405 => x"ee3f7877",
          6406 => x"2e098106",
          6407 => x"9b387552",
          6408 => x"7951ffbf",
          6409 => x"ee3f7951",
          6410 => x"ffbefa3f",
          6411 => x"ab3d0854",
          6412 => x"82b5a808",
          6413 => x"74348058",
          6414 => x"7782b5a8",
          6415 => x"0ca93d0d",
          6416 => x"04f63d0d",
          6417 => x"7c7e715c",
          6418 => x"71723357",
          6419 => x"595a5873",
          6420 => x"a02e0981",
          6421 => x"06a23878",
          6422 => x"33780556",
          6423 => x"77762798",
          6424 => x"38811770",
          6425 => x"5b707133",
          6426 => x"56585573",
          6427 => x"a02e0981",
          6428 => x"06863875",
          6429 => x"7526ea38",
          6430 => x"80547388",
          6431 => x"2982b584",
          6432 => x"05700852",
          6433 => x"55ffbe9d",
          6434 => x"3f82b5a8",
          6435 => x"08537952",
          6436 => x"740851c1",
          6437 => x"9d3f82b5",
          6438 => x"a80880c6",
          6439 => x"38841533",
          6440 => x"5574812e",
          6441 => x"88387482",
          6442 => x"2e8838b6",
          6443 => x"39fce83f",
          6444 => x"ad39811a",
          6445 => x"5a8c3dfc",
          6446 => x"1153f805",
          6447 => x"51ffabf2",
          6448 => x"3f82b5a8",
          6449 => x"08802e9a",
          6450 => x"38ff1b53",
          6451 => x"78527751",
          6452 => x"fdb13f82",
          6453 => x"b5a80881",
          6454 => x"ff065574",
          6455 => x"85387454",
          6456 => x"91398114",
          6457 => x"7081ff06",
          6458 => x"51548274",
          6459 => x"27ff8b38",
          6460 => x"80547382",
          6461 => x"b5a80c8c",
          6462 => x"3d0d04d3",
          6463 => x"3d0db03d",
          6464 => x"08b23d08",
          6465 => x"b43d0859",
          6466 => x"5f5a800b",
          6467 => x"af3d3482",
          6468 => x"b5803382",
          6469 => x"b4fc0855",
          6470 => x"5b7381cb",
          6471 => x"387382b4",
          6472 => x"f8335555",
          6473 => x"73833881",
          6474 => x"5576802e",
          6475 => x"81bc3881",
          6476 => x"70760655",
          6477 => x"5673802e",
          6478 => x"81ad38a8",
          6479 => x"5197c03f",
          6480 => x"82b5a808",
          6481 => x"82b4fc0c",
          6482 => x"82b5a808",
          6483 => x"802e8192",
          6484 => x"38935376",
          6485 => x"5282b5a8",
          6486 => x"085180cc",
          6487 => x"b43f82b5",
          6488 => x"a808802e",
          6489 => x"8c3882ad",
          6490 => x"e051ffb0",
          6491 => x"963f80f7",
          6492 => x"3982b5a8",
          6493 => x"085b82b4",
          6494 => x"fc085380",
          6495 => x"f852903d",
          6496 => x"70525481",
          6497 => x"86f13f82",
          6498 => x"b5a80856",
          6499 => x"82b5a808",
          6500 => x"742e0981",
          6501 => x"0680d038",
          6502 => x"82b5a808",
          6503 => x"51ffbc85",
          6504 => x"3f82b5a8",
          6505 => x"0855800b",
          6506 => x"82b5a808",
          6507 => x"25a93882",
          6508 => x"b5a808ff",
          6509 => x"05701755",
          6510 => x"55807434",
          6511 => x"80537481",
          6512 => x"ff065275",
          6513 => x"51f8c43f",
          6514 => x"811b7081",
          6515 => x"ff065c54",
          6516 => x"937b2783",
          6517 => x"38805b74",
          6518 => x"ff2e0981",
          6519 => x"06ff9738",
          6520 => x"86397582",
          6521 => x"b4f83476",
          6522 => x"8c3882b4",
          6523 => x"fc08802e",
          6524 => x"8438f9d7",
          6525 => x"3f8f3d5d",
          6526 => x"ecd43f82",
          6527 => x"b5a80898",
          6528 => x"2b70982c",
          6529 => x"515978ff",
          6530 => x"2eee3878",
          6531 => x"81ff0682",
          6532 => x"ccd43370",
          6533 => x"982b7098",
          6534 => x"2c82ccd0",
          6535 => x"3370982b",
          6536 => x"70972c71",
          6537 => x"982c0570",
          6538 => x"842982aa",
          6539 => x"b4057008",
          6540 => x"15703351",
          6541 => x"51515159",
          6542 => x"5951595d",
          6543 => x"58815673",
          6544 => x"782e80e9",
          6545 => x"38777427",
          6546 => x"b4387481",
          6547 => x"800a2981",
          6548 => x"ff0a0570",
          6549 => x"982c5155",
          6550 => x"80752480",
          6551 => x"ce387653",
          6552 => x"74527751",
          6553 => x"f6963f82",
          6554 => x"b5a80881",
          6555 => x"ff065473",
          6556 => x"802ed738",
          6557 => x"7482ccd0",
          6558 => x"348156b1",
          6559 => x"39748180",
          6560 => x"0a298180",
          6561 => x"0a057098",
          6562 => x"2c7081ff",
          6563 => x"06565155",
          6564 => x"73952697",
          6565 => x"38765374",
          6566 => x"527751f5",
          6567 => x"df3f82b5",
          6568 => x"a80881ff",
          6569 => x"065473cc",
          6570 => x"38d33980",
          6571 => x"5675802e",
          6572 => x"80ca3881",
          6573 => x"1c557482",
          6574 => x"ccd43474",
          6575 => x"982b7098",
          6576 => x"2c82ccd0",
          6577 => x"3370982b",
          6578 => x"70982c70",
          6579 => x"10117082",
          6580 => x"2b82aab8",
          6581 => x"11335e51",
          6582 => x"51515758",
          6583 => x"51557477",
          6584 => x"2e098106",
          6585 => x"fe923882",
          6586 => x"aabc1408",
          6587 => x"7d0c800b",
          6588 => x"82ccd434",
          6589 => x"800b82cc",
          6590 => x"d0349239",
          6591 => x"7582ccd4",
          6592 => x"347582cc",
          6593 => x"d03478af",
          6594 => x"3d34757d",
          6595 => x"0c7e5473",
          6596 => x"9526fde1",
          6597 => x"38738429",
          6598 => x"8295a405",
          6599 => x"54730804",
          6600 => x"82ccdc33",
          6601 => x"54737e2e",
          6602 => x"fdcb3882",
          6603 => x"ccd83355",
          6604 => x"737527ab",
          6605 => x"3874982b",
          6606 => x"70982c51",
          6607 => x"55737524",
          6608 => x"9e38741a",
          6609 => x"54733381",
          6610 => x"15347481",
          6611 => x"800a2981",
          6612 => x"ff0a0570",
          6613 => x"982c82cc",
          6614 => x"dc335651",
          6615 => x"55df3982",
          6616 => x"ccdc3381",
          6617 => x"11565474",
          6618 => x"82ccdc34",
          6619 => x"731a54ae",
          6620 => x"3d337434",
          6621 => x"82ccd833",
          6622 => x"54737e25",
          6623 => x"89388114",
          6624 => x"547382cc",
          6625 => x"d83482cc",
          6626 => x"dc337081",
          6627 => x"800a2981",
          6628 => x"ff0a0570",
          6629 => x"982c82cc",
          6630 => x"d8335a51",
          6631 => x"56567477",
          6632 => x"25a33874",
          6633 => x"1a703352",
          6634 => x"54ffaef9",
          6635 => x"3f748180",
          6636 => x"0a298180",
          6637 => x"0a057098",
          6638 => x"2c82ccd8",
          6639 => x"33565155",
          6640 => x"737524df",
          6641 => x"3882ccdc",
          6642 => x"3370982b",
          6643 => x"70982c82",
          6644 => x"ccd8335a",
          6645 => x"51565674",
          6646 => x"7725fc99",
          6647 => x"388851ff",
          6648 => x"aec33f74",
          6649 => x"81800a29",
          6650 => x"81800a05",
          6651 => x"70982c82",
          6652 => x"ccd83356",
          6653 => x"51557375",
          6654 => x"24e338fb",
          6655 => x"f839837a",
          6656 => x"34800b81",
          6657 => x"1b3482cc",
          6658 => x"dc538052",
          6659 => x"82a2f051",
          6660 => x"f3b73f81",
          6661 => x"e43982cc",
          6662 => x"dc337081",
          6663 => x"ff065555",
          6664 => x"73802efb",
          6665 => x"d03882cc",
          6666 => x"d833ff05",
          6667 => x"547382cc",
          6668 => x"d834ff15",
          6669 => x"547382cc",
          6670 => x"dc348851",
          6671 => x"ffade63f",
          6672 => x"82ccdc33",
          6673 => x"70982b70",
          6674 => x"982c82cc",
          6675 => x"d8335751",
          6676 => x"56577474",
          6677 => x"25a83874",
          6678 => x"1a548114",
          6679 => x"33743473",
          6680 => x"3351ffad",
          6681 => x"c03f7481",
          6682 => x"800a2981",
          6683 => x"800a0570",
          6684 => x"982c82cc",
          6685 => x"d8335851",
          6686 => x"55757524",
          6687 => x"da38a051",
          6688 => x"ffada23f",
          6689 => x"82ccdc33",
          6690 => x"70982b70",
          6691 => x"982c82cc",
          6692 => x"d8335751",
          6693 => x"56577474",
          6694 => x"24fada38",
          6695 => x"8851ffad",
          6696 => x"843f7481",
          6697 => x"800a2981",
          6698 => x"800a0570",
          6699 => x"982c82cc",
          6700 => x"d8335851",
          6701 => x"55757525",
          6702 => x"e338fab9",
          6703 => x"3982ccd8",
          6704 => x"337a0554",
          6705 => x"8074348a",
          6706 => x"51ffacd9",
          6707 => x"3f82ccd8",
          6708 => x"527951f6",
          6709 => x"ec3f82b5",
          6710 => x"a80881ff",
          6711 => x"06547396",
          6712 => x"3882ccd8",
          6713 => x"33547380",
          6714 => x"2e8f3881",
          6715 => x"53735279",
          6716 => x"51f2983f",
          6717 => x"8439807a",
          6718 => x"34800b82",
          6719 => x"ccdc3480",
          6720 => x"0b82ccd8",
          6721 => x"347982b5",
          6722 => x"a80caf3d",
          6723 => x"0d0482cc",
          6724 => x"dc335473",
          6725 => x"802ef9dd",
          6726 => x"388851ff",
          6727 => x"ac873f82",
          6728 => x"ccdc33ff",
          6729 => x"05547382",
          6730 => x"ccdc3473",
          6731 => x"81ff0654",
          6732 => x"e23982cc",
          6733 => x"dc3382cc",
          6734 => x"d8335555",
          6735 => x"73752ef9",
          6736 => x"b438ff14",
          6737 => x"547382cc",
          6738 => x"d8347498",
          6739 => x"2b70982c",
          6740 => x"7581ff06",
          6741 => x"56515574",
          6742 => x"7425a838",
          6743 => x"741a5481",
          6744 => x"14337434",
          6745 => x"733351ff",
          6746 => x"abbb3f74",
          6747 => x"81800a29",
          6748 => x"81800a05",
          6749 => x"70982c82",
          6750 => x"ccd83358",
          6751 => x"51557575",
          6752 => x"24da38a0",
          6753 => x"51ffab9d",
          6754 => x"3f82ccdc",
          6755 => x"3370982b",
          6756 => x"70982c82",
          6757 => x"ccd83357",
          6758 => x"51565774",
          6759 => x"7424f8d5",
          6760 => x"388851ff",
          6761 => x"aaff3f74",
          6762 => x"81800a29",
          6763 => x"81800a05",
          6764 => x"70982c82",
          6765 => x"ccd83358",
          6766 => x"51557575",
          6767 => x"25e338f8",
          6768 => x"b43982cc",
          6769 => x"dc337081",
          6770 => x"ff0682cc",
          6771 => x"d8335956",
          6772 => x"54747727",
          6773 => x"f89f3881",
          6774 => x"14547382",
          6775 => x"ccdc3474",
          6776 => x"1a703352",
          6777 => x"54ffaabd",
          6778 => x"3f82ccdc",
          6779 => x"337081ff",
          6780 => x"0682ccd8",
          6781 => x"33585654",
          6782 => x"757526db",
          6783 => x"38f7f639",
          6784 => x"82ccdc53",
          6785 => x"805282a2",
          6786 => x"f051efbd",
          6787 => x"3f800b82",
          6788 => x"ccdc3480",
          6789 => x"0b82ccd8",
          6790 => x"34f7da39",
          6791 => x"7ab03882",
          6792 => x"b4f40855",
          6793 => x"74802ea6",
          6794 => x"387451ff",
          6795 => x"b2f73f82",
          6796 => x"b5a80882",
          6797 => x"ccd83482",
          6798 => x"b5a80881",
          6799 => x"ff068105",
          6800 => x"53745279",
          6801 => x"51ffb4bd",
          6802 => x"3f935b81",
          6803 => x"c0397a84",
          6804 => x"2982b4a8",
          6805 => x"05fc1108",
          6806 => x"56547480",
          6807 => x"2ea73874",
          6808 => x"51ffb2c1",
          6809 => x"3f82b5a8",
          6810 => x"0882ccd8",
          6811 => x"3482b5a8",
          6812 => x"0881ff06",
          6813 => x"81055374",
          6814 => x"527951ff",
          6815 => x"b4873fff",
          6816 => x"1b5480fa",
          6817 => x"39730855",
          6818 => x"74802ef6",
          6819 => x"e8387451",
          6820 => x"ffb2923f",
          6821 => x"99397a93",
          6822 => x"2e098106",
          6823 => x"ae3882b4",
          6824 => x"a8085574",
          6825 => x"802ea438",
          6826 => x"7451ffb1",
          6827 => x"f83f82b5",
          6828 => x"a80882cc",
          6829 => x"d83482b5",
          6830 => x"a80881ff",
          6831 => x"06810553",
          6832 => x"74527951",
          6833 => x"ffb3be3f",
          6834 => x"80c3397a",
          6835 => x"842982b4",
          6836 => x"ac057008",
          6837 => x"56547480",
          6838 => x"2eab3874",
          6839 => x"51ffb1c5",
          6840 => x"3f82b5a8",
          6841 => x"0882ccd8",
          6842 => x"3482b5a8",
          6843 => x"0881ff06",
          6844 => x"81055374",
          6845 => x"527951ff",
          6846 => x"b38b3f81",
          6847 => x"1b547381",
          6848 => x"ff065b89",
          6849 => x"397482cc",
          6850 => x"d834747a",
          6851 => x"3482ccdc",
          6852 => x"5382ccd8",
          6853 => x"33527951",
          6854 => x"edaf3ff5",
          6855 => x"d83982cc",
          6856 => x"dc337081",
          6857 => x"ff0682cc",
          6858 => x"d8335956",
          6859 => x"54747727",
          6860 => x"f5c33881",
          6861 => x"14547382",
          6862 => x"ccdc3474",
          6863 => x"1a703352",
          6864 => x"54ffa7e1",
          6865 => x"3ff5ae39",
          6866 => x"82ccdc33",
          6867 => x"5473802e",
          6868 => x"f5a33888",
          6869 => x"51ffa7cd",
          6870 => x"3f82ccdc",
          6871 => x"33ff0554",
          6872 => x"7382ccdc",
          6873 => x"34f58e39",
          6874 => x"f93d0d83",
          6875 => x"dff40b82",
          6876 => x"b5a00c82",
          6877 => x"800b82b5",
          6878 => x"9c239080",
          6879 => x"53805283",
          6880 => x"dff451ff",
          6881 => x"b7803f82",
          6882 => x"b5a00854",
          6883 => x"80587774",
          6884 => x"34815776",
          6885 => x"81153482",
          6886 => x"b5a00854",
          6887 => x"77841534",
          6888 => x"76851534",
          6889 => x"82b5a008",
          6890 => x"54778615",
          6891 => x"34768715",
          6892 => x"3482b5a0",
          6893 => x"0882b59c",
          6894 => x"22ff05fe",
          6895 => x"80800770",
          6896 => x"83ffff06",
          6897 => x"70882a58",
          6898 => x"51555674",
          6899 => x"88173473",
          6900 => x"89173482",
          6901 => x"b59c2270",
          6902 => x"882982b5",
          6903 => x"a00805f8",
          6904 => x"11515555",
          6905 => x"77821534",
          6906 => x"76831534",
          6907 => x"893d0d04",
          6908 => x"ff3d0d73",
          6909 => x"52815184",
          6910 => x"72278f38",
          6911 => x"fb12832a",
          6912 => x"82117083",
          6913 => x"ffff0651",
          6914 => x"51517082",
          6915 => x"b5a80c83",
          6916 => x"3d0d04f9",
          6917 => x"3d0d02a6",
          6918 => x"05220284",
          6919 => x"05aa0522",
          6920 => x"710582b5",
          6921 => x"a0087183",
          6922 => x"2b711174",
          6923 => x"832b7311",
          6924 => x"70338112",
          6925 => x"3371882b",
          6926 => x"0702a405",
          6927 => x"ae052271",
          6928 => x"81ffff06",
          6929 => x"0770882a",
          6930 => x"53515259",
          6931 => x"545b5b57",
          6932 => x"53545571",
          6933 => x"77347081",
          6934 => x"183482b5",
          6935 => x"a0081475",
          6936 => x"882a5254",
          6937 => x"70821534",
          6938 => x"74831534",
          6939 => x"82b5a008",
          6940 => x"70177033",
          6941 => x"81123371",
          6942 => x"882b0770",
          6943 => x"832b8fff",
          6944 => x"f8065152",
          6945 => x"56527105",
          6946 => x"7383ffff",
          6947 => x"0670882a",
          6948 => x"54545171",
          6949 => x"82123472",
          6950 => x"81ff0653",
          6951 => x"72831234",
          6952 => x"82b5a008",
          6953 => x"16567176",
          6954 => x"34728117",
          6955 => x"34893d0d",
          6956 => x"04fb3d0d",
          6957 => x"82b5a008",
          6958 => x"0284059e",
          6959 => x"05227083",
          6960 => x"2b721186",
          6961 => x"11338712",
          6962 => x"33718b2b",
          6963 => x"71832b07",
          6964 => x"585b5952",
          6965 => x"55527205",
          6966 => x"84123385",
          6967 => x"13337188",
          6968 => x"2b077088",
          6969 => x"2a545656",
          6970 => x"52708413",
          6971 => x"34738513",
          6972 => x"3482b5a0",
          6973 => x"08701484",
          6974 => x"11338512",
          6975 => x"33718b2b",
          6976 => x"71832b07",
          6977 => x"56595752",
          6978 => x"72058612",
          6979 => x"33871333",
          6980 => x"71882b07",
          6981 => x"70882a54",
          6982 => x"56565270",
          6983 => x"86133473",
          6984 => x"87133482",
          6985 => x"b5a00813",
          6986 => x"70338112",
          6987 => x"3371882b",
          6988 => x"077081ff",
          6989 => x"ff067088",
          6990 => x"2a535153",
          6991 => x"53537173",
          6992 => x"34708114",
          6993 => x"34873d0d",
          6994 => x"04fa3d0d",
          6995 => x"02a20522",
          6996 => x"82b5a008",
          6997 => x"71832b71",
          6998 => x"11703381",
          6999 => x"12337188",
          7000 => x"2b077088",
          7001 => x"29157033",
          7002 => x"81123371",
          7003 => x"982b7190",
          7004 => x"2b07535f",
          7005 => x"5355525a",
          7006 => x"56575354",
          7007 => x"71802580",
          7008 => x"f6387251",
          7009 => x"feab3f82",
          7010 => x"b5a00870",
          7011 => x"16703381",
          7012 => x"1233718b",
          7013 => x"2b71832b",
          7014 => x"07741170",
          7015 => x"33811233",
          7016 => x"71882b07",
          7017 => x"70832b8f",
          7018 => x"fff80651",
          7019 => x"52545153",
          7020 => x"5a585372",
          7021 => x"0574882a",
          7022 => x"54527282",
          7023 => x"13347383",
          7024 => x"133482b5",
          7025 => x"a0087016",
          7026 => x"70338112",
          7027 => x"33718b2b",
          7028 => x"71832b07",
          7029 => x"56595755",
          7030 => x"72057033",
          7031 => x"81123371",
          7032 => x"882b0770",
          7033 => x"81ffff06",
          7034 => x"70882a57",
          7035 => x"51525852",
          7036 => x"72743471",
          7037 => x"81153488",
          7038 => x"3d0d04fb",
          7039 => x"3d0d82b5",
          7040 => x"a0080284",
          7041 => x"059e0522",
          7042 => x"70832b72",
          7043 => x"11821133",
          7044 => x"83123371",
          7045 => x"8b2b7183",
          7046 => x"2b07595b",
          7047 => x"59525652",
          7048 => x"73057133",
          7049 => x"81133371",
          7050 => x"882b0702",
          7051 => x"8c05a205",
          7052 => x"22710770",
          7053 => x"882a5351",
          7054 => x"53535371",
          7055 => x"73347081",
          7056 => x"143482b5",
          7057 => x"a0087015",
          7058 => x"70338112",
          7059 => x"33718b2b",
          7060 => x"71832b07",
          7061 => x"56595752",
          7062 => x"72058212",
          7063 => x"33831333",
          7064 => x"71882b07",
          7065 => x"70882a54",
          7066 => x"55565270",
          7067 => x"82133472",
          7068 => x"83133482",
          7069 => x"b5a00814",
          7070 => x"82113383",
          7071 => x"12337188",
          7072 => x"2b0782b5",
          7073 => x"a80c5254",
          7074 => x"873d0d04",
          7075 => x"f73d0d7b",
          7076 => x"82b5a008",
          7077 => x"31832a70",
          7078 => x"83ffff06",
          7079 => x"70535753",
          7080 => x"fda73f82",
          7081 => x"b5a00876",
          7082 => x"832b7111",
          7083 => x"82113383",
          7084 => x"1233718b",
          7085 => x"2b71832b",
          7086 => x"07751170",
          7087 => x"33811233",
          7088 => x"71982b71",
          7089 => x"902b0753",
          7090 => x"42405153",
          7091 => x"5b585559",
          7092 => x"54728025",
          7093 => x"8d388280",
          7094 => x"80527551",
          7095 => x"fe9d3f81",
          7096 => x"84398414",
          7097 => x"33851533",
          7098 => x"718b2b71",
          7099 => x"832b0776",
          7100 => x"1179882a",
          7101 => x"53515558",
          7102 => x"55768614",
          7103 => x"347581ff",
          7104 => x"06567587",
          7105 => x"143482b5",
          7106 => x"a0087019",
          7107 => x"84123385",
          7108 => x"13337188",
          7109 => x"2b077088",
          7110 => x"2a54575b",
          7111 => x"56537284",
          7112 => x"16347385",
          7113 => x"163482b5",
          7114 => x"a0081853",
          7115 => x"800b8614",
          7116 => x"34800b87",
          7117 => x"143482b5",
          7118 => x"a0085376",
          7119 => x"84143475",
          7120 => x"85143482",
          7121 => x"b5a00818",
          7122 => x"70338112",
          7123 => x"3371882b",
          7124 => x"07708280",
          7125 => x"80077088",
          7126 => x"2a535155",
          7127 => x"56547474",
          7128 => x"34728115",
          7129 => x"348b3d0d",
          7130 => x"04ff3d0d",
          7131 => x"735282b5",
          7132 => x"a0088438",
          7133 => x"f7f23f71",
          7134 => x"802e8638",
          7135 => x"7151fe8c",
          7136 => x"3f833d0d",
          7137 => x"04f53d0d",
          7138 => x"807e5258",
          7139 => x"f8e23f82",
          7140 => x"b5a80883",
          7141 => x"ffff0682",
          7142 => x"b5a00884",
          7143 => x"11338512",
          7144 => x"3371882b",
          7145 => x"07705f59",
          7146 => x"56585a81",
          7147 => x"ffff5975",
          7148 => x"782e80cb",
          7149 => x"38758829",
          7150 => x"17703381",
          7151 => x"12337188",
          7152 => x"2b077081",
          7153 => x"ffff0679",
          7154 => x"317083ff",
          7155 => x"ff06707f",
          7156 => x"27525351",
          7157 => x"56595577",
          7158 => x"79278a38",
          7159 => x"73802e85",
          7160 => x"3875785a",
          7161 => x"5b841533",
          7162 => x"85163371",
          7163 => x"882b0757",
          7164 => x"5475c238",
          7165 => x"7881ffff",
          7166 => x"2e85387a",
          7167 => x"79595680",
          7168 => x"76832b82",
          7169 => x"b5a00811",
          7170 => x"70338112",
          7171 => x"3371882b",
          7172 => x"077081ff",
          7173 => x"ff065152",
          7174 => x"5a565c55",
          7175 => x"73752e83",
          7176 => x"38815580",
          7177 => x"54797826",
          7178 => x"81cc3874",
          7179 => x"5474802e",
          7180 => x"81c43877",
          7181 => x"7a2e0981",
          7182 => x"06893875",
          7183 => x"51f8f23f",
          7184 => x"81ac3982",
          7185 => x"80805379",
          7186 => x"527551f7",
          7187 => x"c63f82b5",
          7188 => x"a008701c",
          7189 => x"86113387",
          7190 => x"1233718b",
          7191 => x"2b71832b",
          7192 => x"07535a5e",
          7193 => x"5574057a",
          7194 => x"177083ff",
          7195 => x"ff067088",
          7196 => x"2a5c5956",
          7197 => x"54788415",
          7198 => x"347681ff",
          7199 => x"06577685",
          7200 => x"153482b5",
          7201 => x"a0087583",
          7202 => x"2b711172",
          7203 => x"1e861133",
          7204 => x"87123371",
          7205 => x"882b0770",
          7206 => x"882a535b",
          7207 => x"5e535a56",
          7208 => x"54738619",
          7209 => x"34758719",
          7210 => x"3482b5a0",
          7211 => x"08701c84",
          7212 => x"11338512",
          7213 => x"33718b2b",
          7214 => x"71832b07",
          7215 => x"535d5a55",
          7216 => x"74055478",
          7217 => x"86153476",
          7218 => x"87153482",
          7219 => x"b5a00870",
          7220 => x"16711d84",
          7221 => x"11338512",
          7222 => x"3371882b",
          7223 => x"0770882a",
          7224 => x"535a5f52",
          7225 => x"56547384",
          7226 => x"16347585",
          7227 => x"163482b5",
          7228 => x"a0081b84",
          7229 => x"05547382",
          7230 => x"b5a80c8d",
          7231 => x"3d0d04fe",
          7232 => x"3d0d7452",
          7233 => x"82b5a008",
          7234 => x"8438f4dc",
          7235 => x"3f715371",
          7236 => x"802e8b38",
          7237 => x"7151fced",
          7238 => x"3f82b5a8",
          7239 => x"08537282",
          7240 => x"b5a80c84",
          7241 => x"3d0d04ee",
          7242 => x"3d0d6466",
          7243 => x"405c8070",
          7244 => x"424082b5",
          7245 => x"a008602e",
          7246 => x"09810684",
          7247 => x"38f4a93f",
          7248 => x"7b8e387e",
          7249 => x"51ffb83f",
          7250 => x"82b5a808",
          7251 => x"5483c739",
          7252 => x"7e8b387b",
          7253 => x"51fc923f",
          7254 => x"7e5483ba",
          7255 => x"397e51f5",
          7256 => x"8f3f82b5",
          7257 => x"a80883ff",
          7258 => x"ff0682b5",
          7259 => x"a0087d71",
          7260 => x"31832a70",
          7261 => x"83ffff06",
          7262 => x"70832b73",
          7263 => x"11703381",
          7264 => x"12337188",
          7265 => x"2b077075",
          7266 => x"317083ff",
          7267 => x"ff067088",
          7268 => x"29fc0573",
          7269 => x"88291a70",
          7270 => x"33811233",
          7271 => x"71882b07",
          7272 => x"70902b53",
          7273 => x"444e5348",
          7274 => x"41525c54",
          7275 => x"5b415c56",
          7276 => x"5b5b7380",
          7277 => x"258f3876",
          7278 => x"81ffff06",
          7279 => x"75317083",
          7280 => x"ffff0642",
          7281 => x"54821633",
          7282 => x"83173371",
          7283 => x"882b0770",
          7284 => x"88291c70",
          7285 => x"33811233",
          7286 => x"71982b71",
          7287 => x"902b0753",
          7288 => x"47455256",
          7289 => x"54738025",
          7290 => x"8b387875",
          7291 => x"317083ff",
          7292 => x"ff064154",
          7293 => x"777b2781",
          7294 => x"fe386018",
          7295 => x"54737b2e",
          7296 => x"0981068f",
          7297 => x"387851f6",
          7298 => x"c03f7a83",
          7299 => x"ffff0658",
          7300 => x"81e5397f",
          7301 => x"8e387a74",
          7302 => x"24893878",
          7303 => x"51f6aa3f",
          7304 => x"81a5397f",
          7305 => x"18557a75",
          7306 => x"2480c838",
          7307 => x"791d8211",
          7308 => x"33831233",
          7309 => x"71882b07",
          7310 => x"535754f4",
          7311 => x"f43f8052",
          7312 => x"7851f7b7",
          7313 => x"3f82b5a8",
          7314 => x"0883ffff",
          7315 => x"067e547c",
          7316 => x"5370832b",
          7317 => x"82b5a008",
          7318 => x"11840553",
          7319 => x"5559ff9f",
          7320 => x"da3f82b5",
          7321 => x"a0081484",
          7322 => x"057583ff",
          7323 => x"ff06595c",
          7324 => x"81853960",
          7325 => x"15547a74",
          7326 => x"2480d438",
          7327 => x"7851f5c9",
          7328 => x"3f82b5a0",
          7329 => x"081d8211",
          7330 => x"33831233",
          7331 => x"71882b07",
          7332 => x"534354f4",
          7333 => x"9c3f8052",
          7334 => x"7851f6df",
          7335 => x"3f82b5a8",
          7336 => x"0883ffff",
          7337 => x"067e547c",
          7338 => x"5370832b",
          7339 => x"82b5a008",
          7340 => x"11840553",
          7341 => x"5559ff9f",
          7342 => x"823f82b5",
          7343 => x"a0081484",
          7344 => x"05606205",
          7345 => x"19555c73",
          7346 => x"83ffff06",
          7347 => x"58a9397b",
          7348 => x"7f5254f9",
          7349 => x"b03f82b5",
          7350 => x"a8085c82",
          7351 => x"b5a80880",
          7352 => x"2e93387d",
          7353 => x"53735282",
          7354 => x"b5a80851",
          7355 => x"ffa3963f",
          7356 => x"7351f798",
          7357 => x"3f7a587a",
          7358 => x"78279938",
          7359 => x"80537a52",
          7360 => x"7851f28f",
          7361 => x"3f7a1983",
          7362 => x"2b82b5a0",
          7363 => x"08058405",
          7364 => x"51f6f93f",
          7365 => x"7b547382",
          7366 => x"b5a80c94",
          7367 => x"3d0d04fc",
          7368 => x"3d0d7777",
          7369 => x"29705254",
          7370 => x"fbd53f82",
          7371 => x"b5a80855",
          7372 => x"82b5a808",
          7373 => x"802e8e38",
          7374 => x"73538052",
          7375 => x"82b5a808",
          7376 => x"51ffa7c2",
          7377 => x"3f7482b5",
          7378 => x"a80c863d",
          7379 => x"0d04ff3d",
          7380 => x"0d028f05",
          7381 => x"33518152",
          7382 => x"70722687",
          7383 => x"3882b5a4",
          7384 => x"11335271",
          7385 => x"82b5a80c",
          7386 => x"833d0d04",
          7387 => x"fc3d0d02",
          7388 => x"9b053302",
          7389 => x"84059f05",
          7390 => x"33565383",
          7391 => x"51728126",
          7392 => x"80e03872",
          7393 => x"842b87c0",
          7394 => x"928c1153",
          7395 => x"51885474",
          7396 => x"802e8438",
          7397 => x"81885473",
          7398 => x"720c87c0",
          7399 => x"928c1151",
          7400 => x"81710c85",
          7401 => x"0b87c098",
          7402 => x"8c0c7052",
          7403 => x"71087082",
          7404 => x"06515170",
          7405 => x"802e8a38",
          7406 => x"87c0988c",
          7407 => x"085170ec",
          7408 => x"387108fc",
          7409 => x"80800652",
          7410 => x"71923887",
          7411 => x"c0988c08",
          7412 => x"5170802e",
          7413 => x"87387182",
          7414 => x"b5a41434",
          7415 => x"82b5a413",
          7416 => x"33517082",
          7417 => x"b5a80c86",
          7418 => x"3d0d04f3",
          7419 => x"3d0d6062",
          7420 => x"64028c05",
          7421 => x"bf053357",
          7422 => x"40585b83",
          7423 => x"74525afe",
          7424 => x"cd3f82b5",
          7425 => x"a8088106",
          7426 => x"7a545271",
          7427 => x"81be3871",
          7428 => x"7275842b",
          7429 => x"87c09280",
          7430 => x"1187c092",
          7431 => x"8c1287c0",
          7432 => x"92841341",
          7433 => x"5a40575a",
          7434 => x"58850b87",
          7435 => x"c0988c0c",
          7436 => x"767d0c84",
          7437 => x"760c7508",
          7438 => x"70852a70",
          7439 => x"81065153",
          7440 => x"5471802e",
          7441 => x"8e387b08",
          7442 => x"52717b70",
          7443 => x"81055d34",
          7444 => x"81195980",
          7445 => x"74a20653",
          7446 => x"5371732e",
          7447 => x"83388153",
          7448 => x"7883ff26",
          7449 => x"8f387280",
          7450 => x"2e8a3887",
          7451 => x"c0988c08",
          7452 => x"5271c338",
          7453 => x"87c0988c",
          7454 => x"08527180",
          7455 => x"2e873878",
          7456 => x"84802e99",
          7457 => x"3881760c",
          7458 => x"87c0928c",
          7459 => x"15537208",
          7460 => x"70820651",
          7461 => x"5271f738",
          7462 => x"ff1a5a8d",
          7463 => x"39848017",
          7464 => x"81197081",
          7465 => x"ff065a53",
          7466 => x"5779802e",
          7467 => x"903873fc",
          7468 => x"80800652",
          7469 => x"7187387d",
          7470 => x"7826feed",
          7471 => x"3873fc80",
          7472 => x"80065271",
          7473 => x"802e8338",
          7474 => x"81527153",
          7475 => x"7282b5a8",
          7476 => x"0c8f3d0d",
          7477 => x"04f33d0d",
          7478 => x"60626402",
          7479 => x"8c05bf05",
          7480 => x"33574058",
          7481 => x"5b835980",
          7482 => x"745258fc",
          7483 => x"e13f82b5",
          7484 => x"a8088106",
          7485 => x"79545271",
          7486 => x"782e0981",
          7487 => x"0681b138",
          7488 => x"7774842b",
          7489 => x"87c09280",
          7490 => x"1187c092",
          7491 => x"8c1287c0",
          7492 => x"92841340",
          7493 => x"595f565a",
          7494 => x"850b87c0",
          7495 => x"988c0c76",
          7496 => x"7d0c8276",
          7497 => x"0c805875",
          7498 => x"0870842a",
          7499 => x"70810651",
          7500 => x"53547180",
          7501 => x"2e8c387a",
          7502 => x"7081055c",
          7503 => x"337c0c81",
          7504 => x"18587381",
          7505 => x"2a708106",
          7506 => x"51527180",
          7507 => x"2e8a3887",
          7508 => x"c0988c08",
          7509 => x"5271d038",
          7510 => x"87c0988c",
          7511 => x"08527180",
          7512 => x"2e873877",
          7513 => x"84802e99",
          7514 => x"3881760c",
          7515 => x"87c0928c",
          7516 => x"15537208",
          7517 => x"70820651",
          7518 => x"5271f738",
          7519 => x"ff19598d",
          7520 => x"39811a70",
          7521 => x"81ff0684",
          7522 => x"8019595b",
          7523 => x"5278802e",
          7524 => x"903873fc",
          7525 => x"80800652",
          7526 => x"7187387d",
          7527 => x"7a26fef8",
          7528 => x"3873fc80",
          7529 => x"80065271",
          7530 => x"802e8338",
          7531 => x"81527153",
          7532 => x"7282b5a8",
          7533 => x"0c8f3d0d",
          7534 => x"04fa3d0d",
          7535 => x"7a028405",
          7536 => x"a3053302",
          7537 => x"8805a705",
          7538 => x"33715454",
          7539 => x"5657fafe",
          7540 => x"3f82b5a8",
          7541 => x"08810653",
          7542 => x"83547280",
          7543 => x"fe38850b",
          7544 => x"87c0988c",
          7545 => x"0c815671",
          7546 => x"762e80dc",
          7547 => x"38717624",
          7548 => x"93387484",
          7549 => x"2b87c092",
          7550 => x"8c115454",
          7551 => x"71802e8d",
          7552 => x"3880d439",
          7553 => x"71832e80",
          7554 => x"c63880cb",
          7555 => x"39720870",
          7556 => x"812a7081",
          7557 => x"06515152",
          7558 => x"71802e8a",
          7559 => x"3887c098",
          7560 => x"8c085271",
          7561 => x"e83887c0",
          7562 => x"988c0852",
          7563 => x"71963881",
          7564 => x"730c87c0",
          7565 => x"928c1453",
          7566 => x"72087082",
          7567 => x"06515271",
          7568 => x"f7389639",
          7569 => x"80569239",
          7570 => x"88800a77",
          7571 => x"0c853981",
          7572 => x"80770c72",
          7573 => x"56833984",
          7574 => x"56755473",
          7575 => x"82b5a80c",
          7576 => x"883d0d04",
          7577 => x"fe3d0d74",
          7578 => x"81113371",
          7579 => x"3371882b",
          7580 => x"0782b5a8",
          7581 => x"0c535184",
          7582 => x"3d0d04fd",
          7583 => x"3d0d7583",
          7584 => x"11338212",
          7585 => x"3371902b",
          7586 => x"71882b07",
          7587 => x"81143370",
          7588 => x"7207882b",
          7589 => x"75337107",
          7590 => x"82b5a80c",
          7591 => x"52535456",
          7592 => x"5452853d",
          7593 => x"0d04ff3d",
          7594 => x"0d730284",
          7595 => x"05920522",
          7596 => x"52527072",
          7597 => x"70810554",
          7598 => x"3470882a",
          7599 => x"51707234",
          7600 => x"833d0d04",
          7601 => x"ff3d0d73",
          7602 => x"75525270",
          7603 => x"72708105",
          7604 => x"54347088",
          7605 => x"2a517072",
          7606 => x"70810554",
          7607 => x"3470882a",
          7608 => x"51707270",
          7609 => x"81055434",
          7610 => x"70882a51",
          7611 => x"70723483",
          7612 => x"3d0d04fe",
          7613 => x"3d0d7675",
          7614 => x"77545451",
          7615 => x"70802e92",
          7616 => x"38717081",
          7617 => x"05533373",
          7618 => x"70810555",
          7619 => x"34ff1151",
          7620 => x"eb39843d",
          7621 => x"0d04fe3d",
          7622 => x"0d757776",
          7623 => x"54525372",
          7624 => x"72708105",
          7625 => x"5434ff11",
          7626 => x"5170f438",
          7627 => x"843d0d04",
          7628 => x"fc3d0d78",
          7629 => x"77795656",
          7630 => x"53747081",
          7631 => x"05563374",
          7632 => x"70810556",
          7633 => x"33717131",
          7634 => x"ff165652",
          7635 => x"52527280",
          7636 => x"2e863871",
          7637 => x"802ee238",
          7638 => x"7182b5a8",
          7639 => x"0c863d0d",
          7640 => x"04fe3d0d",
          7641 => x"74765451",
          7642 => x"89397173",
          7643 => x"2e8a3881",
          7644 => x"11517033",
          7645 => x"5271f338",
          7646 => x"703382b5",
          7647 => x"a80c843d",
          7648 => x"0d04800b",
          7649 => x"82b5a80c",
          7650 => x"04800b82",
          7651 => x"b5a80c04",
          7652 => x"f73d0d7b",
          7653 => x"56800b83",
          7654 => x"1733565a",
          7655 => x"747a2e80",
          7656 => x"d6388154",
          7657 => x"b0160853",
          7658 => x"b4167053",
          7659 => x"81173352",
          7660 => x"59faa23f",
          7661 => x"82b5a808",
          7662 => x"7a2e0981",
          7663 => x"06b73882",
          7664 => x"b5a80883",
          7665 => x"1734b016",
          7666 => x"0870a418",
          7667 => x"08319c18",
          7668 => x"08595658",
          7669 => x"7477279f",
          7670 => x"38821633",
          7671 => x"5574822e",
          7672 => x"09810693",
          7673 => x"38815476",
          7674 => x"18537852",
          7675 => x"81163351",
          7676 => x"f9e33f83",
          7677 => x"39815a79",
          7678 => x"82b5a80c",
          7679 => x"8b3d0d04",
          7680 => x"fa3d0d78",
          7681 => x"7a565680",
          7682 => x"5774b017",
          7683 => x"082eaf38",
          7684 => x"7551fefc",
          7685 => x"3f82b5a8",
          7686 => x"085782b5",
          7687 => x"a8089f38",
          7688 => x"81547453",
          7689 => x"b4165281",
          7690 => x"163351f7",
          7691 => x"be3f82b5",
          7692 => x"a808802e",
          7693 => x"8538ff55",
          7694 => x"815774b0",
          7695 => x"170c7682",
          7696 => x"b5a80c88",
          7697 => x"3d0d04f8",
          7698 => x"3d0d7a70",
          7699 => x"5257fec0",
          7700 => x"3f82b5a8",
          7701 => x"085882b5",
          7702 => x"a8088191",
          7703 => x"38763355",
          7704 => x"74832e09",
          7705 => x"810680f0",
          7706 => x"38841733",
          7707 => x"5978812e",
          7708 => x"09810680",
          7709 => x"e3388480",
          7710 => x"5382b5a8",
          7711 => x"0852b417",
          7712 => x"705256fd",
          7713 => x"913f82d4",
          7714 => x"d55284b2",
          7715 => x"1751fc96",
          7716 => x"3f848b85",
          7717 => x"a4d25275",
          7718 => x"51fca93f",
          7719 => x"868a85e4",
          7720 => x"f2528498",
          7721 => x"1751fc9c",
          7722 => x"3f901708",
          7723 => x"52849c17",
          7724 => x"51fc913f",
          7725 => x"8c170852",
          7726 => x"84a01751",
          7727 => x"fc863fa0",
          7728 => x"17088105",
          7729 => x"70b0190c",
          7730 => x"79555375",
          7731 => x"52811733",
          7732 => x"51f8823f",
          7733 => x"77841834",
          7734 => x"80538052",
          7735 => x"81173351",
          7736 => x"f9d73f82",
          7737 => x"b5a80880",
          7738 => x"2e833881",
          7739 => x"587782b5",
          7740 => x"a80c8a3d",
          7741 => x"0d04fb3d",
          7742 => x"0d77fe1a",
          7743 => x"981208fe",
          7744 => x"05555654",
          7745 => x"80567473",
          7746 => x"278d388a",
          7747 => x"14227571",
          7748 => x"29ac1608",
          7749 => x"05575375",
          7750 => x"82b5a80c",
          7751 => x"873d0d04",
          7752 => x"f93d0d7a",
          7753 => x"7a700856",
          7754 => x"54578177",
          7755 => x"2781df38",
          7756 => x"76981508",
          7757 => x"2781d738",
          7758 => x"ff743354",
          7759 => x"5872822e",
          7760 => x"80f53872",
          7761 => x"82248938",
          7762 => x"72812e8d",
          7763 => x"3881bf39",
          7764 => x"72832e81",
          7765 => x"8e3881b6",
          7766 => x"3976812a",
          7767 => x"1770892a",
          7768 => x"a4160805",
          7769 => x"53745255",
          7770 => x"fd963f82",
          7771 => x"b5a80881",
          7772 => x"9f387483",
          7773 => x"ff0614b4",
          7774 => x"11338117",
          7775 => x"70892aa4",
          7776 => x"18080555",
          7777 => x"76545757",
          7778 => x"53fcf53f",
          7779 => x"82b5a808",
          7780 => x"80fe3874",
          7781 => x"83ff0614",
          7782 => x"b4113370",
          7783 => x"882b7807",
          7784 => x"79810671",
          7785 => x"842a5c52",
          7786 => x"58515372",
          7787 => x"80e23875",
          7788 => x"9fff0658",
          7789 => x"80da3976",
          7790 => x"882aa415",
          7791 => x"08055273",
          7792 => x"51fcbd3f",
          7793 => x"82b5a808",
          7794 => x"80c63876",
          7795 => x"1083fe06",
          7796 => x"7405b405",
          7797 => x"51f98d3f",
          7798 => x"82b5a808",
          7799 => x"83ffff06",
          7800 => x"58ae3976",
          7801 => x"872aa415",
          7802 => x"08055273",
          7803 => x"51fc913f",
          7804 => x"82b5a808",
          7805 => x"9b387682",
          7806 => x"2b83fc06",
          7807 => x"7405b405",
          7808 => x"51f8f83f",
          7809 => x"82b5a808",
          7810 => x"f00a0658",
          7811 => x"83398158",
          7812 => x"7782b5a8",
          7813 => x"0c893d0d",
          7814 => x"04f83d0d",
          7815 => x"7a7c7e5a",
          7816 => x"58568259",
          7817 => x"81772782",
          7818 => x"9e387698",
          7819 => x"17082782",
          7820 => x"96387533",
          7821 => x"5372792e",
          7822 => x"819d3872",
          7823 => x"79248938",
          7824 => x"72812e8d",
          7825 => x"38828039",
          7826 => x"72832e81",
          7827 => x"b83881f7",
          7828 => x"3976812a",
          7829 => x"1770892a",
          7830 => x"a4180805",
          7831 => x"53765255",
          7832 => x"fb9e3f82",
          7833 => x"b5a80859",
          7834 => x"82b5a808",
          7835 => x"81d93874",
          7836 => x"83ff0616",
          7837 => x"b4058116",
          7838 => x"78810659",
          7839 => x"56547753",
          7840 => x"76802e8f",
          7841 => x"3877842b",
          7842 => x"9ff00674",
          7843 => x"338f0671",
          7844 => x"07515372",
          7845 => x"7434810b",
          7846 => x"83173474",
          7847 => x"892aa417",
          7848 => x"08055275",
          7849 => x"51fad93f",
          7850 => x"82b5a808",
          7851 => x"5982b5a8",
          7852 => x"08819438",
          7853 => x"7483ff06",
          7854 => x"16b40578",
          7855 => x"842a5454",
          7856 => x"768f3877",
          7857 => x"882a7433",
          7858 => x"81f00671",
          7859 => x"8f060751",
          7860 => x"53727434",
          7861 => x"80ec3976",
          7862 => x"882aa417",
          7863 => x"08055275",
          7864 => x"51fa9d3f",
          7865 => x"82b5a808",
          7866 => x"5982b5a8",
          7867 => x"0880d838",
          7868 => x"7783ffff",
          7869 => x"06527610",
          7870 => x"83fe0676",
          7871 => x"05b40551",
          7872 => x"f7a43fbe",
          7873 => x"3976872a",
          7874 => x"a4170805",
          7875 => x"527551f9",
          7876 => x"ef3f82b5",
          7877 => x"a8085982",
          7878 => x"b5a808ab",
          7879 => x"3877f00a",
          7880 => x"0677822b",
          7881 => x"83fc0670",
          7882 => x"18b40570",
          7883 => x"54515454",
          7884 => x"f6c93f82",
          7885 => x"b5a8088f",
          7886 => x"0a067407",
          7887 => x"527251f7",
          7888 => x"833f810b",
          7889 => x"83173478",
          7890 => x"82b5a80c",
          7891 => x"8a3d0d04",
          7892 => x"f83d0d7a",
          7893 => x"7c7e7208",
          7894 => x"59565659",
          7895 => x"817527a4",
          7896 => x"38749817",
          7897 => x"08279d38",
          7898 => x"73802eaa",
          7899 => x"38ff5373",
          7900 => x"527551fd",
          7901 => x"a43f82b5",
          7902 => x"a8085482",
          7903 => x"b5a80880",
          7904 => x"f2389339",
          7905 => x"825480eb",
          7906 => x"39815480",
          7907 => x"e63982b5",
          7908 => x"a8085480",
          7909 => x"de397452",
          7910 => x"7851fb84",
          7911 => x"3f82b5a8",
          7912 => x"085882b5",
          7913 => x"a808802e",
          7914 => x"80c73882",
          7915 => x"b5a80881",
          7916 => x"2ed23882",
          7917 => x"b5a808ff",
          7918 => x"2ecf3880",
          7919 => x"53745275",
          7920 => x"51fcd63f",
          7921 => x"82b5a808",
          7922 => x"c5389816",
          7923 => x"08fe1190",
          7924 => x"18085755",
          7925 => x"57747427",
          7926 => x"90388115",
          7927 => x"90170c84",
          7928 => x"16338107",
          7929 => x"54738417",
          7930 => x"34775576",
          7931 => x"7826ffa6",
          7932 => x"38805473",
          7933 => x"82b5a80c",
          7934 => x"8a3d0d04",
          7935 => x"f63d0d7c",
          7936 => x"7e710859",
          7937 => x"5b5b7995",
          7938 => x"388c1708",
          7939 => x"5877802e",
          7940 => x"88389817",
          7941 => x"087826b2",
          7942 => x"388158ae",
          7943 => x"3979527a",
          7944 => x"51f9fd3f",
          7945 => x"81557482",
          7946 => x"b5a80827",
          7947 => x"82e03882",
          7948 => x"b5a80855",
          7949 => x"82b5a808",
          7950 => x"ff2e82d2",
          7951 => x"38981708",
          7952 => x"82b5a808",
          7953 => x"2682c738",
          7954 => x"79589017",
          7955 => x"08705654",
          7956 => x"73802e82",
          7957 => x"b938777a",
          7958 => x"2e098106",
          7959 => x"80e23881",
          7960 => x"1a569817",
          7961 => x"08762683",
          7962 => x"38825675",
          7963 => x"527a51f9",
          7964 => x"af3f8059",
          7965 => x"82b5a808",
          7966 => x"812e0981",
          7967 => x"06863882",
          7968 => x"b5a80859",
          7969 => x"82b5a808",
          7970 => x"09703070",
          7971 => x"72078025",
          7972 => x"707c0782",
          7973 => x"b5a80854",
          7974 => x"51515555",
          7975 => x"7381ef38",
          7976 => x"82b5a808",
          7977 => x"802e9538",
          7978 => x"8c170854",
          7979 => x"81742790",
          7980 => x"38739818",
          7981 => x"08278938",
          7982 => x"73588539",
          7983 => x"7580db38",
          7984 => x"77568116",
          7985 => x"56981708",
          7986 => x"76268938",
          7987 => x"82567578",
          7988 => x"2681ac38",
          7989 => x"75527a51",
          7990 => x"f8c63f82",
          7991 => x"b5a80880",
          7992 => x"2eb83880",
          7993 => x"5982b5a8",
          7994 => x"08812e09",
          7995 => x"81068638",
          7996 => x"82b5a808",
          7997 => x"5982b5a8",
          7998 => x"08097030",
          7999 => x"70720780",
          8000 => x"25707c07",
          8001 => x"51515555",
          8002 => x"7380f838",
          8003 => x"75782e09",
          8004 => x"8106ffae",
          8005 => x"38735580",
          8006 => x"f539ff53",
          8007 => x"75527651",
          8008 => x"f9f73f82",
          8009 => x"b5a80882",
          8010 => x"b5a80830",
          8011 => x"7082b5a8",
          8012 => x"08078025",
          8013 => x"51555579",
          8014 => x"802e9438",
          8015 => x"73802e8f",
          8016 => x"38755379",
          8017 => x"527651f9",
          8018 => x"d03f82b5",
          8019 => x"a8085574",
          8020 => x"a538758c",
          8021 => x"180c9817",
          8022 => x"08fe0590",
          8023 => x"18085654",
          8024 => x"74742686",
          8025 => x"38ff1590",
          8026 => x"180c8417",
          8027 => x"33810754",
          8028 => x"73841834",
          8029 => x"9739ff56",
          8030 => x"74812e90",
          8031 => x"388c3980",
          8032 => x"558c3982",
          8033 => x"b5a80855",
          8034 => x"85398156",
          8035 => x"75557482",
          8036 => x"b5a80c8c",
          8037 => x"3d0d04f8",
          8038 => x"3d0d7a70",
          8039 => x"5255f3f0",
          8040 => x"3f82b5a8",
          8041 => x"08588156",
          8042 => x"82b5a808",
          8043 => x"80d8387b",
          8044 => x"527451f6",
          8045 => x"c13f82b5",
          8046 => x"a80882b5",
          8047 => x"a808b017",
          8048 => x"0c598480",
          8049 => x"537752b4",
          8050 => x"15705257",
          8051 => x"f2c83f77",
          8052 => x"56843981",
          8053 => x"16568a15",
          8054 => x"22587578",
          8055 => x"27973881",
          8056 => x"54751953",
          8057 => x"76528115",
          8058 => x"3351ede9",
          8059 => x"3f82b5a8",
          8060 => x"08802edf",
          8061 => x"388a1522",
          8062 => x"76327030",
          8063 => x"70720770",
          8064 => x"9f2a5351",
          8065 => x"56567582",
          8066 => x"b5a80c8a",
          8067 => x"3d0d04f8",
          8068 => x"3d0d7a7c",
          8069 => x"71085856",
          8070 => x"5774f080",
          8071 => x"0a2680f1",
          8072 => x"38749f06",
          8073 => x"537280e9",
          8074 => x"38749018",
          8075 => x"0c881708",
          8076 => x"5473aa38",
          8077 => x"75335382",
          8078 => x"73278838",
          8079 => x"a8160854",
          8080 => x"739b3874",
          8081 => x"852a5382",
          8082 => x"0b881722",
          8083 => x"5a587279",
          8084 => x"2780fe38",
          8085 => x"a8160898",
          8086 => x"180c80cd",
          8087 => x"398a1622",
          8088 => x"70892b54",
          8089 => x"58727526",
          8090 => x"b2387352",
          8091 => x"7651f5b0",
          8092 => x"3f82b5a8",
          8093 => x"085482b5",
          8094 => x"a808ff2e",
          8095 => x"bd38810b",
          8096 => x"82b5a808",
          8097 => x"278b3898",
          8098 => x"160882b5",
          8099 => x"a8082685",
          8100 => x"388258bd",
          8101 => x"39747331",
          8102 => x"55cb3973",
          8103 => x"527551f4",
          8104 => x"d53f82b5",
          8105 => x"a8089818",
          8106 => x"0c739418",
          8107 => x"0c981708",
          8108 => x"53825872",
          8109 => x"802e9a38",
          8110 => x"85398158",
          8111 => x"94397489",
          8112 => x"2a139818",
          8113 => x"0c7483ff",
          8114 => x"0616b405",
          8115 => x"9c180c80",
          8116 => x"587782b5",
          8117 => x"a80c8a3d",
          8118 => x"0d04f83d",
          8119 => x"0d7a7008",
          8120 => x"901208a0",
          8121 => x"05595754",
          8122 => x"f0800a77",
          8123 => x"27863880",
          8124 => x"0b98150c",
          8125 => x"98140853",
          8126 => x"84557280",
          8127 => x"2e81cb38",
          8128 => x"7683ff06",
          8129 => x"587781b5",
          8130 => x"38811398",
          8131 => x"150c9414",
          8132 => x"08557492",
          8133 => x"3876852a",
          8134 => x"88172256",
          8135 => x"53747326",
          8136 => x"819b3880",
          8137 => x"c0398a16",
          8138 => x"22ff0577",
          8139 => x"892a0653",
          8140 => x"72818a38",
          8141 => x"74527351",
          8142 => x"f3e63f82",
          8143 => x"b5a80853",
          8144 => x"8255810b",
          8145 => x"82b5a808",
          8146 => x"2780ff38",
          8147 => x"815582b5",
          8148 => x"a808ff2e",
          8149 => x"80f43898",
          8150 => x"160882b5",
          8151 => x"a8082680",
          8152 => x"ca387b8a",
          8153 => x"38779815",
          8154 => x"0c845580",
          8155 => x"dd399414",
          8156 => x"08527351",
          8157 => x"f9863f82",
          8158 => x"b5a80853",
          8159 => x"875582b5",
          8160 => x"a808802e",
          8161 => x"80c43882",
          8162 => x"5582b5a8",
          8163 => x"08812eba",
          8164 => x"38815582",
          8165 => x"b5a808ff",
          8166 => x"2eb03882",
          8167 => x"b5a80852",
          8168 => x"7551fbf3",
          8169 => x"3f82b5a8",
          8170 => x"08a03872",
          8171 => x"94150c72",
          8172 => x"527551f2",
          8173 => x"c13f82b5",
          8174 => x"a8089815",
          8175 => x"0c769015",
          8176 => x"0c7716b4",
          8177 => x"059c150c",
          8178 => x"80557482",
          8179 => x"b5a80c8a",
          8180 => x"3d0d04f7",
          8181 => x"3d0d7b7d",
          8182 => x"71085b5b",
          8183 => x"57805276",
          8184 => x"51fcac3f",
          8185 => x"82b5a808",
          8186 => x"5482b5a8",
          8187 => x"0880ec38",
          8188 => x"82b5a808",
          8189 => x"56981708",
          8190 => x"527851f0",
          8191 => x"833f82b5",
          8192 => x"a8085482",
          8193 => x"b5a80880",
          8194 => x"d23882b5",
          8195 => x"a8089c18",
          8196 => x"08703351",
          8197 => x"54587281",
          8198 => x"e52e0981",
          8199 => x"06833881",
          8200 => x"5882b5a8",
          8201 => x"08557283",
          8202 => x"38815577",
          8203 => x"75075372",
          8204 => x"802e8e38",
          8205 => x"81165675",
          8206 => x"7a2e0981",
          8207 => x"068838a5",
          8208 => x"3982b5a8",
          8209 => x"08568152",
          8210 => x"7651fd8e",
          8211 => x"3f82b5a8",
          8212 => x"085482b5",
          8213 => x"a808802e",
          8214 => x"ff9b3873",
          8215 => x"842e0981",
          8216 => x"06833887",
          8217 => x"547382b5",
          8218 => x"a80c8b3d",
          8219 => x"0d04fd3d",
          8220 => x"0d769a11",
          8221 => x"5254ebec",
          8222 => x"3f82b5a8",
          8223 => x"0883ffff",
          8224 => x"06767033",
          8225 => x"51535371",
          8226 => x"832e0981",
          8227 => x"06903894",
          8228 => x"1451ebd0",
          8229 => x"3f82b5a8",
          8230 => x"08902b73",
          8231 => x"07537282",
          8232 => x"b5a80c85",
          8233 => x"3d0d04fc",
          8234 => x"3d0d7779",
          8235 => x"7083ffff",
          8236 => x"06549a12",
          8237 => x"535555eb",
          8238 => x"ed3f7670",
          8239 => x"33515372",
          8240 => x"832e0981",
          8241 => x"068b3873",
          8242 => x"902a5294",
          8243 => x"1551ebd6",
          8244 => x"3f863d0d",
          8245 => x"04f73d0d",
          8246 => x"7b7d5b55",
          8247 => x"8475085a",
          8248 => x"58981508",
          8249 => x"802e818a",
          8250 => x"38981508",
          8251 => x"527851ee",
          8252 => x"8f3f82b5",
          8253 => x"a8085882",
          8254 => x"b5a80880",
          8255 => x"f5389c15",
          8256 => x"08703355",
          8257 => x"53738638",
          8258 => x"845880e6",
          8259 => x"398b1333",
          8260 => x"70bf0670",
          8261 => x"81ff0658",
          8262 => x"51537286",
          8263 => x"163482b5",
          8264 => x"a8085373",
          8265 => x"81e52e83",
          8266 => x"38815373",
          8267 => x"ae2ea938",
          8268 => x"81707406",
          8269 => x"54577280",
          8270 => x"2e9e3875",
          8271 => x"8f2e9938",
          8272 => x"82b5a808",
          8273 => x"76df0654",
          8274 => x"5472882e",
          8275 => x"09810683",
          8276 => x"38765473",
          8277 => x"7a2ea038",
          8278 => x"80527451",
          8279 => x"fafc3f82",
          8280 => x"b5a80858",
          8281 => x"82b5a808",
          8282 => x"89389815",
          8283 => x"08fefa38",
          8284 => x"8639800b",
          8285 => x"98160c77",
          8286 => x"82b5a80c",
          8287 => x"8b3d0d04",
          8288 => x"fb3d0d77",
          8289 => x"70085754",
          8290 => x"81527351",
          8291 => x"fcc53f82",
          8292 => x"b5a80855",
          8293 => x"82b5a808",
          8294 => x"b4389814",
          8295 => x"08527551",
          8296 => x"ecde3f82",
          8297 => x"b5a80855",
          8298 => x"82b5a808",
          8299 => x"a038a053",
          8300 => x"82b5a808",
          8301 => x"529c1408",
          8302 => x"51eadb3f",
          8303 => x"8b53a014",
          8304 => x"529c1408",
          8305 => x"51eaac3f",
          8306 => x"810b8317",
          8307 => x"347482b5",
          8308 => x"a80c873d",
          8309 => x"0d04fd3d",
          8310 => x"0d757008",
          8311 => x"98120854",
          8312 => x"70535553",
          8313 => x"ec9a3f82",
          8314 => x"b5a8088d",
          8315 => x"389c1308",
          8316 => x"53e57334",
          8317 => x"810b8315",
          8318 => x"34853d0d",
          8319 => x"04fa3d0d",
          8320 => x"787a5757",
          8321 => x"800b8917",
          8322 => x"34981708",
          8323 => x"802e8182",
          8324 => x"38807089",
          8325 => x"18555555",
          8326 => x"9c170814",
          8327 => x"70338116",
          8328 => x"56515271",
          8329 => x"a02ea838",
          8330 => x"71852e09",
          8331 => x"81068438",
          8332 => x"81e55273",
          8333 => x"892e0981",
          8334 => x"068b38ae",
          8335 => x"73708105",
          8336 => x"55348115",
          8337 => x"55717370",
          8338 => x"81055534",
          8339 => x"8115558a",
          8340 => x"7427c538",
          8341 => x"75158805",
          8342 => x"52800b81",
          8343 => x"13349c17",
          8344 => x"08528b12",
          8345 => x"33881734",
          8346 => x"9c17089c",
          8347 => x"115252e8",
          8348 => x"8a3f82b5",
          8349 => x"a808760c",
          8350 => x"961251e7",
          8351 => x"e73f82b5",
          8352 => x"a8088617",
          8353 => x"23981251",
          8354 => x"e7da3f82",
          8355 => x"b5a80884",
          8356 => x"1723883d",
          8357 => x"0d04f33d",
          8358 => x"0d7f7008",
          8359 => x"5e5b8061",
          8360 => x"70335155",
          8361 => x"5573af2e",
          8362 => x"83388155",
          8363 => x"7380dc2e",
          8364 => x"91387480",
          8365 => x"2e8c3894",
          8366 => x"1d08881c",
          8367 => x"0caa3981",
          8368 => x"15418061",
          8369 => x"70335656",
          8370 => x"5673af2e",
          8371 => x"09810683",
          8372 => x"38815673",
          8373 => x"80dc3270",
          8374 => x"30708025",
          8375 => x"78075151",
          8376 => x"5473dc38",
          8377 => x"73881c0c",
          8378 => x"60703351",
          8379 => x"54739f26",
          8380 => x"9638ff80",
          8381 => x"0bab1c34",
          8382 => x"80527a51",
          8383 => x"f6913f82",
          8384 => x"b5a80855",
          8385 => x"85983991",
          8386 => x"3d61a01d",
          8387 => x"5c5a5e8b",
          8388 => x"53a05279",
          8389 => x"51e7ff3f",
          8390 => x"80705957",
          8391 => x"88793355",
          8392 => x"5c73ae2e",
          8393 => x"09810680",
          8394 => x"d4387818",
          8395 => x"7033811a",
          8396 => x"71ae3270",
          8397 => x"30709f2a",
          8398 => x"73822607",
          8399 => x"5151535a",
          8400 => x"5754738c",
          8401 => x"38791754",
          8402 => x"75743481",
          8403 => x"1757db39",
          8404 => x"75af3270",
          8405 => x"30709f2a",
          8406 => x"51515475",
          8407 => x"80dc2e8c",
          8408 => x"3873802e",
          8409 => x"873875a0",
          8410 => x"2682bd38",
          8411 => x"77197e0c",
          8412 => x"a454a076",
          8413 => x"2782bd38",
          8414 => x"a05482b8",
          8415 => x"39781870",
          8416 => x"33811a5a",
          8417 => x"5754a076",
          8418 => x"2781fc38",
          8419 => x"75af3270",
          8420 => x"307780dc",
          8421 => x"32703072",
          8422 => x"80257180",
          8423 => x"25075151",
          8424 => x"56515573",
          8425 => x"802eac38",
          8426 => x"84398118",
          8427 => x"5880781a",
          8428 => x"70335155",
          8429 => x"5573af2e",
          8430 => x"09810683",
          8431 => x"38815573",
          8432 => x"80dc3270",
          8433 => x"30708025",
          8434 => x"77075151",
          8435 => x"5473db38",
          8436 => x"81b53975",
          8437 => x"ae2e0981",
          8438 => x"06833881",
          8439 => x"54767c27",
          8440 => x"74075473",
          8441 => x"802ea238",
          8442 => x"7b8b3270",
          8443 => x"3077ae32",
          8444 => x"70307280",
          8445 => x"25719f2a",
          8446 => x"07535156",
          8447 => x"51557481",
          8448 => x"a7388857",
          8449 => x"8b5cfef5",
          8450 => x"3975982b",
          8451 => x"54738025",
          8452 => x"8c387580",
          8453 => x"ff0682ae",
          8454 => x"f0113357",
          8455 => x"547551e6",
          8456 => x"e13f82b5",
          8457 => x"a808802e",
          8458 => x"b2387818",
          8459 => x"7033811a",
          8460 => x"71545a56",
          8461 => x"54e6d23f",
          8462 => x"82b5a808",
          8463 => x"802e80e8",
          8464 => x"38ff1c54",
          8465 => x"76742780",
          8466 => x"df387917",
          8467 => x"54757434",
          8468 => x"81177a11",
          8469 => x"55577474",
          8470 => x"34a73975",
          8471 => x"5282ae90",
          8472 => x"51e5fe3f",
          8473 => x"82b5a808",
          8474 => x"bf38ff9f",
          8475 => x"16547399",
          8476 => x"268938e0",
          8477 => x"167081ff",
          8478 => x"06575479",
          8479 => x"17547574",
          8480 => x"34811757",
          8481 => x"fdf73977",
          8482 => x"197e0c76",
          8483 => x"802e9938",
          8484 => x"79335473",
          8485 => x"81e52e09",
          8486 => x"81068438",
          8487 => x"857a3484",
          8488 => x"54a07627",
          8489 => x"8f388b39",
          8490 => x"865581f2",
          8491 => x"39845680",
          8492 => x"f3398054",
          8493 => x"738b1b34",
          8494 => x"807b0858",
          8495 => x"527a51f2",
          8496 => x"ce3f82b5",
          8497 => x"a8085682",
          8498 => x"b5a80880",
          8499 => x"d738981b",
          8500 => x"08527651",
          8501 => x"e6aa3f82",
          8502 => x"b5a80856",
          8503 => x"82b5a808",
          8504 => x"80c2389c",
          8505 => x"1b087033",
          8506 => x"55557380",
          8507 => x"2effbe38",
          8508 => x"8b1533bf",
          8509 => x"06547386",
          8510 => x"1c348b15",
          8511 => x"3370832a",
          8512 => x"70810651",
          8513 => x"55587392",
          8514 => x"388b5379",
          8515 => x"527451e4",
          8516 => x"9f3f82b5",
          8517 => x"a808802e",
          8518 => x"8b387552",
          8519 => x"7a51f3ba",
          8520 => x"3fff9f39",
          8521 => x"75ab1c33",
          8522 => x"57557480",
          8523 => x"2ebb3874",
          8524 => x"842e0981",
          8525 => x"0680e738",
          8526 => x"75852a70",
          8527 => x"81067782",
          8528 => x"2a585154",
          8529 => x"73802e96",
          8530 => x"38758106",
          8531 => x"5473802e",
          8532 => x"fbb538ff",
          8533 => x"800bab1c",
          8534 => x"34805580",
          8535 => x"c1397581",
          8536 => x"065473ba",
          8537 => x"388555b6",
          8538 => x"3975822a",
          8539 => x"70810651",
          8540 => x"5473ab38",
          8541 => x"861b3370",
          8542 => x"842a7081",
          8543 => x"06515555",
          8544 => x"73802ee1",
          8545 => x"38901b08",
          8546 => x"83ff061d",
          8547 => x"b405527c",
          8548 => x"51f5db3f",
          8549 => x"82b5a808",
          8550 => x"881c0cfa",
          8551 => x"ea397482",
          8552 => x"b5a80c8f",
          8553 => x"3d0d04f6",
          8554 => x"3d0d7c5b",
          8555 => x"ff7b0870",
          8556 => x"71735559",
          8557 => x"5c555973",
          8558 => x"802e81c6",
          8559 => x"38757081",
          8560 => x"05573370",
          8561 => x"a0265252",
          8562 => x"71ba2e8d",
          8563 => x"3870ee38",
          8564 => x"71ba2e09",
          8565 => x"810681a5",
          8566 => x"387333d0",
          8567 => x"117081ff",
          8568 => x"06515253",
          8569 => x"70892691",
          8570 => x"38821473",
          8571 => x"81ff06d0",
          8572 => x"05565271",
          8573 => x"762e80f7",
          8574 => x"38800b82",
          8575 => x"aee05955",
          8576 => x"77087a55",
          8577 => x"57767081",
          8578 => x"05583374",
          8579 => x"70810556",
          8580 => x"33ff9f12",
          8581 => x"53535370",
          8582 => x"99268938",
          8583 => x"e0137081",
          8584 => x"ff065451",
          8585 => x"ff9f1251",
          8586 => x"70992689",
          8587 => x"38e01270",
          8588 => x"81ff0653",
          8589 => x"51723070",
          8590 => x"9f2a5151",
          8591 => x"72722e09",
          8592 => x"81068538",
          8593 => x"70ffbe38",
          8594 => x"72307477",
          8595 => x"32703070",
          8596 => x"72079f2a",
          8597 => x"739f2a07",
          8598 => x"53545451",
          8599 => x"70802e8f",
          8600 => x"38811584",
          8601 => x"19595583",
          8602 => x"7525ff94",
          8603 => x"388b3974",
          8604 => x"83248638",
          8605 => x"74767c0c",
          8606 => x"59785186",
          8607 => x"3982ccf4",
          8608 => x"33517082",
          8609 => x"b5a80c8c",
          8610 => x"3d0d04fa",
          8611 => x"3d0d7856",
          8612 => x"800b8317",
          8613 => x"34ff0bb0",
          8614 => x"170c7952",
          8615 => x"7551e2e0",
          8616 => x"3f845582",
          8617 => x"b5a80881",
          8618 => x"803884b2",
          8619 => x"1651dfb4",
          8620 => x"3f82b5a8",
          8621 => x"0883ffff",
          8622 => x"06548355",
          8623 => x"7382d4d5",
          8624 => x"2e098106",
          8625 => x"80e33880",
          8626 => x"0bb41733",
          8627 => x"56577481",
          8628 => x"e92e0981",
          8629 => x"06833881",
          8630 => x"577481eb",
          8631 => x"32703070",
          8632 => x"80257907",
          8633 => x"51515473",
          8634 => x"8a387481",
          8635 => x"e82e0981",
          8636 => x"06b53883",
          8637 => x"5382aea0",
          8638 => x"5280ea16",
          8639 => x"51e0b13f",
          8640 => x"82b5a808",
          8641 => x"5582b5a8",
          8642 => x"08802e9d",
          8643 => x"38855382",
          8644 => x"aea45281",
          8645 => x"861651e0",
          8646 => x"973f82b5",
          8647 => x"a8085582",
          8648 => x"b5a80880",
          8649 => x"2e833882",
          8650 => x"557482b5",
          8651 => x"a80c883d",
          8652 => x"0d04f23d",
          8653 => x"0d610284",
          8654 => x"0580cb05",
          8655 => x"33585580",
          8656 => x"750c6051",
          8657 => x"fce13f82",
          8658 => x"b5a80858",
          8659 => x"8b56800b",
          8660 => x"82b5a808",
          8661 => x"2486fc38",
          8662 => x"82b5a808",
          8663 => x"842982cc",
          8664 => x"e0057008",
          8665 => x"55538c56",
          8666 => x"73802e86",
          8667 => x"e6387375",
          8668 => x"0c7681fe",
          8669 => x"06743354",
          8670 => x"5772802e",
          8671 => x"ae388114",
          8672 => x"3351d7ca",
          8673 => x"3f82b5a8",
          8674 => x"0881ff06",
          8675 => x"70810654",
          8676 => x"55729838",
          8677 => x"76802e86",
          8678 => x"b8387482",
          8679 => x"2a708106",
          8680 => x"51538a56",
          8681 => x"7286ac38",
          8682 => x"86a73980",
          8683 => x"74347781",
          8684 => x"15348152",
          8685 => x"81143351",
          8686 => x"d7b23f82",
          8687 => x"b5a80881",
          8688 => x"ff067081",
          8689 => x"06545583",
          8690 => x"56728687",
          8691 => x"3876802e",
          8692 => x"8f387482",
          8693 => x"2a708106",
          8694 => x"51538a56",
          8695 => x"7285f438",
          8696 => x"80705374",
          8697 => x"525bfda3",
          8698 => x"3f82b5a8",
          8699 => x"0881ff06",
          8700 => x"5776822e",
          8701 => x"09810680",
          8702 => x"e2388c3d",
          8703 => x"74565883",
          8704 => x"5683f615",
          8705 => x"33705853",
          8706 => x"72802e8d",
          8707 => x"3883fa15",
          8708 => x"51dce83f",
          8709 => x"82b5a808",
          8710 => x"57767870",
          8711 => x"84055a0c",
          8712 => x"ff169016",
          8713 => x"56567580",
          8714 => x"25d73880",
          8715 => x"0b8d3d54",
          8716 => x"56727084",
          8717 => x"0554085b",
          8718 => x"83577a80",
          8719 => x"2e95387a",
          8720 => x"527351fc",
          8721 => x"c63f82b5",
          8722 => x"a80881ff",
          8723 => x"06578177",
          8724 => x"27893881",
          8725 => x"16568376",
          8726 => x"27d73881",
          8727 => x"5676842e",
          8728 => x"84f1388d",
          8729 => x"56768126",
          8730 => x"84e938bf",
          8731 => x"1451dbf4",
          8732 => x"3f82b5a8",
          8733 => x"0883ffff",
          8734 => x"06537284",
          8735 => x"802e0981",
          8736 => x"0684d038",
          8737 => x"80ca1451",
          8738 => x"dbda3f82",
          8739 => x"b5a80883",
          8740 => x"ffff0658",
          8741 => x"778d3880",
          8742 => x"d81451db",
          8743 => x"de3f82b5",
          8744 => x"a8085877",
          8745 => x"9c150c80",
          8746 => x"c4143382",
          8747 => x"153480c4",
          8748 => x"1433ff11",
          8749 => x"7081ff06",
          8750 => x"5154558d",
          8751 => x"56728126",
          8752 => x"84913874",
          8753 => x"81ff0678",
          8754 => x"712980c1",
          8755 => x"16335259",
          8756 => x"53728a15",
          8757 => x"2372802e",
          8758 => x"8b38ff13",
          8759 => x"73065372",
          8760 => x"802e8638",
          8761 => x"8d5683eb",
          8762 => x"3980c514",
          8763 => x"51daf53f",
          8764 => x"82b5a808",
          8765 => x"5382b5a8",
          8766 => x"08881523",
          8767 => x"728f0657",
          8768 => x"8d567683",
          8769 => x"ce3880c7",
          8770 => x"1451dad8",
          8771 => x"3f82b5a8",
          8772 => x"0883ffff",
          8773 => x"0655748d",
          8774 => x"3880d414",
          8775 => x"51dadc3f",
          8776 => x"82b5a808",
          8777 => x"5580c214",
          8778 => x"51dab93f",
          8779 => x"82b5a808",
          8780 => x"83ffff06",
          8781 => x"538d5672",
          8782 => x"802e8397",
          8783 => x"38881422",
          8784 => x"78147184",
          8785 => x"2a055a5a",
          8786 => x"78752683",
          8787 => x"86388a14",
          8788 => x"22527479",
          8789 => x"3151feff",
          8790 => x"ca3f82b5",
          8791 => x"a8085582",
          8792 => x"b5a80880",
          8793 => x"2e82ec38",
          8794 => x"82b5a808",
          8795 => x"80ffffff",
          8796 => x"f5268338",
          8797 => x"83577483",
          8798 => x"fff52683",
          8799 => x"38825774",
          8800 => x"9ff52685",
          8801 => x"38815789",
          8802 => x"398d5676",
          8803 => x"802e82c3",
          8804 => x"38821570",
          8805 => x"98160c7b",
          8806 => x"a0160c73",
          8807 => x"1c70a417",
          8808 => x"0c7a1dac",
          8809 => x"170c5455",
          8810 => x"76832e09",
          8811 => x"8106af38",
          8812 => x"80de1451",
          8813 => x"d9ae3f82",
          8814 => x"b5a80883",
          8815 => x"ffff0653",
          8816 => x"8d567282",
          8817 => x"8e387982",
          8818 => x"8a3880e0",
          8819 => x"1451d9ab",
          8820 => x"3f82b5a8",
          8821 => x"08a8150c",
          8822 => x"74822b53",
          8823 => x"a2398d56",
          8824 => x"79802e81",
          8825 => x"ee387713",
          8826 => x"a8150c74",
          8827 => x"15537682",
          8828 => x"2e8d3874",
          8829 => x"10157081",
          8830 => x"2a768106",
          8831 => x"05515383",
          8832 => x"ff13892a",
          8833 => x"538d5672",
          8834 => x"9c150826",
          8835 => x"81c538ff",
          8836 => x"0b90150c",
          8837 => x"ff0b8c15",
          8838 => x"0cff800b",
          8839 => x"84153476",
          8840 => x"832e0981",
          8841 => x"06819238",
          8842 => x"80e41451",
          8843 => x"d8b63f82",
          8844 => x"b5a80883",
          8845 => x"ffff0653",
          8846 => x"72812e09",
          8847 => x"810680f9",
          8848 => x"38811b52",
          8849 => x"7351dbb8",
          8850 => x"3f82b5a8",
          8851 => x"0880ea38",
          8852 => x"82b5a808",
          8853 => x"84153484",
          8854 => x"b21451d8",
          8855 => x"873f82b5",
          8856 => x"a80883ff",
          8857 => x"ff065372",
          8858 => x"82d4d52e",
          8859 => x"09810680",
          8860 => x"c838b414",
          8861 => x"51d8843f",
          8862 => x"82b5a808",
          8863 => x"848b85a4",
          8864 => x"d22e0981",
          8865 => x"06b33884",
          8866 => x"981451d7",
          8867 => x"ee3f82b5",
          8868 => x"a808868a",
          8869 => x"85e4f22e",
          8870 => x"0981069d",
          8871 => x"38849c14",
          8872 => x"51d7d83f",
          8873 => x"82b5a808",
          8874 => x"90150c84",
          8875 => x"a01451d7",
          8876 => x"ca3f82b5",
          8877 => x"a8088c15",
          8878 => x"0c767434",
          8879 => x"82ccf022",
          8880 => x"81055372",
          8881 => x"82ccf023",
          8882 => x"72861523",
          8883 => x"800b9415",
          8884 => x"0c805675",
          8885 => x"82b5a80c",
          8886 => x"903d0d04",
          8887 => x"fb3d0d77",
          8888 => x"54895573",
          8889 => x"802eb938",
          8890 => x"73085372",
          8891 => x"802eb138",
          8892 => x"72335271",
          8893 => x"802ea938",
          8894 => x"86132284",
          8895 => x"15225752",
          8896 => x"71762e09",
          8897 => x"81069938",
          8898 => x"81133351",
          8899 => x"d0c03f82",
          8900 => x"b5a80881",
          8901 => x"06527188",
          8902 => x"38717408",
          8903 => x"54558339",
          8904 => x"80537873",
          8905 => x"710c5274",
          8906 => x"82b5a80c",
          8907 => x"873d0d04",
          8908 => x"fa3d0d02",
          8909 => x"ab05337a",
          8910 => x"58893dfc",
          8911 => x"055256f4",
          8912 => x"e63f8b54",
          8913 => x"800b82b5",
          8914 => x"a80824bc",
          8915 => x"3882b5a8",
          8916 => x"08842982",
          8917 => x"cce00570",
          8918 => x"08555573",
          8919 => x"802e8438",
          8920 => x"80743478",
          8921 => x"5473802e",
          8922 => x"84388074",
          8923 => x"3478750c",
          8924 => x"75547580",
          8925 => x"2e923880",
          8926 => x"53893d70",
          8927 => x"53840551",
          8928 => x"f7b03f82",
          8929 => x"b5a80854",
          8930 => x"7382b5a8",
          8931 => x"0c883d0d",
          8932 => x"04eb3d0d",
          8933 => x"67028405",
          8934 => x"80e70533",
          8935 => x"59598954",
          8936 => x"78802e84",
          8937 => x"c83877bf",
          8938 => x"06705498",
          8939 => x"3dd00553",
          8940 => x"993d8405",
          8941 => x"5258f6fa",
          8942 => x"3f82b5a8",
          8943 => x"085582b5",
          8944 => x"a80884a4",
          8945 => x"387a5c68",
          8946 => x"528c3d70",
          8947 => x"5256edc6",
          8948 => x"3f82b5a8",
          8949 => x"085582b5",
          8950 => x"a8089238",
          8951 => x"0280d705",
          8952 => x"3370982b",
          8953 => x"55577380",
          8954 => x"25833886",
          8955 => x"55779c06",
          8956 => x"5473802e",
          8957 => x"81ab3874",
          8958 => x"802e9538",
          8959 => x"74842e09",
          8960 => x"8106aa38",
          8961 => x"7551eaf8",
          8962 => x"3f82b5a8",
          8963 => x"08559e39",
          8964 => x"02b20533",
          8965 => x"91065473",
          8966 => x"81b83877",
          8967 => x"822a7081",
          8968 => x"06515473",
          8969 => x"802e8e38",
          8970 => x"885583bc",
          8971 => x"39778807",
          8972 => x"587483b4",
          8973 => x"3877832a",
          8974 => x"70810651",
          8975 => x"5473802e",
          8976 => x"81af3862",
          8977 => x"527a51e8",
          8978 => x"a53f82b5",
          8979 => x"a8085682",
          8980 => x"88b20a52",
          8981 => x"628e0551",
          8982 => x"d4ea3f62",
          8983 => x"54a00b8b",
          8984 => x"15348053",
          8985 => x"62527a51",
          8986 => x"e8bd3f80",
          8987 => x"52629c05",
          8988 => x"51d4d13f",
          8989 => x"7a54810b",
          8990 => x"83153475",
          8991 => x"802e80f1",
          8992 => x"387ab011",
          8993 => x"08515480",
          8994 => x"53755297",
          8995 => x"3dd40551",
          8996 => x"ddbe3f82",
          8997 => x"b5a80855",
          8998 => x"82b5a808",
          8999 => x"82ca38b7",
          9000 => x"397482c4",
          9001 => x"3802b205",
          9002 => x"3370842a",
          9003 => x"70810651",
          9004 => x"55567380",
          9005 => x"2e863884",
          9006 => x"5582ad39",
          9007 => x"77812a70",
          9008 => x"81065154",
          9009 => x"73802ea9",
          9010 => x"38758106",
          9011 => x"5473802e",
          9012 => x"a0388755",
          9013 => x"82923973",
          9014 => x"527a51d6",
          9015 => x"a33f82b5",
          9016 => x"a8087bff",
          9017 => x"188c120c",
          9018 => x"555582b5",
          9019 => x"a80881f8",
          9020 => x"3877832a",
          9021 => x"70810651",
          9022 => x"5473802e",
          9023 => x"86387780",
          9024 => x"c007587a",
          9025 => x"b01108a0",
          9026 => x"1b0c63a4",
          9027 => x"1b0c6353",
          9028 => x"705257e6",
          9029 => x"d93f82b5",
          9030 => x"a80882b5",
          9031 => x"a808881b",
          9032 => x"0c639c05",
          9033 => x"525ad2d3",
          9034 => x"3f82b5a8",
          9035 => x"0882b5a8",
          9036 => x"088c1b0c",
          9037 => x"777a0c56",
          9038 => x"86172284",
          9039 => x"1a237790",
          9040 => x"1a34800b",
          9041 => x"911a3480",
          9042 => x"0b9c1a0c",
          9043 => x"800b941a",
          9044 => x"0c77852a",
          9045 => x"70810651",
          9046 => x"5473802e",
          9047 => x"818d3882",
          9048 => x"b5a80880",
          9049 => x"2e818438",
          9050 => x"82b5a808",
          9051 => x"941a0c8a",
          9052 => x"17227089",
          9053 => x"2b7b5259",
          9054 => x"57a83976",
          9055 => x"527851d7",
          9056 => x"9f3f82b5",
          9057 => x"a8085782",
          9058 => x"b5a80881",
          9059 => x"26833882",
          9060 => x"5582b5a8",
          9061 => x"08ff2e09",
          9062 => x"81068338",
          9063 => x"79557578",
          9064 => x"31567430",
          9065 => x"70760780",
          9066 => x"25515477",
          9067 => x"76278a38",
          9068 => x"81707506",
          9069 => x"555a73c3",
          9070 => x"3876981a",
          9071 => x"0c74a938",
          9072 => x"7583ff06",
          9073 => x"5473802e",
          9074 => x"a2387652",
          9075 => x"7a51d6a6",
          9076 => x"3f82b5a8",
          9077 => x"08853882",
          9078 => x"558e3975",
          9079 => x"892a82b5",
          9080 => x"a808059c",
          9081 => x"1a0c8439",
          9082 => x"80790c74",
          9083 => x"547382b5",
          9084 => x"a80c973d",
          9085 => x"0d04f23d",
          9086 => x"0d606365",
          9087 => x"6440405d",
          9088 => x"59807e0c",
          9089 => x"903dfc05",
          9090 => x"527851f9",
          9091 => x"cf3f82b5",
          9092 => x"a8085582",
          9093 => x"b5a8088a",
          9094 => x"38911933",
          9095 => x"5574802e",
          9096 => x"86387456",
          9097 => x"82c43990",
          9098 => x"19338106",
          9099 => x"55875674",
          9100 => x"802e82b6",
          9101 => x"38953982",
          9102 => x"0b911a34",
          9103 => x"825682aa",
          9104 => x"39810b91",
          9105 => x"1a348156",
          9106 => x"82a0398c",
          9107 => x"1908941a",
          9108 => x"08315574",
          9109 => x"7c278338",
          9110 => x"745c7b80",
          9111 => x"2e828938",
          9112 => x"94190870",
          9113 => x"83ff0656",
          9114 => x"567481b2",
          9115 => x"387e8a11",
          9116 => x"22ff0577",
          9117 => x"892a065b",
          9118 => x"5579a838",
          9119 => x"75873888",
          9120 => x"1908558f",
          9121 => x"39981908",
          9122 => x"527851d5",
          9123 => x"933f82b5",
          9124 => x"a8085581",
          9125 => x"7527ff9f",
          9126 => x"3874ff2e",
          9127 => x"ffa33874",
          9128 => x"981a0c98",
          9129 => x"1908527e",
          9130 => x"51d4cb3f",
          9131 => x"82b5a808",
          9132 => x"802eff83",
          9133 => x"3882b5a8",
          9134 => x"081a7c89",
          9135 => x"2a595777",
          9136 => x"802e80d6",
          9137 => x"38771a7f",
          9138 => x"8a112258",
          9139 => x"5c557575",
          9140 => x"27853875",
          9141 => x"7a315877",
          9142 => x"5476537c",
          9143 => x"52811b33",
          9144 => x"51ca883f",
          9145 => x"82b5a808",
          9146 => x"fed7387e",
          9147 => x"83113356",
          9148 => x"5674802e",
          9149 => x"9f38b016",
          9150 => x"08773155",
          9151 => x"74782794",
          9152 => x"38848053",
          9153 => x"b41652b0",
          9154 => x"16087731",
          9155 => x"892b7d05",
          9156 => x"51cfe03f",
          9157 => x"77892b56",
          9158 => x"b939769c",
          9159 => x"1a0c9419",
          9160 => x"0883ff06",
          9161 => x"84807131",
          9162 => x"57557b76",
          9163 => x"2783387b",
          9164 => x"569c1908",
          9165 => x"527e51d1",
          9166 => x"c73f82b5",
          9167 => x"a808fe81",
          9168 => x"38755394",
          9169 => x"190883ff",
          9170 => x"061fb405",
          9171 => x"527c51cf",
          9172 => x"a23f7b76",
          9173 => x"317e0817",
          9174 => x"7f0c761e",
          9175 => x"941b0818",
          9176 => x"941c0c5e",
          9177 => x"5cfdf339",
          9178 => x"80567582",
          9179 => x"b5a80c90",
          9180 => x"3d0d04f2",
          9181 => x"3d0d6063",
          9182 => x"65644040",
          9183 => x"5d58807e",
          9184 => x"0c903dfc",
          9185 => x"05527751",
          9186 => x"f6d23f82",
          9187 => x"b5a80855",
          9188 => x"82b5a808",
          9189 => x"8a389118",
          9190 => x"33557480",
          9191 => x"2e863874",
          9192 => x"5683b839",
          9193 => x"90183370",
          9194 => x"812a7081",
          9195 => x"06515656",
          9196 => x"87567480",
          9197 => x"2e83a438",
          9198 => x"9539820b",
          9199 => x"91193482",
          9200 => x"56839839",
          9201 => x"810b9119",
          9202 => x"34815683",
          9203 => x"8e399418",
          9204 => x"087c1156",
          9205 => x"56747627",
          9206 => x"84387509",
          9207 => x"5c7b802e",
          9208 => x"82ec3894",
          9209 => x"18087083",
          9210 => x"ff065656",
          9211 => x"7481fd38",
          9212 => x"7e8a1122",
          9213 => x"ff057789",
          9214 => x"2a065c55",
          9215 => x"7abf3875",
          9216 => x"8c388818",
          9217 => x"0855749c",
          9218 => x"387a5285",
          9219 => x"39981808",
          9220 => x"527751d7",
          9221 => x"e73f82b5",
          9222 => x"a8085582",
          9223 => x"b5a80880",
          9224 => x"2e82ab38",
          9225 => x"74812eff",
          9226 => x"913874ff",
          9227 => x"2eff9538",
          9228 => x"7498190c",
          9229 => x"88180885",
          9230 => x"38748819",
          9231 => x"0c7e55b0",
          9232 => x"15089c19",
          9233 => x"082e0981",
          9234 => x"068d3874",
          9235 => x"51cec13f",
          9236 => x"82b5a808",
          9237 => x"feee3898",
          9238 => x"1808527e",
          9239 => x"51d1973f",
          9240 => x"82b5a808",
          9241 => x"802efed2",
          9242 => x"3882b5a8",
          9243 => x"081b7c89",
          9244 => x"2a5a5778",
          9245 => x"802e80d5",
          9246 => x"38781b7f",
          9247 => x"8a112258",
          9248 => x"5b557575",
          9249 => x"27853875",
          9250 => x"7b315978",
          9251 => x"5476537c",
          9252 => x"52811a33",
          9253 => x"51c8be3f",
          9254 => x"82b5a808",
          9255 => x"fea6387e",
          9256 => x"b0110878",
          9257 => x"31565674",
          9258 => x"79279b38",
          9259 => x"848053b0",
          9260 => x"16087731",
          9261 => x"892b7d05",
          9262 => x"52b41651",
          9263 => x"ccb53f7e",
          9264 => x"55800b83",
          9265 => x"16347889",
          9266 => x"2b5680db",
          9267 => x"398c1808",
          9268 => x"94190826",
          9269 => x"93387e51",
          9270 => x"cdb63f82",
          9271 => x"b5a808fd",
          9272 => x"e3387e77",
          9273 => x"b0120c55",
          9274 => x"769c190c",
          9275 => x"94180883",
          9276 => x"ff068480",
          9277 => x"71315755",
          9278 => x"7b762783",
          9279 => x"387b569c",
          9280 => x"1808527e",
          9281 => x"51cdf93f",
          9282 => x"82b5a808",
          9283 => x"fdb63875",
          9284 => x"537c5294",
          9285 => x"180883ff",
          9286 => x"061fb405",
          9287 => x"51cbd43f",
          9288 => x"7e55810b",
          9289 => x"8316347b",
          9290 => x"76317e08",
          9291 => x"177f0c76",
          9292 => x"1e941a08",
          9293 => x"1870941c",
          9294 => x"0c8c1b08",
          9295 => x"58585e5c",
          9296 => x"74762783",
          9297 => x"38755574",
          9298 => x"8c190cfd",
          9299 => x"90399018",
          9300 => x"3380c007",
          9301 => x"55749019",
          9302 => x"34805675",
          9303 => x"82b5a80c",
          9304 => x"903d0d04",
          9305 => x"f83d0d7a",
          9306 => x"8b3dfc05",
          9307 => x"53705256",
          9308 => x"f2ea3f82",
          9309 => x"b5a80857",
          9310 => x"82b5a808",
          9311 => x"80fb3890",
          9312 => x"16337086",
          9313 => x"2a708106",
          9314 => x"51555573",
          9315 => x"802e80e9",
          9316 => x"38a01608",
          9317 => x"527851cc",
          9318 => x"e73f82b5",
          9319 => x"a8085782",
          9320 => x"b5a80880",
          9321 => x"d438a416",
          9322 => x"088b1133",
          9323 => x"a0075555",
          9324 => x"738b1634",
          9325 => x"88160853",
          9326 => x"74527508",
          9327 => x"51dde83f",
          9328 => x"8c160852",
          9329 => x"9c1551c9",
          9330 => x"fb3f8288",
          9331 => x"b20a5296",
          9332 => x"1551c9f0",
          9333 => x"3f765292",
          9334 => x"1551c9ca",
          9335 => x"3f785481",
          9336 => x"0b831534",
          9337 => x"7851ccdf",
          9338 => x"3f82b5a8",
          9339 => x"08901733",
          9340 => x"81bf0655",
          9341 => x"57739017",
          9342 => x"347682b5",
          9343 => x"a80c8a3d",
          9344 => x"0d04fc3d",
          9345 => x"0d767052",
          9346 => x"54fed93f",
          9347 => x"82b5a808",
          9348 => x"5382b5a8",
          9349 => x"089c3886",
          9350 => x"3dfc0552",
          9351 => x"7351f1bc",
          9352 => x"3f82b5a8",
          9353 => x"085382b5",
          9354 => x"a8088738",
          9355 => x"82b5a808",
          9356 => x"740c7282",
          9357 => x"b5a80c86",
          9358 => x"3d0d04ff",
          9359 => x"3d0d843d",
          9360 => x"51e6e43f",
          9361 => x"8b52800b",
          9362 => x"82b5a808",
          9363 => x"248b3882",
          9364 => x"b5a80882",
          9365 => x"ccf43480",
          9366 => x"527182b5",
          9367 => x"a80c833d",
          9368 => x"0d04ef3d",
          9369 => x"0d805393",
          9370 => x"3dd00552",
          9371 => x"943d51e9",
          9372 => x"c13f82b5",
          9373 => x"a8085582",
          9374 => x"b5a80880",
          9375 => x"e0387658",
          9376 => x"6352933d",
          9377 => x"d40551e0",
          9378 => x"8d3f82b5",
          9379 => x"a8085582",
          9380 => x"b5a808bc",
          9381 => x"380280c7",
          9382 => x"05337098",
          9383 => x"2b555673",
          9384 => x"80258938",
          9385 => x"767a9412",
          9386 => x"0c54b239",
          9387 => x"02a20533",
          9388 => x"70842a70",
          9389 => x"81065155",
          9390 => x"5673802e",
          9391 => x"9e38767f",
          9392 => x"53705254",
          9393 => x"dba83f82",
          9394 => x"b5a80894",
          9395 => x"150c8e39",
          9396 => x"82b5a808",
          9397 => x"842e0981",
          9398 => x"06833885",
          9399 => x"557482b5",
          9400 => x"a80c933d",
          9401 => x"0d04e43d",
          9402 => x"0d6f6f5b",
          9403 => x"5b807a34",
          9404 => x"80539e3d",
          9405 => x"ffb80552",
          9406 => x"9f3d51e8",
          9407 => x"b53f82b5",
          9408 => x"a8085782",
          9409 => x"b5a80882",
          9410 => x"fc387b43",
          9411 => x"7a7c9411",
          9412 => x"08475558",
          9413 => x"64547380",
          9414 => x"2e81ed38",
          9415 => x"a052933d",
          9416 => x"705255d5",
          9417 => x"ea3f82b5",
          9418 => x"a8085782",
          9419 => x"b5a80882",
          9420 => x"d4386852",
          9421 => x"7b51c9c8",
          9422 => x"3f82b5a8",
          9423 => x"085782b5",
          9424 => x"a80882c1",
          9425 => x"3869527b",
          9426 => x"51daa33f",
          9427 => x"82b5a808",
          9428 => x"45765274",
          9429 => x"51d5b83f",
          9430 => x"82b5a808",
          9431 => x"5782b5a8",
          9432 => x"0882a238",
          9433 => x"80527451",
          9434 => x"daeb3f82",
          9435 => x"b5a80857",
          9436 => x"82b5a808",
          9437 => x"a4386952",
          9438 => x"7b51d9f2",
          9439 => x"3f7382b5",
          9440 => x"a8082ea6",
          9441 => x"38765274",
          9442 => x"51d6cf3f",
          9443 => x"82b5a808",
          9444 => x"5782b5a8",
          9445 => x"08802ecc",
          9446 => x"3876842e",
          9447 => x"09810686",
          9448 => x"38825781",
          9449 => x"e0397681",
          9450 => x"dc389e3d",
          9451 => x"ffbc0552",
          9452 => x"7451dcc9",
          9453 => x"3f76903d",
          9454 => x"78118111",
          9455 => x"3351565a",
          9456 => x"5673802e",
          9457 => x"913802b9",
          9458 => x"05558116",
          9459 => x"81167033",
          9460 => x"56565673",
          9461 => x"f5388116",
          9462 => x"54737826",
          9463 => x"81903875",
          9464 => x"802e9938",
          9465 => x"78168105",
          9466 => x"55ff186f",
          9467 => x"11ff18ff",
          9468 => x"18585855",
          9469 => x"58743374",
          9470 => x"3475ee38",
          9471 => x"ff186f11",
          9472 => x"5558af74",
          9473 => x"34fe8d39",
          9474 => x"777b2e09",
          9475 => x"81068a38",
          9476 => x"ff186f11",
          9477 => x"5558af74",
          9478 => x"34800b82",
          9479 => x"ccf43370",
          9480 => x"842982ae",
          9481 => x"e0057008",
          9482 => x"7033525c",
          9483 => x"56565673",
          9484 => x"762e8d38",
          9485 => x"8116701a",
          9486 => x"70335155",
          9487 => x"5673f538",
          9488 => x"82165473",
          9489 => x"7826a738",
          9490 => x"80557476",
          9491 => x"27913874",
          9492 => x"19547333",
          9493 => x"7a708105",
          9494 => x"5c348115",
          9495 => x"55ec39ba",
          9496 => x"7a708105",
          9497 => x"5c3474ff",
          9498 => x"2e098106",
          9499 => x"85389157",
          9500 => x"94396e18",
          9501 => x"81195954",
          9502 => x"73337a70",
          9503 => x"81055c34",
          9504 => x"7a7826ee",
          9505 => x"38807a34",
          9506 => x"7682b5a8",
          9507 => x"0c9e3d0d",
          9508 => x"04f73d0d",
          9509 => x"7b7d8d3d",
          9510 => x"fc055471",
          9511 => x"535755ec",
          9512 => x"bb3f82b5",
          9513 => x"a8085382",
          9514 => x"b5a80882",
          9515 => x"fa389115",
          9516 => x"33537282",
          9517 => x"f2388c15",
          9518 => x"08547376",
          9519 => x"27923890",
          9520 => x"15337081",
          9521 => x"2a708106",
          9522 => x"51545772",
          9523 => x"83387356",
          9524 => x"94150854",
          9525 => x"80709417",
          9526 => x"0c587578",
          9527 => x"2e829738",
          9528 => x"798a1122",
          9529 => x"70892b59",
          9530 => x"51537378",
          9531 => x"2eb73876",
          9532 => x"52ff1651",
          9533 => x"fee8ac3f",
          9534 => x"82b5a808",
          9535 => x"ff157854",
          9536 => x"70535553",
          9537 => x"fee89c3f",
          9538 => x"82b5a808",
          9539 => x"73269638",
          9540 => x"76307075",
          9541 => x"06709418",
          9542 => x"0c777131",
          9543 => x"98180857",
          9544 => x"585153b1",
          9545 => x"39881508",
          9546 => x"5473a638",
          9547 => x"73527451",
          9548 => x"cdca3f82",
          9549 => x"b5a80854",
          9550 => x"82b5a808",
          9551 => x"812e819a",
          9552 => x"3882b5a8",
          9553 => x"08ff2e81",
          9554 => x"9b3882b5",
          9555 => x"a8088816",
          9556 => x"0c739816",
          9557 => x"0c73802e",
          9558 => x"819c3876",
          9559 => x"762780dc",
          9560 => x"38757731",
          9561 => x"94160818",
          9562 => x"94170c90",
          9563 => x"16337081",
          9564 => x"2a708106",
          9565 => x"51555a56",
          9566 => x"72802e9a",
          9567 => x"38735274",
          9568 => x"51ccf93f",
          9569 => x"82b5a808",
          9570 => x"5482b5a8",
          9571 => x"08943882",
          9572 => x"b5a80856",
          9573 => x"a7397352",
          9574 => x"7451c784",
          9575 => x"3f82b5a8",
          9576 => x"085473ff",
          9577 => x"2ebe3881",
          9578 => x"7427af38",
          9579 => x"79537398",
          9580 => x"140827a6",
          9581 => x"38739816",
          9582 => x"0cffa039",
          9583 => x"94150816",
          9584 => x"94160c75",
          9585 => x"83ff0653",
          9586 => x"72802eaa",
          9587 => x"38735279",
          9588 => x"51c6a33f",
          9589 => x"82b5a808",
          9590 => x"9438820b",
          9591 => x"91163482",
          9592 => x"5380c439",
          9593 => x"810b9116",
          9594 => x"348153bb",
          9595 => x"3975892a",
          9596 => x"82b5a808",
          9597 => x"05589415",
          9598 => x"08548c15",
          9599 => x"08742790",
          9600 => x"38738c16",
          9601 => x"0c901533",
          9602 => x"80c00753",
          9603 => x"72901634",
          9604 => x"7383ff06",
          9605 => x"5372802e",
          9606 => x"8c38779c",
          9607 => x"16082e85",
          9608 => x"38779c16",
          9609 => x"0c805372",
          9610 => x"82b5a80c",
          9611 => x"8b3d0d04",
          9612 => x"f93d0d79",
          9613 => x"56895475",
          9614 => x"802e818a",
          9615 => x"38805389",
          9616 => x"3dfc0552",
          9617 => x"8a3d8405",
          9618 => x"51e1e73f",
          9619 => x"82b5a808",
          9620 => x"5582b5a8",
          9621 => x"0880ea38",
          9622 => x"77760c7a",
          9623 => x"527551d8",
          9624 => x"b53f82b5",
          9625 => x"a8085582",
          9626 => x"b5a80880",
          9627 => x"c338ab16",
          9628 => x"3370982b",
          9629 => x"55578074",
          9630 => x"24a23886",
          9631 => x"16337084",
          9632 => x"2a708106",
          9633 => x"51555773",
          9634 => x"802ead38",
          9635 => x"9c160852",
          9636 => x"7751d3da",
          9637 => x"3f82b5a8",
          9638 => x"0888170c",
          9639 => x"77548614",
          9640 => x"22841723",
          9641 => x"74527551",
          9642 => x"cee53f82",
          9643 => x"b5a80855",
          9644 => x"74842e09",
          9645 => x"81068538",
          9646 => x"85558639",
          9647 => x"74802e84",
          9648 => x"3880760c",
          9649 => x"74547382",
          9650 => x"b5a80c89",
          9651 => x"3d0d04fc",
          9652 => x"3d0d7687",
          9653 => x"3dfc0553",
          9654 => x"705253e7",
          9655 => x"ff3f82b5",
          9656 => x"a8088738",
          9657 => x"82b5a808",
          9658 => x"730c863d",
          9659 => x"0d04fb3d",
          9660 => x"0d777989",
          9661 => x"3dfc0554",
          9662 => x"71535654",
          9663 => x"e7de3f82",
          9664 => x"b5a80853",
          9665 => x"82b5a808",
          9666 => x"80df3874",
          9667 => x"933882b5",
          9668 => x"a8085273",
          9669 => x"51cdf83f",
          9670 => x"82b5a808",
          9671 => x"5380ca39",
          9672 => x"82b5a808",
          9673 => x"527351d3",
          9674 => x"ac3f82b5",
          9675 => x"a8085382",
          9676 => x"b5a80884",
          9677 => x"2e098106",
          9678 => x"85388053",
          9679 => x"873982b5",
          9680 => x"a808a638",
          9681 => x"74527351",
          9682 => x"d5b33f72",
          9683 => x"527351cf",
          9684 => x"893f82b5",
          9685 => x"a8088432",
          9686 => x"70307072",
          9687 => x"079f2c70",
          9688 => x"82b5a808",
          9689 => x"06515154",
          9690 => x"547282b5",
          9691 => x"a80c873d",
          9692 => x"0d04ee3d",
          9693 => x"0d655780",
          9694 => x"53893d70",
          9695 => x"53963d52",
          9696 => x"56dfaf3f",
          9697 => x"82b5a808",
          9698 => x"5582b5a8",
          9699 => x"08b23864",
          9700 => x"527551d6",
          9701 => x"813f82b5",
          9702 => x"a8085582",
          9703 => x"b5a808a0",
          9704 => x"380280cb",
          9705 => x"05337098",
          9706 => x"2b555873",
          9707 => x"80258538",
          9708 => x"86558d39",
          9709 => x"76802e88",
          9710 => x"38765275",
          9711 => x"51d4be3f",
          9712 => x"7482b5a8",
          9713 => x"0c943d0d",
          9714 => x"04f03d0d",
          9715 => x"6365555c",
          9716 => x"8053923d",
          9717 => x"ec055293",
          9718 => x"3d51ded6",
          9719 => x"3f82b5a8",
          9720 => x"085b82b5",
          9721 => x"a8088280",
          9722 => x"387c740c",
          9723 => x"73089811",
          9724 => x"08fe1190",
          9725 => x"13085956",
          9726 => x"58557574",
          9727 => x"26913875",
          9728 => x"7c0c81e4",
          9729 => x"39815b81",
          9730 => x"cc39825b",
          9731 => x"81c73982",
          9732 => x"b5a80875",
          9733 => x"33555973",
          9734 => x"812e0981",
          9735 => x"06bf3882",
          9736 => x"755f5776",
          9737 => x"52923df0",
          9738 => x"0551c1f4",
          9739 => x"3f82b5a8",
          9740 => x"08ff2ed1",
          9741 => x"3882b5a8",
          9742 => x"08812ece",
          9743 => x"3882b5a8",
          9744 => x"08307082",
          9745 => x"b5a80807",
          9746 => x"80257a05",
          9747 => x"81197f53",
          9748 => x"595a5498",
          9749 => x"14087726",
          9750 => x"ca3880f9",
          9751 => x"39a41508",
          9752 => x"82b5a808",
          9753 => x"57587598",
          9754 => x"38775281",
          9755 => x"187d5258",
          9756 => x"ffbf8d3f",
          9757 => x"82b5a808",
          9758 => x"5b82b5a8",
          9759 => x"0880d638",
          9760 => x"7c703377",
          9761 => x"12ff1a5d",
          9762 => x"52565474",
          9763 => x"822e0981",
          9764 => x"069e38b4",
          9765 => x"1451ffbb",
          9766 => x"cb3f82b5",
          9767 => x"a80883ff",
          9768 => x"ff067030",
          9769 => x"7080251b",
          9770 => x"8219595b",
          9771 => x"51549b39",
          9772 => x"b41451ff",
          9773 => x"bbc53f82",
          9774 => x"b5a808f0",
          9775 => x"0a067030",
          9776 => x"7080251b",
          9777 => x"8419595b",
          9778 => x"51547583",
          9779 => x"ff067a58",
          9780 => x"5679ff92",
          9781 => x"38787c0c",
          9782 => x"7c799012",
          9783 => x"0c841133",
          9784 => x"81075654",
          9785 => x"74841534",
          9786 => x"7a82b5a8",
          9787 => x"0c923d0d",
          9788 => x"04f93d0d",
          9789 => x"798a3dfc",
          9790 => x"05537052",
          9791 => x"57e3dd3f",
          9792 => x"82b5a808",
          9793 => x"5682b5a8",
          9794 => x"0881a838",
          9795 => x"91173356",
          9796 => x"7581a038",
          9797 => x"90173370",
          9798 => x"812a7081",
          9799 => x"06515555",
          9800 => x"87557380",
          9801 => x"2e818e38",
          9802 => x"94170854",
          9803 => x"738c1808",
          9804 => x"27818038",
          9805 => x"739b3882",
          9806 => x"b5a80853",
          9807 => x"88170852",
          9808 => x"7651c48c",
          9809 => x"3f82b5a8",
          9810 => x"08748819",
          9811 => x"0c5680c9",
          9812 => x"39981708",
          9813 => x"527651ff",
          9814 => x"bfc63f82",
          9815 => x"b5a808ff",
          9816 => x"2e098106",
          9817 => x"83388156",
          9818 => x"82b5a808",
          9819 => x"812e0981",
          9820 => x"06853882",
          9821 => x"56a33975",
          9822 => x"a0387754",
          9823 => x"82b5a808",
          9824 => x"98150827",
          9825 => x"94389817",
          9826 => x"085382b5",
          9827 => x"a8085276",
          9828 => x"51c3bd3f",
          9829 => x"82b5a808",
          9830 => x"56941708",
          9831 => x"8c180c90",
          9832 => x"173380c0",
          9833 => x"07547390",
          9834 => x"18347580",
          9835 => x"2e853875",
          9836 => x"91183475",
          9837 => x"557482b5",
          9838 => x"a80c893d",
          9839 => x"0d04e23d",
          9840 => x"0d8253a0",
          9841 => x"3dffa405",
          9842 => x"52a13d51",
          9843 => x"dae43f82",
          9844 => x"b5a80855",
          9845 => x"82b5a808",
          9846 => x"81f53878",
          9847 => x"45a13d08",
          9848 => x"52953d70",
          9849 => x"5258d1ae",
          9850 => x"3f82b5a8",
          9851 => x"085582b5",
          9852 => x"a80881db",
          9853 => x"380280fb",
          9854 => x"05337085",
          9855 => x"2a708106",
          9856 => x"51555686",
          9857 => x"557381c7",
          9858 => x"3875982b",
          9859 => x"54807424",
          9860 => x"81bd3802",
          9861 => x"80d60533",
          9862 => x"70810658",
          9863 => x"54875576",
          9864 => x"81ad386b",
          9865 => x"527851cc",
          9866 => x"c53f82b5",
          9867 => x"a8087484",
          9868 => x"2a708106",
          9869 => x"51555673",
          9870 => x"802e80d4",
          9871 => x"38785482",
          9872 => x"b5a80894",
          9873 => x"15082e81",
          9874 => x"8638735a",
          9875 => x"82b5a808",
          9876 => x"5c76528a",
          9877 => x"3d705254",
          9878 => x"c7b53f82",
          9879 => x"b5a80855",
          9880 => x"82b5a808",
          9881 => x"80e93882",
          9882 => x"b5a80852",
          9883 => x"7351cce5",
          9884 => x"3f82b5a8",
          9885 => x"085582b5",
          9886 => x"a8088638",
          9887 => x"875580cf",
          9888 => x"3982b5a8",
          9889 => x"08842e88",
          9890 => x"3882b5a8",
          9891 => x"0880c038",
          9892 => x"7751cec2",
          9893 => x"3f82b5a8",
          9894 => x"0882b5a8",
          9895 => x"08307082",
          9896 => x"b5a80807",
          9897 => x"80255155",
          9898 => x"5575802e",
          9899 => x"94387380",
          9900 => x"2e8f3880",
          9901 => x"53755277",
          9902 => x"51c1953f",
          9903 => x"82b5a808",
          9904 => x"55748c38",
          9905 => x"7851ffba",
          9906 => x"fe3f82b5",
          9907 => x"a8085574",
          9908 => x"82b5a80c",
          9909 => x"a03d0d04",
          9910 => x"e93d0d82",
          9911 => x"53993dc0",
          9912 => x"05529a3d",
          9913 => x"51d8cb3f",
          9914 => x"82b5a808",
          9915 => x"5482b5a8",
          9916 => x"0882b038",
          9917 => x"785e6952",
          9918 => x"8e3d7052",
          9919 => x"58cf973f",
          9920 => x"82b5a808",
          9921 => x"5482b5a8",
          9922 => x"08863888",
          9923 => x"54829439",
          9924 => x"82b5a808",
          9925 => x"842e0981",
          9926 => x"06828838",
          9927 => x"0280df05",
          9928 => x"3370852a",
          9929 => x"81065155",
          9930 => x"86547481",
          9931 => x"f638785a",
          9932 => x"74528a3d",
          9933 => x"705257c1",
          9934 => x"c33f82b5",
          9935 => x"a8087555",
          9936 => x"5682b5a8",
          9937 => x"08833887",
          9938 => x"5482b5a8",
          9939 => x"08812e09",
          9940 => x"81068338",
          9941 => x"825482b5",
          9942 => x"a808ff2e",
          9943 => x"09810686",
          9944 => x"38815481",
          9945 => x"b4397381",
          9946 => x"b03882b5",
          9947 => x"a8085278",
          9948 => x"51c4a43f",
          9949 => x"82b5a808",
          9950 => x"5482b5a8",
          9951 => x"08819a38",
          9952 => x"8b53a052",
          9953 => x"b41951ff",
          9954 => x"b78c3f78",
          9955 => x"54ae0bb4",
          9956 => x"15347854",
          9957 => x"900bbf15",
          9958 => x"348288b2",
          9959 => x"0a5280ca",
          9960 => x"1951ffb6",
          9961 => x"9f3f7553",
          9962 => x"78b41153",
          9963 => x"51c9f83f",
          9964 => x"a05378b4",
          9965 => x"115380d4",
          9966 => x"0551ffb6",
          9967 => x"b63f7854",
          9968 => x"ae0b80d5",
          9969 => x"15347f53",
          9970 => x"7880d411",
          9971 => x"5351c9d7",
          9972 => x"3f785481",
          9973 => x"0b831534",
          9974 => x"7751cba4",
          9975 => x"3f82b5a8",
          9976 => x"085482b5",
          9977 => x"a808b238",
          9978 => x"8288b20a",
          9979 => x"52649605",
          9980 => x"51ffb5d0",
          9981 => x"3f755364",
          9982 => x"527851c9",
          9983 => x"aa3f6454",
          9984 => x"900b8b15",
          9985 => x"34785481",
          9986 => x"0b831534",
          9987 => x"7851ffb8",
          9988 => x"b63f82b5",
          9989 => x"a808548b",
          9990 => x"39805375",
          9991 => x"527651ff",
          9992 => x"beae3f73",
          9993 => x"82b5a80c",
          9994 => x"993d0d04",
          9995 => x"da3d0da9",
          9996 => x"3d840551",
          9997 => x"d2f13f82",
          9998 => x"53a83dff",
          9999 => x"840552a9",
         10000 => x"3d51d5ee",
         10001 => x"3f82b5a8",
         10002 => x"085582b5",
         10003 => x"a80882d3",
         10004 => x"38784da9",
         10005 => x"3d08529d",
         10006 => x"3d705258",
         10007 => x"ccb83f82",
         10008 => x"b5a80855",
         10009 => x"82b5a808",
         10010 => x"82b93802",
         10011 => x"819b0533",
         10012 => x"81a00654",
         10013 => x"86557382",
         10014 => x"aa38a053",
         10015 => x"a43d0852",
         10016 => x"a83dff88",
         10017 => x"0551ffb4",
         10018 => x"ea3fac53",
         10019 => x"7752923d",
         10020 => x"705254ff",
         10021 => x"b4dd3faa",
         10022 => x"3d085273",
         10023 => x"51cbf73f",
         10024 => x"82b5a808",
         10025 => x"5582b5a8",
         10026 => x"08953863",
         10027 => x"6f2e0981",
         10028 => x"06883865",
         10029 => x"a23d082e",
         10030 => x"92388855",
         10031 => x"81e53982",
         10032 => x"b5a80884",
         10033 => x"2e098106",
         10034 => x"81b83873",
         10035 => x"51c9b13f",
         10036 => x"82b5a808",
         10037 => x"5582b5a8",
         10038 => x"0881c838",
         10039 => x"68569353",
         10040 => x"a83dff95",
         10041 => x"05528d16",
         10042 => x"51ffb487",
         10043 => x"3f02af05",
         10044 => x"338b1734",
         10045 => x"8b163370",
         10046 => x"842a7081",
         10047 => x"06515555",
         10048 => x"73893874",
         10049 => x"a0075473",
         10050 => x"8b173478",
         10051 => x"54810b83",
         10052 => x"15348b16",
         10053 => x"3370842a",
         10054 => x"70810651",
         10055 => x"55557380",
         10056 => x"2e80e538",
         10057 => x"6e642e80",
         10058 => x"df387552",
         10059 => x"7851c6be",
         10060 => x"3f82b5a8",
         10061 => x"08527851",
         10062 => x"ffb7bb3f",
         10063 => x"825582b5",
         10064 => x"a808802e",
         10065 => x"80dd3882",
         10066 => x"b5a80852",
         10067 => x"7851ffb5",
         10068 => x"af3f82b5",
         10069 => x"a8087980",
         10070 => x"d4115858",
         10071 => x"5582b5a8",
         10072 => x"0880c038",
         10073 => x"81163354",
         10074 => x"73ae2e09",
         10075 => x"81069938",
         10076 => x"63537552",
         10077 => x"7651c6af",
         10078 => x"3f785481",
         10079 => x"0b831534",
         10080 => x"873982b5",
         10081 => x"a8089c38",
         10082 => x"7751c8ca",
         10083 => x"3f82b5a8",
         10084 => x"085582b5",
         10085 => x"a8088c38",
         10086 => x"7851ffb5",
         10087 => x"aa3f82b5",
         10088 => x"a8085574",
         10089 => x"82b5a80c",
         10090 => x"a83d0d04",
         10091 => x"ed3d0d02",
         10092 => x"80db0533",
         10093 => x"02840580",
         10094 => x"df053357",
         10095 => x"57825395",
         10096 => x"3dd00552",
         10097 => x"963d51d2",
         10098 => x"e93f82b5",
         10099 => x"a8085582",
         10100 => x"b5a80880",
         10101 => x"cf38785a",
         10102 => x"6552953d",
         10103 => x"d40551c9",
         10104 => x"b53f82b5",
         10105 => x"a8085582",
         10106 => x"b5a808b8",
         10107 => x"380280cf",
         10108 => x"053381a0",
         10109 => x"06548655",
         10110 => x"73aa3875",
         10111 => x"a7066171",
         10112 => x"098b1233",
         10113 => x"71067a74",
         10114 => x"06075157",
         10115 => x"5556748b",
         10116 => x"15347854",
         10117 => x"810b8315",
         10118 => x"347851ff",
         10119 => x"b4a93f82",
         10120 => x"b5a80855",
         10121 => x"7482b5a8",
         10122 => x"0c953d0d",
         10123 => x"04ef3d0d",
         10124 => x"64568253",
         10125 => x"933dd005",
         10126 => x"52943d51",
         10127 => x"d1f43f82",
         10128 => x"b5a80855",
         10129 => x"82b5a808",
         10130 => x"80cb3876",
         10131 => x"58635293",
         10132 => x"3dd40551",
         10133 => x"c8c03f82",
         10134 => x"b5a80855",
         10135 => x"82b5a808",
         10136 => x"b4380280",
         10137 => x"c7053381",
         10138 => x"a0065486",
         10139 => x"5573a638",
         10140 => x"84162286",
         10141 => x"17227190",
         10142 => x"2b075354",
         10143 => x"961f51ff",
         10144 => x"b0c23f76",
         10145 => x"54810b83",
         10146 => x"15347651",
         10147 => x"ffb3b83f",
         10148 => x"82b5a808",
         10149 => x"557482b5",
         10150 => x"a80c933d",
         10151 => x"0d04ea3d",
         10152 => x"0d696b5c",
         10153 => x"5a805398",
         10154 => x"3dd00552",
         10155 => x"993d51d1",
         10156 => x"813f82b5",
         10157 => x"a80882b5",
         10158 => x"a8083070",
         10159 => x"82b5a808",
         10160 => x"07802551",
         10161 => x"55577980",
         10162 => x"2e818538",
         10163 => x"81707506",
         10164 => x"55557380",
         10165 => x"2e80f938",
         10166 => x"7b5d805f",
         10167 => x"80528d3d",
         10168 => x"705254ff",
         10169 => x"bea93f82",
         10170 => x"b5a80857",
         10171 => x"82b5a808",
         10172 => x"80d13874",
         10173 => x"527351c3",
         10174 => x"dc3f82b5",
         10175 => x"a8085782",
         10176 => x"b5a808bf",
         10177 => x"3882b5a8",
         10178 => x"0882b5a8",
         10179 => x"08655b59",
         10180 => x"56781881",
         10181 => x"197b1856",
         10182 => x"59557433",
         10183 => x"74348116",
         10184 => x"568a7827",
         10185 => x"ec388b56",
         10186 => x"751a5480",
         10187 => x"74347580",
         10188 => x"2e9e38ff",
         10189 => x"16701b70",
         10190 => x"33515556",
         10191 => x"73a02ee8",
         10192 => x"388e3976",
         10193 => x"842e0981",
         10194 => x"06863880",
         10195 => x"7a348057",
         10196 => x"76307078",
         10197 => x"07802551",
         10198 => x"547a802e",
         10199 => x"80c13873",
         10200 => x"802ebc38",
         10201 => x"7ba01108",
         10202 => x"5351ffb1",
         10203 => x"933f82b5",
         10204 => x"a8085782",
         10205 => x"b5a808a7",
         10206 => x"387b7033",
         10207 => x"555580c3",
         10208 => x"5673832e",
         10209 => x"8b3880e4",
         10210 => x"5673842e",
         10211 => x"8338a756",
         10212 => x"7515b405",
         10213 => x"51ffade3",
         10214 => x"3f82b5a8",
         10215 => x"087b0c76",
         10216 => x"82b5a80c",
         10217 => x"983d0d04",
         10218 => x"e63d0d82",
         10219 => x"539c3dff",
         10220 => x"b805529d",
         10221 => x"3d51cefa",
         10222 => x"3f82b5a8",
         10223 => x"0882b5a8",
         10224 => x"08565482",
         10225 => x"b5a80883",
         10226 => x"98388b53",
         10227 => x"a0528b3d",
         10228 => x"705259ff",
         10229 => x"aec03f73",
         10230 => x"6d703370",
         10231 => x"81ff0652",
         10232 => x"5755579f",
         10233 => x"742781bc",
         10234 => x"38785874",
         10235 => x"81ff066d",
         10236 => x"81054e70",
         10237 => x"5255ffaf",
         10238 => x"893f82b5",
         10239 => x"a808802e",
         10240 => x"a5386c70",
         10241 => x"33705357",
         10242 => x"54ffaefd",
         10243 => x"3f82b5a8",
         10244 => x"08802e8d",
         10245 => x"3874882b",
         10246 => x"76076d81",
         10247 => x"054e5586",
         10248 => x"3982b5a8",
         10249 => x"0855ff9f",
         10250 => x"157083ff",
         10251 => x"ff065154",
         10252 => x"7399268a",
         10253 => x"38e01570",
         10254 => x"83ffff06",
         10255 => x"565480ff",
         10256 => x"75278738",
         10257 => x"82adf015",
         10258 => x"33557480",
         10259 => x"2ea33874",
         10260 => x"5282aff0",
         10261 => x"51ffae89",
         10262 => x"3f82b5a8",
         10263 => x"08933881",
         10264 => x"ff752788",
         10265 => x"38768926",
         10266 => x"88388b39",
         10267 => x"8a772786",
         10268 => x"38865581",
         10269 => x"ec3981ff",
         10270 => x"75278f38",
         10271 => x"74882a54",
         10272 => x"73787081",
         10273 => x"055a3481",
         10274 => x"17577478",
         10275 => x"7081055a",
         10276 => x"3481176d",
         10277 => x"70337081",
         10278 => x"ff065257",
         10279 => x"5557739f",
         10280 => x"26fec838",
         10281 => x"8b3d3354",
         10282 => x"86557381",
         10283 => x"e52e81b1",
         10284 => x"3876802e",
         10285 => x"993802a7",
         10286 => x"05557615",
         10287 => x"70335154",
         10288 => x"73a02e09",
         10289 => x"81068738",
         10290 => x"ff175776",
         10291 => x"ed387941",
         10292 => x"80438052",
         10293 => x"913d7052",
         10294 => x"55ffbab3",
         10295 => x"3f82b5a8",
         10296 => x"085482b5",
         10297 => x"a80880f7",
         10298 => x"38815274",
         10299 => x"51ffbfe5",
         10300 => x"3f82b5a8",
         10301 => x"085482b5",
         10302 => x"a8088d38",
         10303 => x"7680c438",
         10304 => x"6754e574",
         10305 => x"3480c639",
         10306 => x"82b5a808",
         10307 => x"842e0981",
         10308 => x"0680cc38",
         10309 => x"80547674",
         10310 => x"2e80c438",
         10311 => x"81527451",
         10312 => x"ffbdb03f",
         10313 => x"82b5a808",
         10314 => x"5482b5a8",
         10315 => x"08b138a0",
         10316 => x"5382b5a8",
         10317 => x"08526751",
         10318 => x"ffabdb3f",
         10319 => x"6754880b",
         10320 => x"8b15348b",
         10321 => x"53785267",
         10322 => x"51ffaba7",
         10323 => x"3f795481",
         10324 => x"0b831534",
         10325 => x"7951ffad",
         10326 => x"ee3f82b5",
         10327 => x"a8085473",
         10328 => x"557482b5",
         10329 => x"a80c9c3d",
         10330 => x"0d04f23d",
         10331 => x"0d606202",
         10332 => x"880580cb",
         10333 => x"0533933d",
         10334 => x"fc055572",
         10335 => x"54405e5a",
         10336 => x"d2da3f82",
         10337 => x"b5a80858",
         10338 => x"82b5a808",
         10339 => x"82bd3891",
         10340 => x"1a335877",
         10341 => x"82b5387c",
         10342 => x"802e9738",
         10343 => x"8c1a0859",
         10344 => x"78903890",
         10345 => x"1a337081",
         10346 => x"2a708106",
         10347 => x"51555573",
         10348 => x"90388754",
         10349 => x"82973982",
         10350 => x"58829039",
         10351 => x"8158828b",
         10352 => x"397e8a11",
         10353 => x"2270892b",
         10354 => x"70557f54",
         10355 => x"565656fe",
         10356 => x"ced13fff",
         10357 => x"147d0670",
         10358 => x"30707207",
         10359 => x"9f2a82b5",
         10360 => x"a808058c",
         10361 => x"19087c40",
         10362 => x"5a5d5555",
         10363 => x"81772788",
         10364 => x"38981608",
         10365 => x"77268338",
         10366 => x"82577677",
         10367 => x"56598056",
         10368 => x"74527951",
         10369 => x"ffae993f",
         10370 => x"81157f55",
         10371 => x"55981408",
         10372 => x"75268338",
         10373 => x"825582b5",
         10374 => x"a808812e",
         10375 => x"ff993882",
         10376 => x"b5a808ff",
         10377 => x"2eff9538",
         10378 => x"82b5a808",
         10379 => x"8e388116",
         10380 => x"56757b2e",
         10381 => x"09810687",
         10382 => x"38933974",
         10383 => x"59805674",
         10384 => x"772e0981",
         10385 => x"06ffb938",
         10386 => x"875880ff",
         10387 => x"397d802e",
         10388 => x"ba38787b",
         10389 => x"55557a80",
         10390 => x"2eb43881",
         10391 => x"15567381",
         10392 => x"2e098106",
         10393 => x"8338ff56",
         10394 => x"75537452",
         10395 => x"7e51ffaf",
         10396 => x"a83f82b5",
         10397 => x"a8085882",
         10398 => x"b5a80880",
         10399 => x"ce387481",
         10400 => x"16ff1656",
         10401 => x"565c73d3",
         10402 => x"388439ff",
         10403 => x"195c7e7c",
         10404 => x"8c120c55",
         10405 => x"7d802eb3",
         10406 => x"3878881b",
         10407 => x"0c7c8c1b",
         10408 => x"0c901a33",
         10409 => x"80c00754",
         10410 => x"73901b34",
         10411 => x"981508fe",
         10412 => x"05901608",
         10413 => x"57547574",
         10414 => x"26913875",
         10415 => x"7b319016",
         10416 => x"0c841533",
         10417 => x"81075473",
         10418 => x"84163477",
         10419 => x"547382b5",
         10420 => x"a80c903d",
         10421 => x"0d04e93d",
         10422 => x"0d6b6d02",
         10423 => x"880580eb",
         10424 => x"05339d3d",
         10425 => x"545a5c59",
         10426 => x"c5bd3f8b",
         10427 => x"56800b82",
         10428 => x"b5a80824",
         10429 => x"8bf83882",
         10430 => x"b5a80884",
         10431 => x"2982cce0",
         10432 => x"05700851",
         10433 => x"5574802e",
         10434 => x"84388075",
         10435 => x"3482b5a8",
         10436 => x"0881ff06",
         10437 => x"5f81527e",
         10438 => x"51ffa0d0",
         10439 => x"3f82b5a8",
         10440 => x"0881ff06",
         10441 => x"70810656",
         10442 => x"57835674",
         10443 => x"8bc03876",
         10444 => x"822a7081",
         10445 => x"0651558a",
         10446 => x"56748bb2",
         10447 => x"38993dfc",
         10448 => x"05538352",
         10449 => x"7e51ffa4",
         10450 => x"f03f82b5",
         10451 => x"a8089938",
         10452 => x"67557480",
         10453 => x"2e923874",
         10454 => x"82808026",
         10455 => x"8b38ff15",
         10456 => x"75065574",
         10457 => x"802e8338",
         10458 => x"81487880",
         10459 => x"2e873884",
         10460 => x"80792692",
         10461 => x"38788180",
         10462 => x"0a268b38",
         10463 => x"ff197906",
         10464 => x"5574802e",
         10465 => x"86389356",
         10466 => x"8ae43978",
         10467 => x"892a6e89",
         10468 => x"2a70892b",
         10469 => x"77594843",
         10470 => x"597a8338",
         10471 => x"81566130",
         10472 => x"70802577",
         10473 => x"07515591",
         10474 => x"56748ac2",
         10475 => x"38993df8",
         10476 => x"05538152",
         10477 => x"7e51ffa4",
         10478 => x"803f8156",
         10479 => x"82b5a808",
         10480 => x"8aac3877",
         10481 => x"832a7077",
         10482 => x"0682b5a8",
         10483 => x"08435645",
         10484 => x"748338bf",
         10485 => x"4166558e",
         10486 => x"56607526",
         10487 => x"8a903874",
         10488 => x"61317048",
         10489 => x"5580ff75",
         10490 => x"278a8338",
         10491 => x"93567881",
         10492 => x"802689fa",
         10493 => x"3877812a",
         10494 => x"70810656",
         10495 => x"4374802e",
         10496 => x"95387787",
         10497 => x"06557482",
         10498 => x"2e838d38",
         10499 => x"77810655",
         10500 => x"74802e83",
         10501 => x"83387781",
         10502 => x"06559356",
         10503 => x"825e7480",
         10504 => x"2e89cb38",
         10505 => x"785a7d83",
         10506 => x"2e098106",
         10507 => x"80e13878",
         10508 => x"ae386691",
         10509 => x"2a57810b",
         10510 => x"82b09422",
         10511 => x"565a7480",
         10512 => x"2e9d3874",
         10513 => x"77269838",
         10514 => x"82b09456",
         10515 => x"79108217",
         10516 => x"70225757",
         10517 => x"5a74802e",
         10518 => x"86387675",
         10519 => x"27ee3879",
         10520 => x"526651fe",
         10521 => x"c9bd3f82",
         10522 => x"b5a80884",
         10523 => x"29848705",
         10524 => x"70892a5e",
         10525 => x"55a05c80",
         10526 => x"0b82b5a8",
         10527 => x"08fc808a",
         10528 => x"055644fd",
         10529 => x"fff00a75",
         10530 => x"2780ec38",
         10531 => x"88d33978",
         10532 => x"ae38668c",
         10533 => x"2a57810b",
         10534 => x"82b08422",
         10535 => x"565a7480",
         10536 => x"2e9d3874",
         10537 => x"77269838",
         10538 => x"82b08456",
         10539 => x"79108217",
         10540 => x"70225757",
         10541 => x"5a74802e",
         10542 => x"86387675",
         10543 => x"27ee3879",
         10544 => x"526651fe",
         10545 => x"c8dd3f82",
         10546 => x"b5a80810",
         10547 => x"84055782",
         10548 => x"b5a8089f",
         10549 => x"f5269638",
         10550 => x"810b82b5",
         10551 => x"a8081082",
         10552 => x"b5a80805",
         10553 => x"7111722a",
         10554 => x"83055956",
         10555 => x"5e83ff17",
         10556 => x"892a5d81",
         10557 => x"5ca04460",
         10558 => x"1c7d1165",
         10559 => x"05697012",
         10560 => x"ff057130",
         10561 => x"70720674",
         10562 => x"315c5259",
         10563 => x"5759407d",
         10564 => x"832e0981",
         10565 => x"06893876",
         10566 => x"1c601841",
         10567 => x"5c843976",
         10568 => x"1d5d7990",
         10569 => x"29187062",
         10570 => x"31685851",
         10571 => x"55747626",
         10572 => x"87af3875",
         10573 => x"7c317d31",
         10574 => x"7a537065",
         10575 => x"315255fe",
         10576 => x"c7e13f82",
         10577 => x"b5a80858",
         10578 => x"7d832e09",
         10579 => x"81069b38",
         10580 => x"82b5a808",
         10581 => x"83fff526",
         10582 => x"80dd3878",
         10583 => x"87833879",
         10584 => x"812a5978",
         10585 => x"fdbe3886",
         10586 => x"f8397d82",
         10587 => x"2e098106",
         10588 => x"80c53883",
         10589 => x"fff50b82",
         10590 => x"b5a80827",
         10591 => x"a038788f",
         10592 => x"38791a55",
         10593 => x"7480c026",
         10594 => x"86387459",
         10595 => x"fd963962",
         10596 => x"81065574",
         10597 => x"802e8f38",
         10598 => x"835efd88",
         10599 => x"3982b5a8",
         10600 => x"089ff526",
         10601 => x"92387886",
         10602 => x"b838791a",
         10603 => x"59818079",
         10604 => x"27fcf138",
         10605 => x"86ab3980",
         10606 => x"557d812e",
         10607 => x"09810683",
         10608 => x"387d559f",
         10609 => x"f578278b",
         10610 => x"38748106",
         10611 => x"558e5674",
         10612 => x"869c3884",
         10613 => x"80538052",
         10614 => x"7a51ffa2",
         10615 => x"b93f8b53",
         10616 => x"82aeac52",
         10617 => x"7a51ffa2",
         10618 => x"8a3f8480",
         10619 => x"528b1b51",
         10620 => x"ffa1b33f",
         10621 => x"798d1c34",
         10622 => x"7b83ffff",
         10623 => x"06528e1b",
         10624 => x"51ffa1a2",
         10625 => x"3f810b90",
         10626 => x"1c347d83",
         10627 => x"32703070",
         10628 => x"962a8480",
         10629 => x"06545155",
         10630 => x"911b51ff",
         10631 => x"a1883f66",
         10632 => x"557483ff",
         10633 => x"ff269038",
         10634 => x"7483ffff",
         10635 => x"0652931b",
         10636 => x"51ffa0f2",
         10637 => x"3f8a3974",
         10638 => x"52a01b51",
         10639 => x"ffa1853f",
         10640 => x"f80b951c",
         10641 => x"34bf5298",
         10642 => x"1b51ffa0",
         10643 => x"d93f81ff",
         10644 => x"529a1b51",
         10645 => x"ffa0cf3f",
         10646 => x"60529c1b",
         10647 => x"51ffa0e4",
         10648 => x"3f7d832e",
         10649 => x"09810680",
         10650 => x"cb388288",
         10651 => x"b20a5280",
         10652 => x"c31b51ff",
         10653 => x"a0ce3f7c",
         10654 => x"52a41b51",
         10655 => x"ffa0c53f",
         10656 => x"8252ac1b",
         10657 => x"51ffa0bc",
         10658 => x"3f8152b0",
         10659 => x"1b51ffa0",
         10660 => x"953f8652",
         10661 => x"b21b51ff",
         10662 => x"a08c3fff",
         10663 => x"800b80c0",
         10664 => x"1c34a90b",
         10665 => x"80c21c34",
         10666 => x"935382ae",
         10667 => x"b85280c7",
         10668 => x"1b51ae39",
         10669 => x"8288b20a",
         10670 => x"52a71b51",
         10671 => x"ffa0853f",
         10672 => x"7c83ffff",
         10673 => x"0652961b",
         10674 => x"51ff9fda",
         10675 => x"3fff800b",
         10676 => x"a41c34a9",
         10677 => x"0ba61c34",
         10678 => x"935382ae",
         10679 => x"cc52ab1b",
         10680 => x"51ffa08f",
         10681 => x"3f82d4d5",
         10682 => x"5283fe1b",
         10683 => x"705259ff",
         10684 => x"9fb43f81",
         10685 => x"5460537a",
         10686 => x"527e51ff",
         10687 => x"9bd73f81",
         10688 => x"5682b5a8",
         10689 => x"0883e738",
         10690 => x"7d832e09",
         10691 => x"810680ee",
         10692 => x"38755460",
         10693 => x"8605537a",
         10694 => x"527e51ff",
         10695 => x"9bb73f84",
         10696 => x"80538052",
         10697 => x"7a51ff9f",
         10698 => x"ed3f848b",
         10699 => x"85a4d252",
         10700 => x"7a51ff9f",
         10701 => x"8f3f868a",
         10702 => x"85e4f252",
         10703 => x"83e41b51",
         10704 => x"ff9f813f",
         10705 => x"ff185283",
         10706 => x"e81b51ff",
         10707 => x"9ef63f82",
         10708 => x"5283ec1b",
         10709 => x"51ff9eec",
         10710 => x"3f82d4d5",
         10711 => x"527851ff",
         10712 => x"9ec43f75",
         10713 => x"54608705",
         10714 => x"537a527e",
         10715 => x"51ff9ae5",
         10716 => x"3f755460",
         10717 => x"16537a52",
         10718 => x"7e51ff9a",
         10719 => x"d83f6553",
         10720 => x"80527a51",
         10721 => x"ff9f8f3f",
         10722 => x"7f568058",
         10723 => x"7d832e09",
         10724 => x"81069a38",
         10725 => x"f8527a51",
         10726 => x"ff9ea93f",
         10727 => x"ff52841b",
         10728 => x"51ff9ea0",
         10729 => x"3ff00a52",
         10730 => x"881b5191",
         10731 => x"3987ffff",
         10732 => x"f8557d81",
         10733 => x"2e8338f8",
         10734 => x"5574527a",
         10735 => x"51ff9e84",
         10736 => x"3f7c5561",
         10737 => x"57746226",
         10738 => x"83387457",
         10739 => x"76547553",
         10740 => x"7a527e51",
         10741 => x"ff99fe3f",
         10742 => x"82b5a808",
         10743 => x"82873884",
         10744 => x"805382b5",
         10745 => x"a808527a",
         10746 => x"51ff9eaa",
         10747 => x"3f761675",
         10748 => x"78315656",
         10749 => x"74cd3881",
         10750 => x"18587780",
         10751 => x"2eff8d38",
         10752 => x"79557d83",
         10753 => x"2e833863",
         10754 => x"55615774",
         10755 => x"62268338",
         10756 => x"74577654",
         10757 => x"75537a52",
         10758 => x"7e51ff99",
         10759 => x"b83f82b5",
         10760 => x"a80881c1",
         10761 => x"38761675",
         10762 => x"78315656",
         10763 => x"74db388c",
         10764 => x"567d832e",
         10765 => x"93388656",
         10766 => x"6683ffff",
         10767 => x"268a3884",
         10768 => x"567d822e",
         10769 => x"83388156",
         10770 => x"64810658",
         10771 => x"7780fe38",
         10772 => x"84805377",
         10773 => x"527a51ff",
         10774 => x"9dbc3f82",
         10775 => x"d4d55278",
         10776 => x"51ff9cc2",
         10777 => x"3f83be1b",
         10778 => x"55777534",
         10779 => x"810b8116",
         10780 => x"34810b82",
         10781 => x"16347783",
         10782 => x"16347584",
         10783 => x"16346067",
         10784 => x"055680fd",
         10785 => x"c1527551",
         10786 => x"fec1983f",
         10787 => x"fe0b8516",
         10788 => x"3482b5a8",
         10789 => x"08822abf",
         10790 => x"07567586",
         10791 => x"163482b5",
         10792 => x"a8088716",
         10793 => x"34605283",
         10794 => x"c61b51ff",
         10795 => x"9c963f66",
         10796 => x"5283ca1b",
         10797 => x"51ff9c8c",
         10798 => x"3f815477",
         10799 => x"537a527e",
         10800 => x"51ff9891",
         10801 => x"3f815682",
         10802 => x"b5a808a2",
         10803 => x"38805380",
         10804 => x"527e51ff",
         10805 => x"99e33f81",
         10806 => x"5682b5a8",
         10807 => x"08903889",
         10808 => x"398e568a",
         10809 => x"39815686",
         10810 => x"3982b5a8",
         10811 => x"08567582",
         10812 => x"b5a80c99",
         10813 => x"3d0d04f5",
         10814 => x"3d0d7d60",
         10815 => x"5b598079",
         10816 => x"60ff055a",
         10817 => x"57577678",
         10818 => x"25b4388d",
         10819 => x"3df81155",
         10820 => x"558153fc",
         10821 => x"15527951",
         10822 => x"c9dc3f7a",
         10823 => x"812e0981",
         10824 => x"069c388c",
         10825 => x"3d335574",
         10826 => x"8d2edb38",
         10827 => x"74767081",
         10828 => x"05583481",
         10829 => x"1757748a",
         10830 => x"2e098106",
         10831 => x"c9388076",
         10832 => x"34785576",
         10833 => x"83387655",
         10834 => x"7482b5a8",
         10835 => x"0c8d3d0d",
         10836 => x"04f73d0d",
         10837 => x"7b028405",
         10838 => x"b3053359",
         10839 => x"57778a2e",
         10840 => x"09810687",
         10841 => x"388d5276",
         10842 => x"51e73f84",
         10843 => x"17085680",
         10844 => x"7624be38",
         10845 => x"88170877",
         10846 => x"178c0556",
         10847 => x"59777534",
         10848 => x"811656bb",
         10849 => x"7625a138",
         10850 => x"8b3dfc05",
         10851 => x"5475538c",
         10852 => x"17527608",
         10853 => x"51cbdc3f",
         10854 => x"79763270",
         10855 => x"30707207",
         10856 => x"9f2a7030",
         10857 => x"53515656",
         10858 => x"7584180c",
         10859 => x"81198818",
         10860 => x"0c8b3d0d",
         10861 => x"04f93d0d",
         10862 => x"79841108",
         10863 => x"56568075",
         10864 => x"24a73889",
         10865 => x"3dfc0554",
         10866 => x"74538c16",
         10867 => x"52750851",
         10868 => x"cba13f82",
         10869 => x"b5a80891",
         10870 => x"38841608",
         10871 => x"782e0981",
         10872 => x"06873888",
         10873 => x"16085583",
         10874 => x"39ff5574",
         10875 => x"82b5a80c",
         10876 => x"893d0d04",
         10877 => x"fd3d0d75",
         10878 => x"5480cc53",
         10879 => x"80527351",
         10880 => x"ff9a933f",
         10881 => x"76740c85",
         10882 => x"3d0d04ea",
         10883 => x"3d0d0280",
         10884 => x"e305336a",
         10885 => x"53863d70",
         10886 => x"535454d8",
         10887 => x"3f735272",
         10888 => x"51feae3f",
         10889 => x"7251ff8d",
         10890 => x"3f983d0d",
         10891 => x"04000000",
         10892 => x"00ffffff",
         10893 => x"ff00ffff",
         10894 => x"ffff00ff",
         10895 => x"ffffff00",
         10896 => x"00002ba8",
         10897 => x"00002b2c",
         10898 => x"00002b33",
         10899 => x"00002b3a",
         10900 => x"00002b41",
         10901 => x"00002b48",
         10902 => x"00002b4f",
         10903 => x"00002b56",
         10904 => x"00002b5d",
         10905 => x"00002b64",
         10906 => x"00002b6b",
         10907 => x"00002b72",
         10908 => x"00002b78",
         10909 => x"00002b7e",
         10910 => x"00002b84",
         10911 => x"00002b8a",
         10912 => x"00002b90",
         10913 => x"00002b96",
         10914 => x"00002b9c",
         10915 => x"00002ba2",
         10916 => x"0000413b",
         10917 => x"00004141",
         10918 => x"00004147",
         10919 => x"0000414d",
         10920 => x"00004153",
         10921 => x"00004720",
         10922 => x"00004816",
         10923 => x"0000490e",
         10924 => x"00004b48",
         10925 => x"000047fe",
         10926 => x"000045f5",
         10927 => x"000049c2",
         10928 => x"00004b1e",
         10929 => x"00004a00",
         10930 => x"00004a96",
         10931 => x"00004a1c",
         10932 => x"000048bd",
         10933 => x"000045f5",
         10934 => x"0000490e",
         10935 => x"00004932",
         10936 => x"000049c2",
         10937 => x"000045f5",
         10938 => x"000045f5",
         10939 => x"00004a1c",
         10940 => x"00004a96",
         10941 => x"00004b1e",
         10942 => x"00004b48",
         10943 => x"00000e2f",
         10944 => x"00001718",
         10945 => x"00001718",
         10946 => x"00000e5e",
         10947 => x"00001718",
         10948 => x"00001718",
         10949 => x"00001718",
         10950 => x"00001718",
         10951 => x"00001718",
         10952 => x"00001718",
         10953 => x"00001718",
         10954 => x"00000e1b",
         10955 => x"00001718",
         10956 => x"00000e46",
         10957 => x"00000e76",
         10958 => x"00001718",
         10959 => x"00001718",
         10960 => x"00001718",
         10961 => x"00001718",
         10962 => x"00001718",
         10963 => x"00001718",
         10964 => x"00001718",
         10965 => x"00001718",
         10966 => x"00001718",
         10967 => x"00001718",
         10968 => x"00001718",
         10969 => x"00001718",
         10970 => x"00001718",
         10971 => x"00001718",
         10972 => x"00001718",
         10973 => x"00001718",
         10974 => x"00001718",
         10975 => x"00001718",
         10976 => x"00001718",
         10977 => x"00001718",
         10978 => x"00001718",
         10979 => x"00001718",
         10980 => x"00001718",
         10981 => x"00001718",
         10982 => x"00001718",
         10983 => x"00001718",
         10984 => x"00001718",
         10985 => x"00001718",
         10986 => x"00001718",
         10987 => x"00001718",
         10988 => x"00001718",
         10989 => x"00001718",
         10990 => x"00001718",
         10991 => x"00001718",
         10992 => x"00001718",
         10993 => x"00001718",
         10994 => x"00000fa6",
         10995 => x"00001718",
         10996 => x"00001718",
         10997 => x"00001718",
         10998 => x"00001718",
         10999 => x"00001114",
         11000 => x"00001718",
         11001 => x"00001718",
         11002 => x"00001718",
         11003 => x"00001718",
         11004 => x"00001718",
         11005 => x"00001718",
         11006 => x"00001718",
         11007 => x"00001718",
         11008 => x"00001718",
         11009 => x"00001718",
         11010 => x"00000ed6",
         11011 => x"0000103d",
         11012 => x"00000ead",
         11013 => x"00000ead",
         11014 => x"00000ead",
         11015 => x"00001718",
         11016 => x"0000103d",
         11017 => x"00001718",
         11018 => x"00001718",
         11019 => x"00000e96",
         11020 => x"00001718",
         11021 => x"00001718",
         11022 => x"000010ea",
         11023 => x"000010f5",
         11024 => x"00001718",
         11025 => x"00001718",
         11026 => x"00000f0f",
         11027 => x"00001718",
         11028 => x"0000111d",
         11029 => x"00001718",
         11030 => x"00001718",
         11031 => x"00001114",
         11032 => x"64696e69",
         11033 => x"74000000",
         11034 => x"64696f63",
         11035 => x"746c0000",
         11036 => x"66696e69",
         11037 => x"74000000",
         11038 => x"666c6f61",
         11039 => x"64000000",
         11040 => x"66657865",
         11041 => x"63000000",
         11042 => x"6d636c65",
         11043 => x"61720000",
         11044 => x"6d636f70",
         11045 => x"79000000",
         11046 => x"6d646966",
         11047 => x"66000000",
         11048 => x"6d64756d",
         11049 => x"70000000",
         11050 => x"6d656200",
         11051 => x"6d656800",
         11052 => x"6d657700",
         11053 => x"68696400",
         11054 => x"68696500",
         11055 => x"68666400",
         11056 => x"68666500",
         11057 => x"63616c6c",
         11058 => x"00000000",
         11059 => x"6a6d7000",
         11060 => x"72657374",
         11061 => x"61727400",
         11062 => x"72657365",
         11063 => x"74000000",
         11064 => x"696e666f",
         11065 => x"00000000",
         11066 => x"74657374",
         11067 => x"00000000",
         11068 => x"74626173",
         11069 => x"69630000",
         11070 => x"6d626173",
         11071 => x"69630000",
         11072 => x"6b696c6f",
         11073 => x"00000000",
         11074 => x"65640000",
         11075 => x"4469736b",
         11076 => x"20457272",
         11077 => x"6f720a00",
         11078 => x"496e7465",
         11079 => x"726e616c",
         11080 => x"20657272",
         11081 => x"6f722e0a",
         11082 => x"00000000",
         11083 => x"4469736b",
         11084 => x"206e6f74",
         11085 => x"20726561",
         11086 => x"64792e0a",
         11087 => x"00000000",
         11088 => x"4e6f2066",
         11089 => x"696c6520",
         11090 => x"666f756e",
         11091 => x"642e0a00",
         11092 => x"4e6f2070",
         11093 => x"61746820",
         11094 => x"666f756e",
         11095 => x"642e0a00",
         11096 => x"496e7661",
         11097 => x"6c696420",
         11098 => x"66696c65",
         11099 => x"6e616d65",
         11100 => x"2e0a0000",
         11101 => x"41636365",
         11102 => x"73732064",
         11103 => x"656e6965",
         11104 => x"642e0a00",
         11105 => x"46696c65",
         11106 => x"20616c72",
         11107 => x"65616479",
         11108 => x"20657869",
         11109 => x"7374732e",
         11110 => x"0a000000",
         11111 => x"46696c65",
         11112 => x"2068616e",
         11113 => x"646c6520",
         11114 => x"696e7661",
         11115 => x"6c69642e",
         11116 => x"0a000000",
         11117 => x"53442069",
         11118 => x"73207772",
         11119 => x"69746520",
         11120 => x"70726f74",
         11121 => x"65637465",
         11122 => x"642e0a00",
         11123 => x"44726976",
         11124 => x"65206e75",
         11125 => x"6d626572",
         11126 => x"20697320",
         11127 => x"696e7661",
         11128 => x"6c69642e",
         11129 => x"0a000000",
         11130 => x"4469736b",
         11131 => x"206e6f74",
         11132 => x"20656e61",
         11133 => x"626c6564",
         11134 => x"2e0a0000",
         11135 => x"4e6f2063",
         11136 => x"6f6d7061",
         11137 => x"7469626c",
         11138 => x"65206669",
         11139 => x"6c657379",
         11140 => x"7374656d",
         11141 => x"20666f75",
         11142 => x"6e64206f",
         11143 => x"6e206469",
         11144 => x"736b2e0a",
         11145 => x"00000000",
         11146 => x"466f726d",
         11147 => x"61742061",
         11148 => x"626f7274",
         11149 => x"65642e0a",
         11150 => x"00000000",
         11151 => x"54696d65",
         11152 => x"6f75742c",
         11153 => x"206f7065",
         11154 => x"72617469",
         11155 => x"6f6e2063",
         11156 => x"616e6365",
         11157 => x"6c6c6564",
         11158 => x"2e0a0000",
         11159 => x"46696c65",
         11160 => x"20697320",
         11161 => x"6c6f636b",
         11162 => x"65642e0a",
         11163 => x"00000000",
         11164 => x"496e7375",
         11165 => x"66666963",
         11166 => x"69656e74",
         11167 => x"206d656d",
         11168 => x"6f72792e",
         11169 => x"0a000000",
         11170 => x"546f6f20",
         11171 => x"6d616e79",
         11172 => x"206f7065",
         11173 => x"6e206669",
         11174 => x"6c65732e",
         11175 => x"0a000000",
         11176 => x"50617261",
         11177 => x"6d657465",
         11178 => x"72732069",
         11179 => x"6e636f72",
         11180 => x"72656374",
         11181 => x"2e0a0000",
         11182 => x"53756363",
         11183 => x"6573732e",
         11184 => x"0a000000",
         11185 => x"556e6b6e",
         11186 => x"6f776e20",
         11187 => x"6572726f",
         11188 => x"722e0a00",
         11189 => x"0a256c75",
         11190 => x"20627974",
         11191 => x"65732025",
         11192 => x"73206174",
         11193 => x"20256c75",
         11194 => x"20627974",
         11195 => x"65732f73",
         11196 => x"65632e0a",
         11197 => x"00000000",
         11198 => x"72656164",
         11199 => x"00000000",
         11200 => x"25303858",
         11201 => x"00000000",
         11202 => x"3a202000",
         11203 => x"25303458",
         11204 => x"00000000",
         11205 => x"20202020",
         11206 => x"20202020",
         11207 => x"00000000",
         11208 => x"25303258",
         11209 => x"00000000",
         11210 => x"20200000",
         11211 => x"207c0000",
         11212 => x"7c0d0a00",
         11213 => x"7a4f5300",
         11214 => x"0a2a2a20",
         11215 => x"25732028",
         11216 => x"00000000",
         11217 => x"30322f30",
         11218 => x"352f3230",
         11219 => x"32300000",
         11220 => x"76312e30",
         11221 => x"32000000",
         11222 => x"205a5055",
         11223 => x"2c207265",
         11224 => x"76202530",
         11225 => x"32782920",
         11226 => x"25732025",
         11227 => x"73202a2a",
         11228 => x"0a0a0000",
         11229 => x"5a505520",
         11230 => x"496e7465",
         11231 => x"72727570",
         11232 => x"74204861",
         11233 => x"6e646c65",
         11234 => x"720a0000",
         11235 => x"54696d65",
         11236 => x"7220696e",
         11237 => x"74657272",
         11238 => x"7570740a",
         11239 => x"00000000",
         11240 => x"50533220",
         11241 => x"696e7465",
         11242 => x"72727570",
         11243 => x"740a0000",
         11244 => x"494f4354",
         11245 => x"4c205244",
         11246 => x"20696e74",
         11247 => x"65727275",
         11248 => x"70740a00",
         11249 => x"494f4354",
         11250 => x"4c205752",
         11251 => x"20696e74",
         11252 => x"65727275",
         11253 => x"70740a00",
         11254 => x"55415254",
         11255 => x"30205258",
         11256 => x"20696e74",
         11257 => x"65727275",
         11258 => x"70740a00",
         11259 => x"55415254",
         11260 => x"30205458",
         11261 => x"20696e74",
         11262 => x"65727275",
         11263 => x"70740a00",
         11264 => x"55415254",
         11265 => x"31205258",
         11266 => x"20696e74",
         11267 => x"65727275",
         11268 => x"70740a00",
         11269 => x"55415254",
         11270 => x"31205458",
         11271 => x"20696e74",
         11272 => x"65727275",
         11273 => x"70740a00",
         11274 => x"53657474",
         11275 => x"696e6720",
         11276 => x"75702074",
         11277 => x"696d6572",
         11278 => x"2e2e2e0a",
         11279 => x"00000000",
         11280 => x"456e6162",
         11281 => x"6c696e67",
         11282 => x"2074696d",
         11283 => x"65722e2e",
         11284 => x"2e0a0000",
         11285 => x"6175746f",
         11286 => x"65786563",
         11287 => x"2e626174",
         11288 => x"00000000",
         11289 => x"7a4f532e",
         11290 => x"68737400",
         11291 => x"303a0000",
         11292 => x"4661696c",
         11293 => x"65642074",
         11294 => x"6f20696e",
         11295 => x"69746961",
         11296 => x"6c697365",
         11297 => x"20736420",
         11298 => x"63617264",
         11299 => x"20302c20",
         11300 => x"706c6561",
         11301 => x"73652069",
         11302 => x"6e697420",
         11303 => x"6d616e75",
         11304 => x"616c6c79",
         11305 => x"2e000000",
         11306 => x"2a200000",
         11307 => x"436c6561",
         11308 => x"72696e67",
         11309 => x"2e2e2e2e",
         11310 => x"00000000",
         11311 => x"436f7079",
         11312 => x"696e672e",
         11313 => x"2e2e0000",
         11314 => x"436f6d70",
         11315 => x"6172696e",
         11316 => x"672e2e2e",
         11317 => x"00000000",
         11318 => x"2530386c",
         11319 => x"78282530",
         11320 => x"3878292d",
         11321 => x"3e253038",
         11322 => x"6c782825",
         11323 => x"30387829",
         11324 => x"0a000000",
         11325 => x"44756d70",
         11326 => x"204d656d",
         11327 => x"6f72790a",
         11328 => x"00000000",
         11329 => x"0a436f6d",
         11330 => x"706c6574",
         11331 => x"652e0a00",
         11332 => x"25303858",
         11333 => x"20253032",
         11334 => x"582d0000",
         11335 => x"3f3f3f0a",
         11336 => x"00000000",
         11337 => x"25303858",
         11338 => x"20253034",
         11339 => x"582d0000",
         11340 => x"25303858",
         11341 => x"20253038",
         11342 => x"582d0000",
         11343 => x"45786563",
         11344 => x"7574696e",
         11345 => x"6720636f",
         11346 => x"64652040",
         11347 => x"20253038",
         11348 => x"78202e2e",
         11349 => x"2e0a0000",
         11350 => x"43616c6c",
         11351 => x"696e6720",
         11352 => x"636f6465",
         11353 => x"20402025",
         11354 => x"30387820",
         11355 => x"2e2e2e0a",
         11356 => x"00000000",
         11357 => x"43616c6c",
         11358 => x"20726574",
         11359 => x"75726e65",
         11360 => x"6420636f",
         11361 => x"64652028",
         11362 => x"2564292e",
         11363 => x"0a000000",
         11364 => x"52657374",
         11365 => x"61727469",
         11366 => x"6e672061",
         11367 => x"70706c69",
         11368 => x"63617469",
         11369 => x"6f6e2e2e",
         11370 => x"2e0a0000",
         11371 => x"436f6c64",
         11372 => x"20726562",
         11373 => x"6f6f7469",
         11374 => x"6e672e2e",
         11375 => x"2e0a0000",
         11376 => x"5a505500",
         11377 => x"62696e00",
         11378 => x"25643a5c",
         11379 => x"25735c25",
         11380 => x"732e2573",
         11381 => x"00000000",
         11382 => x"25643a5c",
         11383 => x"25735c25",
         11384 => x"73000000",
         11385 => x"25643a5c",
         11386 => x"25730000",
         11387 => x"42616420",
         11388 => x"636f6d6d",
         11389 => x"616e642e",
         11390 => x"00000000",
         11391 => x"48454c4c",
         11392 => x"4f203120",
         11393 => x"46524f4d",
         11394 => x"20505249",
         11395 => x"4e544600",
         11396 => x"48454c4c",
         11397 => x"4f203220",
         11398 => x"46524f4d",
         11399 => x"20505249",
         11400 => x"4e544600",
         11401 => x"52756e6e",
         11402 => x"696e672e",
         11403 => x"2e2e0a00",
         11404 => x"456e6162",
         11405 => x"6c696e67",
         11406 => x"20696e74",
         11407 => x"65727275",
         11408 => x"7074732e",
         11409 => x"2e2e0a00",
         11410 => x"25642f25",
         11411 => x"642f2564",
         11412 => x"2025643a",
         11413 => x"25643a25",
         11414 => x"642e2564",
         11415 => x"25640a00",
         11416 => x"536f4320",
         11417 => x"436f6e66",
         11418 => x"69677572",
         11419 => x"6174696f",
         11420 => x"6e000000",
         11421 => x"20286672",
         11422 => x"6f6d2053",
         11423 => x"6f432063",
         11424 => x"6f6e6669",
         11425 => x"67290000",
         11426 => x"3a0a4465",
         11427 => x"76696365",
         11428 => x"7320696d",
         11429 => x"706c656d",
         11430 => x"656e7465",
         11431 => x"643a0a00",
         11432 => x"20202020",
         11433 => x"57422053",
         11434 => x"4452414d",
         11435 => x"20202825",
         11436 => x"3038583a",
         11437 => x"25303858",
         11438 => x"292e0a00",
         11439 => x"20202020",
         11440 => x"53445241",
         11441 => x"4d202020",
         11442 => x"20202825",
         11443 => x"3038583a",
         11444 => x"25303858",
         11445 => x"292e0a00",
         11446 => x"20202020",
         11447 => x"494e534e",
         11448 => x"20425241",
         11449 => x"4d202825",
         11450 => x"3038583a",
         11451 => x"25303858",
         11452 => x"292e0a00",
         11453 => x"20202020",
         11454 => x"4252414d",
         11455 => x"20202020",
         11456 => x"20202825",
         11457 => x"3038583a",
         11458 => x"25303858",
         11459 => x"292e0a00",
         11460 => x"20202020",
         11461 => x"52414d20",
         11462 => x"20202020",
         11463 => x"20202825",
         11464 => x"3038583a",
         11465 => x"25303858",
         11466 => x"292e0a00",
         11467 => x"20202020",
         11468 => x"53442043",
         11469 => x"41524420",
         11470 => x"20202844",
         11471 => x"65766963",
         11472 => x"6573203d",
         11473 => x"25303264",
         11474 => x"292e0a00",
         11475 => x"20202020",
         11476 => x"54494d45",
         11477 => x"52312020",
         11478 => x"20202854",
         11479 => x"696d6572",
         11480 => x"7320203d",
         11481 => x"25303264",
         11482 => x"292e0a00",
         11483 => x"20202020",
         11484 => x"494e5452",
         11485 => x"20435452",
         11486 => x"4c202843",
         11487 => x"68616e6e",
         11488 => x"656c733d",
         11489 => x"25303264",
         11490 => x"292e0a00",
         11491 => x"20202020",
         11492 => x"57495348",
         11493 => x"424f4e45",
         11494 => x"20425553",
         11495 => x"0a000000",
         11496 => x"20202020",
         11497 => x"57422049",
         11498 => x"32430a00",
         11499 => x"20202020",
         11500 => x"494f4354",
         11501 => x"4c0a0000",
         11502 => x"20202020",
         11503 => x"5053320a",
         11504 => x"00000000",
         11505 => x"20202020",
         11506 => x"5350490a",
         11507 => x"00000000",
         11508 => x"41646472",
         11509 => x"65737365",
         11510 => x"733a0a00",
         11511 => x"20202020",
         11512 => x"43505520",
         11513 => x"52657365",
         11514 => x"74205665",
         11515 => x"63746f72",
         11516 => x"20416464",
         11517 => x"72657373",
         11518 => x"203d2025",
         11519 => x"3038580a",
         11520 => x"00000000",
         11521 => x"20202020",
         11522 => x"43505520",
         11523 => x"4d656d6f",
         11524 => x"72792053",
         11525 => x"74617274",
         11526 => x"20416464",
         11527 => x"72657373",
         11528 => x"203d2025",
         11529 => x"3038580a",
         11530 => x"00000000",
         11531 => x"20202020",
         11532 => x"53746163",
         11533 => x"6b205374",
         11534 => x"61727420",
         11535 => x"41646472",
         11536 => x"65737320",
         11537 => x"20202020",
         11538 => x"203d2025",
         11539 => x"3038580a",
         11540 => x"00000000",
         11541 => x"4d697363",
         11542 => x"3a0a0000",
         11543 => x"20202020",
         11544 => x"5a505520",
         11545 => x"49642020",
         11546 => x"20202020",
         11547 => x"20202020",
         11548 => x"20202020",
         11549 => x"20202020",
         11550 => x"203d2025",
         11551 => x"3034580a",
         11552 => x"00000000",
         11553 => x"20202020",
         11554 => x"53797374",
         11555 => x"656d2043",
         11556 => x"6c6f636b",
         11557 => x"20467265",
         11558 => x"71202020",
         11559 => x"20202020",
         11560 => x"203d2025",
         11561 => x"642e2530",
         11562 => x"34644d48",
         11563 => x"7a0a0000",
         11564 => x"20202020",
         11565 => x"53445241",
         11566 => x"4d20436c",
         11567 => x"6f636b20",
         11568 => x"46726571",
         11569 => x"20202020",
         11570 => x"20202020",
         11571 => x"203d2025",
         11572 => x"642e2530",
         11573 => x"34644d48",
         11574 => x"7a0a0000",
         11575 => x"20202020",
         11576 => x"57697368",
         11577 => x"626f6e65",
         11578 => x"20534452",
         11579 => x"414d2043",
         11580 => x"6c6f636b",
         11581 => x"20467265",
         11582 => x"713d2025",
         11583 => x"642e2530",
         11584 => x"34644d48",
         11585 => x"7a0a0000",
         11586 => x"536d616c",
         11587 => x"6c000000",
         11588 => x"4d656469",
         11589 => x"756d0000",
         11590 => x"466c6578",
         11591 => x"00000000",
         11592 => x"45564f00",
         11593 => x"45564f6d",
         11594 => x"696e0000",
         11595 => x"556e6b6e",
         11596 => x"6f776e00",
         11597 => x"00009690",
         11598 => x"01000000",
         11599 => x"00000002",
         11600 => x"0000968c",
         11601 => x"01000000",
         11602 => x"00000003",
         11603 => x"00009688",
         11604 => x"01000000",
         11605 => x"00000004",
         11606 => x"00009684",
         11607 => x"01000000",
         11608 => x"00000005",
         11609 => x"00009680",
         11610 => x"01000000",
         11611 => x"00000006",
         11612 => x"0000967c",
         11613 => x"01000000",
         11614 => x"00000007",
         11615 => x"00009678",
         11616 => x"01000000",
         11617 => x"00000001",
         11618 => x"00009674",
         11619 => x"01000000",
         11620 => x"00000008",
         11621 => x"00009670",
         11622 => x"01000000",
         11623 => x"0000000b",
         11624 => x"0000966c",
         11625 => x"01000000",
         11626 => x"00000009",
         11627 => x"00009668",
         11628 => x"01000000",
         11629 => x"0000000a",
         11630 => x"00009664",
         11631 => x"04000000",
         11632 => x"0000000d",
         11633 => x"00009660",
         11634 => x"04000000",
         11635 => x"0000000c",
         11636 => x"0000965c",
         11637 => x"04000000",
         11638 => x"0000000e",
         11639 => x"00009658",
         11640 => x"03000000",
         11641 => x"0000000f",
         11642 => x"00009654",
         11643 => x"04000000",
         11644 => x"0000000f",
         11645 => x"00009650",
         11646 => x"04000000",
         11647 => x"00000010",
         11648 => x"0000964c",
         11649 => x"04000000",
         11650 => x"00000011",
         11651 => x"00009648",
         11652 => x"03000000",
         11653 => x"00000012",
         11654 => x"00009644",
         11655 => x"03000000",
         11656 => x"00000013",
         11657 => x"00009640",
         11658 => x"03000000",
         11659 => x"00000014",
         11660 => x"0000963c",
         11661 => x"03000000",
         11662 => x"00000015",
         11663 => x"1b5b4400",
         11664 => x"1b5b4300",
         11665 => x"1b5b4200",
         11666 => x"1b5b4100",
         11667 => x"1b5b367e",
         11668 => x"1b5b357e",
         11669 => x"1b5b347e",
         11670 => x"1b304600",
         11671 => x"1b5b337e",
         11672 => x"1b5b327e",
         11673 => x"1b5b317e",
         11674 => x"10000000",
         11675 => x"0e000000",
         11676 => x"0d000000",
         11677 => x"0b000000",
         11678 => x"08000000",
         11679 => x"06000000",
         11680 => x"05000000",
         11681 => x"04000000",
         11682 => x"03000000",
         11683 => x"02000000",
         11684 => x"01000000",
         11685 => x"68697374",
         11686 => x"6f727900",
         11687 => x"68697374",
         11688 => x"00000000",
         11689 => x"21000000",
         11690 => x"25303464",
         11691 => x"20202573",
         11692 => x"0a000000",
         11693 => x"4661696c",
         11694 => x"65642074",
         11695 => x"6f207265",
         11696 => x"73657420",
         11697 => x"74686520",
         11698 => x"68697374",
         11699 => x"6f727920",
         11700 => x"66696c65",
         11701 => x"20746f20",
         11702 => x"454f462e",
         11703 => x"0a000000",
         11704 => x"43616e6e",
         11705 => x"6f74206f",
         11706 => x"70656e2f",
         11707 => x"63726561",
         11708 => x"74652068",
         11709 => x"6973746f",
         11710 => x"72792066",
         11711 => x"696c652c",
         11712 => x"20646973",
         11713 => x"61626c69",
         11714 => x"6e672e00",
         11715 => x"53440000",
         11716 => x"222a2b2c",
         11717 => x"3a3b3c3d",
         11718 => x"3e3f5b5d",
         11719 => x"7c7f0000",
         11720 => x"46415400",
         11721 => x"46415433",
         11722 => x"32000000",
         11723 => x"ebfe904d",
         11724 => x"53444f53",
         11725 => x"352e3000",
         11726 => x"4e4f204e",
         11727 => x"414d4520",
         11728 => x"20202046",
         11729 => x"41543332",
         11730 => x"20202000",
         11731 => x"4e4f204e",
         11732 => x"414d4520",
         11733 => x"20202046",
         11734 => x"41542020",
         11735 => x"20202000",
         11736 => x"0000970c",
         11737 => x"00000000",
         11738 => x"00000000",
         11739 => x"00000000",
         11740 => x"809a4541",
         11741 => x"8e418f80",
         11742 => x"45454549",
         11743 => x"49498e8f",
         11744 => x"9092924f",
         11745 => x"994f5555",
         11746 => x"59999a9b",
         11747 => x"9c9d9e9f",
         11748 => x"41494f55",
         11749 => x"a5a5a6a7",
         11750 => x"a8a9aaab",
         11751 => x"acadaeaf",
         11752 => x"b0b1b2b3",
         11753 => x"b4b5b6b7",
         11754 => x"b8b9babb",
         11755 => x"bcbdbebf",
         11756 => x"c0c1c2c3",
         11757 => x"c4c5c6c7",
         11758 => x"c8c9cacb",
         11759 => x"cccdcecf",
         11760 => x"d0d1d2d3",
         11761 => x"d4d5d6d7",
         11762 => x"d8d9dadb",
         11763 => x"dcdddedf",
         11764 => x"e0e1e2e3",
         11765 => x"e4e5e6e7",
         11766 => x"e8e9eaeb",
         11767 => x"ecedeeef",
         11768 => x"f0f1f2f3",
         11769 => x"f4f5f6f7",
         11770 => x"f8f9fafb",
         11771 => x"fcfdfeff",
         11772 => x"2b2e2c3b",
         11773 => x"3d5b5d2f",
         11774 => x"5c222a3a",
         11775 => x"3c3e3f7c",
         11776 => x"7f000000",
         11777 => x"00010004",
         11778 => x"00100040",
         11779 => x"01000200",
         11780 => x"00000000",
         11781 => x"00010002",
         11782 => x"00040008",
         11783 => x"00100020",
         11784 => x"00000000",
         11785 => x"00000000",
         11786 => x"00008c60",
         11787 => x"01020100",
         11788 => x"00000000",
         11789 => x"00000000",
         11790 => x"00008c68",
         11791 => x"01040100",
         11792 => x"00000000",
         11793 => x"00000000",
         11794 => x"00008c70",
         11795 => x"01140300",
         11796 => x"00000000",
         11797 => x"00000000",
         11798 => x"00008c78",
         11799 => x"012b0300",
         11800 => x"00000000",
         11801 => x"00000000",
         11802 => x"00008c80",
         11803 => x"01300300",
         11804 => x"00000000",
         11805 => x"00000000",
         11806 => x"00008c88",
         11807 => x"013c0400",
         11808 => x"00000000",
         11809 => x"00000000",
         11810 => x"00008c90",
         11811 => x"013d0400",
         11812 => x"00000000",
         11813 => x"00000000",
         11814 => x"00008c98",
         11815 => x"013f0400",
         11816 => x"00000000",
         11817 => x"00000000",
         11818 => x"00008ca0",
         11819 => x"01400400",
         11820 => x"00000000",
         11821 => x"00000000",
         11822 => x"00008ca8",
         11823 => x"01410400",
         11824 => x"00000000",
         11825 => x"00000000",
         11826 => x"00008cac",
         11827 => x"01420400",
         11828 => x"00000000",
         11829 => x"00000000",
         11830 => x"00008cb0",
         11831 => x"01430400",
         11832 => x"00000000",
         11833 => x"00000000",
         11834 => x"00008cb4",
         11835 => x"01500500",
         11836 => x"00000000",
         11837 => x"00000000",
         11838 => x"00008cb8",
         11839 => x"01510500",
         11840 => x"00000000",
         11841 => x"00000000",
         11842 => x"00008cbc",
         11843 => x"01540500",
         11844 => x"00000000",
         11845 => x"00000000",
         11846 => x"00008cc0",
         11847 => x"01550500",
         11848 => x"00000000",
         11849 => x"00000000",
         11850 => x"00008cc4",
         11851 => x"01790700",
         11852 => x"00000000",
         11853 => x"00000000",
         11854 => x"00008ccc",
         11855 => x"01780700",
         11856 => x"00000000",
         11857 => x"00000000",
         11858 => x"00008cd0",
         11859 => x"01820800",
         11860 => x"00000000",
         11861 => x"00000000",
         11862 => x"00008cd8",
         11863 => x"01830800",
         11864 => x"00000000",
         11865 => x"00000000",
         11866 => x"00008ce0",
         11867 => x"01850800",
         11868 => x"00000000",
         11869 => x"00000000",
         11870 => x"00008ce8",
         11871 => x"01870800",
         11872 => x"00000000",
         11873 => x"00000000",
         11874 => x"00008cf0",
         11875 => x"018c0900",
         11876 => x"00000000",
         11877 => x"00000000",
         11878 => x"00008cf8",
         11879 => x"018d0900",
         11880 => x"00000000",
         11881 => x"00000000",
         11882 => x"00008d00",
         11883 => x"018e0900",
         11884 => x"00000000",
         11885 => x"00000000",
         11886 => x"00008d08",
         11887 => x"018f0900",
         11888 => x"00000000",
         11889 => x"00000000",
         11890 => x"00000000",
         11891 => x"00000000",
         11892 => x"00007fff",
         11893 => x"00000000",
         11894 => x"00007fff",
         11895 => x"00010000",
         11896 => x"00007fff",
         11897 => x"00010000",
         11898 => x"00810000",
         11899 => x"01000000",
         11900 => x"017fffff",
         11901 => x"00000000",
         11902 => x"00000000",
         11903 => x"00007800",
         11904 => x"00000000",
         11905 => x"05f5e100",
         11906 => x"05f5e100",
         11907 => x"05f5e100",
         11908 => x"00000000",
         11909 => x"01010101",
         11910 => x"01010101",
         11911 => x"01011001",
         11912 => x"01000000",
         11913 => x"00000000",
         11914 => x"00000000",
         11915 => x"00000000",
         11916 => x"00000000",
         11917 => x"00000000",
         11918 => x"00000000",
         11919 => x"00000000",
         11920 => x"00000000",
         11921 => x"00000000",
         11922 => x"00000000",
         11923 => x"00000000",
         11924 => x"00000000",
         11925 => x"00000000",
         11926 => x"00000000",
         11927 => x"00000000",
         11928 => x"00000000",
         11929 => x"00000000",
         11930 => x"00000000",
         11931 => x"00000000",
         11932 => x"00000000",
         11933 => x"00000000",
         11934 => x"00000000",
         11935 => x"00000000",
         11936 => x"00000000",
         11937 => x"00009694",
         11938 => x"01000000",
         11939 => x"0000969c",
         11940 => x"01000000",
         11941 => x"000096a4",
         11942 => x"02000000",
         11943 => x"00000000",
         11944 => x"00000000",
         11945 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

