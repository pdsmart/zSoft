-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b0b93",
          2049 => x"99040000",
          2050 => x"00000000",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b92",
          2121 => x"fd040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b92e0",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b81e8",
          2210 => x"b4738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"92e50400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b80eb",
          2219 => x"b62d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b80ed",
          2227 => x"f22d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"94040b0b",
          2317 => x"0b8ca404",
          2318 => x"0b0b0b8c",
          2319 => x"b4040b0b",
          2320 => x"0b8cc404",
          2321 => x"0b0b0b8c",
          2322 => x"d4040b0b",
          2323 => x"0b8ce404",
          2324 => x"0b0b0b8c",
          2325 => x"f4040b0b",
          2326 => x"0b8d8404",
          2327 => x"0b0b0b8d",
          2328 => x"94040b0b",
          2329 => x"0b8da404",
          2330 => x"0b0b0b8d",
          2331 => x"b4040b0b",
          2332 => x"0b8dc404",
          2333 => x"0b0b0b8d",
          2334 => x"d4040b0b",
          2335 => x"0b8de404",
          2336 => x"0b0b0b8d",
          2337 => x"f4040b0b",
          2338 => x"0b8e8304",
          2339 => x"0b0b0b8e",
          2340 => x"92040b0b",
          2341 => x"0b8ea104",
          2342 => x"0b0b0b8e",
          2343 => x"b1040b0b",
          2344 => x"0b8ec104",
          2345 => x"0b0b0b8e",
          2346 => x"d1040b0b",
          2347 => x"0b8ee104",
          2348 => x"0b0b0b8e",
          2349 => x"f1040b0b",
          2350 => x"0b8f8104",
          2351 => x"0b0b0b8f",
          2352 => x"91040b0b",
          2353 => x"0b8fa104",
          2354 => x"0b0b0b8f",
          2355 => x"b1040b0b",
          2356 => x"0b8fc104",
          2357 => x"0b0b0b8f",
          2358 => x"d1040b0b",
          2359 => x"0b8fe104",
          2360 => x"0b0b0b8f",
          2361 => x"f1040b0b",
          2362 => x"0b908104",
          2363 => x"0b0b0b90",
          2364 => x"91040b0b",
          2365 => x"0b90a104",
          2366 => x"0b0b0b90",
          2367 => x"b1040b0b",
          2368 => x"0b90c104",
          2369 => x"0b0b0b90",
          2370 => x"d1040b0b",
          2371 => x"0b90e104",
          2372 => x"0b0b0b90",
          2373 => x"f1040b0b",
          2374 => x"0b918104",
          2375 => x"0b0b0b91",
          2376 => x"91040b0b",
          2377 => x"0b91a104",
          2378 => x"0b0b0b91",
          2379 => x"b1040b0b",
          2380 => x"0b91c104",
          2381 => x"0b0b0b91",
          2382 => x"d1040b0b",
          2383 => x"0b91e104",
          2384 => x"0b0b0b91",
          2385 => x"f1040b0b",
          2386 => x"0b928104",
          2387 => x"0b0b0b92",
          2388 => x"90040b0b",
          2389 => x"0b929f04",
          2390 => x"0b0b0b92",
          2391 => x"ae04ffff",
          2392 => x"ffffffff",
          2393 => x"ffffffff",
          2394 => x"ffffffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"048287d8",
          2434 => x"0cbe972d",
          2435 => x"8287d808",
          2436 => x"82a09004",
          2437 => x"8287d80c",
          2438 => x"80cbc32d",
          2439 => x"8287d808",
          2440 => x"82a09004",
          2441 => x"8287d80c",
          2442 => x"80cc822d",
          2443 => x"8287d808",
          2444 => x"82a09004",
          2445 => x"8287d80c",
          2446 => x"80cca02d",
          2447 => x"8287d808",
          2448 => x"82a09004",
          2449 => x"8287d80c",
          2450 => x"80d2de2d",
          2451 => x"8287d808",
          2452 => x"82a09004",
          2453 => x"8287d80c",
          2454 => x"80d3dc2d",
          2455 => x"8287d808",
          2456 => x"82a09004",
          2457 => x"8287d80c",
          2458 => x"80ccc32d",
          2459 => x"8287d808",
          2460 => x"82a09004",
          2461 => x"8287d80c",
          2462 => x"80d3f92d",
          2463 => x"8287d808",
          2464 => x"82a09004",
          2465 => x"8287d80c",
          2466 => x"80d5eb2d",
          2467 => x"8287d808",
          2468 => x"82a09004",
          2469 => x"8287d80c",
          2470 => x"80d2842d",
          2471 => x"8287d808",
          2472 => x"82a09004",
          2473 => x"8287d80c",
          2474 => x"80ccf52d",
          2475 => x"8287d808",
          2476 => x"82a09004",
          2477 => x"8287d80c",
          2478 => x"80d29a2d",
          2479 => x"8287d808",
          2480 => x"82a09004",
          2481 => x"8287d80c",
          2482 => x"80d2be2d",
          2483 => x"8287d808",
          2484 => x"82a09004",
          2485 => x"8287d80c",
          2486 => x"80c0a02d",
          2487 => x"8287d808",
          2488 => x"82a09004",
          2489 => x"8287d80c",
          2490 => x"80c0ef2d",
          2491 => x"8287d808",
          2492 => x"82a09004",
          2493 => x"8287d80c",
          2494 => x"b8d32d82",
          2495 => x"87d80882",
          2496 => x"a0900482",
          2497 => x"87d80cba",
          2498 => x"ca2d8287",
          2499 => x"d80882a0",
          2500 => x"90048287",
          2501 => x"d80cbbfd",
          2502 => x"2d8287d8",
          2503 => x"0882a090",
          2504 => x"048287d8",
          2505 => x"0c81ab97",
          2506 => x"2d8287d8",
          2507 => x"0882a090",
          2508 => x"048287d8",
          2509 => x"0c81b888",
          2510 => x"2d8287d8",
          2511 => x"0882a090",
          2512 => x"048287d8",
          2513 => x"0c81affc",
          2514 => x"2d8287d8",
          2515 => x"0882a090",
          2516 => x"048287d8",
          2517 => x"0c81b2f9",
          2518 => x"2d8287d8",
          2519 => x"0882a090",
          2520 => x"048287d8",
          2521 => x"0c81bd97",
          2522 => x"2d8287d8",
          2523 => x"0882a090",
          2524 => x"048287d8",
          2525 => x"0c81c5f7",
          2526 => x"2d8287d8",
          2527 => x"0882a090",
          2528 => x"048287d8",
          2529 => x"0c81b6ea",
          2530 => x"2d8287d8",
          2531 => x"0882a090",
          2532 => x"048287d8",
          2533 => x"0c81c0b6",
          2534 => x"2d8287d8",
          2535 => x"0882a090",
          2536 => x"048287d8",
          2537 => x"0c81c1d5",
          2538 => x"2d8287d8",
          2539 => x"0882a090",
          2540 => x"048287d8",
          2541 => x"0c81c1f4",
          2542 => x"2d8287d8",
          2543 => x"0882a090",
          2544 => x"048287d8",
          2545 => x"0c81c9de",
          2546 => x"2d8287d8",
          2547 => x"0882a090",
          2548 => x"048287d8",
          2549 => x"0c81c7c4",
          2550 => x"2d8287d8",
          2551 => x"0882a090",
          2552 => x"048287d8",
          2553 => x"0c81ccb2",
          2554 => x"2d8287d8",
          2555 => x"0882a090",
          2556 => x"048287d8",
          2557 => x"0c81c2f8",
          2558 => x"2d8287d8",
          2559 => x"0882a090",
          2560 => x"048287d8",
          2561 => x"0c81cfb2",
          2562 => x"2d8287d8",
          2563 => x"0882a090",
          2564 => x"048287d8",
          2565 => x"0c81d0b3",
          2566 => x"2d8287d8",
          2567 => x"0882a090",
          2568 => x"048287d8",
          2569 => x"0c81b8e8",
          2570 => x"2d8287d8",
          2571 => x"0882a090",
          2572 => x"048287d8",
          2573 => x"0c81b8c1",
          2574 => x"2d8287d8",
          2575 => x"0882a090",
          2576 => x"048287d8",
          2577 => x"0c81b9ec",
          2578 => x"2d8287d8",
          2579 => x"0882a090",
          2580 => x"048287d8",
          2581 => x"0c81c3cf",
          2582 => x"2d8287d8",
          2583 => x"0882a090",
          2584 => x"048287d8",
          2585 => x"0c81d1a4",
          2586 => x"2d8287d8",
          2587 => x"0882a090",
          2588 => x"048287d8",
          2589 => x"0c81d3ae",
          2590 => x"2d8287d8",
          2591 => x"0882a090",
          2592 => x"048287d8",
          2593 => x"0c81d6f0",
          2594 => x"2d8287d8",
          2595 => x"0882a090",
          2596 => x"048287d8",
          2597 => x"0c81aab6",
          2598 => x"2d8287d8",
          2599 => x"0882a090",
          2600 => x"048287d8",
          2601 => x"0c81d9dc",
          2602 => x"2d8287d8",
          2603 => x"0882a090",
          2604 => x"048287d8",
          2605 => x"0c81e891",
          2606 => x"2d8287d8",
          2607 => x"0882a090",
          2608 => x"048287d8",
          2609 => x"0c81e5fd",
          2610 => x"2d8287d8",
          2611 => x"0882a090",
          2612 => x"048287d8",
          2613 => x"0c80fbf2",
          2614 => x"2d8287d8",
          2615 => x"0882a090",
          2616 => x"048287d8",
          2617 => x"0c80fddc",
          2618 => x"2d8287d8",
          2619 => x"0882a090",
          2620 => x"048287d8",
          2621 => x"0c80ffc0",
          2622 => x"2d8287d8",
          2623 => x"0882a090",
          2624 => x"048287d8",
          2625 => x"0cb8fc2d",
          2626 => x"8287d808",
          2627 => x"82a09004",
          2628 => x"8287d80c",
          2629 => x"baa02d82",
          2630 => x"87d80882",
          2631 => x"a0900482",
          2632 => x"87d80cbd",
          2633 => x"8d2d8287",
          2634 => x"d80882a0",
          2635 => x"90048287",
          2636 => x"d80c9af4",
          2637 => x"2d8287d8",
          2638 => x"0882a090",
          2639 => x"043c0400",
          2640 => x"00101010",
          2641 => x"10101010",
          2642 => x"10101010",
          2643 => x"10101010",
          2644 => x"10101010",
          2645 => x"10101010",
          2646 => x"10101010",
          2647 => x"10101010",
          2648 => x"53510400",
          2649 => x"007381ff",
          2650 => x"06738306",
          2651 => x"09810583",
          2652 => x"05101010",
          2653 => x"2b0772fc",
          2654 => x"060c5151",
          2655 => x"04727280",
          2656 => x"728106ff",
          2657 => x"05097206",
          2658 => x"05711052",
          2659 => x"720a100a",
          2660 => x"5372ed38",
          2661 => x"51515351",
          2662 => x"048287cc",
          2663 => x"70829f88",
          2664 => x"278e3880",
          2665 => x"71708405",
          2666 => x"530c0b0b",
          2667 => x"0b939c04",
          2668 => x"8c8151b7",
          2669 => x"ad040082",
          2670 => x"87d80802",
          2671 => x"8287d80c",
          2672 => x"fe3d0d82",
          2673 => x"87d80888",
          2674 => x"05088287",
          2675 => x"d808fc05",
          2676 => x"0c8287d8",
          2677 => x"08fc0508",
          2678 => x"52713382",
          2679 => x"87d808fc",
          2680 => x"05088105",
          2681 => x"8287d808",
          2682 => x"fc050c70",
          2683 => x"81ff0651",
          2684 => x"5170802e",
          2685 => x"8338da39",
          2686 => x"8287d808",
          2687 => x"fc0508ff",
          2688 => x"058287d8",
          2689 => x"08fc050c",
          2690 => x"8287d808",
          2691 => x"fc050882",
          2692 => x"87d80888",
          2693 => x"05083170",
          2694 => x"8287cc0c",
          2695 => x"51843d0d",
          2696 => x"8287d80c",
          2697 => x"048287d8",
          2698 => x"08028287",
          2699 => x"d80cfe3d",
          2700 => x"0d8287d8",
          2701 => x"08880508",
          2702 => x"8287d808",
          2703 => x"fc050c82",
          2704 => x"87d8088c",
          2705 => x"05085271",
          2706 => x"338287d8",
          2707 => x"088c0508",
          2708 => x"81058287",
          2709 => x"d8088c05",
          2710 => x"0c8287d8",
          2711 => x"08fc0508",
          2712 => x"53517072",
          2713 => x"348287d8",
          2714 => x"08fc0508",
          2715 => x"81058287",
          2716 => x"d808fc05",
          2717 => x"0c7081ff",
          2718 => x"06517080",
          2719 => x"2e8438ff",
          2720 => x"be398287",
          2721 => x"d8088805",
          2722 => x"08708287",
          2723 => x"cc0c5184",
          2724 => x"3d0d8287",
          2725 => x"d80c0482",
          2726 => x"87d80802",
          2727 => x"8287d80c",
          2728 => x"fd3d0d82",
          2729 => x"87d80888",
          2730 => x"05088287",
          2731 => x"d808fc05",
          2732 => x"0c8287d8",
          2733 => x"088c0508",
          2734 => x"8287d808",
          2735 => x"f8050c82",
          2736 => x"87d80890",
          2737 => x"0508802e",
          2738 => x"80e53882",
          2739 => x"87d80890",
          2740 => x"05088105",
          2741 => x"8287d808",
          2742 => x"90050c82",
          2743 => x"87d80890",
          2744 => x"0508ff05",
          2745 => x"8287d808",
          2746 => x"90050c82",
          2747 => x"87d80890",
          2748 => x"0508802e",
          2749 => x"ba388287",
          2750 => x"d808f805",
          2751 => x"08517033",
          2752 => x"8287d808",
          2753 => x"f8050881",
          2754 => x"058287d8",
          2755 => x"08f8050c",
          2756 => x"8287d808",
          2757 => x"fc050852",
          2758 => x"52717134",
          2759 => x"8287d808",
          2760 => x"fc050881",
          2761 => x"058287d8",
          2762 => x"08fc050c",
          2763 => x"ffad3982",
          2764 => x"87d80888",
          2765 => x"05087082",
          2766 => x"87cc0c51",
          2767 => x"853d0d82",
          2768 => x"87d80c04",
          2769 => x"8287d808",
          2770 => x"028287d8",
          2771 => x"0cfd3d0d",
          2772 => x"8287d808",
          2773 => x"90050880",
          2774 => x"2e81f438",
          2775 => x"8287d808",
          2776 => x"8c050852",
          2777 => x"71338287",
          2778 => x"d8088c05",
          2779 => x"08810582",
          2780 => x"87d8088c",
          2781 => x"050c8287",
          2782 => x"d8088805",
          2783 => x"08703372",
          2784 => x"81ff0653",
          2785 => x"54545171",
          2786 => x"712e8438",
          2787 => x"80ce3982",
          2788 => x"87d80888",
          2789 => x"05085271",
          2790 => x"338287d8",
          2791 => x"08880508",
          2792 => x"81058287",
          2793 => x"d8088805",
          2794 => x"0c7081ff",
          2795 => x"06515170",
          2796 => x"8d38800b",
          2797 => x"8287d808",
          2798 => x"fc050c81",
          2799 => x"9b398287",
          2800 => x"d8089005",
          2801 => x"08ff0582",
          2802 => x"87d80890",
          2803 => x"050c8287",
          2804 => x"d8089005",
          2805 => x"08802e84",
          2806 => x"38ff8139",
          2807 => x"8287d808",
          2808 => x"90050880",
          2809 => x"2e80e838",
          2810 => x"8287d808",
          2811 => x"88050870",
          2812 => x"33525370",
          2813 => x"8d38ff0b",
          2814 => x"8287d808",
          2815 => x"fc050c80",
          2816 => x"d7398287",
          2817 => x"d8088c05",
          2818 => x"08ff0582",
          2819 => x"87d8088c",
          2820 => x"050c8287",
          2821 => x"d8088c05",
          2822 => x"08703352",
          2823 => x"52708c38",
          2824 => x"810b8287",
          2825 => x"d808fc05",
          2826 => x"0cae3982",
          2827 => x"87d80888",
          2828 => x"05087033",
          2829 => x"8287d808",
          2830 => x"8c050870",
          2831 => x"33727131",
          2832 => x"708287d8",
          2833 => x"08fc050c",
          2834 => x"53555252",
          2835 => x"538a3980",
          2836 => x"0b8287d8",
          2837 => x"08fc050c",
          2838 => x"8287d808",
          2839 => x"fc050882",
          2840 => x"87cc0c85",
          2841 => x"3d0d8287",
          2842 => x"d80c0482",
          2843 => x"87d80802",
          2844 => x"8287d80c",
          2845 => x"fe3d0d82",
          2846 => x"87d80888",
          2847 => x"05088287",
          2848 => x"d808fc05",
          2849 => x"0c8287d8",
          2850 => x"08900508",
          2851 => x"802e80d4",
          2852 => x"388287d8",
          2853 => x"08900508",
          2854 => x"81058287",
          2855 => x"d8089005",
          2856 => x"0c8287d8",
          2857 => x"08900508",
          2858 => x"ff058287",
          2859 => x"d8089005",
          2860 => x"0c8287d8",
          2861 => x"08900508",
          2862 => x"802ea938",
          2863 => x"8287d808",
          2864 => x"8c050851",
          2865 => x"708287d8",
          2866 => x"08fc0508",
          2867 => x"52527171",
          2868 => x"348287d8",
          2869 => x"08fc0508",
          2870 => x"81058287",
          2871 => x"d808fc05",
          2872 => x"0cffbe39",
          2873 => x"8287d808",
          2874 => x"88050870",
          2875 => x"8287cc0c",
          2876 => x"51843d0d",
          2877 => x"8287d80c",
          2878 => x"04f93d0d",
          2879 => x"79700870",
          2880 => x"56565874",
          2881 => x"802e80e3",
          2882 => x"38953975",
          2883 => x"0851f9a7",
          2884 => x"3f8287cc",
          2885 => x"0815780c",
          2886 => x"85163354",
          2887 => x"80cd3974",
          2888 => x"335473a0",
          2889 => x"2e098106",
          2890 => x"86388115",
          2891 => x"55f13980",
          2892 => x"57769029",
          2893 => x"8282cc05",
          2894 => x"70085256",
          2895 => x"f8f93f82",
          2896 => x"87cc0853",
          2897 => x"74527508",
          2898 => x"51fbf93f",
          2899 => x"8287cc08",
          2900 => x"8b388416",
          2901 => x"33547381",
          2902 => x"2effb038",
          2903 => x"81177081",
          2904 => x"ff065854",
          2905 => x"997727c9",
          2906 => x"38ff5473",
          2907 => x"8287cc0c",
          2908 => x"893d0d04",
          2909 => x"ff3d0d73",
          2910 => x"52719326",
          2911 => x"818e3871",
          2912 => x"842981e8",
          2913 => x"c4055271",
          2914 => x"080481eb",
          2915 => x"ac518180",
          2916 => x"3981ebb8",
          2917 => x"5180f939",
          2918 => x"81ebcc51",
          2919 => x"80f23981",
          2920 => x"ebe05180",
          2921 => x"eb3981eb",
          2922 => x"f05180e4",
          2923 => x"3981ec80",
          2924 => x"5180dd39",
          2925 => x"81ec9451",
          2926 => x"80d63981",
          2927 => x"eca45180",
          2928 => x"cf3981ec",
          2929 => x"bc5180c8",
          2930 => x"3981ecd4",
          2931 => x"5180c139",
          2932 => x"81ecec51",
          2933 => x"bb3981ed",
          2934 => x"8851b539",
          2935 => x"81ed9c51",
          2936 => x"af3981ed",
          2937 => x"c851a939",
          2938 => x"81eddc51",
          2939 => x"a33981ed",
          2940 => x"fc519d39",
          2941 => x"81ee9051",
          2942 => x"973981ee",
          2943 => x"a8519139",
          2944 => x"81eec051",
          2945 => x"8b3981ee",
          2946 => x"d8518539",
          2947 => x"81eee451",
          2948 => x"b08e3f83",
          2949 => x"3d0d04fb",
          2950 => x"3d0d7779",
          2951 => x"56567487",
          2952 => x"e7268a38",
          2953 => x"74527587",
          2954 => x"e8295191",
          2955 => x"3987e852",
          2956 => x"745180cf",
          2957 => x"b63f8287",
          2958 => x"cc085275",
          2959 => x"5180cfab",
          2960 => x"3f8287cc",
          2961 => x"08547953",
          2962 => x"755281ee",
          2963 => x"f451b5b4",
          2964 => x"3f873d0d",
          2965 => x"04ec3d0d",
          2966 => x"66028405",
          2967 => x"80e30533",
          2968 => x"5b578068",
          2969 => x"7830707a",
          2970 => x"07732551",
          2971 => x"57595978",
          2972 => x"567787ff",
          2973 => x"26833881",
          2974 => x"56747607",
          2975 => x"7081ff06",
          2976 => x"51559356",
          2977 => x"74818238",
          2978 => x"81537652",
          2979 => x"8c3d7052",
          2980 => x"56818e83",
          2981 => x"3f8287cc",
          2982 => x"08578287",
          2983 => x"cc08b938",
          2984 => x"8287cc08",
          2985 => x"87c09888",
          2986 => x"0c8287cc",
          2987 => x"0859963d",
          2988 => x"d4055484",
          2989 => x"80537752",
          2990 => x"75518192",
          2991 => x"bf3f8287",
          2992 => x"cc085782",
          2993 => x"87cc0890",
          2994 => x"387a5574",
          2995 => x"802e8938",
          2996 => x"74197519",
          2997 => x"5959d739",
          2998 => x"963dd805",
          2999 => x"51819aa8",
          3000 => x"3f763070",
          3001 => x"78078025",
          3002 => x"7b30709f",
          3003 => x"2a720651",
          3004 => x"57515674",
          3005 => x"802e9038",
          3006 => x"81ef9853",
          3007 => x"87c09888",
          3008 => x"08527851",
          3009 => x"fe913f76",
          3010 => x"56758287",
          3011 => x"cc0c963d",
          3012 => x"0d04f93d",
          3013 => x"0d7b0284",
          3014 => x"05b30533",
          3015 => x"5758ff57",
          3016 => x"80537a52",
          3017 => x"7951fead",
          3018 => x"3f8287cc",
          3019 => x"08a43875",
          3020 => x"802e8838",
          3021 => x"75812e98",
          3022 => x"38983960",
          3023 => x"557f5482",
          3024 => x"87cc537e",
          3025 => x"527d5177",
          3026 => x"2d8287cc",
          3027 => x"08578339",
          3028 => x"77047682",
          3029 => x"87cc0c89",
          3030 => x"3d0d04f3",
          3031 => x"3d0d7f61",
          3032 => x"63028c05",
          3033 => x"80cf0533",
          3034 => x"73731568",
          3035 => x"415f5c5c",
          3036 => x"5e5e5e7a",
          3037 => x"5281efa0",
          3038 => x"51b3893f",
          3039 => x"81efa851",
          3040 => x"ad9e3f80",
          3041 => x"55747927",
          3042 => x"80f4387b",
          3043 => x"902e8938",
          3044 => x"7ba02ea4",
          3045 => x"3880c139",
          3046 => x"74185372",
          3047 => x"7a278d38",
          3048 => x"72225281",
          3049 => x"efac51b2",
          3050 => x"db3f8839",
          3051 => x"81efb851",
          3052 => x"acee3f82",
          3053 => x"1555bf39",
          3054 => x"74185372",
          3055 => x"7a278d38",
          3056 => x"72085281",
          3057 => x"efa051b2",
          3058 => x"bb3f8839",
          3059 => x"81efb451",
          3060 => x"acce3f84",
          3061 => x"15559f39",
          3062 => x"74185372",
          3063 => x"7a278d38",
          3064 => x"72335281",
          3065 => x"efc051b2",
          3066 => x"9b3f8839",
          3067 => x"81efc851",
          3068 => x"acae3f81",
          3069 => x"1555a051",
          3070 => x"abc93fff",
          3071 => x"883981ef",
          3072 => x"cc51ac9c",
          3073 => x"3f805574",
          3074 => x"7927bb38",
          3075 => x"74187033",
          3076 => x"55538056",
          3077 => x"727a2783",
          3078 => x"38815680",
          3079 => x"539f7427",
          3080 => x"83388153",
          3081 => x"75730670",
          3082 => x"81ff0651",
          3083 => x"5372802e",
          3084 => x"8b387380",
          3085 => x"fe268538",
          3086 => x"73518339",
          3087 => x"a051ab83",
          3088 => x"3f811555",
          3089 => x"c23981ef",
          3090 => x"d051abd4",
          3091 => x"3f781879",
          3092 => x"1c5c58a0",
          3093 => x"9a3f8287",
          3094 => x"cc08982b",
          3095 => x"70982c51",
          3096 => x"5776a02e",
          3097 => x"098106aa",
          3098 => x"38a0843f",
          3099 => x"8287cc08",
          3100 => x"982b7098",
          3101 => x"2c70a032",
          3102 => x"7030729b",
          3103 => x"32703070",
          3104 => x"72077375",
          3105 => x"07065158",
          3106 => x"58595751",
          3107 => x"57807324",
          3108 => x"d838769b",
          3109 => x"2e098106",
          3110 => x"85388053",
          3111 => x"8c397c1e",
          3112 => x"53727826",
          3113 => x"fdcd38ff",
          3114 => x"53728287",
          3115 => x"cc0c8f3d",
          3116 => x"0d04fc3d",
          3117 => x"0d029b05",
          3118 => x"3381efd4",
          3119 => x"5381efdc",
          3120 => x"5255b0c0",
          3121 => x"3f8286a4",
          3122 => x"2251a8dc",
          3123 => x"3f81efe8",
          3124 => x"5481eff4",
          3125 => x"538286a5",
          3126 => x"335281ef",
          3127 => x"fc51b0a4",
          3128 => x"3f74802e",
          3129 => x"8438a4a9",
          3130 => x"3f863d0d",
          3131 => x"04fe3d0d",
          3132 => x"87c09680",
          3133 => x"0853a9b9",
          3134 => x"3f81519b",
          3135 => x"903f81f0",
          3136 => x"98519d83",
          3137 => x"3f80519b",
          3138 => x"843f7281",
          3139 => x"2a708106",
          3140 => x"51527180",
          3141 => x"2e923881",
          3142 => x"519af23f",
          3143 => x"81f0b451",
          3144 => x"9ce53f80",
          3145 => x"519ae63f",
          3146 => x"72822a70",
          3147 => x"81065152",
          3148 => x"71802e92",
          3149 => x"3881519a",
          3150 => x"d43f81f0",
          3151 => x"c8519cc7",
          3152 => x"3f80519a",
          3153 => x"c83f7283",
          3154 => x"2a708106",
          3155 => x"51527180",
          3156 => x"2e923881",
          3157 => x"519ab63f",
          3158 => x"81f0d851",
          3159 => x"9ca93f80",
          3160 => x"519aaa3f",
          3161 => x"72842a70",
          3162 => x"81065152",
          3163 => x"71802e92",
          3164 => x"3881519a",
          3165 => x"983f81f0",
          3166 => x"ec519c8b",
          3167 => x"3f80519a",
          3168 => x"8c3f7285",
          3169 => x"2a708106",
          3170 => x"51527180",
          3171 => x"2e923881",
          3172 => x"5199fa3f",
          3173 => x"81f18051",
          3174 => x"9bed3f80",
          3175 => x"5199ee3f",
          3176 => x"72862a70",
          3177 => x"81065152",
          3178 => x"71802e92",
          3179 => x"38815199",
          3180 => x"dc3f81f1",
          3181 => x"94519bcf",
          3182 => x"3f805199",
          3183 => x"d03f7287",
          3184 => x"2a708106",
          3185 => x"51527180",
          3186 => x"2e923881",
          3187 => x"5199be3f",
          3188 => x"81f1a851",
          3189 => x"9bb13f80",
          3190 => x"5199b23f",
          3191 => x"72882a70",
          3192 => x"81065152",
          3193 => x"71802e92",
          3194 => x"38815199",
          3195 => x"a03f81f1",
          3196 => x"bc519b93",
          3197 => x"3f805199",
          3198 => x"943fa7bd",
          3199 => x"3f843d0d",
          3200 => x"04fb3d0d",
          3201 => x"77028405",
          3202 => x"a3053370",
          3203 => x"55565680",
          3204 => x"527551f4",
          3205 => x"d63f0b0b",
          3206 => x"8282c833",
          3207 => x"5473a938",
          3208 => x"815381f1",
          3209 => x"fc52829e",
          3210 => x"ac518186",
          3211 => x"ea3f8287",
          3212 => x"cc083070",
          3213 => x"8287cc08",
          3214 => x"07802582",
          3215 => x"71315151",
          3216 => x"54730b0b",
          3217 => x"8282c834",
          3218 => x"0b0b8282",
          3219 => x"c8335473",
          3220 => x"812e0981",
          3221 => x"06af3882",
          3222 => x"9eac5374",
          3223 => x"52755181",
          3224 => x"c19b3f82",
          3225 => x"87cc0880",
          3226 => x"2e8b3882",
          3227 => x"87cc0851",
          3228 => x"a7ae3f91",
          3229 => x"39829eac",
          3230 => x"5181938c",
          3231 => x"3f820b0b",
          3232 => x"0b8282c8",
          3233 => x"340b0b82",
          3234 => x"82c83354",
          3235 => x"73822e09",
          3236 => x"81068c38",
          3237 => x"81f28c53",
          3238 => x"74527551",
          3239 => x"b9ba3f80",
          3240 => x"0b8287cc",
          3241 => x"0c873d0d",
          3242 => x"04ce3d0d",
          3243 => x"80707182",
          3244 => x"9ea80c5f",
          3245 => x"5d81527c",
          3246 => x"5180d5b7",
          3247 => x"3f8287cc",
          3248 => x"0881ff06",
          3249 => x"59787d2e",
          3250 => x"098106a1",
          3251 => x"3881f298",
          3252 => x"52963d70",
          3253 => x"5259acc2",
          3254 => x"3f7c5378",
          3255 => x"528288d8",
          3256 => x"518184d2",
          3257 => x"3f8287cc",
          3258 => x"087d2e88",
          3259 => x"3881f29c",
          3260 => x"5191b439",
          3261 => x"81705f5d",
          3262 => x"81f2d451",
          3263 => x"a6a23f96",
          3264 => x"3d70465a",
          3265 => x"80f85279",
          3266 => x"51fdf63f",
          3267 => x"b43dff84",
          3268 => x"0551f3e5",
          3269 => x"3f8287cc",
          3270 => x"08902b70",
          3271 => x"902c5159",
          3272 => x"7880c12e",
          3273 => x"89d13878",
          3274 => x"80c12480",
          3275 => x"d93878ab",
          3276 => x"2e83b838",
          3277 => x"78ab24a4",
          3278 => x"3878822e",
          3279 => x"81b33878",
          3280 => x"82248a38",
          3281 => x"78802eff",
          3282 => x"af388ee1",
          3283 => x"3978842e",
          3284 => x"82833878",
          3285 => x"942e82ad",
          3286 => x"388ed239",
          3287 => x"78bd2e84",
          3288 => x"fa3878bd",
          3289 => x"24903878",
          3290 => x"b02e83a5",
          3291 => x"3878bc2e",
          3292 => x"8483388e",
          3293 => x"b83978bf",
          3294 => x"2e85c138",
          3295 => x"7880c02e",
          3296 => x"86b7388e",
          3297 => x"a8397880",
          3298 => x"d52e8d88",
          3299 => x"387880d5",
          3300 => x"24b03878",
          3301 => x"80d02e8c",
          3302 => x"c1387880",
          3303 => x"d0249238",
          3304 => x"7880c22e",
          3305 => x"89f23878",
          3306 => x"80c32e8b",
          3307 => x"94388dfd",
          3308 => x"397880d1",
          3309 => x"2e8cb238",
          3310 => x"7880d42e",
          3311 => x"8cba388d",
          3312 => x"ec397881",
          3313 => x"822e8dc6",
          3314 => x"38788182",
          3315 => x"24923878",
          3316 => x"80f82e8c",
          3317 => x"db387880",
          3318 => x"f92e8cf7",
          3319 => x"388dce39",
          3320 => x"7881832e",
          3321 => x"8db53878",
          3322 => x"81852e8d",
          3323 => x"ba388dbd",
          3324 => x"39b43dff",
          3325 => x"801153ff",
          3326 => x"840551ab",
          3327 => x"fc3f8287",
          3328 => x"cc088838",
          3329 => x"81f2d851",
          3330 => x"8f9d39b4",
          3331 => x"3dfefc11",
          3332 => x"53ff8405",
          3333 => x"51abe23f",
          3334 => x"8287cc08",
          3335 => x"802e8838",
          3336 => x"81632583",
          3337 => x"38804302",
          3338 => x"80cb0533",
          3339 => x"520280cf",
          3340 => x"05335180",
          3341 => x"d2bd3f82",
          3342 => x"87cc0881",
          3343 => x"ff065978",
          3344 => x"8d3881f2",
          3345 => x"e851a3d8",
          3346 => x"3f815efd",
          3347 => x"ab3981f2",
          3348 => x"f851879d",
          3349 => x"39b43dff",
          3350 => x"801153ff",
          3351 => x"840551ab",
          3352 => x"983f8287",
          3353 => x"cc08802e",
          3354 => x"fd8e3880",
          3355 => x"53805202",
          3356 => x"80cf0533",
          3357 => x"5180d6c8",
          3358 => x"3f8287cc",
          3359 => x"085281f3",
          3360 => x"90518c84",
          3361 => x"39b43dff",
          3362 => x"801153ff",
          3363 => x"840551aa",
          3364 => x"e83f8287",
          3365 => x"cc08802e",
          3366 => x"87386389",
          3367 => x"26fcd938",
          3368 => x"b43dfefc",
          3369 => x"1153ff84",
          3370 => x"0551aacd",
          3371 => x"3f8287cc",
          3372 => x"08863882",
          3373 => x"87cc0843",
          3374 => x"635381f3",
          3375 => x"98527951",
          3376 => x"a8d83f02",
          3377 => x"80cb0533",
          3378 => x"53795263",
          3379 => x"84b42982",
          3380 => x"88d80551",
          3381 => x"8180df3f",
          3382 => x"8287cc08",
          3383 => x"818c3881",
          3384 => x"f2e851a2",
          3385 => x"bb3f815d",
          3386 => x"fc8e39b4",
          3387 => x"3dff8405",
          3388 => x"518f893f",
          3389 => x"8287cc08",
          3390 => x"b53dff84",
          3391 => x"05525b90",
          3392 => x"9f3f8153",
          3393 => x"8287cc08",
          3394 => x"527a51f2",
          3395 => x"c83f80d1",
          3396 => x"39b43dff",
          3397 => x"8405518e",
          3398 => x"e33f8287",
          3399 => x"cc08b53d",
          3400 => x"ff840552",
          3401 => x"5b8ff93f",
          3402 => x"8287cc08",
          3403 => x"b53dff84",
          3404 => x"05525a8f",
          3405 => x"eb3f8287",
          3406 => x"cc08b53d",
          3407 => x"ff840552",
          3408 => x"598fdd3f",
          3409 => x"8285f058",
          3410 => x"8287dc57",
          3411 => x"80568055",
          3412 => x"8287cc08",
          3413 => x"81ff0654",
          3414 => x"78537952",
          3415 => x"7a51f3b2",
          3416 => x"3f8287cc",
          3417 => x"08802efb",
          3418 => x"8f388287",
          3419 => x"cc0851f0",
          3420 => x"833ffb84",
          3421 => x"39b43dff",
          3422 => x"801153ff",
          3423 => x"840551a8",
          3424 => x"f83f8287",
          3425 => x"cc08802e",
          3426 => x"faee38b4",
          3427 => x"3dfefc11",
          3428 => x"53ff8405",
          3429 => x"51a8e23f",
          3430 => x"8287cc08",
          3431 => x"802efad8",
          3432 => x"38b43dfe",
          3433 => x"f81153ff",
          3434 => x"840551a8",
          3435 => x"cc3f8287",
          3436 => x"cc088638",
          3437 => x"8287cc08",
          3438 => x"4281f39c",
          3439 => x"51a0e13f",
          3440 => x"63635c5a",
          3441 => x"797b2781",
          3442 => x"e9386159",
          3443 => x"787a7084",
          3444 => x"055c0c7a",
          3445 => x"7a26f538",
          3446 => x"81d839b4",
          3447 => x"3dff8011",
          3448 => x"53ff8405",
          3449 => x"51a8923f",
          3450 => x"8287cc08",
          3451 => x"802efa88",
          3452 => x"38b43dfe",
          3453 => x"fc1153ff",
          3454 => x"840551a7",
          3455 => x"fc3f8287",
          3456 => x"cc08802e",
          3457 => x"f9f238b4",
          3458 => x"3dfef811",
          3459 => x"53ff8405",
          3460 => x"51a7e63f",
          3461 => x"8287cc08",
          3462 => x"802ef9dc",
          3463 => x"3881f3ac",
          3464 => x"519ffd3f",
          3465 => x"635a7963",
          3466 => x"27818738",
          3467 => x"61597970",
          3468 => x"81055b33",
          3469 => x"79346181",
          3470 => x"0542eb39",
          3471 => x"b43dff80",
          3472 => x"1153ff84",
          3473 => x"0551a7b1",
          3474 => x"3f8287cc",
          3475 => x"08802ef9",
          3476 => x"a738b43d",
          3477 => x"fefc1153",
          3478 => x"ff840551",
          3479 => x"a79b3f82",
          3480 => x"87cc0880",
          3481 => x"2ef99138",
          3482 => x"b43dfef8",
          3483 => x"1153ff84",
          3484 => x"0551a785",
          3485 => x"3f8287cc",
          3486 => x"08802ef8",
          3487 => x"fb3881f3",
          3488 => x"b8519f9c",
          3489 => x"3f635a79",
          3490 => x"6327a738",
          3491 => x"6170337b",
          3492 => x"335e5a5b",
          3493 => x"787c2e91",
          3494 => x"3878557a",
          3495 => x"54793353",
          3496 => x"795281f3",
          3497 => x"c851a4dc",
          3498 => x"3f811a62",
          3499 => x"8105435a",
          3500 => x"d63981f2",
          3501 => x"e45182b9",
          3502 => x"39b43dff",
          3503 => x"801153ff",
          3504 => x"840551a6",
          3505 => x"b43f8287",
          3506 => x"cc0880df",
          3507 => x"388286b8",
          3508 => x"33597880",
          3509 => x"2e893882",
          3510 => x"85f00844",
          3511 => x"80cd3982",
          3512 => x"86b93359",
          3513 => x"78802e88",
          3514 => x"388285f8",
          3515 => x"0844bc39",
          3516 => x"8286ba33",
          3517 => x"5978802e",
          3518 => x"88388286",
          3519 => x"800844ab",
          3520 => x"398286bb",
          3521 => x"33597880",
          3522 => x"2e883882",
          3523 => x"86880844",
          3524 => x"9a398286",
          3525 => x"b6335978",
          3526 => x"802e8838",
          3527 => x"82869008",
          3528 => x"44893982",
          3529 => x"86a008fc",
          3530 => x"800544b4",
          3531 => x"3dfefc11",
          3532 => x"53ff8405",
          3533 => x"51a5c23f",
          3534 => x"8287cc08",
          3535 => x"80de3882",
          3536 => x"86b83359",
          3537 => x"78802e89",
          3538 => x"388285f4",
          3539 => x"084380cc",
          3540 => x"398286b9",
          3541 => x"33597880",
          3542 => x"2e883882",
          3543 => x"85fc0843",
          3544 => x"bb398286",
          3545 => x"ba335978",
          3546 => x"802e8838",
          3547 => x"82868408",
          3548 => x"43aa3982",
          3549 => x"86bb3359",
          3550 => x"78802e88",
          3551 => x"3882868c",
          3552 => x"08439939",
          3553 => x"8286b633",
          3554 => x"5978802e",
          3555 => x"88388286",
          3556 => x"94084388",
          3557 => x"398286a0",
          3558 => x"08880543",
          3559 => x"b43dfef8",
          3560 => x"1153ff84",
          3561 => x"0551a4d1",
          3562 => x"3f8287cc",
          3563 => x"08802ea7",
          3564 => x"3880625c",
          3565 => x"5c7a882e",
          3566 => x"8338815c",
          3567 => x"7a903270",
          3568 => x"30707207",
          3569 => x"9f2a707f",
          3570 => x"0651515a",
          3571 => x"5a78802e",
          3572 => x"88387aa0",
          3573 => x"2e833888",
          3574 => x"4281f3e4",
          3575 => x"519cc13f",
          3576 => x"a0556354",
          3577 => x"61536252",
          3578 => x"6351eeef",
          3579 => x"3f81f3f4",
          3580 => x"519cad3f",
          3581 => x"f68239b4",
          3582 => x"3dff8011",
          3583 => x"53ff8405",
          3584 => x"51a3f63f",
          3585 => x"8287cc08",
          3586 => x"802ef5ec",
          3587 => x"38b43dfe",
          3588 => x"fc1153ff",
          3589 => x"840551a3",
          3590 => x"e03f8287",
          3591 => x"cc08802e",
          3592 => x"a4386359",
          3593 => x"0280cb05",
          3594 => x"33793463",
          3595 => x"810544b4",
          3596 => x"3dfefc11",
          3597 => x"53ff8405",
          3598 => x"51a3be3f",
          3599 => x"8287cc08",
          3600 => x"e138f5b4",
          3601 => x"39637033",
          3602 => x"545281f4",
          3603 => x"8051a1b4",
          3604 => x"3f80f852",
          3605 => x"7951a286",
          3606 => x"3f794579",
          3607 => x"335978ae",
          3608 => x"2ef59538",
          3609 => x"9f79279f",
          3610 => x"38b43dfe",
          3611 => x"fc1153ff",
          3612 => x"840551a3",
          3613 => x"843f8287",
          3614 => x"cc08802e",
          3615 => x"91386359",
          3616 => x"0280cb05",
          3617 => x"33793463",
          3618 => x"810544ff",
          3619 => x"b83981f4",
          3620 => x"8c519b8c",
          3621 => x"3fffae39",
          3622 => x"b43dfef4",
          3623 => x"1153ff84",
          3624 => x"0551a4c7",
          3625 => x"3f8287cc",
          3626 => x"08802ef4",
          3627 => x"cb38b43d",
          3628 => x"fef01153",
          3629 => x"ff840551",
          3630 => x"a4b13f82",
          3631 => x"87cc0880",
          3632 => x"2ea53860",
          3633 => x"5902be05",
          3634 => x"22797082",
          3635 => x"055b2378",
          3636 => x"41b43dfe",
          3637 => x"f01153ff",
          3638 => x"840551a4",
          3639 => x"8e3f8287",
          3640 => x"cc08e038",
          3641 => x"f4923960",
          3642 => x"70225452",
          3643 => x"81f49451",
          3644 => x"a0923f80",
          3645 => x"f8527951",
          3646 => x"a0e43f79",
          3647 => x"45793359",
          3648 => x"78ae2ef3",
          3649 => x"f338789f",
          3650 => x"26873860",
          3651 => x"820541d7",
          3652 => x"39b43dfe",
          3653 => x"f01153ff",
          3654 => x"840551a3",
          3655 => x"ce3f8287",
          3656 => x"cc08802e",
          3657 => x"92386059",
          3658 => x"02be0522",
          3659 => x"79708205",
          3660 => x"5b237841",
          3661 => x"ffb13981",
          3662 => x"f48c5199",
          3663 => x"e33fffa7",
          3664 => x"39b43dfe",
          3665 => x"f41153ff",
          3666 => x"840551a3",
          3667 => x"9e3f8287",
          3668 => x"cc08802e",
          3669 => x"f3a238b4",
          3670 => x"3dfef011",
          3671 => x"53ff8405",
          3672 => x"51a3883f",
          3673 => x"8287cc08",
          3674 => x"802ea038",
          3675 => x"6060710c",
          3676 => x"59608405",
          3677 => x"41b43dfe",
          3678 => x"f01153ff",
          3679 => x"840551a2",
          3680 => x"ea3f8287",
          3681 => x"cc08e538",
          3682 => x"f2ee3960",
          3683 => x"70085452",
          3684 => x"81f4a051",
          3685 => x"9eee3f80",
          3686 => x"f8527951",
          3687 => x"9fc03f79",
          3688 => x"45793359",
          3689 => x"78ae2ef2",
          3690 => x"cf389f79",
          3691 => x"279b38b4",
          3692 => x"3dfef011",
          3693 => x"53ff8405",
          3694 => x"51a2b03f",
          3695 => x"8287cc08",
          3696 => x"802e8d38",
          3697 => x"6060710c",
          3698 => x"59608405",
          3699 => x"41ffbc39",
          3700 => x"81f48c51",
          3701 => x"98ca3fff",
          3702 => x"b23981f4",
          3703 => x"ac5198c0",
          3704 => x"3f825197",
          3705 => x"a73ff290",
          3706 => x"3981f4c4",
          3707 => x"5198b13f",
          3708 => x"a25196fc",
          3709 => x"3ff28139",
          3710 => x"81f4dc51",
          3711 => x"98a23f84",
          3712 => x"80810b87",
          3713 => x"c094840c",
          3714 => x"8480810b",
          3715 => x"87c09494",
          3716 => x"0cf1e539",
          3717 => x"81f4f051",
          3718 => x"98863f8c",
          3719 => x"80830b87",
          3720 => x"c094840c",
          3721 => x"8c80830b",
          3722 => x"87c09494",
          3723 => x"0cf1c939",
          3724 => x"b43dff80",
          3725 => x"1153ff84",
          3726 => x"05519fbd",
          3727 => x"3f8287cc",
          3728 => x"08802ef1",
          3729 => x"b3386352",
          3730 => x"81f58451",
          3731 => x"9db63f63",
          3732 => x"597804b4",
          3733 => x"3dff8011",
          3734 => x"53ff8405",
          3735 => x"519f9a3f",
          3736 => x"8287cc08",
          3737 => x"802ef190",
          3738 => x"38635281",
          3739 => x"f5a0519d",
          3740 => x"933f6359",
          3741 => x"782d8287",
          3742 => x"cc08802e",
          3743 => x"f0fa3882",
          3744 => x"87cc0852",
          3745 => x"81f5bc51",
          3746 => x"9cfa3ff0",
          3747 => x"eb3981f5",
          3748 => x"d851978c",
          3749 => x"3fde823f",
          3750 => x"f0de3981",
          3751 => x"f5f45196",
          3752 => x"ff3f8059",
          3753 => x"ffab3990",
          3754 => x"e83ff0cc",
          3755 => x"39794579",
          3756 => x"33597880",
          3757 => x"2ef0c138",
          3758 => x"7d7d0659",
          3759 => x"78802e81",
          3760 => x"ce38b43d",
          3761 => x"ff840551",
          3762 => x"83b23f82",
          3763 => x"87cc085b",
          3764 => x"815c7b82",
          3765 => x"2eb1387b",
          3766 => x"82248938",
          3767 => x"7b812e8c",
          3768 => x"3880ca39",
          3769 => x"7b832eae",
          3770 => x"3880c239",
          3771 => x"81f68856",
          3772 => x"7a5581f6",
          3773 => x"8c548053",
          3774 => x"81f69052",
          3775 => x"b43dffb0",
          3776 => x"05519c96",
          3777 => x"3fb83981",
          3778 => x"f6b052b4",
          3779 => x"3dffb005",
          3780 => x"519c873f",
          3781 => x"a9397a55",
          3782 => x"81f68c54",
          3783 => x"805381f6",
          3784 => x"a052b43d",
          3785 => x"ffb00551",
          3786 => x"9bf03f92",
          3787 => x"397a5480",
          3788 => x"5381f6ac",
          3789 => x"52b43dff",
          3790 => x"b005519b",
          3791 => x"dd3f8285",
          3792 => x"f0588287",
          3793 => x"dc578056",
          3794 => x"64558054",
          3795 => x"82a08053",
          3796 => x"82a08052",
          3797 => x"b43dffb0",
          3798 => x"0551e7b6",
          3799 => x"3f8287cc",
          3800 => x"088287cc",
          3801 => x"08097030",
          3802 => x"70720780",
          3803 => x"25515b5b",
          3804 => x"5f805a7b",
          3805 => x"83268338",
          3806 => x"815a787a",
          3807 => x"06597880",
          3808 => x"2e8d3881",
          3809 => x"1c7081ff",
          3810 => x"065d597b",
          3811 => x"fec4387d",
          3812 => x"81327d81",
          3813 => x"32075978",
          3814 => x"8a387eff",
          3815 => x"2e098106",
          3816 => x"eed63881",
          3817 => x"f6b4519a",
          3818 => x"db3feecc",
          3819 => x"39fc3d0d",
          3820 => x"800b8287",
          3821 => x"dc3487c0",
          3822 => x"948c7008",
          3823 => x"54558784",
          3824 => x"80527251",
          3825 => x"b4a53f82",
          3826 => x"87cc0890",
          3827 => x"2b750855",
          3828 => x"53878480",
          3829 => x"527351b4",
          3830 => x"923f7282",
          3831 => x"87cc0807",
          3832 => x"750c87c0",
          3833 => x"949c7008",
          3834 => x"54558784",
          3835 => x"80527251",
          3836 => x"b3f93f82",
          3837 => x"87cc0890",
          3838 => x"2b750855",
          3839 => x"53878480",
          3840 => x"527351b3",
          3841 => x"e63f7282",
          3842 => x"87cc0807",
          3843 => x"750c8c80",
          3844 => x"830b87c0",
          3845 => x"94840c8c",
          3846 => x"80830b87",
          3847 => x"c094940c",
          3848 => x"bda50b82",
          3849 => x"9ed40c80",
          3850 => x"c0a00b82",
          3851 => x"9ed80c89",
          3852 => x"943f92fd",
          3853 => x"3f81f6c4",
          3854 => x"5193e53f",
          3855 => x"81f6d051",
          3856 => x"93de3fa1",
          3857 => x"ed5192a3",
          3858 => x"3f8151e8",
          3859 => x"e53fecd9",
          3860 => x"3f8004fe",
          3861 => x"3d0d8052",
          3862 => x"83537188",
          3863 => x"2b5287c0",
          3864 => x"3f8287cc",
          3865 => x"0881ff06",
          3866 => x"7207ff14",
          3867 => x"54527280",
          3868 => x"25e83871",
          3869 => x"8287cc0c",
          3870 => x"843d0d04",
          3871 => x"fc3d0d76",
          3872 => x"70085455",
          3873 => x"80735254",
          3874 => x"72742e81",
          3875 => x"8a387233",
          3876 => x"5170a02e",
          3877 => x"09810686",
          3878 => x"38811353",
          3879 => x"f1397233",
          3880 => x"5170a22e",
          3881 => x"09810686",
          3882 => x"38811353",
          3883 => x"81547252",
          3884 => x"73812e09",
          3885 => x"81069f38",
          3886 => x"84398112",
          3887 => x"52807233",
          3888 => x"525470a2",
          3889 => x"2e833881",
          3890 => x"5470802e",
          3891 => x"9d3873ea",
          3892 => x"38983981",
          3893 => x"12528072",
          3894 => x"33525470",
          3895 => x"a02e8338",
          3896 => x"81547080",
          3897 => x"2e843873",
          3898 => x"ea388072",
          3899 => x"33525470",
          3900 => x"a02e0981",
          3901 => x"06833881",
          3902 => x"5470a232",
          3903 => x"70307080",
          3904 => x"25760751",
          3905 => x"51517080",
          3906 => x"2e883880",
          3907 => x"72708105",
          3908 => x"54347175",
          3909 => x"0c725170",
          3910 => x"8287cc0c",
          3911 => x"863d0d04",
          3912 => x"fc3d0d76",
          3913 => x"53720880",
          3914 => x"2e913886",
          3915 => x"3dfc0552",
          3916 => x"72519bb7",
          3917 => x"3f8287cc",
          3918 => x"08853880",
          3919 => x"53833974",
          3920 => x"53728287",
          3921 => x"cc0c863d",
          3922 => x"0d04fc3d",
          3923 => x"0d768211",
          3924 => x"33ff0552",
          3925 => x"53815270",
          3926 => x"8b268198",
          3927 => x"38831333",
          3928 => x"ff055182",
          3929 => x"52709e26",
          3930 => x"818a3884",
          3931 => x"13335183",
          3932 => x"52709726",
          3933 => x"80fe3885",
          3934 => x"13335184",
          3935 => x"5270bb26",
          3936 => x"80f23886",
          3937 => x"13335185",
          3938 => x"5270bb26",
          3939 => x"80e63888",
          3940 => x"13225586",
          3941 => x"527487e7",
          3942 => x"2680d938",
          3943 => x"8a132254",
          3944 => x"87527387",
          3945 => x"e72680cc",
          3946 => x"38810b87",
          3947 => x"c0989c0c",
          3948 => x"722287c0",
          3949 => x"98bc0c82",
          3950 => x"133387c0",
          3951 => x"98b80c83",
          3952 => x"133387c0",
          3953 => x"98b40c84",
          3954 => x"133387c0",
          3955 => x"98b00c85",
          3956 => x"133387c0",
          3957 => x"98ac0c86",
          3958 => x"133387c0",
          3959 => x"98a80c74",
          3960 => x"87c098a4",
          3961 => x"0c7387c0",
          3962 => x"98a00c80",
          3963 => x"0b87c098",
          3964 => x"9c0c8052",
          3965 => x"718287cc",
          3966 => x"0c863d0d",
          3967 => x"04f33d0d",
          3968 => x"7f5b87c0",
          3969 => x"989c5d81",
          3970 => x"7d0c87c0",
          3971 => x"98bc085e",
          3972 => x"7d7b2387",
          3973 => x"c098b808",
          3974 => x"5a79821c",
          3975 => x"3487c098",
          3976 => x"b4085a79",
          3977 => x"831c3487",
          3978 => x"c098b008",
          3979 => x"5a79841c",
          3980 => x"3487c098",
          3981 => x"ac085a79",
          3982 => x"851c3487",
          3983 => x"c098a808",
          3984 => x"5a79861c",
          3985 => x"3487c098",
          3986 => x"a4085c7b",
          3987 => x"881c2387",
          3988 => x"c098a008",
          3989 => x"5a798a1c",
          3990 => x"23807d0c",
          3991 => x"7983ffff",
          3992 => x"06597b83",
          3993 => x"ffff0658",
          3994 => x"861b3357",
          3995 => x"851b3356",
          3996 => x"841b3355",
          3997 => x"831b3354",
          3998 => x"821b3353",
          3999 => x"7d83ffff",
          4000 => x"065281f6",
          4001 => x"e85194fc",
          4002 => x"3f8f3d0d",
          4003 => x"04ff3d0d",
          4004 => x"028f0533",
          4005 => x"7030709f",
          4006 => x"2a515252",
          4007 => x"708285ec",
          4008 => x"34833d0d",
          4009 => x"04fb3d0d",
          4010 => x"778285ec",
          4011 => x"337081ff",
          4012 => x"06575556",
          4013 => x"87c09484",
          4014 => x"5174802e",
          4015 => x"863887c0",
          4016 => x"94945170",
          4017 => x"0870962a",
          4018 => x"70810653",
          4019 => x"54527080",
          4020 => x"2e8c3871",
          4021 => x"912a7081",
          4022 => x"06515170",
          4023 => x"d7387281",
          4024 => x"32708106",
          4025 => x"51517080",
          4026 => x"2e8d3871",
          4027 => x"932a7081",
          4028 => x"06515170",
          4029 => x"ffbe3873",
          4030 => x"81ff0651",
          4031 => x"87c09480",
          4032 => x"5270802e",
          4033 => x"863887c0",
          4034 => x"94905275",
          4035 => x"720c7582",
          4036 => x"87cc0c87",
          4037 => x"3d0d04fb",
          4038 => x"3d0d029f",
          4039 => x"05338285",
          4040 => x"ec337081",
          4041 => x"ff065755",
          4042 => x"5687c094",
          4043 => x"84517480",
          4044 => x"2e863887",
          4045 => x"c0949451",
          4046 => x"70087096",
          4047 => x"2a708106",
          4048 => x"53545270",
          4049 => x"802e8c38",
          4050 => x"71912a70",
          4051 => x"81065151",
          4052 => x"70d73872",
          4053 => x"81327081",
          4054 => x"06515170",
          4055 => x"802e8d38",
          4056 => x"71932a70",
          4057 => x"81065151",
          4058 => x"70ffbe38",
          4059 => x"7381ff06",
          4060 => x"5187c094",
          4061 => x"80527080",
          4062 => x"2e863887",
          4063 => x"c0949052",
          4064 => x"75720c87",
          4065 => x"3d0d04f9",
          4066 => x"3d0d7954",
          4067 => x"80743370",
          4068 => x"81ff0653",
          4069 => x"53577077",
          4070 => x"2e80fc38",
          4071 => x"7181ff06",
          4072 => x"81158285",
          4073 => x"ec337081",
          4074 => x"ff065957",
          4075 => x"555887c0",
          4076 => x"94845175",
          4077 => x"802e8638",
          4078 => x"87c09494",
          4079 => x"51700870",
          4080 => x"962a7081",
          4081 => x"06535452",
          4082 => x"70802e8c",
          4083 => x"3871912a",
          4084 => x"70810651",
          4085 => x"5170d738",
          4086 => x"72813270",
          4087 => x"81065151",
          4088 => x"70802e8d",
          4089 => x"3871932a",
          4090 => x"70810651",
          4091 => x"5170ffbe",
          4092 => x"387481ff",
          4093 => x"065187c0",
          4094 => x"94805270",
          4095 => x"802e8638",
          4096 => x"87c09490",
          4097 => x"5277720c",
          4098 => x"81177433",
          4099 => x"7081ff06",
          4100 => x"53535770",
          4101 => x"ff863876",
          4102 => x"8287cc0c",
          4103 => x"893d0d04",
          4104 => x"fe3d0d82",
          4105 => x"85ec3370",
          4106 => x"81ff0654",
          4107 => x"5287c094",
          4108 => x"84517280",
          4109 => x"2e863887",
          4110 => x"c0949451",
          4111 => x"70087082",
          4112 => x"2a708106",
          4113 => x"51515170",
          4114 => x"802ee238",
          4115 => x"7181ff06",
          4116 => x"5187c094",
          4117 => x"80527080",
          4118 => x"2e863887",
          4119 => x"c0949052",
          4120 => x"71087081",
          4121 => x"ff068287",
          4122 => x"cc0c5184",
          4123 => x"3d0d04fe",
          4124 => x"3d0d8285",
          4125 => x"ec337081",
          4126 => x"ff065253",
          4127 => x"87c09484",
          4128 => x"5270802e",
          4129 => x"863887c0",
          4130 => x"94945271",
          4131 => x"0870822a",
          4132 => x"70810651",
          4133 => x"5151ff52",
          4134 => x"70802ea0",
          4135 => x"387281ff",
          4136 => x"065187c0",
          4137 => x"94805270",
          4138 => x"802e8638",
          4139 => x"87c09490",
          4140 => x"52710870",
          4141 => x"982b7098",
          4142 => x"2c515351",
          4143 => x"718287cc",
          4144 => x"0c843d0d",
          4145 => x"04ff3d0d",
          4146 => x"87c09e80",
          4147 => x"08709c2a",
          4148 => x"8a065151",
          4149 => x"70802e84",
          4150 => x"b43887c0",
          4151 => x"9ea40882",
          4152 => x"85f00c87",
          4153 => x"c09ea808",
          4154 => x"8285f40c",
          4155 => x"87c09e94",
          4156 => x"088285f8",
          4157 => x"0c87c09e",
          4158 => x"98088285",
          4159 => x"fc0c87c0",
          4160 => x"9e9c0882",
          4161 => x"86800c87",
          4162 => x"c09ea008",
          4163 => x"8286840c",
          4164 => x"87c09eac",
          4165 => x"08828688",
          4166 => x"0c87c09e",
          4167 => x"b0088286",
          4168 => x"8c0c87c0",
          4169 => x"9eb40882",
          4170 => x"86900c87",
          4171 => x"c09eb808",
          4172 => x"8286940c",
          4173 => x"87c09ebc",
          4174 => x"08828698",
          4175 => x"0c87c09e",
          4176 => x"c0088286",
          4177 => x"9c0c87c0",
          4178 => x"9ec40882",
          4179 => x"86a00c87",
          4180 => x"c09e8008",
          4181 => x"51708286",
          4182 => x"a42387c0",
          4183 => x"9e840882",
          4184 => x"86a80c87",
          4185 => x"c09e8808",
          4186 => x"8286ac0c",
          4187 => x"87c09e8c",
          4188 => x"088286b0",
          4189 => x"0c810b82",
          4190 => x"86b43480",
          4191 => x"0b87c09e",
          4192 => x"90087084",
          4193 => x"800a0651",
          4194 => x"52527080",
          4195 => x"2e833881",
          4196 => x"52718286",
          4197 => x"b534800b",
          4198 => x"87c09e90",
          4199 => x"08708880",
          4200 => x"0a065152",
          4201 => x"5270802e",
          4202 => x"83388152",
          4203 => x"718286b6",
          4204 => x"34800b87",
          4205 => x"c09e9008",
          4206 => x"7090800a",
          4207 => x"06515252",
          4208 => x"70802e83",
          4209 => x"38815271",
          4210 => x"8286b734",
          4211 => x"800b87c0",
          4212 => x"9e900870",
          4213 => x"88808006",
          4214 => x"51525270",
          4215 => x"802e8338",
          4216 => x"81527182",
          4217 => x"86b83480",
          4218 => x"0b87c09e",
          4219 => x"900870a0",
          4220 => x"80800651",
          4221 => x"52527080",
          4222 => x"2e833881",
          4223 => x"52718286",
          4224 => x"b934800b",
          4225 => x"87c09e90",
          4226 => x"08709080",
          4227 => x"80065152",
          4228 => x"5270802e",
          4229 => x"83388152",
          4230 => x"718286ba",
          4231 => x"34800b87",
          4232 => x"c09e9008",
          4233 => x"70848080",
          4234 => x"06515252",
          4235 => x"70802e83",
          4236 => x"38815271",
          4237 => x"8286bb34",
          4238 => x"800b87c0",
          4239 => x"9e900870",
          4240 => x"82808006",
          4241 => x"51525270",
          4242 => x"802e8338",
          4243 => x"81527182",
          4244 => x"86bc3480",
          4245 => x"0b87c09e",
          4246 => x"90087081",
          4247 => x"80800651",
          4248 => x"52527080",
          4249 => x"2e833881",
          4250 => x"52718286",
          4251 => x"bd34800b",
          4252 => x"87c09e90",
          4253 => x"087080c0",
          4254 => x"80065152",
          4255 => x"5270802e",
          4256 => x"83388152",
          4257 => x"718286be",
          4258 => x"34800b87",
          4259 => x"c09e9008",
          4260 => x"70a08006",
          4261 => x"51525270",
          4262 => x"802e8338",
          4263 => x"81527182",
          4264 => x"86bf3487",
          4265 => x"c09e9008",
          4266 => x"70988006",
          4267 => x"708a2a51",
          4268 => x"51517082",
          4269 => x"86c03480",
          4270 => x"0b87c09e",
          4271 => x"90087084",
          4272 => x"80065152",
          4273 => x"5270802e",
          4274 => x"83388152",
          4275 => x"718286c1",
          4276 => x"3487c09e",
          4277 => x"90087083",
          4278 => x"f0067084",
          4279 => x"2a515151",
          4280 => x"708286c2",
          4281 => x"34800b87",
          4282 => x"c09e9008",
          4283 => x"70880651",
          4284 => x"52527080",
          4285 => x"2e833881",
          4286 => x"52718286",
          4287 => x"c33487c0",
          4288 => x"9e900870",
          4289 => x"87065151",
          4290 => x"708286c4",
          4291 => x"34833d0d",
          4292 => x"04fb3d0d",
          4293 => x"81f78051",
          4294 => x"86863f82",
          4295 => x"86b43354",
          4296 => x"73802e88",
          4297 => x"3881f794",
          4298 => x"5185f53f",
          4299 => x"81f7a851",
          4300 => x"85ee3f82",
          4301 => x"86b63354",
          4302 => x"73802e93",
          4303 => x"38828690",
          4304 => x"08828694",
          4305 => x"08115452",
          4306 => x"81f7c051",
          4307 => x"8bb63f82",
          4308 => x"86bb3354",
          4309 => x"73802e93",
          4310 => x"38828688",
          4311 => x"0882868c",
          4312 => x"08115452",
          4313 => x"81f7dc51",
          4314 => x"8b9a3f82",
          4315 => x"86b83354",
          4316 => x"73802e93",
          4317 => x"388285f0",
          4318 => x"088285f4",
          4319 => x"08115452",
          4320 => x"81f7f851",
          4321 => x"8afe3f82",
          4322 => x"86b93354",
          4323 => x"73802e93",
          4324 => x"388285f8",
          4325 => x"088285fc",
          4326 => x"08115452",
          4327 => x"81f89451",
          4328 => x"8ae23f82",
          4329 => x"86ba3354",
          4330 => x"73802e93",
          4331 => x"38828680",
          4332 => x"08828684",
          4333 => x"08115452",
          4334 => x"81f8b051",
          4335 => x"8ac63f82",
          4336 => x"86bf3354",
          4337 => x"73802e8d",
          4338 => x"388286c0",
          4339 => x"335281f8",
          4340 => x"cc518ab0",
          4341 => x"3f8286c3",
          4342 => x"33547380",
          4343 => x"2e8d3882",
          4344 => x"86c43352",
          4345 => x"81f8ec51",
          4346 => x"8a9a3f82",
          4347 => x"86c13354",
          4348 => x"73802e8d",
          4349 => x"388286c2",
          4350 => x"335281f9",
          4351 => x"8c518a84",
          4352 => x"3f8286b5",
          4353 => x"33547380",
          4354 => x"2e883881",
          4355 => x"f9ac5184",
          4356 => x"8f3f8286",
          4357 => x"b7335473",
          4358 => x"802e8838",
          4359 => x"81f9c051",
          4360 => x"83fe3f82",
          4361 => x"86bc3354",
          4362 => x"73802e88",
          4363 => x"3881f9cc",
          4364 => x"5183ed3f",
          4365 => x"8286bd33",
          4366 => x"5473802e",
          4367 => x"883881f9",
          4368 => x"d85183dc",
          4369 => x"3f8286be",
          4370 => x"33547380",
          4371 => x"2e883881",
          4372 => x"f9e45183",
          4373 => x"cb3f81f9",
          4374 => x"f05183c4",
          4375 => x"3f828698",
          4376 => x"085281f9",
          4377 => x"fc51899c",
          4378 => x"3f82869c",
          4379 => x"085281fa",
          4380 => x"a4518990",
          4381 => x"3f8286a0",
          4382 => x"085281fa",
          4383 => x"cc518984",
          4384 => x"3f81faf4",
          4385 => x"5183993f",
          4386 => x"8286a422",
          4387 => x"5281fafc",
          4388 => x"5188f13f",
          4389 => x"8286a808",
          4390 => x"56bd84c0",
          4391 => x"527551a2",
          4392 => x"ca3f8287",
          4393 => x"cc08bd84",
          4394 => x"c0297671",
          4395 => x"31545482",
          4396 => x"87cc0852",
          4397 => x"81fba451",
          4398 => x"88ca3f82",
          4399 => x"86bb3354",
          4400 => x"73802ea8",
          4401 => x"388286ac",
          4402 => x"0856bd84",
          4403 => x"c0527551",
          4404 => x"a2993f82",
          4405 => x"87cc08bd",
          4406 => x"84c02976",
          4407 => x"71315454",
          4408 => x"8287cc08",
          4409 => x"5281fbd0",
          4410 => x"5188993f",
          4411 => x"8286b633",
          4412 => x"5473802e",
          4413 => x"a8388286",
          4414 => x"b00856bd",
          4415 => x"84c05275",
          4416 => x"51a1e83f",
          4417 => x"8287cc08",
          4418 => x"bd84c029",
          4419 => x"76713154",
          4420 => x"548287cc",
          4421 => x"085281fb",
          4422 => x"fc5187e8",
          4423 => x"3f81f2e4",
          4424 => x"5181fd3f",
          4425 => x"873d0d04",
          4426 => x"fe3d0d02",
          4427 => x"920533ff",
          4428 => x"05527184",
          4429 => x"26aa3871",
          4430 => x"842981e9",
          4431 => x"94055271",
          4432 => x"080481fc",
          4433 => x"a8519d39",
          4434 => x"81fcb051",
          4435 => x"973981fc",
          4436 => x"b8519139",
          4437 => x"81fcc051",
          4438 => x"8b3981fc",
          4439 => x"c4518539",
          4440 => x"81fccc51",
          4441 => x"81ba3f84",
          4442 => x"3d0d0471",
          4443 => x"88800c04",
          4444 => x"ff3d0d87",
          4445 => x"c0968470",
          4446 => x"08525280",
          4447 => x"720c7074",
          4448 => x"07708286",
          4449 => x"c80c720c",
          4450 => x"833d0d04",
          4451 => x"ff3d0d87",
          4452 => x"c0968470",
          4453 => x"088286c8",
          4454 => x"0c528072",
          4455 => x"0c730970",
          4456 => x"8286c808",
          4457 => x"06708286",
          4458 => x"c80c730c",
          4459 => x"51833d0d",
          4460 => x"04800b87",
          4461 => x"c096840c",
          4462 => x"048286c8",
          4463 => x"0887c096",
          4464 => x"840c04fe",
          4465 => x"3d0d0293",
          4466 => x"05335372",
          4467 => x"8a2e0981",
          4468 => x"0685388d",
          4469 => x"51ed3f82",
          4470 => x"9edc0852",
          4471 => x"71802e90",
          4472 => x"38727234",
          4473 => x"829edc08",
          4474 => x"8105829e",
          4475 => x"dc0c8f39",
          4476 => x"829ed408",
          4477 => x"5271802e",
          4478 => x"85387251",
          4479 => x"712d843d",
          4480 => x"0d04fe3d",
          4481 => x"0d029705",
          4482 => x"33829ed4",
          4483 => x"0876829e",
          4484 => x"d40c5451",
          4485 => x"ffad3f72",
          4486 => x"829ed40c",
          4487 => x"843d0d04",
          4488 => x"fd3d0d75",
          4489 => x"54733370",
          4490 => x"81ff0653",
          4491 => x"5371802e",
          4492 => x"8e387281",
          4493 => x"ff065181",
          4494 => x"1454ff87",
          4495 => x"3fe73985",
          4496 => x"3d0d04fc",
          4497 => x"3d0d7782",
          4498 => x"9ed40878",
          4499 => x"829ed40c",
          4500 => x"56547333",
          4501 => x"7081ff06",
          4502 => x"53537180",
          4503 => x"2e8e3872",
          4504 => x"81ff0651",
          4505 => x"811454fe",
          4506 => x"da3fe739",
          4507 => x"74829ed4",
          4508 => x"0c863d0d",
          4509 => x"04ec3d0d",
          4510 => x"66685959",
          4511 => x"78708105",
          4512 => x"5a335675",
          4513 => x"802e84f8",
          4514 => x"3875a52e",
          4515 => x"09810682",
          4516 => x"de388070",
          4517 => x"7a708105",
          4518 => x"5c33585b",
          4519 => x"5b75b02e",
          4520 => x"09810685",
          4521 => x"38815a8b",
          4522 => x"3975ad2e",
          4523 => x"0981068a",
          4524 => x"38825a78",
          4525 => x"7081055a",
          4526 => x"335675aa",
          4527 => x"2e098106",
          4528 => x"92387784",
          4529 => x"1971087b",
          4530 => x"7081055d",
          4531 => x"33595d59",
          4532 => x"539d39d0",
          4533 => x"16537289",
          4534 => x"2695387a",
          4535 => x"88297b10",
          4536 => x"057605d0",
          4537 => x"05797081",
          4538 => x"055b3357",
          4539 => x"5be53975",
          4540 => x"80ec3270",
          4541 => x"30707207",
          4542 => x"80257880",
          4543 => x"cc327030",
          4544 => x"70720780",
          4545 => x"25730753",
          4546 => x"54585155",
          4547 => x"5373802e",
          4548 => x"8c387984",
          4549 => x"07797081",
          4550 => x"055b3357",
          4551 => x"5a75802e",
          4552 => x"83de3875",
          4553 => x"5480e076",
          4554 => x"278938e0",
          4555 => x"167081ff",
          4556 => x"06555373",
          4557 => x"80cf2e81",
          4558 => x"aa387380",
          4559 => x"cf24a238",
          4560 => x"7380c32e",
          4561 => x"818e3873",
          4562 => x"80c3248b",
          4563 => x"387380c2",
          4564 => x"2e818c38",
          4565 => x"81993973",
          4566 => x"80c42e81",
          4567 => x"8a38818f",
          4568 => x"397380d5",
          4569 => x"2e818038",
          4570 => x"7380d524",
          4571 => x"8a387380",
          4572 => x"d32e8e38",
          4573 => x"80f93973",
          4574 => x"80d82e80",
          4575 => x"ee3880ef",
          4576 => x"39778419",
          4577 => x"71085659",
          4578 => x"53807433",
          4579 => x"54557275",
          4580 => x"2e8d3881",
          4581 => x"15701570",
          4582 => x"33515455",
          4583 => x"72f53879",
          4584 => x"812a5690",
          4585 => x"39748116",
          4586 => x"5653727b",
          4587 => x"278f38a0",
          4588 => x"51fc903f",
          4589 => x"75810653",
          4590 => x"72802ee9",
          4591 => x"387351fc",
          4592 => x"df3f7481",
          4593 => x"16565372",
          4594 => x"7b27fdb0",
          4595 => x"38a051fb",
          4596 => x"f23fef39",
          4597 => x"77841983",
          4598 => x"12335359",
          4599 => x"53933982",
          4600 => x"5c953988",
          4601 => x"5c91398a",
          4602 => x"5c8d3990",
          4603 => x"5c893975",
          4604 => x"51fbd03f",
          4605 => x"fd863979",
          4606 => x"822a7081",
          4607 => x"06515372",
          4608 => x"802e8838",
          4609 => x"77841959",
          4610 => x"53863984",
          4611 => x"18785458",
          4612 => x"72087480",
          4613 => x"c4327030",
          4614 => x"70720780",
          4615 => x"25515555",
          4616 => x"55748025",
          4617 => x"8d387280",
          4618 => x"2e883874",
          4619 => x"307a9007",
          4620 => x"5b55800b",
          4621 => x"8f3d5e57",
          4622 => x"7b527451",
          4623 => x"9dd43f82",
          4624 => x"87cc0881",
          4625 => x"ff067c53",
          4626 => x"7552549b",
          4627 => x"9e3f8287",
          4628 => x"cc085589",
          4629 => x"74279238",
          4630 => x"a7145375",
          4631 => x"80f82e84",
          4632 => x"38871453",
          4633 => x"7281ff06",
          4634 => x"54b01453",
          4635 => x"727d7081",
          4636 => x"055f3481",
          4637 => x"17753070",
          4638 => x"77079f2a",
          4639 => x"51545776",
          4640 => x"9f268538",
          4641 => x"72ffb138",
          4642 => x"79842a70",
          4643 => x"81065153",
          4644 => x"72802e8e",
          4645 => x"38963d77",
          4646 => x"05e00553",
          4647 => x"ad733481",
          4648 => x"1757767a",
          4649 => x"81065455",
          4650 => x"b0547283",
          4651 => x"38a05479",
          4652 => x"812a7081",
          4653 => x"06545672",
          4654 => x"9f388117",
          4655 => x"55767b27",
          4656 => x"97387351",
          4657 => x"f9fd3f75",
          4658 => x"81065372",
          4659 => x"8b387481",
          4660 => x"1656537a",
          4661 => x"7326eb38",
          4662 => x"963d7705",
          4663 => x"e00553ff",
          4664 => x"17ff1470",
          4665 => x"33535457",
          4666 => x"f9d93f76",
          4667 => x"f2387481",
          4668 => x"16565372",
          4669 => x"7b27fb84",
          4670 => x"38a051f9",
          4671 => x"c63fef39",
          4672 => x"963d0d04",
          4673 => x"fd3d0d86",
          4674 => x"3d707084",
          4675 => x"05520855",
          4676 => x"527351fa",
          4677 => x"e03f853d",
          4678 => x"0d04fe3d",
          4679 => x"0d74829e",
          4680 => x"dc0c853d",
          4681 => x"88055275",
          4682 => x"51faca3f",
          4683 => x"829edc08",
          4684 => x"53807334",
          4685 => x"800b829e",
          4686 => x"dc0c843d",
          4687 => x"0d04fd3d",
          4688 => x"0d829ed4",
          4689 => x"0876829e",
          4690 => x"d40c873d",
          4691 => x"88055377",
          4692 => x"5253faa1",
          4693 => x"3f72829e",
          4694 => x"d40c853d",
          4695 => x"0d04fb3d",
          4696 => x"0d777982",
          4697 => x"9ed80870",
          4698 => x"56545755",
          4699 => x"80547180",
          4700 => x"2e80e038",
          4701 => x"829ed808",
          4702 => x"52712d82",
          4703 => x"87cc0881",
          4704 => x"ff065372",
          4705 => x"802e80cb",
          4706 => x"38728d2e",
          4707 => x"b9387288",
          4708 => x"32703070",
          4709 => x"80255151",
          4710 => x"5273802e",
          4711 => x"8b387180",
          4712 => x"2e8638ff",
          4713 => x"14549739",
          4714 => x"9f7325c8",
          4715 => x"38ff1652",
          4716 => x"737225c0",
          4717 => x"38741452",
          4718 => x"72723481",
          4719 => x"14547251",
          4720 => x"f8813fff",
          4721 => x"af397315",
          4722 => x"52807234",
          4723 => x"8a51f7f3",
          4724 => x"3f815372",
          4725 => x"8287cc0c",
          4726 => x"873d0d04",
          4727 => x"fe3d0d82",
          4728 => x"9ed80875",
          4729 => x"829ed80c",
          4730 => x"77537652",
          4731 => x"53feef3f",
          4732 => x"72829ed8",
          4733 => x"0c843d0d",
          4734 => x"04f83d0d",
          4735 => x"7a7c5a56",
          4736 => x"80707a0c",
          4737 => x"58750870",
          4738 => x"33555373",
          4739 => x"a02e0981",
          4740 => x"06873881",
          4741 => x"13760ced",
          4742 => x"3973ad2e",
          4743 => x"0981068e",
          4744 => x"38817608",
          4745 => x"11770c76",
          4746 => x"08703356",
          4747 => x"545873b0",
          4748 => x"2e098106",
          4749 => x"80c23875",
          4750 => x"08810576",
          4751 => x"0c750870",
          4752 => x"33555373",
          4753 => x"80e22e8b",
          4754 => x"38905773",
          4755 => x"80f82e85",
          4756 => x"388f3982",
          4757 => x"57811376",
          4758 => x"0c750870",
          4759 => x"335553ac",
          4760 => x"398155a0",
          4761 => x"742780fa",
          4762 => x"38d01453",
          4763 => x"80558857",
          4764 => x"89732798",
          4765 => x"3880eb39",
          4766 => x"d0145380",
          4767 => x"55728926",
          4768 => x"80e03886",
          4769 => x"39805580",
          4770 => x"d9398a57",
          4771 => x"8055a074",
          4772 => x"2780c238",
          4773 => x"80e07427",
          4774 => x"8938e014",
          4775 => x"7081ff06",
          4776 => x"5553d014",
          4777 => x"7081ff06",
          4778 => x"55539074",
          4779 => x"278e38f9",
          4780 => x"147081ff",
          4781 => x"06555389",
          4782 => x"7427ca38",
          4783 => x"737727c5",
          4784 => x"38747729",
          4785 => x"14760881",
          4786 => x"05770c76",
          4787 => x"08703356",
          4788 => x"5455ffba",
          4789 => x"3977802e",
          4790 => x"84387430",
          4791 => x"5574790c",
          4792 => x"81557482",
          4793 => x"87cc0c8a",
          4794 => x"3d0d04f8",
          4795 => x"3d0d7a7c",
          4796 => x"5a568070",
          4797 => x"7a0c5875",
          4798 => x"08703355",
          4799 => x"5373a02e",
          4800 => x"09810687",
          4801 => x"38811376",
          4802 => x"0ced3973",
          4803 => x"ad2e0981",
          4804 => x"068e3881",
          4805 => x"76081177",
          4806 => x"0c760870",
          4807 => x"33565458",
          4808 => x"73b02e09",
          4809 => x"810680c2",
          4810 => x"38750881",
          4811 => x"05760c75",
          4812 => x"08703355",
          4813 => x"537380e2",
          4814 => x"2e8b3890",
          4815 => x"577380f8",
          4816 => x"2e85388f",
          4817 => x"39825781",
          4818 => x"13760c75",
          4819 => x"08703355",
          4820 => x"53ac3981",
          4821 => x"55a07427",
          4822 => x"80fa38d0",
          4823 => x"14538055",
          4824 => x"88578973",
          4825 => x"27983880",
          4826 => x"eb39d014",
          4827 => x"53805572",
          4828 => x"892680e0",
          4829 => x"38863980",
          4830 => x"5580d939",
          4831 => x"8a578055",
          4832 => x"a0742780",
          4833 => x"c23880e0",
          4834 => x"74278938",
          4835 => x"e0147081",
          4836 => x"ff065553",
          4837 => x"d0147081",
          4838 => x"ff065553",
          4839 => x"9074278e",
          4840 => x"38f91470",
          4841 => x"81ff0655",
          4842 => x"53897427",
          4843 => x"ca387377",
          4844 => x"27c53874",
          4845 => x"77291476",
          4846 => x"08810577",
          4847 => x"0c760870",
          4848 => x"33565455",
          4849 => x"ffba3977",
          4850 => x"802e8438",
          4851 => x"74305574",
          4852 => x"790c8155",
          4853 => x"748287cc",
          4854 => x"0c8a3d0d",
          4855 => x"04fd3d0d",
          4856 => x"76982b70",
          4857 => x"982c7998",
          4858 => x"2b70982c",
          4859 => x"72101370",
          4860 => x"822b5153",
          4861 => x"51545151",
          4862 => x"800b81fc",
          4863 => x"d8123355",
          4864 => x"53717425",
          4865 => x"9c3881fc",
          4866 => x"d4110812",
          4867 => x"02840597",
          4868 => x"05337133",
          4869 => x"52525270",
          4870 => x"722e0981",
          4871 => x"06833881",
          4872 => x"53728287",
          4873 => x"cc0c853d",
          4874 => x"0d04fc3d",
          4875 => x"0d780284",
          4876 => x"059f0533",
          4877 => x"71335455",
          4878 => x"5371802e",
          4879 => x"9f388851",
          4880 => x"f3813fa0",
          4881 => x"51f2fc3f",
          4882 => x"8851f2f7",
          4883 => x"3f7233ff",
          4884 => x"05527173",
          4885 => x"347181ff",
          4886 => x"0652de39",
          4887 => x"7651f3c0",
          4888 => x"3f737334",
          4889 => x"863d0d04",
          4890 => x"f63d0d7c",
          4891 => x"028405b7",
          4892 => x"05330288",
          4893 => x"05bb0533",
          4894 => x"8287a433",
          4895 => x"70842982",
          4896 => x"86cc0570",
          4897 => x"08515959",
          4898 => x"5a585974",
          4899 => x"802e8638",
          4900 => x"74519e83",
          4901 => x"3f8287a4",
          4902 => x"33708429",
          4903 => x"8286cc05",
          4904 => x"81197054",
          4905 => x"58565aa1",
          4906 => x"843f8287",
          4907 => x"cc08750c",
          4908 => x"8287a433",
          4909 => x"70842982",
          4910 => x"86cc0570",
          4911 => x"0851565a",
          4912 => x"74802ea7",
          4913 => x"38755378",
          4914 => x"527451ff",
          4915 => x"bbc93f82",
          4916 => x"87a43381",
          4917 => x"05557482",
          4918 => x"87a43474",
          4919 => x"81ff0655",
          4920 => x"93752787",
          4921 => x"38800b82",
          4922 => x"87a43477",
          4923 => x"802eb638",
          4924 => x"8287a008",
          4925 => x"5675802e",
          4926 => x"ac388287",
          4927 => x"9c335574",
          4928 => x"a4388c3d",
          4929 => x"fc055476",
          4930 => x"53785275",
          4931 => x"5180d8e9",
          4932 => x"3f8287a0",
          4933 => x"08528a51",
          4934 => x"818df63f",
          4935 => x"8287a008",
          4936 => x"5180dcc6",
          4937 => x"3f8c3d0d",
          4938 => x"04fd3d0d",
          4939 => x"8286cc53",
          4940 => x"93547208",
          4941 => x"5271802e",
          4942 => x"89387151",
          4943 => x"9cd93f80",
          4944 => x"730cff14",
          4945 => x"84145454",
          4946 => x"738025e6",
          4947 => x"38800b82",
          4948 => x"87a43482",
          4949 => x"87a00852",
          4950 => x"71802e95",
          4951 => x"38715180",
          4952 => x"dda63f82",
          4953 => x"87a00851",
          4954 => x"9cad3f80",
          4955 => x"0b8287a0",
          4956 => x"0c853d0d",
          4957 => x"04dc3d0d",
          4958 => x"81578052",
          4959 => x"8287a008",
          4960 => x"5180e293",
          4961 => x"3f8287cc",
          4962 => x"0880d238",
          4963 => x"8287a008",
          4964 => x"5380f852",
          4965 => x"883d7052",
          4966 => x"56818ae1",
          4967 => x"3f8287cc",
          4968 => x"08802eb9",
          4969 => x"387551ff",
          4970 => x"b88d3f82",
          4971 => x"87cc0855",
          4972 => x"800b8287",
          4973 => x"cc08259c",
          4974 => x"388287cc",
          4975 => x"08ff0570",
          4976 => x"17555580",
          4977 => x"74347553",
          4978 => x"76528117",
          4979 => x"81ffc852",
          4980 => x"57f6b13f",
          4981 => x"74ff2e09",
          4982 => x"8106ffb0",
          4983 => x"38a63d0d",
          4984 => x"04d93d0d",
          4985 => x"aa3d08ad",
          4986 => x"3d085a5a",
          4987 => x"81705858",
          4988 => x"80528287",
          4989 => x"a0085180",
          4990 => x"e19d3f82",
          4991 => x"87cc0881",
          4992 => x"9438ff0b",
          4993 => x"8287a008",
          4994 => x"545580f8",
          4995 => x"528b3d70",
          4996 => x"52568189",
          4997 => x"e83f8287",
          4998 => x"cc08802e",
          4999 => x"a5387551",
          5000 => x"ffb7943f",
          5001 => x"8287cc08",
          5002 => x"81185855",
          5003 => x"800b8287",
          5004 => x"cc08258e",
          5005 => x"388287cc",
          5006 => x"08ff0570",
          5007 => x"17555580",
          5008 => x"74347409",
          5009 => x"70307072",
          5010 => x"079f2a51",
          5011 => x"55557877",
          5012 => x"2e853873",
          5013 => x"ffac3882",
          5014 => x"87a0088c",
          5015 => x"11085351",
          5016 => x"80e0b43f",
          5017 => x"8287cc08",
          5018 => x"802e8838",
          5019 => x"81ffd451",
          5020 => x"efae3f78",
          5021 => x"772e0981",
          5022 => x"069b3875",
          5023 => x"527951ff",
          5024 => x"b7a33f79",
          5025 => x"51ffb6af",
          5026 => x"3fab3d08",
          5027 => x"548287cc",
          5028 => x"08743480",
          5029 => x"58778287",
          5030 => x"cc0ca93d",
          5031 => x"0d04f63d",
          5032 => x"0d7c7e71",
          5033 => x"5c717233",
          5034 => x"57595a58",
          5035 => x"73a02e09",
          5036 => x"8106a238",
          5037 => x"78337805",
          5038 => x"56777627",
          5039 => x"98388117",
          5040 => x"705b7071",
          5041 => x"33565855",
          5042 => x"73a02e09",
          5043 => x"81068638",
          5044 => x"757526ea",
          5045 => x"38805473",
          5046 => x"88298287",
          5047 => x"a8057008",
          5048 => x"5255ffb5",
          5049 => x"d23f8287",
          5050 => x"cc085379",
          5051 => x"52740851",
          5052 => x"ffb8d13f",
          5053 => x"8287cc08",
          5054 => x"80c53884",
          5055 => x"15335574",
          5056 => x"812e8838",
          5057 => x"74822e88",
          5058 => x"38b539fc",
          5059 => x"e83fac39",
          5060 => x"811a5a8c",
          5061 => x"3dfc1153",
          5062 => x"f80551f5",
          5063 => x"dc3f8287",
          5064 => x"cc08802e",
          5065 => x"9a38ff1b",
          5066 => x"53785277",
          5067 => x"51fdb23f",
          5068 => x"8287cc08",
          5069 => x"81ff0655",
          5070 => x"74853874",
          5071 => x"54913981",
          5072 => x"147081ff",
          5073 => x"06515482",
          5074 => x"7427ff8b",
          5075 => x"38805473",
          5076 => x"8287cc0c",
          5077 => x"8c3d0d04",
          5078 => x"d33d0db0",
          5079 => x"3d08b23d",
          5080 => x"08b43d08",
          5081 => x"595f5a80",
          5082 => x"0baf3d34",
          5083 => x"8287a433",
          5084 => x"8287a008",
          5085 => x"555b7381",
          5086 => x"ca387382",
          5087 => x"879c3355",
          5088 => x"55738338",
          5089 => x"81557680",
          5090 => x"2e81bb38",
          5091 => x"81707606",
          5092 => x"55567380",
          5093 => x"2e81ac38",
          5094 => x"a8519b91",
          5095 => x"3f8287cc",
          5096 => x"088287a0",
          5097 => x"0c8287cc",
          5098 => x"08802e81",
          5099 => x"91389353",
          5100 => x"76528287",
          5101 => x"cc085180",
          5102 => x"cbdd3f82",
          5103 => x"87cc0880",
          5104 => x"2e8b3882",
          5105 => x"808051f2",
          5106 => x"bb3f80f7",
          5107 => x"398287cc",
          5108 => x"085b8287",
          5109 => x"a0085380",
          5110 => x"f852903d",
          5111 => x"70525481",
          5112 => x"869b3f82",
          5113 => x"87cc0856",
          5114 => x"8287cc08",
          5115 => x"742e0981",
          5116 => x"0680d038",
          5117 => x"8287cc08",
          5118 => x"51ffb3bb",
          5119 => x"3f8287cc",
          5120 => x"0855800b",
          5121 => x"8287cc08",
          5122 => x"25a93882",
          5123 => x"87cc08ff",
          5124 => x"05701755",
          5125 => x"55807434",
          5126 => x"80537481",
          5127 => x"ff065275",
          5128 => x"51f8c53f",
          5129 => x"811b7081",
          5130 => x"ff065c54",
          5131 => x"937b2783",
          5132 => x"38805b74",
          5133 => x"ff2e0981",
          5134 => x"06ff9738",
          5135 => x"86397582",
          5136 => x"879c3476",
          5137 => x"8c388287",
          5138 => x"a008802e",
          5139 => x"8438f9d9",
          5140 => x"3f8f3d5d",
          5141 => x"e0993f82",
          5142 => x"87cc0898",
          5143 => x"2b70982c",
          5144 => x"515978ff",
          5145 => x"2eee3878",
          5146 => x"81ff0682",
          5147 => x"9ee43370",
          5148 => x"982b7098",
          5149 => x"2c829ee0",
          5150 => x"3370982b",
          5151 => x"70972c71",
          5152 => x"982c0570",
          5153 => x"842981fc",
          5154 => x"d4057008",
          5155 => x"15703351",
          5156 => x"51515159",
          5157 => x"5951595d",
          5158 => x"58815673",
          5159 => x"782e80e9",
          5160 => x"38777427",
          5161 => x"b4387481",
          5162 => x"800a2981",
          5163 => x"ff0a0570",
          5164 => x"982c5155",
          5165 => x"80752480",
          5166 => x"ce387653",
          5167 => x"74527751",
          5168 => x"f69b3f82",
          5169 => x"87cc0881",
          5170 => x"ff065473",
          5171 => x"802ed738",
          5172 => x"74829ee0",
          5173 => x"348156b1",
          5174 => x"39748180",
          5175 => x"0a298180",
          5176 => x"0a057098",
          5177 => x"2c7081ff",
          5178 => x"06565155",
          5179 => x"73952697",
          5180 => x"38765374",
          5181 => x"527751f5",
          5182 => x"e43f8287",
          5183 => x"cc0881ff",
          5184 => x"065473cc",
          5185 => x"38d33980",
          5186 => x"5675802e",
          5187 => x"80ca3881",
          5188 => x"1c557482",
          5189 => x"9ee43474",
          5190 => x"982b7098",
          5191 => x"2c829ee0",
          5192 => x"3370982b",
          5193 => x"70982c70",
          5194 => x"10117082",
          5195 => x"2b81fcd8",
          5196 => x"11335e51",
          5197 => x"51515758",
          5198 => x"51557477",
          5199 => x"2e098106",
          5200 => x"fe923881",
          5201 => x"fcdc1408",
          5202 => x"7d0c800b",
          5203 => x"829ee434",
          5204 => x"800b829e",
          5205 => x"e0349239",
          5206 => x"75829ee4",
          5207 => x"3475829e",
          5208 => x"e03478af",
          5209 => x"3d34757d",
          5210 => x"0c7e5473",
          5211 => x"9526fde1",
          5212 => x"38738429",
          5213 => x"81e9a805",
          5214 => x"54730804",
          5215 => x"829eec33",
          5216 => x"54737e2e",
          5217 => x"fdcb3882",
          5218 => x"9ee83355",
          5219 => x"737527ab",
          5220 => x"3874982b",
          5221 => x"70982c51",
          5222 => x"55737524",
          5223 => x"9e38741a",
          5224 => x"54733381",
          5225 => x"15347481",
          5226 => x"800a2981",
          5227 => x"ff0a0570",
          5228 => x"982c829e",
          5229 => x"ec335651",
          5230 => x"55df3982",
          5231 => x"9eec3381",
          5232 => x"11565474",
          5233 => x"829eec34",
          5234 => x"731a54ae",
          5235 => x"3d337434",
          5236 => x"829ee833",
          5237 => x"54737e25",
          5238 => x"89388114",
          5239 => x"5473829e",
          5240 => x"e834829e",
          5241 => x"ec337081",
          5242 => x"800a2981",
          5243 => x"ff0a0570",
          5244 => x"982c829e",
          5245 => x"e8335a51",
          5246 => x"56567477",
          5247 => x"25a23874",
          5248 => x"1a703352",
          5249 => x"54e7bc3f",
          5250 => x"7481800a",
          5251 => x"2981800a",
          5252 => x"0570982c",
          5253 => x"829ee833",
          5254 => x"56515573",
          5255 => x"7524e038",
          5256 => x"829eec33",
          5257 => x"70982b70",
          5258 => x"982c829e",
          5259 => x"e8335a51",
          5260 => x"56567477",
          5261 => x"25fc9a38",
          5262 => x"8851e787",
          5263 => x"3f748180",
          5264 => x"0a298180",
          5265 => x"0a057098",
          5266 => x"2c829ee8",
          5267 => x"33565155",
          5268 => x"737524e4",
          5269 => x"38fbfa39",
          5270 => x"837a3480",
          5271 => x"0b811b34",
          5272 => x"829eec53",
          5273 => x"805281f5",
          5274 => x"b851f3be",
          5275 => x"3f81df39",
          5276 => x"829eec33",
          5277 => x"7081ff06",
          5278 => x"55557380",
          5279 => x"2efbd238",
          5280 => x"829ee833",
          5281 => x"ff055473",
          5282 => x"829ee834",
          5283 => x"ff155473",
          5284 => x"829eec34",
          5285 => x"8851e6ab",
          5286 => x"3f829eec",
          5287 => x"3370982b",
          5288 => x"70982c82",
          5289 => x"9ee83357",
          5290 => x"51565774",
          5291 => x"7425a738",
          5292 => x"741a5481",
          5293 => x"14337434",
          5294 => x"733351e6",
          5295 => x"863f7481",
          5296 => x"800a2981",
          5297 => x"800a0570",
          5298 => x"982c829e",
          5299 => x"e8335851",
          5300 => x"55757524",
          5301 => x"db38a051",
          5302 => x"e5e93f82",
          5303 => x"9eec3370",
          5304 => x"982b7098",
          5305 => x"2c829ee8",
          5306 => x"33575156",
          5307 => x"57747424",
          5308 => x"fadf3888",
          5309 => x"51e5cc3f",
          5310 => x"7481800a",
          5311 => x"2981800a",
          5312 => x"0570982c",
          5313 => x"829ee833",
          5314 => x"58515575",
          5315 => x"7525e438",
          5316 => x"fabf3982",
          5317 => x"9ee8337a",
          5318 => x"05548074",
          5319 => x"348a51e5",
          5320 => x"a23f829e",
          5321 => x"e8527951",
          5322 => x"f6f43f82",
          5323 => x"87cc0881",
          5324 => x"ff065473",
          5325 => x"9638829e",
          5326 => x"e8335473",
          5327 => x"802e8f38",
          5328 => x"81537352",
          5329 => x"7951f2a0",
          5330 => x"3f843980",
          5331 => x"7a34800b",
          5332 => x"829eec34",
          5333 => x"800b829e",
          5334 => x"e8347982",
          5335 => x"87cc0caf",
          5336 => x"3d0d0482",
          5337 => x"9eec3354",
          5338 => x"73802ef9",
          5339 => x"e4388851",
          5340 => x"e4d13f82",
          5341 => x"9eec33ff",
          5342 => x"05547382",
          5343 => x"9eec3473",
          5344 => x"81ff0654",
          5345 => x"e339829e",
          5346 => x"ec33829e",
          5347 => x"e8335555",
          5348 => x"73752ef9",
          5349 => x"bc38ff14",
          5350 => x"5473829e",
          5351 => x"e8347498",
          5352 => x"2b70982c",
          5353 => x"7581ff06",
          5354 => x"56515574",
          5355 => x"7425a738",
          5356 => x"741a5481",
          5357 => x"14337434",
          5358 => x"733351e4",
          5359 => x"863f7481",
          5360 => x"800a2981",
          5361 => x"800a0570",
          5362 => x"982c829e",
          5363 => x"e8335851",
          5364 => x"55757524",
          5365 => x"db38a051",
          5366 => x"e3e93f82",
          5367 => x"9eec3370",
          5368 => x"982b7098",
          5369 => x"2c829ee8",
          5370 => x"33575156",
          5371 => x"57747424",
          5372 => x"f8df3888",
          5373 => x"51e3cc3f",
          5374 => x"7481800a",
          5375 => x"2981800a",
          5376 => x"0570982c",
          5377 => x"829ee833",
          5378 => x"58515575",
          5379 => x"7525e438",
          5380 => x"f8bf3982",
          5381 => x"9eec3370",
          5382 => x"81ff0682",
          5383 => x"9ee83359",
          5384 => x"56547477",
          5385 => x"27f8aa38",
          5386 => x"81145473",
          5387 => x"829eec34",
          5388 => x"741a7033",
          5389 => x"5254e38b",
          5390 => x"3f829eec",
          5391 => x"337081ff",
          5392 => x"06829ee8",
          5393 => x"33585654",
          5394 => x"757526dc",
          5395 => x"38f88239",
          5396 => x"829eec53",
          5397 => x"805281f5",
          5398 => x"b851efce",
          5399 => x"3f800b82",
          5400 => x"9eec3480",
          5401 => x"0b829ee8",
          5402 => x"34f7e639",
          5403 => x"7ab03882",
          5404 => x"87980855",
          5405 => x"74802ea6",
          5406 => x"387451ff",
          5407 => x"aab93f82",
          5408 => x"87cc0882",
          5409 => x"9ee83482",
          5410 => x"87cc0881",
          5411 => x"ff068105",
          5412 => x"53745279",
          5413 => x"51ffabff",
          5414 => x"3f935b81",
          5415 => x"c0397a84",
          5416 => x"298286cc",
          5417 => x"05fc1108",
          5418 => x"56547480",
          5419 => x"2ea73874",
          5420 => x"51ffaa83",
          5421 => x"3f8287cc",
          5422 => x"08829ee8",
          5423 => x"348287cc",
          5424 => x"0881ff06",
          5425 => x"81055374",
          5426 => x"527951ff",
          5427 => x"abc93fff",
          5428 => x"1b5480fa",
          5429 => x"39730855",
          5430 => x"74802ef6",
          5431 => x"f4387451",
          5432 => x"ffa9d43f",
          5433 => x"99397a93",
          5434 => x"2e098106",
          5435 => x"ae388286",
          5436 => x"cc085574",
          5437 => x"802ea438",
          5438 => x"7451ffa9",
          5439 => x"ba3f8287",
          5440 => x"cc08829e",
          5441 => x"e8348287",
          5442 => x"cc0881ff",
          5443 => x"06810553",
          5444 => x"74527951",
          5445 => x"ffab803f",
          5446 => x"80c3397a",
          5447 => x"84298286",
          5448 => x"d0057008",
          5449 => x"56547480",
          5450 => x"2eab3874",
          5451 => x"51ffa987",
          5452 => x"3f8287cc",
          5453 => x"08829ee8",
          5454 => x"348287cc",
          5455 => x"0881ff06",
          5456 => x"81055374",
          5457 => x"527951ff",
          5458 => x"aacd3f81",
          5459 => x"1b547381",
          5460 => x"ff065b89",
          5461 => x"3974829e",
          5462 => x"e834747a",
          5463 => x"34829eec",
          5464 => x"53829ee8",
          5465 => x"33527951",
          5466 => x"edc03ff5",
          5467 => x"e439829e",
          5468 => x"ec337081",
          5469 => x"ff06829e",
          5470 => x"e8335956",
          5471 => x"54747727",
          5472 => x"f5cf3881",
          5473 => x"14547382",
          5474 => x"9eec3474",
          5475 => x"1a703352",
          5476 => x"54e0b03f",
          5477 => x"f5bb3982",
          5478 => x"9eec3354",
          5479 => x"73802ef5",
          5480 => x"b0388851",
          5481 => x"e09d3f82",
          5482 => x"9eec33ff",
          5483 => x"05547382",
          5484 => x"9eec34f5",
          5485 => x"9c39fb3d",
          5486 => x"0d779f2c",
          5487 => x"799f2c79",
          5488 => x"9f2c7a32",
          5489 => x"7073317c",
          5490 => x"9f2c7d32",
          5491 => x"74743271",
          5492 => x"75315855",
          5493 => x"59545557",
          5494 => x"54913f82",
          5495 => x"87cc0874",
          5496 => x"32743182",
          5497 => x"87cc0c87",
          5498 => x"3d0d04fa",
          5499 => x"3d0d787a",
          5500 => x"5855a052",
          5501 => x"76802e8b",
          5502 => x"38765180",
          5503 => x"f53f8287",
          5504 => x"cc0852e0",
          5505 => x"12537480",
          5506 => x"2e8d3874",
          5507 => x"5180e33f",
          5508 => x"718287cc",
          5509 => x"08315380",
          5510 => x"52729f26",
          5511 => x"80cb3874",
          5512 => x"52729f2e",
          5513 => x"80c33881",
          5514 => x"1375712a",
          5515 => x"a0723177",
          5516 => x"712b5854",
          5517 => x"55538056",
          5518 => x"72762ea8",
          5519 => x"38731075",
          5520 => x"9f2a0775",
          5521 => x"10770778",
          5522 => x"7231ff11",
          5523 => x"9f2c7081",
          5524 => x"067b7206",
          5525 => x"757131ff",
          5526 => x"1a5a5652",
          5527 => x"5a515456",
          5528 => x"5472da38",
          5529 => x"74107607",
          5530 => x"52718287",
          5531 => x"cc0c883d",
          5532 => x"0d04fd3d",
          5533 => x"0d7570fc",
          5534 => x"80800670",
          5535 => x"30707207",
          5536 => x"80257084",
          5537 => x"2b907131",
          5538 => x"75712a56",
          5539 => x"527483fe",
          5540 => x"80067030",
          5541 => x"70802583",
          5542 => x"2b887131",
          5543 => x"78712a59",
          5544 => x"52730577",
          5545 => x"81f00670",
          5546 => x"30708025",
          5547 => x"822b8471",
          5548 => x"317b712a",
          5549 => x"5c527305",
          5550 => x"7a8c0670",
          5551 => x"30708025",
          5552 => x"10827131",
          5553 => x"7e712a70",
          5554 => x"812a8132",
          5555 => x"70810670",
          5556 => x"30827431",
          5557 => x"06751905",
          5558 => x"8287cc0c",
          5559 => x"51525f52",
          5560 => x"41515253",
          5561 => x"51525351",
          5562 => x"52535153",
          5563 => x"5452853d",
          5564 => x"0d04fd3d",
          5565 => x"0d757770",
          5566 => x"54715354",
          5567 => x"54fdb73f",
          5568 => x"8287cc08",
          5569 => x"73297471",
          5570 => x"318287cc",
          5571 => x"0c53853d",
          5572 => x"0d04fa3d",
          5573 => x"0d787a57",
          5574 => x"55a05275",
          5575 => x"802e8b38",
          5576 => x"7551fece",
          5577 => x"3f8287cc",
          5578 => x"0852e012",
          5579 => x"5374802e",
          5580 => x"8d387451",
          5581 => x"febc3f71",
          5582 => x"8287cc08",
          5583 => x"31537452",
          5584 => x"729f2680",
          5585 => x"c8388052",
          5586 => x"729f2e80",
          5587 => x"c0388113",
          5588 => x"75712aa0",
          5589 => x"72317771",
          5590 => x"2b585455",
          5591 => x"53805772",
          5592 => x"772ea838",
          5593 => x"7310759f",
          5594 => x"2a077510",
          5595 => x"78077772",
          5596 => x"31ff119f",
          5597 => x"2c708106",
          5598 => x"7a720675",
          5599 => x"7131ff1a",
          5600 => x"5a56525b",
          5601 => x"51545654",
          5602 => x"72da3873",
          5603 => x"52718287",
          5604 => x"cc0c883d",
          5605 => x"0d04f93d",
          5606 => x"0d83c080",
          5607 => x"0b8287c4",
          5608 => x"0c84800b",
          5609 => x"8287c023",
          5610 => x"a0805380",
          5611 => x"5283c080",
          5612 => x"51ffa9b7",
          5613 => x"3f8287c4",
          5614 => x"08548058",
          5615 => x"77743481",
          5616 => x"57768115",
          5617 => x"348287c4",
          5618 => x"08547784",
          5619 => x"15347685",
          5620 => x"15348287",
          5621 => x"c4085477",
          5622 => x"86153476",
          5623 => x"87153482",
          5624 => x"87c40882",
          5625 => x"87c022ff",
          5626 => x"05fe8080",
          5627 => x"077083ff",
          5628 => x"ff067088",
          5629 => x"2a585155",
          5630 => x"56748817",
          5631 => x"34738917",
          5632 => x"348287c0",
          5633 => x"22708829",
          5634 => x"8287c408",
          5635 => x"05f81151",
          5636 => x"55557782",
          5637 => x"15347683",
          5638 => x"1534893d",
          5639 => x"0d04ff3d",
          5640 => x"0d735281",
          5641 => x"51847227",
          5642 => x"8f38fb12",
          5643 => x"832a8211",
          5644 => x"7083ffff",
          5645 => x"06515151",
          5646 => x"708287cc",
          5647 => x"0c833d0d",
          5648 => x"04f93d0d",
          5649 => x"02a60522",
          5650 => x"028405aa",
          5651 => x"05227105",
          5652 => x"8287c408",
          5653 => x"71832b71",
          5654 => x"1174832b",
          5655 => x"73117033",
          5656 => x"81123371",
          5657 => x"882b0702",
          5658 => x"a405ae05",
          5659 => x"227181ff",
          5660 => x"ff060770",
          5661 => x"882a5351",
          5662 => x"5259545b",
          5663 => x"5b575354",
          5664 => x"55717734",
          5665 => x"70811834",
          5666 => x"8287c408",
          5667 => x"1475882a",
          5668 => x"52547082",
          5669 => x"15347483",
          5670 => x"15348287",
          5671 => x"c4087017",
          5672 => x"70338112",
          5673 => x"3371882b",
          5674 => x"0770832b",
          5675 => x"8ffff806",
          5676 => x"51525652",
          5677 => x"71057383",
          5678 => x"ffff0670",
          5679 => x"882a5454",
          5680 => x"51718212",
          5681 => x"347281ff",
          5682 => x"06537283",
          5683 => x"12348287",
          5684 => x"c4081656",
          5685 => x"71763472",
          5686 => x"81173489",
          5687 => x"3d0d04fb",
          5688 => x"3d0d8287",
          5689 => x"c4080284",
          5690 => x"059e0522",
          5691 => x"70832b72",
          5692 => x"11861133",
          5693 => x"87123371",
          5694 => x"8b2b7183",
          5695 => x"2b07585b",
          5696 => x"59525552",
          5697 => x"72058412",
          5698 => x"33851333",
          5699 => x"71882b07",
          5700 => x"70882a54",
          5701 => x"56565270",
          5702 => x"84133473",
          5703 => x"85133482",
          5704 => x"87c40870",
          5705 => x"14841133",
          5706 => x"85123371",
          5707 => x"8b2b7183",
          5708 => x"2b075659",
          5709 => x"57527205",
          5710 => x"86123387",
          5711 => x"13337188",
          5712 => x"2b077088",
          5713 => x"2a545656",
          5714 => x"52708613",
          5715 => x"34738713",
          5716 => x"348287c4",
          5717 => x"08137033",
          5718 => x"81123371",
          5719 => x"882b0770",
          5720 => x"81ffff06",
          5721 => x"70882a53",
          5722 => x"51535353",
          5723 => x"71733470",
          5724 => x"81143487",
          5725 => x"3d0d04fa",
          5726 => x"3d0d02a2",
          5727 => x"05228287",
          5728 => x"c4087183",
          5729 => x"2b711170",
          5730 => x"33811233",
          5731 => x"71882b07",
          5732 => x"70882915",
          5733 => x"70338112",
          5734 => x"3371982b",
          5735 => x"71902b07",
          5736 => x"535f5355",
          5737 => x"525a5657",
          5738 => x"53547180",
          5739 => x"2580f638",
          5740 => x"7251feab",
          5741 => x"3f8287c4",
          5742 => x"08701670",
          5743 => x"33811233",
          5744 => x"718b2b71",
          5745 => x"832b0774",
          5746 => x"11703381",
          5747 => x"12337188",
          5748 => x"2b077083",
          5749 => x"2b8ffff8",
          5750 => x"06515254",
          5751 => x"51535a58",
          5752 => x"53720574",
          5753 => x"882a5452",
          5754 => x"72821334",
          5755 => x"73831334",
          5756 => x"8287c408",
          5757 => x"70167033",
          5758 => x"81123371",
          5759 => x"8b2b7183",
          5760 => x"2b075659",
          5761 => x"57557205",
          5762 => x"70338112",
          5763 => x"3371882b",
          5764 => x"077081ff",
          5765 => x"ff067088",
          5766 => x"2a575152",
          5767 => x"58527274",
          5768 => x"34718115",
          5769 => x"34883d0d",
          5770 => x"04fb3d0d",
          5771 => x"8287c408",
          5772 => x"0284059e",
          5773 => x"05227083",
          5774 => x"2b721182",
          5775 => x"11338312",
          5776 => x"33718b2b",
          5777 => x"71832b07",
          5778 => x"595b5952",
          5779 => x"56527305",
          5780 => x"71338113",
          5781 => x"3371882b",
          5782 => x"07028c05",
          5783 => x"a2052271",
          5784 => x"0770882a",
          5785 => x"53515353",
          5786 => x"53717334",
          5787 => x"70811434",
          5788 => x"8287c408",
          5789 => x"70157033",
          5790 => x"81123371",
          5791 => x"8b2b7183",
          5792 => x"2b075659",
          5793 => x"57527205",
          5794 => x"82123383",
          5795 => x"13337188",
          5796 => x"2b077088",
          5797 => x"2a545556",
          5798 => x"52708213",
          5799 => x"34728313",
          5800 => x"348287c4",
          5801 => x"08148211",
          5802 => x"33831233",
          5803 => x"71882b07",
          5804 => x"8287cc0c",
          5805 => x"5254873d",
          5806 => x"0d04f73d",
          5807 => x"0d7b8287",
          5808 => x"c4083183",
          5809 => x"2a7083ff",
          5810 => x"ff067053",
          5811 => x"5753fda7",
          5812 => x"3f8287c4",
          5813 => x"0876832b",
          5814 => x"71118211",
          5815 => x"33831233",
          5816 => x"718b2b71",
          5817 => x"832b0775",
          5818 => x"11703381",
          5819 => x"12337198",
          5820 => x"2b71902b",
          5821 => x"07534240",
          5822 => x"51535b58",
          5823 => x"55595472",
          5824 => x"80258d38",
          5825 => x"82808052",
          5826 => x"7551fe9d",
          5827 => x"3f818439",
          5828 => x"84143385",
          5829 => x"1533718b",
          5830 => x"2b71832b",
          5831 => x"07761179",
          5832 => x"882a5351",
          5833 => x"55585576",
          5834 => x"86143475",
          5835 => x"81ff0656",
          5836 => x"75871434",
          5837 => x"8287c408",
          5838 => x"70198412",
          5839 => x"33851333",
          5840 => x"71882b07",
          5841 => x"70882a54",
          5842 => x"575b5653",
          5843 => x"72841634",
          5844 => x"73851634",
          5845 => x"8287c408",
          5846 => x"1853800b",
          5847 => x"86143480",
          5848 => x"0b871434",
          5849 => x"8287c408",
          5850 => x"53768414",
          5851 => x"34758514",
          5852 => x"348287c4",
          5853 => x"08187033",
          5854 => x"81123371",
          5855 => x"882b0770",
          5856 => x"82808007",
          5857 => x"70882a53",
          5858 => x"51555654",
          5859 => x"74743472",
          5860 => x"8115348b",
          5861 => x"3d0d04ff",
          5862 => x"3d0d7352",
          5863 => x"8287c408",
          5864 => x"8438f7f2",
          5865 => x"3f71802e",
          5866 => x"86387151",
          5867 => x"fe8c3f83",
          5868 => x"3d0d04f5",
          5869 => x"3d0d807e",
          5870 => x"5258f8e2",
          5871 => x"3f8287cc",
          5872 => x"0883ffff",
          5873 => x"068287c4",
          5874 => x"08841133",
          5875 => x"85123371",
          5876 => x"882b0770",
          5877 => x"5f595658",
          5878 => x"5a81ffff",
          5879 => x"5975782e",
          5880 => x"80cb3875",
          5881 => x"88291770",
          5882 => x"33811233",
          5883 => x"71882b07",
          5884 => x"7081ffff",
          5885 => x"06793170",
          5886 => x"83ffff06",
          5887 => x"707f2752",
          5888 => x"53515659",
          5889 => x"55777927",
          5890 => x"8a387380",
          5891 => x"2e853875",
          5892 => x"785a5b84",
          5893 => x"15338516",
          5894 => x"3371882b",
          5895 => x"07575475",
          5896 => x"c2387881",
          5897 => x"ffff2e85",
          5898 => x"387a7959",
          5899 => x"56807683",
          5900 => x"2b8287c4",
          5901 => x"08117033",
          5902 => x"81123371",
          5903 => x"882b0770",
          5904 => x"81ffff06",
          5905 => x"51525a56",
          5906 => x"5c557375",
          5907 => x"2e833881",
          5908 => x"55805479",
          5909 => x"782681cc",
          5910 => x"38745474",
          5911 => x"802e81c4",
          5912 => x"38777a2e",
          5913 => x"09810689",
          5914 => x"387551f8",
          5915 => x"f23f81ac",
          5916 => x"39828080",
          5917 => x"53795275",
          5918 => x"51f7c63f",
          5919 => x"8287c408",
          5920 => x"701c8611",
          5921 => x"33871233",
          5922 => x"718b2b71",
          5923 => x"832b0753",
          5924 => x"5a5e5574",
          5925 => x"057a1770",
          5926 => x"83ffff06",
          5927 => x"70882a5c",
          5928 => x"59565478",
          5929 => x"84153476",
          5930 => x"81ff0657",
          5931 => x"76851534",
          5932 => x"8287c408",
          5933 => x"75832b71",
          5934 => x"11721e86",
          5935 => x"11338712",
          5936 => x"3371882b",
          5937 => x"0770882a",
          5938 => x"535b5e53",
          5939 => x"5a565473",
          5940 => x"86193475",
          5941 => x"87193482",
          5942 => x"87c40870",
          5943 => x"1c841133",
          5944 => x"85123371",
          5945 => x"8b2b7183",
          5946 => x"2b07535d",
          5947 => x"5a557405",
          5948 => x"54788615",
          5949 => x"34768715",
          5950 => x"348287c4",
          5951 => x"08701671",
          5952 => x"1d841133",
          5953 => x"85123371",
          5954 => x"882b0770",
          5955 => x"882a535a",
          5956 => x"5f525654",
          5957 => x"73841634",
          5958 => x"75851634",
          5959 => x"8287c408",
          5960 => x"1b840554",
          5961 => x"738287cc",
          5962 => x"0c8d3d0d",
          5963 => x"04fe3d0d",
          5964 => x"74528287",
          5965 => x"c4088438",
          5966 => x"f4dc3f71",
          5967 => x"5371802e",
          5968 => x"8b387151",
          5969 => x"fced3f82",
          5970 => x"87cc0853",
          5971 => x"728287cc",
          5972 => x"0c843d0d",
          5973 => x"04ff3d0d",
          5974 => x"028f0533",
          5975 => x"51815270",
          5976 => x"72268738",
          5977 => x"8287c811",
          5978 => x"33527182",
          5979 => x"87cc0c83",
          5980 => x"3d0d04fc",
          5981 => x"3d0d029b",
          5982 => x"05330284",
          5983 => x"059f0533",
          5984 => x"56538351",
          5985 => x"72812680",
          5986 => x"e0387284",
          5987 => x"2b87c092",
          5988 => x"8c115351",
          5989 => x"88547480",
          5990 => x"2e843881",
          5991 => x"88547372",
          5992 => x"0c87c092",
          5993 => x"8c115181",
          5994 => x"710c850b",
          5995 => x"87c0988c",
          5996 => x"0c705271",
          5997 => x"08708206",
          5998 => x"51517080",
          5999 => x"2e8a3887",
          6000 => x"c0988c08",
          6001 => x"5170ec38",
          6002 => x"7108fc80",
          6003 => x"80065271",
          6004 => x"923887c0",
          6005 => x"988c0851",
          6006 => x"70802e87",
          6007 => x"38718287",
          6008 => x"c8143482",
          6009 => x"87c81333",
          6010 => x"51708287",
          6011 => x"cc0c863d",
          6012 => x"0d04f33d",
          6013 => x"0d606264",
          6014 => x"028c05bf",
          6015 => x"05335740",
          6016 => x"585b8374",
          6017 => x"525afecd",
          6018 => x"3f8287cc",
          6019 => x"0881067a",
          6020 => x"54527181",
          6021 => x"be387172",
          6022 => x"75842b87",
          6023 => x"c0928011",
          6024 => x"87c0928c",
          6025 => x"1287c092",
          6026 => x"8413415a",
          6027 => x"40575a58",
          6028 => x"850b87c0",
          6029 => x"988c0c76",
          6030 => x"7d0c8476",
          6031 => x"0c750870",
          6032 => x"852a7081",
          6033 => x"06515354",
          6034 => x"71802e8e",
          6035 => x"387b0852",
          6036 => x"717b7081",
          6037 => x"055d3481",
          6038 => x"19598074",
          6039 => x"a2065353",
          6040 => x"71732e83",
          6041 => x"38815378",
          6042 => x"83ff268f",
          6043 => x"3872802e",
          6044 => x"8a3887c0",
          6045 => x"988c0852",
          6046 => x"71c33887",
          6047 => x"c0988c08",
          6048 => x"5271802e",
          6049 => x"87387884",
          6050 => x"802e9938",
          6051 => x"81760c87",
          6052 => x"c0928c15",
          6053 => x"53720870",
          6054 => x"82065152",
          6055 => x"71f738ff",
          6056 => x"1a5a8d39",
          6057 => x"84801781",
          6058 => x"197081ff",
          6059 => x"065a5357",
          6060 => x"79802e90",
          6061 => x"3873fc80",
          6062 => x"80065271",
          6063 => x"87387d78",
          6064 => x"26feed38",
          6065 => x"73fc8080",
          6066 => x"06527180",
          6067 => x"2e833881",
          6068 => x"52715372",
          6069 => x"8287cc0c",
          6070 => x"8f3d0d04",
          6071 => x"f33d0d60",
          6072 => x"6264028c",
          6073 => x"05bf0533",
          6074 => x"5740585b",
          6075 => x"83598074",
          6076 => x"5258fce1",
          6077 => x"3f8287cc",
          6078 => x"08810679",
          6079 => x"54527178",
          6080 => x"2e098106",
          6081 => x"81b13877",
          6082 => x"74842b87",
          6083 => x"c0928011",
          6084 => x"87c0928c",
          6085 => x"1287c092",
          6086 => x"84134059",
          6087 => x"5f565a85",
          6088 => x"0b87c098",
          6089 => x"8c0c767d",
          6090 => x"0c82760c",
          6091 => x"80587508",
          6092 => x"70842a70",
          6093 => x"81065153",
          6094 => x"5471802e",
          6095 => x"8c387a70",
          6096 => x"81055c33",
          6097 => x"7c0c8118",
          6098 => x"5873812a",
          6099 => x"70810651",
          6100 => x"5271802e",
          6101 => x"8a3887c0",
          6102 => x"988c0852",
          6103 => x"71d03887",
          6104 => x"c0988c08",
          6105 => x"5271802e",
          6106 => x"87387784",
          6107 => x"802e9938",
          6108 => x"81760c87",
          6109 => x"c0928c15",
          6110 => x"53720870",
          6111 => x"82065152",
          6112 => x"71f738ff",
          6113 => x"19598d39",
          6114 => x"811a7081",
          6115 => x"ff068480",
          6116 => x"19595b52",
          6117 => x"78802e90",
          6118 => x"3873fc80",
          6119 => x"80065271",
          6120 => x"87387d7a",
          6121 => x"26fef838",
          6122 => x"73fc8080",
          6123 => x"06527180",
          6124 => x"2e833881",
          6125 => x"52715372",
          6126 => x"8287cc0c",
          6127 => x"8f3d0d04",
          6128 => x"fa3d0d7a",
          6129 => x"028405a3",
          6130 => x"05330288",
          6131 => x"05a70533",
          6132 => x"71545456",
          6133 => x"57fafe3f",
          6134 => x"8287cc08",
          6135 => x"81065383",
          6136 => x"547280fe",
          6137 => x"38850b87",
          6138 => x"c0988c0c",
          6139 => x"81567176",
          6140 => x"2e80dc38",
          6141 => x"71762493",
          6142 => x"3874842b",
          6143 => x"87c0928c",
          6144 => x"11545471",
          6145 => x"802e8d38",
          6146 => x"80d43971",
          6147 => x"832e80c6",
          6148 => x"3880cb39",
          6149 => x"72087081",
          6150 => x"2a708106",
          6151 => x"51515271",
          6152 => x"802e8a38",
          6153 => x"87c0988c",
          6154 => x"085271e8",
          6155 => x"3887c098",
          6156 => x"8c085271",
          6157 => x"96388173",
          6158 => x"0c87c092",
          6159 => x"8c145372",
          6160 => x"08708206",
          6161 => x"515271f7",
          6162 => x"38963980",
          6163 => x"56923988",
          6164 => x"800a770c",
          6165 => x"85398180",
          6166 => x"770c7256",
          6167 => x"83398456",
          6168 => x"75547382",
          6169 => x"87cc0c88",
          6170 => x"3d0d04fe",
          6171 => x"3d0d7481",
          6172 => x"11337133",
          6173 => x"71882b07",
          6174 => x"8287cc0c",
          6175 => x"5351843d",
          6176 => x"0d04fd3d",
          6177 => x"0d758311",
          6178 => x"33821233",
          6179 => x"71902b71",
          6180 => x"882b0781",
          6181 => x"14337072",
          6182 => x"07882b75",
          6183 => x"33710782",
          6184 => x"87cc0c52",
          6185 => x"53545654",
          6186 => x"52853d0d",
          6187 => x"04ff3d0d",
          6188 => x"73028405",
          6189 => x"92052252",
          6190 => x"52707270",
          6191 => x"81055434",
          6192 => x"70882a51",
          6193 => x"70723483",
          6194 => x"3d0d04ff",
          6195 => x"3d0d7375",
          6196 => x"52527072",
          6197 => x"70810554",
          6198 => x"3470882a",
          6199 => x"51707270",
          6200 => x"81055434",
          6201 => x"70882a51",
          6202 => x"70727081",
          6203 => x"05543470",
          6204 => x"882a5170",
          6205 => x"7234833d",
          6206 => x"0d04fe3d",
          6207 => x"0d767577",
          6208 => x"54545170",
          6209 => x"802e9238",
          6210 => x"71708105",
          6211 => x"53337370",
          6212 => x"81055534",
          6213 => x"ff1151eb",
          6214 => x"39843d0d",
          6215 => x"04fe3d0d",
          6216 => x"75777654",
          6217 => x"52537272",
          6218 => x"70810554",
          6219 => x"34ff1151",
          6220 => x"70f43884",
          6221 => x"3d0d04fc",
          6222 => x"3d0d7877",
          6223 => x"79565653",
          6224 => x"74708105",
          6225 => x"56337470",
          6226 => x"81055633",
          6227 => x"717131ff",
          6228 => x"16565252",
          6229 => x"5272802e",
          6230 => x"86387180",
          6231 => x"2ee23871",
          6232 => x"8287cc0c",
          6233 => x"863d0d04",
          6234 => x"fe3d0d74",
          6235 => x"76545189",
          6236 => x"3971732e",
          6237 => x"8a388111",
          6238 => x"51703352",
          6239 => x"71f33870",
          6240 => x"338287cc",
          6241 => x"0c843d0d",
          6242 => x"04800b82",
          6243 => x"87cc0c04",
          6244 => x"800b8287",
          6245 => x"cc0c04f7",
          6246 => x"3d0d7b56",
          6247 => x"800b8317",
          6248 => x"33565a74",
          6249 => x"7a2e80d6",
          6250 => x"388154b0",
          6251 => x"160853b4",
          6252 => x"16705381",
          6253 => x"17335259",
          6254 => x"faa23f82",
          6255 => x"87cc087a",
          6256 => x"2e098106",
          6257 => x"b7388287",
          6258 => x"cc088317",
          6259 => x"34b01608",
          6260 => x"70a41808",
          6261 => x"319c1808",
          6262 => x"59565874",
          6263 => x"77279f38",
          6264 => x"82163355",
          6265 => x"74822e09",
          6266 => x"81069338",
          6267 => x"81547618",
          6268 => x"53785281",
          6269 => x"163351f9",
          6270 => x"e33f8339",
          6271 => x"815a7982",
          6272 => x"87cc0c8b",
          6273 => x"3d0d04fa",
          6274 => x"3d0d787a",
          6275 => x"56568057",
          6276 => x"74b01708",
          6277 => x"2eaf3875",
          6278 => x"51fefc3f",
          6279 => x"8287cc08",
          6280 => x"578287cc",
          6281 => x"089f3881",
          6282 => x"547453b4",
          6283 => x"16528116",
          6284 => x"3351f7be",
          6285 => x"3f8287cc",
          6286 => x"08802e85",
          6287 => x"38ff5581",
          6288 => x"5774b017",
          6289 => x"0c768287",
          6290 => x"cc0c883d",
          6291 => x"0d04f83d",
          6292 => x"0d7a7052",
          6293 => x"57fec03f",
          6294 => x"8287cc08",
          6295 => x"588287cc",
          6296 => x"08819138",
          6297 => x"76335574",
          6298 => x"832e0981",
          6299 => x"0680f038",
          6300 => x"84173359",
          6301 => x"78812e09",
          6302 => x"810680e3",
          6303 => x"38848053",
          6304 => x"8287cc08",
          6305 => x"52b41770",
          6306 => x"5256fd91",
          6307 => x"3f82d4d5",
          6308 => x"5284b217",
          6309 => x"51fc963f",
          6310 => x"848b85a4",
          6311 => x"d2527551",
          6312 => x"fca93f86",
          6313 => x"8a85e4f2",
          6314 => x"52849817",
          6315 => x"51fc9c3f",
          6316 => x"90170852",
          6317 => x"849c1751",
          6318 => x"fc913f8c",
          6319 => x"17085284",
          6320 => x"a01751fc",
          6321 => x"863fa017",
          6322 => x"08810570",
          6323 => x"b0190c79",
          6324 => x"55537552",
          6325 => x"81173351",
          6326 => x"f8823f77",
          6327 => x"84183480",
          6328 => x"53805281",
          6329 => x"173351f9",
          6330 => x"d73f8287",
          6331 => x"cc08802e",
          6332 => x"83388158",
          6333 => x"778287cc",
          6334 => x"0c8a3d0d",
          6335 => x"04fb3d0d",
          6336 => x"77fe1a98",
          6337 => x"1208fe05",
          6338 => x"55565480",
          6339 => x"56747327",
          6340 => x"8d388a14",
          6341 => x"22757129",
          6342 => x"ac160805",
          6343 => x"57537582",
          6344 => x"87cc0c87",
          6345 => x"3d0d04f9",
          6346 => x"3d0d7a7a",
          6347 => x"70085654",
          6348 => x"57817727",
          6349 => x"81df3876",
          6350 => x"98150827",
          6351 => x"81d738ff",
          6352 => x"74335458",
          6353 => x"72822e80",
          6354 => x"f5387282",
          6355 => x"24893872",
          6356 => x"812e8d38",
          6357 => x"81bf3972",
          6358 => x"832e818e",
          6359 => x"3881b639",
          6360 => x"76812a17",
          6361 => x"70892aa4",
          6362 => x"16080553",
          6363 => x"745255fd",
          6364 => x"963f8287",
          6365 => x"cc08819f",
          6366 => x"387483ff",
          6367 => x"0614b411",
          6368 => x"33811770",
          6369 => x"892aa418",
          6370 => x"08055576",
          6371 => x"54575753",
          6372 => x"fcf53f82",
          6373 => x"87cc0880",
          6374 => x"fe387483",
          6375 => x"ff0614b4",
          6376 => x"11337088",
          6377 => x"2b780779",
          6378 => x"81067184",
          6379 => x"2a5c5258",
          6380 => x"51537280",
          6381 => x"e238759f",
          6382 => x"ff065880",
          6383 => x"da397688",
          6384 => x"2aa41508",
          6385 => x"05527351",
          6386 => x"fcbd3f82",
          6387 => x"87cc0880",
          6388 => x"c6387610",
          6389 => x"83fe0674",
          6390 => x"05b40551",
          6391 => x"f98d3f82",
          6392 => x"87cc0883",
          6393 => x"ffff0658",
          6394 => x"ae397687",
          6395 => x"2aa41508",
          6396 => x"05527351",
          6397 => x"fc913f82",
          6398 => x"87cc089b",
          6399 => x"3876822b",
          6400 => x"83fc0674",
          6401 => x"05b40551",
          6402 => x"f8f83f82",
          6403 => x"87cc08f0",
          6404 => x"0a065883",
          6405 => x"39815877",
          6406 => x"8287cc0c",
          6407 => x"893d0d04",
          6408 => x"f83d0d7a",
          6409 => x"7c7e5a58",
          6410 => x"56825981",
          6411 => x"7727829e",
          6412 => x"38769817",
          6413 => x"08278296",
          6414 => x"38753353",
          6415 => x"72792e81",
          6416 => x"9d387279",
          6417 => x"24893872",
          6418 => x"812e8d38",
          6419 => x"82803972",
          6420 => x"832e81b8",
          6421 => x"3881f739",
          6422 => x"76812a17",
          6423 => x"70892aa4",
          6424 => x"18080553",
          6425 => x"765255fb",
          6426 => x"9e3f8287",
          6427 => x"cc085982",
          6428 => x"87cc0881",
          6429 => x"d9387483",
          6430 => x"ff0616b4",
          6431 => x"05811678",
          6432 => x"81065956",
          6433 => x"54775376",
          6434 => x"802e8f38",
          6435 => x"77842b9f",
          6436 => x"f0067433",
          6437 => x"8f067107",
          6438 => x"51537274",
          6439 => x"34810b83",
          6440 => x"17347489",
          6441 => x"2aa41708",
          6442 => x"05527551",
          6443 => x"fad93f82",
          6444 => x"87cc0859",
          6445 => x"8287cc08",
          6446 => x"81943874",
          6447 => x"83ff0616",
          6448 => x"b4057884",
          6449 => x"2a545476",
          6450 => x"8f387788",
          6451 => x"2a743381",
          6452 => x"f006718f",
          6453 => x"06075153",
          6454 => x"72743480",
          6455 => x"ec397688",
          6456 => x"2aa41708",
          6457 => x"05527551",
          6458 => x"fa9d3f82",
          6459 => x"87cc0859",
          6460 => x"8287cc08",
          6461 => x"80d83877",
          6462 => x"83ffff06",
          6463 => x"52761083",
          6464 => x"fe067605",
          6465 => x"b40551f7",
          6466 => x"a43fbe39",
          6467 => x"76872aa4",
          6468 => x"17080552",
          6469 => x"7551f9ef",
          6470 => x"3f8287cc",
          6471 => x"08598287",
          6472 => x"cc08ab38",
          6473 => x"77f00a06",
          6474 => x"77822b83",
          6475 => x"fc067018",
          6476 => x"b4057054",
          6477 => x"515454f6",
          6478 => x"c93f8287",
          6479 => x"cc088f0a",
          6480 => x"06740752",
          6481 => x"7251f783",
          6482 => x"3f810b83",
          6483 => x"17347882",
          6484 => x"87cc0c8a",
          6485 => x"3d0d04f8",
          6486 => x"3d0d7a7c",
          6487 => x"7e720859",
          6488 => x"56565981",
          6489 => x"7527a438",
          6490 => x"74981708",
          6491 => x"279d3873",
          6492 => x"802eaa38",
          6493 => x"ff537352",
          6494 => x"7551fda4",
          6495 => x"3f8287cc",
          6496 => x"08548287",
          6497 => x"cc0880f2",
          6498 => x"38933982",
          6499 => x"5480eb39",
          6500 => x"815480e6",
          6501 => x"398287cc",
          6502 => x"085480de",
          6503 => x"39745278",
          6504 => x"51fb843f",
          6505 => x"8287cc08",
          6506 => x"588287cc",
          6507 => x"08802e80",
          6508 => x"c7388287",
          6509 => x"cc08812e",
          6510 => x"d2388287",
          6511 => x"cc08ff2e",
          6512 => x"cf388053",
          6513 => x"74527551",
          6514 => x"fcd63f82",
          6515 => x"87cc08c5",
          6516 => x"38981608",
          6517 => x"fe119018",
          6518 => x"08575557",
          6519 => x"74742790",
          6520 => x"38811590",
          6521 => x"170c8416",
          6522 => x"33810754",
          6523 => x"73841734",
          6524 => x"77557678",
          6525 => x"26ffa638",
          6526 => x"80547382",
          6527 => x"87cc0c8a",
          6528 => x"3d0d04f6",
          6529 => x"3d0d7c7e",
          6530 => x"7108595b",
          6531 => x"5b799538",
          6532 => x"8c170858",
          6533 => x"77802e88",
          6534 => x"38981708",
          6535 => x"7826b238",
          6536 => x"8158ae39",
          6537 => x"79527a51",
          6538 => x"f9fd3f81",
          6539 => x"55748287",
          6540 => x"cc082782",
          6541 => x"e0388287",
          6542 => x"cc085582",
          6543 => x"87cc08ff",
          6544 => x"2e82d238",
          6545 => x"98170882",
          6546 => x"87cc0826",
          6547 => x"82c73879",
          6548 => x"58901708",
          6549 => x"70565473",
          6550 => x"802e82b9",
          6551 => x"38777a2e",
          6552 => x"09810680",
          6553 => x"e238811a",
          6554 => x"56981708",
          6555 => x"76268338",
          6556 => x"82567552",
          6557 => x"7a51f9af",
          6558 => x"3f805982",
          6559 => x"87cc0881",
          6560 => x"2e098106",
          6561 => x"86388287",
          6562 => x"cc085982",
          6563 => x"87cc0809",
          6564 => x"70307072",
          6565 => x"07802570",
          6566 => x"7c078287",
          6567 => x"cc085451",
          6568 => x"51555573",
          6569 => x"81ef3882",
          6570 => x"87cc0880",
          6571 => x"2e95388c",
          6572 => x"17085481",
          6573 => x"74279038",
          6574 => x"73981808",
          6575 => x"27893873",
          6576 => x"58853975",
          6577 => x"80db3877",
          6578 => x"56811656",
          6579 => x"98170876",
          6580 => x"26893882",
          6581 => x"56757826",
          6582 => x"81ac3875",
          6583 => x"527a51f8",
          6584 => x"c63f8287",
          6585 => x"cc08802e",
          6586 => x"b8388059",
          6587 => x"8287cc08",
          6588 => x"812e0981",
          6589 => x"06863882",
          6590 => x"87cc0859",
          6591 => x"8287cc08",
          6592 => x"09703070",
          6593 => x"72078025",
          6594 => x"707c0751",
          6595 => x"51555573",
          6596 => x"80f83875",
          6597 => x"782e0981",
          6598 => x"06ffae38",
          6599 => x"735580f5",
          6600 => x"39ff5375",
          6601 => x"527651f9",
          6602 => x"f73f8287",
          6603 => x"cc088287",
          6604 => x"cc083070",
          6605 => x"8287cc08",
          6606 => x"07802551",
          6607 => x"55557980",
          6608 => x"2e943873",
          6609 => x"802e8f38",
          6610 => x"75537952",
          6611 => x"7651f9d0",
          6612 => x"3f8287cc",
          6613 => x"085574a5",
          6614 => x"38758c18",
          6615 => x"0c981708",
          6616 => x"fe059018",
          6617 => x"08565474",
          6618 => x"74268638",
          6619 => x"ff159018",
          6620 => x"0c841733",
          6621 => x"81075473",
          6622 => x"84183497",
          6623 => x"39ff5674",
          6624 => x"812e9038",
          6625 => x"8c398055",
          6626 => x"8c398287",
          6627 => x"cc085585",
          6628 => x"39815675",
          6629 => x"55748287",
          6630 => x"cc0c8c3d",
          6631 => x"0d04f83d",
          6632 => x"0d7a7052",
          6633 => x"55f3f03f",
          6634 => x"8287cc08",
          6635 => x"58815682",
          6636 => x"87cc0880",
          6637 => x"d8387b52",
          6638 => x"7451f6c1",
          6639 => x"3f8287cc",
          6640 => x"088287cc",
          6641 => x"08b0170c",
          6642 => x"59848053",
          6643 => x"7752b415",
          6644 => x"705257f2",
          6645 => x"c83f7756",
          6646 => x"84398116",
          6647 => x"568a1522",
          6648 => x"58757827",
          6649 => x"97388154",
          6650 => x"75195376",
          6651 => x"52811533",
          6652 => x"51ede93f",
          6653 => x"8287cc08",
          6654 => x"802edf38",
          6655 => x"8a152276",
          6656 => x"32703070",
          6657 => x"7207709f",
          6658 => x"2a535156",
          6659 => x"56758287",
          6660 => x"cc0c8a3d",
          6661 => x"0d04f83d",
          6662 => x"0d7a7c71",
          6663 => x"08585657",
          6664 => x"74f0800a",
          6665 => x"2680f138",
          6666 => x"749f0653",
          6667 => x"7280e938",
          6668 => x"7490180c",
          6669 => x"88170854",
          6670 => x"73aa3875",
          6671 => x"33538273",
          6672 => x"278838a8",
          6673 => x"16085473",
          6674 => x"9b387485",
          6675 => x"2a53820b",
          6676 => x"8817225a",
          6677 => x"58727927",
          6678 => x"80fe38a8",
          6679 => x"16089818",
          6680 => x"0c80cd39",
          6681 => x"8a162270",
          6682 => x"892b5458",
          6683 => x"727526b2",
          6684 => x"38735276",
          6685 => x"51f5b03f",
          6686 => x"8287cc08",
          6687 => x"548287cc",
          6688 => x"08ff2ebd",
          6689 => x"38810b82",
          6690 => x"87cc0827",
          6691 => x"8b389816",
          6692 => x"088287cc",
          6693 => x"08268538",
          6694 => x"8258bd39",
          6695 => x"74733155",
          6696 => x"cb397352",
          6697 => x"7551f4d5",
          6698 => x"3f8287cc",
          6699 => x"0898180c",
          6700 => x"7394180c",
          6701 => x"98170853",
          6702 => x"82587280",
          6703 => x"2e9a3885",
          6704 => x"39815894",
          6705 => x"3974892a",
          6706 => x"1398180c",
          6707 => x"7483ff06",
          6708 => x"16b4059c",
          6709 => x"180c8058",
          6710 => x"778287cc",
          6711 => x"0c8a3d0d",
          6712 => x"04f83d0d",
          6713 => x"7a700890",
          6714 => x"1208a005",
          6715 => x"595754f0",
          6716 => x"800a7727",
          6717 => x"8638800b",
          6718 => x"98150c98",
          6719 => x"14085384",
          6720 => x"5572802e",
          6721 => x"81cb3876",
          6722 => x"83ff0658",
          6723 => x"7781b538",
          6724 => x"81139815",
          6725 => x"0c941408",
          6726 => x"55749238",
          6727 => x"76852a88",
          6728 => x"17225653",
          6729 => x"74732681",
          6730 => x"9b3880c0",
          6731 => x"398a1622",
          6732 => x"ff057789",
          6733 => x"2a065372",
          6734 => x"818a3874",
          6735 => x"527351f3",
          6736 => x"e63f8287",
          6737 => x"cc085382",
          6738 => x"55810b82",
          6739 => x"87cc0827",
          6740 => x"80ff3881",
          6741 => x"558287cc",
          6742 => x"08ff2e80",
          6743 => x"f4389816",
          6744 => x"088287cc",
          6745 => x"082680ca",
          6746 => x"387b8a38",
          6747 => x"7798150c",
          6748 => x"845580dd",
          6749 => x"39941408",
          6750 => x"527351f9",
          6751 => x"863f8287",
          6752 => x"cc085387",
          6753 => x"558287cc",
          6754 => x"08802e80",
          6755 => x"c4388255",
          6756 => x"8287cc08",
          6757 => x"812eba38",
          6758 => x"81558287",
          6759 => x"cc08ff2e",
          6760 => x"b0388287",
          6761 => x"cc085275",
          6762 => x"51fbf33f",
          6763 => x"8287cc08",
          6764 => x"a0387294",
          6765 => x"150c7252",
          6766 => x"7551f2c1",
          6767 => x"3f8287cc",
          6768 => x"0898150c",
          6769 => x"7690150c",
          6770 => x"7716b405",
          6771 => x"9c150c80",
          6772 => x"55748287",
          6773 => x"cc0c8a3d",
          6774 => x"0d04f73d",
          6775 => x"0d7b7d71",
          6776 => x"085b5b57",
          6777 => x"80527651",
          6778 => x"fcac3f82",
          6779 => x"87cc0854",
          6780 => x"8287cc08",
          6781 => x"80ec3882",
          6782 => x"87cc0856",
          6783 => x"98170852",
          6784 => x"7851f083",
          6785 => x"3f8287cc",
          6786 => x"08548287",
          6787 => x"cc0880d2",
          6788 => x"388287cc",
          6789 => x"089c1808",
          6790 => x"70335154",
          6791 => x"587281e5",
          6792 => x"2e098106",
          6793 => x"83388158",
          6794 => x"8287cc08",
          6795 => x"55728338",
          6796 => x"81557775",
          6797 => x"07537280",
          6798 => x"2e8e3881",
          6799 => x"1656757a",
          6800 => x"2e098106",
          6801 => x"8838a539",
          6802 => x"8287cc08",
          6803 => x"56815276",
          6804 => x"51fd8e3f",
          6805 => x"8287cc08",
          6806 => x"548287cc",
          6807 => x"08802eff",
          6808 => x"9b387384",
          6809 => x"2e098106",
          6810 => x"83388754",
          6811 => x"738287cc",
          6812 => x"0c8b3d0d",
          6813 => x"04fd3d0d",
          6814 => x"769a1152",
          6815 => x"54ebec3f",
          6816 => x"8287cc08",
          6817 => x"83ffff06",
          6818 => x"76703351",
          6819 => x"53537183",
          6820 => x"2e098106",
          6821 => x"90389414",
          6822 => x"51ebd03f",
          6823 => x"8287cc08",
          6824 => x"902b7307",
          6825 => x"53728287",
          6826 => x"cc0c853d",
          6827 => x"0d04fc3d",
          6828 => x"0d777970",
          6829 => x"83ffff06",
          6830 => x"549a1253",
          6831 => x"5555ebed",
          6832 => x"3f767033",
          6833 => x"51537283",
          6834 => x"2e098106",
          6835 => x"8b387390",
          6836 => x"2a529415",
          6837 => x"51ebd63f",
          6838 => x"863d0d04",
          6839 => x"f73d0d7b",
          6840 => x"7d5b5584",
          6841 => x"75085a58",
          6842 => x"98150880",
          6843 => x"2e818a38",
          6844 => x"98150852",
          6845 => x"7851ee8f",
          6846 => x"3f8287cc",
          6847 => x"08588287",
          6848 => x"cc0880f5",
          6849 => x"389c1508",
          6850 => x"70335553",
          6851 => x"73863884",
          6852 => x"5880e639",
          6853 => x"8b133370",
          6854 => x"bf067081",
          6855 => x"ff065851",
          6856 => x"53728616",
          6857 => x"348287cc",
          6858 => x"08537381",
          6859 => x"e52e8338",
          6860 => x"815373ae",
          6861 => x"2ea93881",
          6862 => x"70740654",
          6863 => x"5772802e",
          6864 => x"9e38758f",
          6865 => x"2e993882",
          6866 => x"87cc0876",
          6867 => x"df065454",
          6868 => x"72882e09",
          6869 => x"81068338",
          6870 => x"7654737a",
          6871 => x"2ea03880",
          6872 => x"527451fa",
          6873 => x"fc3f8287",
          6874 => x"cc085882",
          6875 => x"87cc0889",
          6876 => x"38981508",
          6877 => x"fefa3886",
          6878 => x"39800b98",
          6879 => x"160c7782",
          6880 => x"87cc0c8b",
          6881 => x"3d0d04fb",
          6882 => x"3d0d7770",
          6883 => x"08575481",
          6884 => x"527351fc",
          6885 => x"c53f8287",
          6886 => x"cc085582",
          6887 => x"87cc08b4",
          6888 => x"38981408",
          6889 => x"527551ec",
          6890 => x"de3f8287",
          6891 => x"cc085582",
          6892 => x"87cc08a0",
          6893 => x"38a05382",
          6894 => x"87cc0852",
          6895 => x"9c140851",
          6896 => x"eadb3f8b",
          6897 => x"53a01452",
          6898 => x"9c140851",
          6899 => x"eaac3f81",
          6900 => x"0b831734",
          6901 => x"748287cc",
          6902 => x"0c873d0d",
          6903 => x"04fd3d0d",
          6904 => x"75700898",
          6905 => x"12085470",
          6906 => x"535553ec",
          6907 => x"9a3f8287",
          6908 => x"cc088d38",
          6909 => x"9c130853",
          6910 => x"e5733481",
          6911 => x"0b831534",
          6912 => x"853d0d04",
          6913 => x"fa3d0d78",
          6914 => x"7a575780",
          6915 => x"0b891734",
          6916 => x"98170880",
          6917 => x"2e818238",
          6918 => x"80708918",
          6919 => x"5555559c",
          6920 => x"17081470",
          6921 => x"33811656",
          6922 => x"515271a0",
          6923 => x"2ea83871",
          6924 => x"852e0981",
          6925 => x"06843881",
          6926 => x"e5527389",
          6927 => x"2e098106",
          6928 => x"8b38ae73",
          6929 => x"70810555",
          6930 => x"34811555",
          6931 => x"71737081",
          6932 => x"05553481",
          6933 => x"15558a74",
          6934 => x"27c53875",
          6935 => x"15880552",
          6936 => x"800b8113",
          6937 => x"349c1708",
          6938 => x"528b1233",
          6939 => x"8817349c",
          6940 => x"17089c11",
          6941 => x"5252e88a",
          6942 => x"3f8287cc",
          6943 => x"08760c96",
          6944 => x"1251e7e7",
          6945 => x"3f8287cc",
          6946 => x"08861723",
          6947 => x"981251e7",
          6948 => x"da3f8287",
          6949 => x"cc088417",
          6950 => x"23883d0d",
          6951 => x"04f33d0d",
          6952 => x"7f70085e",
          6953 => x"5b806170",
          6954 => x"33515555",
          6955 => x"73af2e83",
          6956 => x"38815573",
          6957 => x"80dc2e91",
          6958 => x"3874802e",
          6959 => x"8c38941d",
          6960 => x"08881c0c",
          6961 => x"aa398115",
          6962 => x"41806170",
          6963 => x"33565656",
          6964 => x"73af2e09",
          6965 => x"81068338",
          6966 => x"81567380",
          6967 => x"dc327030",
          6968 => x"70802578",
          6969 => x"07515154",
          6970 => x"73dc3873",
          6971 => x"881c0c60",
          6972 => x"70335154",
          6973 => x"739f2696",
          6974 => x"38ff800b",
          6975 => x"ab1c3480",
          6976 => x"527a51f6",
          6977 => x"913f8287",
          6978 => x"cc085585",
          6979 => x"9839913d",
          6980 => x"61a01d5c",
          6981 => x"5a5e8b53",
          6982 => x"a0527951",
          6983 => x"e7ff3f80",
          6984 => x"70595788",
          6985 => x"7933555c",
          6986 => x"73ae2e09",
          6987 => x"810680d4",
          6988 => x"38781870",
          6989 => x"33811a71",
          6990 => x"ae327030",
          6991 => x"709f2a73",
          6992 => x"82260751",
          6993 => x"51535a57",
          6994 => x"54738c38",
          6995 => x"79175475",
          6996 => x"74348117",
          6997 => x"57db3975",
          6998 => x"af327030",
          6999 => x"709f2a51",
          7000 => x"51547580",
          7001 => x"dc2e8c38",
          7002 => x"73802e87",
          7003 => x"3875a026",
          7004 => x"82bd3877",
          7005 => x"197e0ca4",
          7006 => x"54a07627",
          7007 => x"82bd38a0",
          7008 => x"5482b839",
          7009 => x"78187033",
          7010 => x"811a5a57",
          7011 => x"54a07627",
          7012 => x"81fc3875",
          7013 => x"af327030",
          7014 => x"7780dc32",
          7015 => x"70307280",
          7016 => x"25718025",
          7017 => x"07515156",
          7018 => x"51557380",
          7019 => x"2eac3884",
          7020 => x"39811858",
          7021 => x"80781a70",
          7022 => x"33515555",
          7023 => x"73af2e09",
          7024 => x"81068338",
          7025 => x"81557380",
          7026 => x"dc327030",
          7027 => x"70802577",
          7028 => x"07515154",
          7029 => x"73db3881",
          7030 => x"b53975ae",
          7031 => x"2e098106",
          7032 => x"83388154",
          7033 => x"767c2774",
          7034 => x"07547380",
          7035 => x"2ea2387b",
          7036 => x"8b327030",
          7037 => x"77ae3270",
          7038 => x"30728025",
          7039 => x"719f2a07",
          7040 => x"53515651",
          7041 => x"557481a7",
          7042 => x"3888578b",
          7043 => x"5cfef539",
          7044 => x"75982b54",
          7045 => x"7380258c",
          7046 => x"387580ff",
          7047 => x"06828194",
          7048 => x"11335754",
          7049 => x"7551e6e1",
          7050 => x"3f8287cc",
          7051 => x"08802eb2",
          7052 => x"38781870",
          7053 => x"33811a71",
          7054 => x"545a5654",
          7055 => x"e6d23f82",
          7056 => x"87cc0880",
          7057 => x"2e80e838",
          7058 => x"ff1c5476",
          7059 => x"742780df",
          7060 => x"38791754",
          7061 => x"75743481",
          7062 => x"177a1155",
          7063 => x"57747434",
          7064 => x"a7397552",
          7065 => x"8280b451",
          7066 => x"e5fe3f82",
          7067 => x"87cc08bf",
          7068 => x"38ff9f16",
          7069 => x"54739926",
          7070 => x"8938e016",
          7071 => x"7081ff06",
          7072 => x"57547917",
          7073 => x"54757434",
          7074 => x"811757fd",
          7075 => x"f7397719",
          7076 => x"7e0c7680",
          7077 => x"2e993879",
          7078 => x"33547381",
          7079 => x"e52e0981",
          7080 => x"06843885",
          7081 => x"7a348454",
          7082 => x"a076278f",
          7083 => x"388b3986",
          7084 => x"5581f239",
          7085 => x"845680f3",
          7086 => x"39805473",
          7087 => x"8b1b3480",
          7088 => x"7b085852",
          7089 => x"7a51f2ce",
          7090 => x"3f8287cc",
          7091 => x"08568287",
          7092 => x"cc0880d7",
          7093 => x"38981b08",
          7094 => x"527651e6",
          7095 => x"aa3f8287",
          7096 => x"cc085682",
          7097 => x"87cc0880",
          7098 => x"c2389c1b",
          7099 => x"08703355",
          7100 => x"5573802e",
          7101 => x"ffbe388b",
          7102 => x"1533bf06",
          7103 => x"5473861c",
          7104 => x"348b1533",
          7105 => x"70832a70",
          7106 => x"81065155",
          7107 => x"58739238",
          7108 => x"8b537952",
          7109 => x"7451e49f",
          7110 => x"3f8287cc",
          7111 => x"08802e8b",
          7112 => x"3875527a",
          7113 => x"51f3ba3f",
          7114 => x"ff9f3975",
          7115 => x"ab1c3357",
          7116 => x"5574802e",
          7117 => x"bb387484",
          7118 => x"2e098106",
          7119 => x"80e73875",
          7120 => x"852a7081",
          7121 => x"0677822a",
          7122 => x"58515473",
          7123 => x"802e9638",
          7124 => x"75810654",
          7125 => x"73802efb",
          7126 => x"b538ff80",
          7127 => x"0bab1c34",
          7128 => x"805580c1",
          7129 => x"39758106",
          7130 => x"5473ba38",
          7131 => x"8555b639",
          7132 => x"75822a70",
          7133 => x"81065154",
          7134 => x"73ab3886",
          7135 => x"1b337084",
          7136 => x"2a708106",
          7137 => x"51555573",
          7138 => x"802ee138",
          7139 => x"901b0883",
          7140 => x"ff061db4",
          7141 => x"05527c51",
          7142 => x"f5db3f82",
          7143 => x"87cc0888",
          7144 => x"1c0cfaea",
          7145 => x"39748287",
          7146 => x"cc0c8f3d",
          7147 => x"0d04f63d",
          7148 => x"0d7c5bff",
          7149 => x"7b087071",
          7150 => x"7355595c",
          7151 => x"55597380",
          7152 => x"2e81c638",
          7153 => x"75708105",
          7154 => x"573370a0",
          7155 => x"26525271",
          7156 => x"ba2e8d38",
          7157 => x"70ee3871",
          7158 => x"ba2e0981",
          7159 => x"0681a538",
          7160 => x"7333d011",
          7161 => x"7081ff06",
          7162 => x"51525370",
          7163 => x"89269138",
          7164 => x"82147381",
          7165 => x"ff06d005",
          7166 => x"56527176",
          7167 => x"2e80f738",
          7168 => x"800b8281",
          7169 => x"84595577",
          7170 => x"087a5557",
          7171 => x"76708105",
          7172 => x"58337470",
          7173 => x"81055633",
          7174 => x"ff9f1253",
          7175 => x"53537099",
          7176 => x"268938e0",
          7177 => x"137081ff",
          7178 => x"065451ff",
          7179 => x"9f125170",
          7180 => x"99268938",
          7181 => x"e0127081",
          7182 => x"ff065351",
          7183 => x"7230709f",
          7184 => x"2a515172",
          7185 => x"722e0981",
          7186 => x"06853870",
          7187 => x"ffbe3872",
          7188 => x"30747732",
          7189 => x"70307072",
          7190 => x"079f2a73",
          7191 => x"9f2a0753",
          7192 => x"54545170",
          7193 => x"802e8f38",
          7194 => x"81158419",
          7195 => x"59558375",
          7196 => x"25ff9438",
          7197 => x"8b397483",
          7198 => x"24863874",
          7199 => x"767c0c59",
          7200 => x"78518639",
          7201 => x"829f8433",
          7202 => x"51708287",
          7203 => x"cc0c8c3d",
          7204 => x"0d04fa3d",
          7205 => x"0d785680",
          7206 => x"0b831734",
          7207 => x"ff0bb017",
          7208 => x"0c795275",
          7209 => x"51e2e03f",
          7210 => x"84558287",
          7211 => x"cc088180",
          7212 => x"3884b216",
          7213 => x"51dfb43f",
          7214 => x"8287cc08",
          7215 => x"83ffff06",
          7216 => x"54835573",
          7217 => x"82d4d52e",
          7218 => x"09810680",
          7219 => x"e338800b",
          7220 => x"b4173356",
          7221 => x"577481e9",
          7222 => x"2e098106",
          7223 => x"83388157",
          7224 => x"7481eb32",
          7225 => x"70307080",
          7226 => x"25790751",
          7227 => x"5154738a",
          7228 => x"387481e8",
          7229 => x"2e098106",
          7230 => x"b5388353",
          7231 => x"8280c452",
          7232 => x"80ea1651",
          7233 => x"e0b13f82",
          7234 => x"87cc0855",
          7235 => x"8287cc08",
          7236 => x"802e9d38",
          7237 => x"85538280",
          7238 => x"c8528186",
          7239 => x"1651e097",
          7240 => x"3f8287cc",
          7241 => x"08558287",
          7242 => x"cc08802e",
          7243 => x"83388255",
          7244 => x"748287cc",
          7245 => x"0c883d0d",
          7246 => x"04f23d0d",
          7247 => x"61028405",
          7248 => x"80cb0533",
          7249 => x"58558075",
          7250 => x"0c6051fc",
          7251 => x"e13f8287",
          7252 => x"cc08588b",
          7253 => x"56800b82",
          7254 => x"87cc0824",
          7255 => x"86fb3882",
          7256 => x"87cc0884",
          7257 => x"29829ef0",
          7258 => x"05700855",
          7259 => x"538c5673",
          7260 => x"802e86e5",
          7261 => x"3873750c",
          7262 => x"7681fe06",
          7263 => x"74335457",
          7264 => x"72802eae",
          7265 => x"38811433",
          7266 => x"51d7ca3f",
          7267 => x"8287cc08",
          7268 => x"81ff0670",
          7269 => x"81065455",
          7270 => x"72983876",
          7271 => x"802e86b7",
          7272 => x"3874822a",
          7273 => x"70810651",
          7274 => x"538a5672",
          7275 => x"86ab3886",
          7276 => x"a6398074",
          7277 => x"34778115",
          7278 => x"34815281",
          7279 => x"143351d7",
          7280 => x"b23f8287",
          7281 => x"cc0881ff",
          7282 => x"06708106",
          7283 => x"54558356",
          7284 => x"72868638",
          7285 => x"76802e8f",
          7286 => x"3874822a",
          7287 => x"70810651",
          7288 => x"538a5672",
          7289 => x"85f33880",
          7290 => x"70537452",
          7291 => x"5bfda33f",
          7292 => x"8287cc08",
          7293 => x"81ff0657",
          7294 => x"76822e09",
          7295 => x"810680e2",
          7296 => x"388c3d74",
          7297 => x"56588356",
          7298 => x"83f61533",
          7299 => x"70585372",
          7300 => x"802e8d38",
          7301 => x"83fa1551",
          7302 => x"dce83f82",
          7303 => x"87cc0857",
          7304 => x"76787084",
          7305 => x"055a0cff",
          7306 => x"16901656",
          7307 => x"56758025",
          7308 => x"d738800b",
          7309 => x"8d3d5456",
          7310 => x"72708405",
          7311 => x"54085b83",
          7312 => x"577a802e",
          7313 => x"95387a52",
          7314 => x"7351fcc6",
          7315 => x"3f8287cc",
          7316 => x"0881ff06",
          7317 => x"57817727",
          7318 => x"89388116",
          7319 => x"56837627",
          7320 => x"d7388156",
          7321 => x"76842e84",
          7322 => x"f0388d56",
          7323 => x"76812684",
          7324 => x"e838bf14",
          7325 => x"51dbf43f",
          7326 => x"8287cc08",
          7327 => x"83ffff06",
          7328 => x"53728480",
          7329 => x"2e098106",
          7330 => x"84cf3880",
          7331 => x"ca1451db",
          7332 => x"da3f8287",
          7333 => x"cc0883ff",
          7334 => x"ff065877",
          7335 => x"8d3880d8",
          7336 => x"1451dbde",
          7337 => x"3f8287cc",
          7338 => x"0858779c",
          7339 => x"150c80c4",
          7340 => x"14338215",
          7341 => x"3480c414",
          7342 => x"33ff1170",
          7343 => x"81ff0651",
          7344 => x"54558d56",
          7345 => x"72812684",
          7346 => x"90387481",
          7347 => x"ff067871",
          7348 => x"2980c116",
          7349 => x"33525953",
          7350 => x"728a1523",
          7351 => x"72802e8b",
          7352 => x"38ff1373",
          7353 => x"06537280",
          7354 => x"2e86388d",
          7355 => x"5683ea39",
          7356 => x"80c51451",
          7357 => x"daf53f82",
          7358 => x"87cc0853",
          7359 => x"8287cc08",
          7360 => x"88152372",
          7361 => x"8f06578d",
          7362 => x"567683cd",
          7363 => x"3880c714",
          7364 => x"51dad83f",
          7365 => x"8287cc08",
          7366 => x"83ffff06",
          7367 => x"55748d38",
          7368 => x"80d41451",
          7369 => x"dadc3f82",
          7370 => x"87cc0855",
          7371 => x"80c21451",
          7372 => x"dab93f82",
          7373 => x"87cc0883",
          7374 => x"ffff0653",
          7375 => x"8d567280",
          7376 => x"2e839638",
          7377 => x"88142278",
          7378 => x"1471842a",
          7379 => x"055a5a78",
          7380 => x"75268385",
          7381 => x"388a1422",
          7382 => x"52747931",
          7383 => x"51c58c3f",
          7384 => x"8287cc08",
          7385 => x"558287cc",
          7386 => x"08802e82",
          7387 => x"ec388287",
          7388 => x"cc0880ff",
          7389 => x"fffff526",
          7390 => x"83388357",
          7391 => x"7483fff5",
          7392 => x"26833882",
          7393 => x"57749ff5",
          7394 => x"26853881",
          7395 => x"5789398d",
          7396 => x"5676802e",
          7397 => x"82c33882",
          7398 => x"15709816",
          7399 => x"0c7ba016",
          7400 => x"0c731c70",
          7401 => x"a4170c7a",
          7402 => x"1dac170c",
          7403 => x"54557683",
          7404 => x"2e098106",
          7405 => x"af3880de",
          7406 => x"1451d9af",
          7407 => x"3f8287cc",
          7408 => x"0883ffff",
          7409 => x"06538d56",
          7410 => x"72828e38",
          7411 => x"79828a38",
          7412 => x"80e01451",
          7413 => x"d9ac3f82",
          7414 => x"87cc08a8",
          7415 => x"150c7482",
          7416 => x"2b53a239",
          7417 => x"8d567980",
          7418 => x"2e81ee38",
          7419 => x"7713a815",
          7420 => x"0c741553",
          7421 => x"76822e8d",
          7422 => x"38741015",
          7423 => x"70812a76",
          7424 => x"81060551",
          7425 => x"5383ff13",
          7426 => x"892a538d",
          7427 => x"56729c15",
          7428 => x"082681c5",
          7429 => x"38ff0b90",
          7430 => x"150cff0b",
          7431 => x"8c150cff",
          7432 => x"800b8415",
          7433 => x"3476832e",
          7434 => x"09810681",
          7435 => x"923880e4",
          7436 => x"1451d8b7",
          7437 => x"3f8287cc",
          7438 => x"0883ffff",
          7439 => x"06537281",
          7440 => x"2e098106",
          7441 => x"80f93881",
          7442 => x"1b527351",
          7443 => x"dbb93f82",
          7444 => x"87cc0880",
          7445 => x"ea388287",
          7446 => x"cc088415",
          7447 => x"3484b214",
          7448 => x"51d8883f",
          7449 => x"8287cc08",
          7450 => x"83ffff06",
          7451 => x"537282d4",
          7452 => x"d52e0981",
          7453 => x"0680c838",
          7454 => x"b41451d8",
          7455 => x"853f8287",
          7456 => x"cc08848b",
          7457 => x"85a4d22e",
          7458 => x"098106b3",
          7459 => x"38849814",
          7460 => x"51d7ef3f",
          7461 => x"8287cc08",
          7462 => x"868a85e4",
          7463 => x"f22e0981",
          7464 => x"069d3884",
          7465 => x"9c1451d7",
          7466 => x"d93f8287",
          7467 => x"cc089015",
          7468 => x"0c84a014",
          7469 => x"51d7cb3f",
          7470 => x"8287cc08",
          7471 => x"8c150c76",
          7472 => x"7434829f",
          7473 => x"80228105",
          7474 => x"5372829f",
          7475 => x"80237286",
          7476 => x"1523800b",
          7477 => x"94150c80",
          7478 => x"56758287",
          7479 => x"cc0c903d",
          7480 => x"0d04fb3d",
          7481 => x"0d775489",
          7482 => x"5573802e",
          7483 => x"b9387308",
          7484 => x"5372802e",
          7485 => x"b1387233",
          7486 => x"5271802e",
          7487 => x"a9388613",
          7488 => x"22841522",
          7489 => x"57527176",
          7490 => x"2e098106",
          7491 => x"99388113",
          7492 => x"3351d0c1",
          7493 => x"3f8287cc",
          7494 => x"08810652",
          7495 => x"71883871",
          7496 => x"74085455",
          7497 => x"83398053",
          7498 => x"7873710c",
          7499 => x"52748287",
          7500 => x"cc0c873d",
          7501 => x"0d04fa3d",
          7502 => x"0d02ab05",
          7503 => x"337a5889",
          7504 => x"3dfc0552",
          7505 => x"56f4e73f",
          7506 => x"8b54800b",
          7507 => x"8287cc08",
          7508 => x"24bc3882",
          7509 => x"87cc0884",
          7510 => x"29829ef0",
          7511 => x"05700855",
          7512 => x"5573802e",
          7513 => x"84388074",
          7514 => x"34785473",
          7515 => x"802e8438",
          7516 => x"80743478",
          7517 => x"750c7554",
          7518 => x"75802e92",
          7519 => x"38805389",
          7520 => x"3d705384",
          7521 => x"0551f7b1",
          7522 => x"3f8287cc",
          7523 => x"08547382",
          7524 => x"87cc0c88",
          7525 => x"3d0d04eb",
          7526 => x"3d0d6702",
          7527 => x"840580e7",
          7528 => x"05335959",
          7529 => x"89547880",
          7530 => x"2e84c838",
          7531 => x"77bf0670",
          7532 => x"54983dd0",
          7533 => x"0553993d",
          7534 => x"84055258",
          7535 => x"f6fb3f82",
          7536 => x"87cc0855",
          7537 => x"8287cc08",
          7538 => x"84a4387a",
          7539 => x"5c68528c",
          7540 => x"3d705256",
          7541 => x"edc73f82",
          7542 => x"87cc0855",
          7543 => x"8287cc08",
          7544 => x"92380280",
          7545 => x"d7053370",
          7546 => x"982b5557",
          7547 => x"73802583",
          7548 => x"38865577",
          7549 => x"9c065473",
          7550 => x"802e81ab",
          7551 => x"3874802e",
          7552 => x"95387484",
          7553 => x"2e098106",
          7554 => x"aa387551",
          7555 => x"eaf93f82",
          7556 => x"87cc0855",
          7557 => x"9e3902b2",
          7558 => x"05339106",
          7559 => x"547381b8",
          7560 => x"3877822a",
          7561 => x"70810651",
          7562 => x"5473802e",
          7563 => x"8e388855",
          7564 => x"83bc3977",
          7565 => x"88075874",
          7566 => x"83b43877",
          7567 => x"832a7081",
          7568 => x"06515473",
          7569 => x"802e81af",
          7570 => x"3862527a",
          7571 => x"51e8a63f",
          7572 => x"8287cc08",
          7573 => x"568288b2",
          7574 => x"0a52628e",
          7575 => x"0551d4eb",
          7576 => x"3f6254a0",
          7577 => x"0b8b1534",
          7578 => x"80536252",
          7579 => x"7a51e8be",
          7580 => x"3f805262",
          7581 => x"9c0551d4",
          7582 => x"d23f7a54",
          7583 => x"810b8315",
          7584 => x"3475802e",
          7585 => x"80f1387a",
          7586 => x"b0110851",
          7587 => x"54805375",
          7588 => x"52973dd4",
          7589 => x"0551ddbf",
          7590 => x"3f8287cc",
          7591 => x"08558287",
          7592 => x"cc0882ca",
          7593 => x"38b73974",
          7594 => x"82c43802",
          7595 => x"b2053370",
          7596 => x"842a7081",
          7597 => x"06515556",
          7598 => x"73802e86",
          7599 => x"38845582",
          7600 => x"ad397781",
          7601 => x"2a708106",
          7602 => x"51547380",
          7603 => x"2ea93875",
          7604 => x"81065473",
          7605 => x"802ea038",
          7606 => x"87558292",
          7607 => x"3973527a",
          7608 => x"51d6a43f",
          7609 => x"8287cc08",
          7610 => x"7bff188c",
          7611 => x"120c5555",
          7612 => x"8287cc08",
          7613 => x"81f83877",
          7614 => x"832a7081",
          7615 => x"06515473",
          7616 => x"802e8638",
          7617 => x"7780c007",
          7618 => x"587ab011",
          7619 => x"08a01b0c",
          7620 => x"63a41b0c",
          7621 => x"63537052",
          7622 => x"57e6da3f",
          7623 => x"8287cc08",
          7624 => x"8287cc08",
          7625 => x"881b0c63",
          7626 => x"9c05525a",
          7627 => x"d2d43f82",
          7628 => x"87cc0882",
          7629 => x"87cc088c",
          7630 => x"1b0c777a",
          7631 => x"0c568617",
          7632 => x"22841a23",
          7633 => x"77901a34",
          7634 => x"800b911a",
          7635 => x"34800b9c",
          7636 => x"1a0c800b",
          7637 => x"941a0c77",
          7638 => x"852a7081",
          7639 => x"06515473",
          7640 => x"802e818d",
          7641 => x"388287cc",
          7642 => x"08802e81",
          7643 => x"84388287",
          7644 => x"cc08941a",
          7645 => x"0c8a1722",
          7646 => x"70892b7b",
          7647 => x"525957a8",
          7648 => x"39765278",
          7649 => x"51d7a03f",
          7650 => x"8287cc08",
          7651 => x"578287cc",
          7652 => x"08812683",
          7653 => x"38825582",
          7654 => x"87cc08ff",
          7655 => x"2e098106",
          7656 => x"83387955",
          7657 => x"75783156",
          7658 => x"74307076",
          7659 => x"07802551",
          7660 => x"54777627",
          7661 => x"8a388170",
          7662 => x"7506555a",
          7663 => x"73c33876",
          7664 => x"981a0c74",
          7665 => x"a9387583",
          7666 => x"ff065473",
          7667 => x"802ea238",
          7668 => x"76527a51",
          7669 => x"d6a73f82",
          7670 => x"87cc0885",
          7671 => x"3882558e",
          7672 => x"3975892a",
          7673 => x"8287cc08",
          7674 => x"059c1a0c",
          7675 => x"84398079",
          7676 => x"0c745473",
          7677 => x"8287cc0c",
          7678 => x"973d0d04",
          7679 => x"f23d0d60",
          7680 => x"63656440",
          7681 => x"405d5980",
          7682 => x"7e0c903d",
          7683 => x"fc055278",
          7684 => x"51f9cf3f",
          7685 => x"8287cc08",
          7686 => x"558287cc",
          7687 => x"088a3891",
          7688 => x"19335574",
          7689 => x"802e8638",
          7690 => x"745682c4",
          7691 => x"39901933",
          7692 => x"81065587",
          7693 => x"5674802e",
          7694 => x"82b63895",
          7695 => x"39820b91",
          7696 => x"1a348256",
          7697 => x"82aa3981",
          7698 => x"0b911a34",
          7699 => x"815682a0",
          7700 => x"398c1908",
          7701 => x"941a0831",
          7702 => x"55747c27",
          7703 => x"8338745c",
          7704 => x"7b802e82",
          7705 => x"89389419",
          7706 => x"087083ff",
          7707 => x"06565674",
          7708 => x"81b2387e",
          7709 => x"8a1122ff",
          7710 => x"0577892a",
          7711 => x"065b5579",
          7712 => x"a8387587",
          7713 => x"38881908",
          7714 => x"558f3998",
          7715 => x"19085278",
          7716 => x"51d5943f",
          7717 => x"8287cc08",
          7718 => x"55817527",
          7719 => x"ff9f3874",
          7720 => x"ff2effa3",
          7721 => x"3874981a",
          7722 => x"0c981908",
          7723 => x"527e51d4",
          7724 => x"cc3f8287",
          7725 => x"cc08802e",
          7726 => x"ff833882",
          7727 => x"87cc081a",
          7728 => x"7c892a59",
          7729 => x"5777802e",
          7730 => x"80d63877",
          7731 => x"1a7f8a11",
          7732 => x"22585c55",
          7733 => x"75752785",
          7734 => x"38757a31",
          7735 => x"58775476",
          7736 => x"537c5281",
          7737 => x"1b3351ca",
          7738 => x"893f8287",
          7739 => x"cc08fed7",
          7740 => x"387e8311",
          7741 => x"33565674",
          7742 => x"802e9f38",
          7743 => x"b0160877",
          7744 => x"31557478",
          7745 => x"27943884",
          7746 => x"8053b416",
          7747 => x"52b01608",
          7748 => x"7731892b",
          7749 => x"7d0551cf",
          7750 => x"e13f7789",
          7751 => x"2b56b939",
          7752 => x"769c1a0c",
          7753 => x"94190883",
          7754 => x"ff068480",
          7755 => x"71315755",
          7756 => x"7b762783",
          7757 => x"387b569c",
          7758 => x"1908527e",
          7759 => x"51d1c83f",
          7760 => x"8287cc08",
          7761 => x"fe813875",
          7762 => x"53941908",
          7763 => x"83ff061f",
          7764 => x"b405527c",
          7765 => x"51cfa33f",
          7766 => x"7b76317e",
          7767 => x"08177f0c",
          7768 => x"761e941b",
          7769 => x"0818941c",
          7770 => x"0c5e5cfd",
          7771 => x"f3398056",
          7772 => x"758287cc",
          7773 => x"0c903d0d",
          7774 => x"04f23d0d",
          7775 => x"60636564",
          7776 => x"40405d58",
          7777 => x"807e0c90",
          7778 => x"3dfc0552",
          7779 => x"7751f6d2",
          7780 => x"3f8287cc",
          7781 => x"08558287",
          7782 => x"cc088a38",
          7783 => x"91183355",
          7784 => x"74802e86",
          7785 => x"38745683",
          7786 => x"b8399018",
          7787 => x"3370812a",
          7788 => x"70810651",
          7789 => x"56568756",
          7790 => x"74802e83",
          7791 => x"a4389539",
          7792 => x"820b9119",
          7793 => x"34825683",
          7794 => x"9839810b",
          7795 => x"91193481",
          7796 => x"56838e39",
          7797 => x"9418087c",
          7798 => x"11565674",
          7799 => x"76278438",
          7800 => x"75095c7b",
          7801 => x"802e82ec",
          7802 => x"38941808",
          7803 => x"7083ff06",
          7804 => x"56567481",
          7805 => x"fd387e8a",
          7806 => x"1122ff05",
          7807 => x"77892a06",
          7808 => x"5c557abf",
          7809 => x"38758c38",
          7810 => x"88180855",
          7811 => x"749c387a",
          7812 => x"52853998",
          7813 => x"18085277",
          7814 => x"51d7e83f",
          7815 => x"8287cc08",
          7816 => x"558287cc",
          7817 => x"08802e82",
          7818 => x"ab387481",
          7819 => x"2eff9138",
          7820 => x"74ff2eff",
          7821 => x"95387498",
          7822 => x"190c8818",
          7823 => x"08853874",
          7824 => x"88190c7e",
          7825 => x"55b01508",
          7826 => x"9c19082e",
          7827 => x"0981068d",
          7828 => x"387451ce",
          7829 => x"c23f8287",
          7830 => x"cc08feee",
          7831 => x"38981808",
          7832 => x"527e51d1",
          7833 => x"983f8287",
          7834 => x"cc08802e",
          7835 => x"fed23882",
          7836 => x"87cc081b",
          7837 => x"7c892a5a",
          7838 => x"5778802e",
          7839 => x"80d53878",
          7840 => x"1b7f8a11",
          7841 => x"22585b55",
          7842 => x"75752785",
          7843 => x"38757b31",
          7844 => x"59785476",
          7845 => x"537c5281",
          7846 => x"1a3351c8",
          7847 => x"bf3f8287",
          7848 => x"cc08fea6",
          7849 => x"387eb011",
          7850 => x"08783156",
          7851 => x"56747927",
          7852 => x"9b388480",
          7853 => x"53b01608",
          7854 => x"7731892b",
          7855 => x"7d0552b4",
          7856 => x"1651ccb6",
          7857 => x"3f7e5580",
          7858 => x"0b831634",
          7859 => x"78892b56",
          7860 => x"80db398c",
          7861 => x"18089419",
          7862 => x"08269338",
          7863 => x"7e51cdb7",
          7864 => x"3f8287cc",
          7865 => x"08fde338",
          7866 => x"7e77b012",
          7867 => x"0c55769c",
          7868 => x"190c9418",
          7869 => x"0883ff06",
          7870 => x"84807131",
          7871 => x"57557b76",
          7872 => x"2783387b",
          7873 => x"569c1808",
          7874 => x"527e51cd",
          7875 => x"fa3f8287",
          7876 => x"cc08fdb6",
          7877 => x"3875537c",
          7878 => x"52941808",
          7879 => x"83ff061f",
          7880 => x"b40551cb",
          7881 => x"d53f7e55",
          7882 => x"810b8316",
          7883 => x"347b7631",
          7884 => x"7e08177f",
          7885 => x"0c761e94",
          7886 => x"1a081870",
          7887 => x"941c0c8c",
          7888 => x"1b085858",
          7889 => x"5e5c7476",
          7890 => x"27833875",
          7891 => x"55748c19",
          7892 => x"0cfd9039",
          7893 => x"90183380",
          7894 => x"c0075574",
          7895 => x"90193480",
          7896 => x"56758287",
          7897 => x"cc0c903d",
          7898 => x"0d04f83d",
          7899 => x"0d7a8b3d",
          7900 => x"fc055370",
          7901 => x"5256f2ea",
          7902 => x"3f8287cc",
          7903 => x"08578287",
          7904 => x"cc0880fb",
          7905 => x"38901633",
          7906 => x"70862a70",
          7907 => x"81065155",
          7908 => x"5573802e",
          7909 => x"80e938a0",
          7910 => x"16085278",
          7911 => x"51cce83f",
          7912 => x"8287cc08",
          7913 => x"578287cc",
          7914 => x"0880d438",
          7915 => x"a416088b",
          7916 => x"1133a007",
          7917 => x"5555738b",
          7918 => x"16348816",
          7919 => x"08537452",
          7920 => x"750851dd",
          7921 => x"e93f8c16",
          7922 => x"08529c15",
          7923 => x"51c9fc3f",
          7924 => x"8288b20a",
          7925 => x"52961551",
          7926 => x"c9f13f76",
          7927 => x"52921551",
          7928 => x"c9cb3f78",
          7929 => x"54810b83",
          7930 => x"15347851",
          7931 => x"cce03f82",
          7932 => x"87cc0890",
          7933 => x"173381bf",
          7934 => x"06555773",
          7935 => x"90173476",
          7936 => x"8287cc0c",
          7937 => x"8a3d0d04",
          7938 => x"fc3d0d76",
          7939 => x"705254fe",
          7940 => x"d93f8287",
          7941 => x"cc085382",
          7942 => x"87cc089c",
          7943 => x"38863dfc",
          7944 => x"05527351",
          7945 => x"f1bc3f82",
          7946 => x"87cc0853",
          7947 => x"8287cc08",
          7948 => x"87388287",
          7949 => x"cc08740c",
          7950 => x"728287cc",
          7951 => x"0c863d0d",
          7952 => x"04ff3d0d",
          7953 => x"843d51e6",
          7954 => x"e53f8b52",
          7955 => x"800b8287",
          7956 => x"cc08248b",
          7957 => x"388287cc",
          7958 => x"08829f84",
          7959 => x"34805271",
          7960 => x"8287cc0c",
          7961 => x"833d0d04",
          7962 => x"ef3d0d80",
          7963 => x"53933dd0",
          7964 => x"0552943d",
          7965 => x"51e9c23f",
          7966 => x"8287cc08",
          7967 => x"558287cc",
          7968 => x"0880e038",
          7969 => x"76586352",
          7970 => x"933dd405",
          7971 => x"51e08e3f",
          7972 => x"8287cc08",
          7973 => x"558287cc",
          7974 => x"08bc3802",
          7975 => x"80c70533",
          7976 => x"70982b55",
          7977 => x"56738025",
          7978 => x"8938767a",
          7979 => x"94120c54",
          7980 => x"b23902a2",
          7981 => x"05337084",
          7982 => x"2a708106",
          7983 => x"51555673",
          7984 => x"802e9e38",
          7985 => x"767f5370",
          7986 => x"5254dba9",
          7987 => x"3f8287cc",
          7988 => x"0894150c",
          7989 => x"8e398287",
          7990 => x"cc08842e",
          7991 => x"09810683",
          7992 => x"38855574",
          7993 => x"8287cc0c",
          7994 => x"933d0d04",
          7995 => x"e43d0d6f",
          7996 => x"6f5b5b80",
          7997 => x"7a348053",
          7998 => x"9e3dffb8",
          7999 => x"05529f3d",
          8000 => x"51e8b63f",
          8001 => x"8287cc08",
          8002 => x"578287cc",
          8003 => x"0882fc38",
          8004 => x"7b437a7c",
          8005 => x"94110847",
          8006 => x"55586454",
          8007 => x"73802e81",
          8008 => x"ed38a052",
          8009 => x"933d7052",
          8010 => x"55d5eb3f",
          8011 => x"8287cc08",
          8012 => x"578287cc",
          8013 => x"0882d438",
          8014 => x"68527b51",
          8015 => x"c9c93f82",
          8016 => x"87cc0857",
          8017 => x"8287cc08",
          8018 => x"82c13869",
          8019 => x"527b51da",
          8020 => x"a43f8287",
          8021 => x"cc084576",
          8022 => x"527451d5",
          8023 => x"b93f8287",
          8024 => x"cc085782",
          8025 => x"87cc0882",
          8026 => x"a2388052",
          8027 => x"7451daec",
          8028 => x"3f8287cc",
          8029 => x"08578287",
          8030 => x"cc08a438",
          8031 => x"69527b51",
          8032 => x"d9f33f73",
          8033 => x"8287cc08",
          8034 => x"2ea63876",
          8035 => x"527451d6",
          8036 => x"d03f8287",
          8037 => x"cc085782",
          8038 => x"87cc0880",
          8039 => x"2ecc3876",
          8040 => x"842e0981",
          8041 => x"06863882",
          8042 => x"5781e039",
          8043 => x"7681dc38",
          8044 => x"9e3dffbc",
          8045 => x"05527451",
          8046 => x"dcca3f76",
          8047 => x"903d7811",
          8048 => x"81113351",
          8049 => x"565a5673",
          8050 => x"802e9138",
          8051 => x"02b90555",
          8052 => x"81168116",
          8053 => x"70335656",
          8054 => x"5673f538",
          8055 => x"81165473",
          8056 => x"78268190",
          8057 => x"3875802e",
          8058 => x"99387816",
          8059 => x"810555ff",
          8060 => x"186f11ff",
          8061 => x"18ff1858",
          8062 => x"58555874",
          8063 => x"33743475",
          8064 => x"ee38ff18",
          8065 => x"6f115558",
          8066 => x"af7434fe",
          8067 => x"8d39777b",
          8068 => x"2e098106",
          8069 => x"8a38ff18",
          8070 => x"6f115558",
          8071 => x"af743480",
          8072 => x"0b829f84",
          8073 => x"33708429",
          8074 => x"82818405",
          8075 => x"70087033",
          8076 => x"525c5656",
          8077 => x"5673762e",
          8078 => x"8d388116",
          8079 => x"701a7033",
          8080 => x"51555673",
          8081 => x"f5388216",
          8082 => x"54737826",
          8083 => x"a7388055",
          8084 => x"74762791",
          8085 => x"38741954",
          8086 => x"73337a70",
          8087 => x"81055c34",
          8088 => x"811555ec",
          8089 => x"39ba7a70",
          8090 => x"81055c34",
          8091 => x"74ff2e09",
          8092 => x"81068538",
          8093 => x"91579439",
          8094 => x"6e188119",
          8095 => x"59547333",
          8096 => x"7a708105",
          8097 => x"5c347a78",
          8098 => x"26ee3880",
          8099 => x"7a347682",
          8100 => x"87cc0c9e",
          8101 => x"3d0d04f7",
          8102 => x"3d0d7b7d",
          8103 => x"8d3dfc05",
          8104 => x"54715357",
          8105 => x"55ecbb3f",
          8106 => x"8287cc08",
          8107 => x"538287cc",
          8108 => x"0882fa38",
          8109 => x"91153353",
          8110 => x"7282f238",
          8111 => x"8c150854",
          8112 => x"73762792",
          8113 => x"38901533",
          8114 => x"70812a70",
          8115 => x"81065154",
          8116 => x"57728338",
          8117 => x"73569415",
          8118 => x"08548070",
          8119 => x"94170c58",
          8120 => x"75782e82",
          8121 => x"9738798a",
          8122 => x"11227089",
          8123 => x"2b595153",
          8124 => x"73782eb7",
          8125 => x"387652ff",
          8126 => x"1651ffad",
          8127 => x"ee3f8287",
          8128 => x"cc08ff15",
          8129 => x"78547053",
          8130 => x"5553ffad",
          8131 => x"de3f8287",
          8132 => x"cc087326",
          8133 => x"96387630",
          8134 => x"70750670",
          8135 => x"94180c77",
          8136 => x"71319818",
          8137 => x"08575851",
          8138 => x"53b13988",
          8139 => x"15085473",
          8140 => x"a6387352",
          8141 => x"7451cdcb",
          8142 => x"3f8287cc",
          8143 => x"08548287",
          8144 => x"cc08812e",
          8145 => x"819a3882",
          8146 => x"87cc08ff",
          8147 => x"2e819b38",
          8148 => x"8287cc08",
          8149 => x"88160c73",
          8150 => x"98160c73",
          8151 => x"802e819c",
          8152 => x"38767627",
          8153 => x"80dc3875",
          8154 => x"77319416",
          8155 => x"08189417",
          8156 => x"0c901633",
          8157 => x"70812a70",
          8158 => x"81065155",
          8159 => x"5a567280",
          8160 => x"2e9a3873",
          8161 => x"527451cc",
          8162 => x"fa3f8287",
          8163 => x"cc085482",
          8164 => x"87cc0894",
          8165 => x"388287cc",
          8166 => x"0856a739",
          8167 => x"73527451",
          8168 => x"c7853f82",
          8169 => x"87cc0854",
          8170 => x"73ff2ebe",
          8171 => x"38817427",
          8172 => x"af387953",
          8173 => x"73981408",
          8174 => x"27a63873",
          8175 => x"98160cff",
          8176 => x"a0399415",
          8177 => x"08169416",
          8178 => x"0c7583ff",
          8179 => x"06537280",
          8180 => x"2eaa3873",
          8181 => x"527951c6",
          8182 => x"a43f8287",
          8183 => x"cc089438",
          8184 => x"820b9116",
          8185 => x"34825380",
          8186 => x"c439810b",
          8187 => x"91163481",
          8188 => x"53bb3975",
          8189 => x"892a8287",
          8190 => x"cc080558",
          8191 => x"94150854",
          8192 => x"8c150874",
          8193 => x"27903873",
          8194 => x"8c160c90",
          8195 => x"153380c0",
          8196 => x"07537290",
          8197 => x"16347383",
          8198 => x"ff065372",
          8199 => x"802e8c38",
          8200 => x"779c1608",
          8201 => x"2e853877",
          8202 => x"9c160c80",
          8203 => x"53728287",
          8204 => x"cc0c8b3d",
          8205 => x"0d04f93d",
          8206 => x"0d795689",
          8207 => x"5475802e",
          8208 => x"818a3880",
          8209 => x"53893dfc",
          8210 => x"05528a3d",
          8211 => x"840551e1",
          8212 => x"e83f8287",
          8213 => x"cc085582",
          8214 => x"87cc0880",
          8215 => x"ea387776",
          8216 => x"0c7a5275",
          8217 => x"51d8b63f",
          8218 => x"8287cc08",
          8219 => x"558287cc",
          8220 => x"0880c338",
          8221 => x"ab163370",
          8222 => x"982b5557",
          8223 => x"807424a2",
          8224 => x"38861633",
          8225 => x"70842a70",
          8226 => x"81065155",
          8227 => x"5773802e",
          8228 => x"ad389c16",
          8229 => x"08527751",
          8230 => x"d3db3f82",
          8231 => x"87cc0888",
          8232 => x"170c7754",
          8233 => x"86142284",
          8234 => x"17237452",
          8235 => x"7551cee6",
          8236 => x"3f8287cc",
          8237 => x"08557484",
          8238 => x"2e098106",
          8239 => x"85388555",
          8240 => x"86397480",
          8241 => x"2e843880",
          8242 => x"760c7454",
          8243 => x"738287cc",
          8244 => x"0c893d0d",
          8245 => x"04fc3d0d",
          8246 => x"76873dfc",
          8247 => x"05537052",
          8248 => x"53e7ff3f",
          8249 => x"8287cc08",
          8250 => x"87388287",
          8251 => x"cc08730c",
          8252 => x"863d0d04",
          8253 => x"fb3d0d77",
          8254 => x"79893dfc",
          8255 => x"05547153",
          8256 => x"5654e7de",
          8257 => x"3f8287cc",
          8258 => x"08538287",
          8259 => x"cc0880df",
          8260 => x"38749338",
          8261 => x"8287cc08",
          8262 => x"527351cd",
          8263 => x"f93f8287",
          8264 => x"cc085380",
          8265 => x"ca398287",
          8266 => x"cc085273",
          8267 => x"51d3ad3f",
          8268 => x"8287cc08",
          8269 => x"538287cc",
          8270 => x"08842e09",
          8271 => x"81068538",
          8272 => x"80538739",
          8273 => x"8287cc08",
          8274 => x"a6387452",
          8275 => x"7351d5b4",
          8276 => x"3f725273",
          8277 => x"51cf8a3f",
          8278 => x"8287cc08",
          8279 => x"84327030",
          8280 => x"7072079f",
          8281 => x"2c708287",
          8282 => x"cc080651",
          8283 => x"51545472",
          8284 => x"8287cc0c",
          8285 => x"873d0d04",
          8286 => x"ee3d0d65",
          8287 => x"57805389",
          8288 => x"3d705396",
          8289 => x"3d5256df",
          8290 => x"b03f8287",
          8291 => x"cc085582",
          8292 => x"87cc08b2",
          8293 => x"38645275",
          8294 => x"51d6823f",
          8295 => x"8287cc08",
          8296 => x"558287cc",
          8297 => x"08a03802",
          8298 => x"80cb0533",
          8299 => x"70982b55",
          8300 => x"58738025",
          8301 => x"85388655",
          8302 => x"8d397680",
          8303 => x"2e883876",
          8304 => x"527551d4",
          8305 => x"bf3f7482",
          8306 => x"87cc0c94",
          8307 => x"3d0d04f0",
          8308 => x"3d0d6365",
          8309 => x"555c8053",
          8310 => x"923dec05",
          8311 => x"52933d51",
          8312 => x"ded73f82",
          8313 => x"87cc085b",
          8314 => x"8287cc08",
          8315 => x"8280387c",
          8316 => x"740c7308",
          8317 => x"981108fe",
          8318 => x"11901308",
          8319 => x"59565855",
          8320 => x"75742691",
          8321 => x"38757c0c",
          8322 => x"81e43981",
          8323 => x"5b81cc39",
          8324 => x"825b81c7",
          8325 => x"398287cc",
          8326 => x"08753355",
          8327 => x"5973812e",
          8328 => x"098106bf",
          8329 => x"3882755f",
          8330 => x"57765292",
          8331 => x"3df00551",
          8332 => x"c1f53f82",
          8333 => x"87cc08ff",
          8334 => x"2ed13882",
          8335 => x"87cc0881",
          8336 => x"2ece3882",
          8337 => x"87cc0830",
          8338 => x"708287cc",
          8339 => x"08078025",
          8340 => x"7a058119",
          8341 => x"7f53595a",
          8342 => x"54981408",
          8343 => x"7726ca38",
          8344 => x"80f939a4",
          8345 => x"15088287",
          8346 => x"cc085758",
          8347 => x"75983877",
          8348 => x"5281187d",
          8349 => x"5258ffbf",
          8350 => x"8e3f8287",
          8351 => x"cc085b82",
          8352 => x"87cc0880",
          8353 => x"d6387c70",
          8354 => x"337712ff",
          8355 => x"1a5d5256",
          8356 => x"5474822e",
          8357 => x"0981069e",
          8358 => x"38b41451",
          8359 => x"ffbbcc3f",
          8360 => x"8287cc08",
          8361 => x"83ffff06",
          8362 => x"70307080",
          8363 => x"251b8219",
          8364 => x"595b5154",
          8365 => x"9b39b414",
          8366 => x"51ffbbc6",
          8367 => x"3f8287cc",
          8368 => x"08f00a06",
          8369 => x"70307080",
          8370 => x"251b8419",
          8371 => x"595b5154",
          8372 => x"7583ff06",
          8373 => x"7a585679",
          8374 => x"ff923878",
          8375 => x"7c0c7c79",
          8376 => x"90120c84",
          8377 => x"11338107",
          8378 => x"56547484",
          8379 => x"15347a82",
          8380 => x"87cc0c92",
          8381 => x"3d0d04f9",
          8382 => x"3d0d798a",
          8383 => x"3dfc0553",
          8384 => x"705257e3",
          8385 => x"dd3f8287",
          8386 => x"cc085682",
          8387 => x"87cc0881",
          8388 => x"a8389117",
          8389 => x"33567581",
          8390 => x"a0389017",
          8391 => x"3370812a",
          8392 => x"70810651",
          8393 => x"55558755",
          8394 => x"73802e81",
          8395 => x"8e389417",
          8396 => x"0854738c",
          8397 => x"18082781",
          8398 => x"8038739b",
          8399 => x"388287cc",
          8400 => x"08538817",
          8401 => x"08527651",
          8402 => x"c48d3f82",
          8403 => x"87cc0874",
          8404 => x"88190c56",
          8405 => x"80c93998",
          8406 => x"17085276",
          8407 => x"51ffbfc7",
          8408 => x"3f8287cc",
          8409 => x"08ff2e09",
          8410 => x"81068338",
          8411 => x"81568287",
          8412 => x"cc08812e",
          8413 => x"09810685",
          8414 => x"388256a3",
          8415 => x"3975a038",
          8416 => x"77548287",
          8417 => x"cc089815",
          8418 => x"08279438",
          8419 => x"98170853",
          8420 => x"8287cc08",
          8421 => x"527651c3",
          8422 => x"be3f8287",
          8423 => x"cc085694",
          8424 => x"17088c18",
          8425 => x"0c901733",
          8426 => x"80c00754",
          8427 => x"73901834",
          8428 => x"75802e85",
          8429 => x"38759118",
          8430 => x"34755574",
          8431 => x"8287cc0c",
          8432 => x"893d0d04",
          8433 => x"e23d0d82",
          8434 => x"53a03dff",
          8435 => x"a40552a1",
          8436 => x"3d51dae5",
          8437 => x"3f8287cc",
          8438 => x"08558287",
          8439 => x"cc0881f5",
          8440 => x"387845a1",
          8441 => x"3d085295",
          8442 => x"3d705258",
          8443 => x"d1af3f82",
          8444 => x"87cc0855",
          8445 => x"8287cc08",
          8446 => x"81db3802",
          8447 => x"80fb0533",
          8448 => x"70852a70",
          8449 => x"81065155",
          8450 => x"56865573",
          8451 => x"81c73875",
          8452 => x"982b5480",
          8453 => x"742481bd",
          8454 => x"380280d6",
          8455 => x"05337081",
          8456 => x"06585487",
          8457 => x"557681ad",
          8458 => x"386b5278",
          8459 => x"51ccc63f",
          8460 => x"8287cc08",
          8461 => x"74842a70",
          8462 => x"81065155",
          8463 => x"5673802e",
          8464 => x"80d43878",
          8465 => x"548287cc",
          8466 => x"08941508",
          8467 => x"2e818638",
          8468 => x"735a8287",
          8469 => x"cc085c76",
          8470 => x"528a3d70",
          8471 => x"5254c7b6",
          8472 => x"3f8287cc",
          8473 => x"08558287",
          8474 => x"cc0880e9",
          8475 => x"388287cc",
          8476 => x"08527351",
          8477 => x"cce63f82",
          8478 => x"87cc0855",
          8479 => x"8287cc08",
          8480 => x"86388755",
          8481 => x"80cf3982",
          8482 => x"87cc0884",
          8483 => x"2e883882",
          8484 => x"87cc0880",
          8485 => x"c0387751",
          8486 => x"cec33f82",
          8487 => x"87cc0882",
          8488 => x"87cc0830",
          8489 => x"708287cc",
          8490 => x"08078025",
          8491 => x"51555575",
          8492 => x"802e9438",
          8493 => x"73802e8f",
          8494 => x"38805375",
          8495 => x"527751c1",
          8496 => x"963f8287",
          8497 => x"cc085574",
          8498 => x"8c387851",
          8499 => x"ffbaff3f",
          8500 => x"8287cc08",
          8501 => x"55748287",
          8502 => x"cc0ca03d",
          8503 => x"0d04e93d",
          8504 => x"0d825399",
          8505 => x"3dc00552",
          8506 => x"9a3d51d8",
          8507 => x"cc3f8287",
          8508 => x"cc085482",
          8509 => x"87cc0882",
          8510 => x"b038785e",
          8511 => x"69528e3d",
          8512 => x"705258cf",
          8513 => x"983f8287",
          8514 => x"cc085482",
          8515 => x"87cc0886",
          8516 => x"38885482",
          8517 => x"94398287",
          8518 => x"cc08842e",
          8519 => x"09810682",
          8520 => x"88380280",
          8521 => x"df053370",
          8522 => x"852a8106",
          8523 => x"51558654",
          8524 => x"7481f638",
          8525 => x"785a7452",
          8526 => x"8a3d7052",
          8527 => x"57c1c43f",
          8528 => x"8287cc08",
          8529 => x"75555682",
          8530 => x"87cc0883",
          8531 => x"38875482",
          8532 => x"87cc0881",
          8533 => x"2e098106",
          8534 => x"83388254",
          8535 => x"8287cc08",
          8536 => x"ff2e0981",
          8537 => x"06863881",
          8538 => x"5481b439",
          8539 => x"7381b038",
          8540 => x"8287cc08",
          8541 => x"527851c4",
          8542 => x"a53f8287",
          8543 => x"cc085482",
          8544 => x"87cc0881",
          8545 => x"9a388b53",
          8546 => x"a052b419",
          8547 => x"51ffb78d",
          8548 => x"3f7854ae",
          8549 => x"0bb41534",
          8550 => x"7854900b",
          8551 => x"bf153482",
          8552 => x"88b20a52",
          8553 => x"80ca1951",
          8554 => x"ffb6a03f",
          8555 => x"755378b4",
          8556 => x"115351c9",
          8557 => x"f93fa053",
          8558 => x"78b41153",
          8559 => x"80d40551",
          8560 => x"ffb6b73f",
          8561 => x"7854ae0b",
          8562 => x"80d51534",
          8563 => x"7f537880",
          8564 => x"d4115351",
          8565 => x"c9d83f78",
          8566 => x"54810b83",
          8567 => x"15347751",
          8568 => x"cba53f82",
          8569 => x"87cc0854",
          8570 => x"8287cc08",
          8571 => x"b2388288",
          8572 => x"b20a5264",
          8573 => x"960551ff",
          8574 => x"b5d13f75",
          8575 => x"53645278",
          8576 => x"51c9ab3f",
          8577 => x"6454900b",
          8578 => x"8b153478",
          8579 => x"54810b83",
          8580 => x"15347851",
          8581 => x"ffb8b73f",
          8582 => x"8287cc08",
          8583 => x"548b3980",
          8584 => x"53755276",
          8585 => x"51ffbeaf",
          8586 => x"3f738287",
          8587 => x"cc0c993d",
          8588 => x"0d04da3d",
          8589 => x"0da93d84",
          8590 => x"0551d2f2",
          8591 => x"3f8253a8",
          8592 => x"3dff8405",
          8593 => x"52a93d51",
          8594 => x"d5ef3f82",
          8595 => x"87cc0855",
          8596 => x"8287cc08",
          8597 => x"82d33878",
          8598 => x"4da93d08",
          8599 => x"529d3d70",
          8600 => x"5258ccb9",
          8601 => x"3f8287cc",
          8602 => x"08558287",
          8603 => x"cc0882b9",
          8604 => x"3802819b",
          8605 => x"053381a0",
          8606 => x"06548655",
          8607 => x"7382aa38",
          8608 => x"a053a43d",
          8609 => x"0852a83d",
          8610 => x"ff880551",
          8611 => x"ffb4eb3f",
          8612 => x"ac537752",
          8613 => x"923d7052",
          8614 => x"54ffb4de",
          8615 => x"3faa3d08",
          8616 => x"527351cb",
          8617 => x"f83f8287",
          8618 => x"cc085582",
          8619 => x"87cc0895",
          8620 => x"38636f2e",
          8621 => x"09810688",
          8622 => x"3865a23d",
          8623 => x"082e9238",
          8624 => x"885581e5",
          8625 => x"398287cc",
          8626 => x"08842e09",
          8627 => x"810681b8",
          8628 => x"387351c9",
          8629 => x"b23f8287",
          8630 => x"cc085582",
          8631 => x"87cc0881",
          8632 => x"c8386856",
          8633 => x"9353a83d",
          8634 => x"ff950552",
          8635 => x"8d1651ff",
          8636 => x"b4883f02",
          8637 => x"af05338b",
          8638 => x"17348b16",
          8639 => x"3370842a",
          8640 => x"70810651",
          8641 => x"55557389",
          8642 => x"3874a007",
          8643 => x"54738b17",
          8644 => x"34785481",
          8645 => x"0b831534",
          8646 => x"8b163370",
          8647 => x"842a7081",
          8648 => x"06515555",
          8649 => x"73802e80",
          8650 => x"e5386e64",
          8651 => x"2e80df38",
          8652 => x"75527851",
          8653 => x"c6bf3f82",
          8654 => x"87cc0852",
          8655 => x"7851ffb7",
          8656 => x"bc3f8255",
          8657 => x"8287cc08",
          8658 => x"802e80dd",
          8659 => x"388287cc",
          8660 => x"08527851",
          8661 => x"ffb5b03f",
          8662 => x"8287cc08",
          8663 => x"7980d411",
          8664 => x"58585582",
          8665 => x"87cc0880",
          8666 => x"c0388116",
          8667 => x"335473ae",
          8668 => x"2e098106",
          8669 => x"99386353",
          8670 => x"75527651",
          8671 => x"c6b03f78",
          8672 => x"54810b83",
          8673 => x"15348739",
          8674 => x"8287cc08",
          8675 => x"9c387751",
          8676 => x"c8cb3f82",
          8677 => x"87cc0855",
          8678 => x"8287cc08",
          8679 => x"8c387851",
          8680 => x"ffb5ab3f",
          8681 => x"8287cc08",
          8682 => x"55748287",
          8683 => x"cc0ca83d",
          8684 => x"0d04ed3d",
          8685 => x"0d0280db",
          8686 => x"05330284",
          8687 => x"0580df05",
          8688 => x"33575782",
          8689 => x"53953dd0",
          8690 => x"0552963d",
          8691 => x"51d2ea3f",
          8692 => x"8287cc08",
          8693 => x"558287cc",
          8694 => x"0880cf38",
          8695 => x"785a6552",
          8696 => x"953dd405",
          8697 => x"51c9b63f",
          8698 => x"8287cc08",
          8699 => x"558287cc",
          8700 => x"08b83802",
          8701 => x"80cf0533",
          8702 => x"81a00654",
          8703 => x"865573aa",
          8704 => x"3875a706",
          8705 => x"6171098b",
          8706 => x"12337106",
          8707 => x"7a740607",
          8708 => x"51575556",
          8709 => x"748b1534",
          8710 => x"7854810b",
          8711 => x"83153478",
          8712 => x"51ffb4aa",
          8713 => x"3f8287cc",
          8714 => x"08557482",
          8715 => x"87cc0c95",
          8716 => x"3d0d04ef",
          8717 => x"3d0d6456",
          8718 => x"8253933d",
          8719 => x"d0055294",
          8720 => x"3d51d1f5",
          8721 => x"3f8287cc",
          8722 => x"08558287",
          8723 => x"cc0880cb",
          8724 => x"38765863",
          8725 => x"52933dd4",
          8726 => x"0551c8c1",
          8727 => x"3f8287cc",
          8728 => x"08558287",
          8729 => x"cc08b438",
          8730 => x"0280c705",
          8731 => x"3381a006",
          8732 => x"54865573",
          8733 => x"a6388416",
          8734 => x"22861722",
          8735 => x"71902b07",
          8736 => x"5354961f",
          8737 => x"51ffb0c3",
          8738 => x"3f765481",
          8739 => x"0b831534",
          8740 => x"7651ffb3",
          8741 => x"b93f8287",
          8742 => x"cc085574",
          8743 => x"8287cc0c",
          8744 => x"933d0d04",
          8745 => x"ea3d0d69",
          8746 => x"6b5c5a80",
          8747 => x"53983dd0",
          8748 => x"0552993d",
          8749 => x"51d1823f",
          8750 => x"8287cc08",
          8751 => x"8287cc08",
          8752 => x"30708287",
          8753 => x"cc080780",
          8754 => x"25515557",
          8755 => x"79802e81",
          8756 => x"85388170",
          8757 => x"75065555",
          8758 => x"73802e80",
          8759 => x"f9387b5d",
          8760 => x"805f8052",
          8761 => x"8d3d7052",
          8762 => x"54ffbeaa",
          8763 => x"3f8287cc",
          8764 => x"08578287",
          8765 => x"cc0880d1",
          8766 => x"38745273",
          8767 => x"51c3dd3f",
          8768 => x"8287cc08",
          8769 => x"578287cc",
          8770 => x"08bf3882",
          8771 => x"87cc0882",
          8772 => x"87cc0865",
          8773 => x"5b595678",
          8774 => x"1881197b",
          8775 => x"18565955",
          8776 => x"74337434",
          8777 => x"8116568a",
          8778 => x"7827ec38",
          8779 => x"8b56751a",
          8780 => x"54807434",
          8781 => x"75802e9e",
          8782 => x"38ff1670",
          8783 => x"1b703351",
          8784 => x"555673a0",
          8785 => x"2ee8388e",
          8786 => x"3976842e",
          8787 => x"09810686",
          8788 => x"38807a34",
          8789 => x"80577630",
          8790 => x"70780780",
          8791 => x"2551547a",
          8792 => x"802e80c1",
          8793 => x"3873802e",
          8794 => x"bc387ba0",
          8795 => x"11085351",
          8796 => x"ffb1943f",
          8797 => x"8287cc08",
          8798 => x"578287cc",
          8799 => x"08a7387b",
          8800 => x"70335555",
          8801 => x"80c35673",
          8802 => x"832e8b38",
          8803 => x"80e45673",
          8804 => x"842e8338",
          8805 => x"a7567515",
          8806 => x"b40551ff",
          8807 => x"ade43f82",
          8808 => x"87cc087b",
          8809 => x"0c768287",
          8810 => x"cc0c983d",
          8811 => x"0d04e63d",
          8812 => x"0d82539c",
          8813 => x"3dffb805",
          8814 => x"529d3d51",
          8815 => x"cefb3f82",
          8816 => x"87cc0882",
          8817 => x"87cc0856",
          8818 => x"548287cc",
          8819 => x"08839838",
          8820 => x"8b53a052",
          8821 => x"8b3d7052",
          8822 => x"59ffaec1",
          8823 => x"3f736d70",
          8824 => x"337081ff",
          8825 => x"06525755",
          8826 => x"579f7427",
          8827 => x"81bc3878",
          8828 => x"587481ff",
          8829 => x"066d8105",
          8830 => x"4e705255",
          8831 => x"ffaf8a3f",
          8832 => x"8287cc08",
          8833 => x"802ea538",
          8834 => x"6c703370",
          8835 => x"535754ff",
          8836 => x"aefe3f82",
          8837 => x"87cc0880",
          8838 => x"2e8d3874",
          8839 => x"882b7607",
          8840 => x"6d81054e",
          8841 => x"55863982",
          8842 => x"87cc0855",
          8843 => x"ff9f1570",
          8844 => x"83ffff06",
          8845 => x"51547399",
          8846 => x"268a38e0",
          8847 => x"157083ff",
          8848 => x"ff065654",
          8849 => x"80ff7527",
          8850 => x"87388280",
          8851 => x"94153355",
          8852 => x"74802ea3",
          8853 => x"38745282",
          8854 => x"829451ff",
          8855 => x"ae8a3f82",
          8856 => x"87cc0893",
          8857 => x"3881ff75",
          8858 => x"27883876",
          8859 => x"89268838",
          8860 => x"8b398a77",
          8861 => x"27863886",
          8862 => x"5581ec39",
          8863 => x"81ff7527",
          8864 => x"8f387488",
          8865 => x"2a547378",
          8866 => x"7081055a",
          8867 => x"34811757",
          8868 => x"74787081",
          8869 => x"055a3481",
          8870 => x"176d7033",
          8871 => x"7081ff06",
          8872 => x"52575557",
          8873 => x"739f26fe",
          8874 => x"c8388b3d",
          8875 => x"33548655",
          8876 => x"7381e52e",
          8877 => x"81b13876",
          8878 => x"802e9938",
          8879 => x"02a70555",
          8880 => x"76157033",
          8881 => x"515473a0",
          8882 => x"2e098106",
          8883 => x"8738ff17",
          8884 => x"5776ed38",
          8885 => x"79418043",
          8886 => x"8052913d",
          8887 => x"705255ff",
          8888 => x"bab43f82",
          8889 => x"87cc0854",
          8890 => x"8287cc08",
          8891 => x"80f73881",
          8892 => x"527451ff",
          8893 => x"bfe63f82",
          8894 => x"87cc0854",
          8895 => x"8287cc08",
          8896 => x"8d387680",
          8897 => x"c4386754",
          8898 => x"e5743480",
          8899 => x"c6398287",
          8900 => x"cc08842e",
          8901 => x"09810680",
          8902 => x"cc388054",
          8903 => x"76742e80",
          8904 => x"c4388152",
          8905 => x"7451ffbd",
          8906 => x"b13f8287",
          8907 => x"cc085482",
          8908 => x"87cc08b1",
          8909 => x"38a05382",
          8910 => x"87cc0852",
          8911 => x"6751ffab",
          8912 => x"dc3f6754",
          8913 => x"880b8b15",
          8914 => x"348b5378",
          8915 => x"526751ff",
          8916 => x"aba83f79",
          8917 => x"54810b83",
          8918 => x"15347951",
          8919 => x"ffadef3f",
          8920 => x"8287cc08",
          8921 => x"54735574",
          8922 => x"8287cc0c",
          8923 => x"9c3d0d04",
          8924 => x"f23d0d60",
          8925 => x"62028805",
          8926 => x"80cb0533",
          8927 => x"933dfc05",
          8928 => x"55725440",
          8929 => x"5e5ad2da",
          8930 => x"3f8287cc",
          8931 => x"08588287",
          8932 => x"cc0882bd",
          8933 => x"38911a33",
          8934 => x"587782b5",
          8935 => x"387c802e",
          8936 => x"97388c1a",
          8937 => x"08597890",
          8938 => x"38901a33",
          8939 => x"70812a70",
          8940 => x"81065155",
          8941 => x"55739038",
          8942 => x"87548297",
          8943 => x"39825882",
          8944 => x"90398158",
          8945 => x"828b397e",
          8946 => x"8a112270",
          8947 => x"892b7055",
          8948 => x"7f545656",
          8949 => x"56ff9493",
          8950 => x"3fff147d",
          8951 => x"06703070",
          8952 => x"72079f2a",
          8953 => x"8287cc08",
          8954 => x"058c1908",
          8955 => x"7c405a5d",
          8956 => x"55558177",
          8957 => x"27883898",
          8958 => x"16087726",
          8959 => x"83388257",
          8960 => x"76775659",
          8961 => x"80567452",
          8962 => x"7951ffae",
          8963 => x"9a3f8115",
          8964 => x"7f555598",
          8965 => x"14087526",
          8966 => x"83388255",
          8967 => x"8287cc08",
          8968 => x"812eff99",
          8969 => x"388287cc",
          8970 => x"08ff2eff",
          8971 => x"95388287",
          8972 => x"cc088e38",
          8973 => x"81165675",
          8974 => x"7b2e0981",
          8975 => x"06873893",
          8976 => x"39745980",
          8977 => x"5674772e",
          8978 => x"098106ff",
          8979 => x"b9388758",
          8980 => x"80ff397d",
          8981 => x"802eba38",
          8982 => x"787b5555",
          8983 => x"7a802eb4",
          8984 => x"38811556",
          8985 => x"73812e09",
          8986 => x"81068338",
          8987 => x"ff567553",
          8988 => x"74527e51",
          8989 => x"ffafa93f",
          8990 => x"8287cc08",
          8991 => x"588287cc",
          8992 => x"0880ce38",
          8993 => x"748116ff",
          8994 => x"1656565c",
          8995 => x"73d33884",
          8996 => x"39ff195c",
          8997 => x"7e7c8c12",
          8998 => x"0c557d80",
          8999 => x"2eb33878",
          9000 => x"881b0c7c",
          9001 => x"8c1b0c90",
          9002 => x"1a3380c0",
          9003 => x"07547390",
          9004 => x"1b349815",
          9005 => x"08fe0590",
          9006 => x"16085754",
          9007 => x"75742691",
          9008 => x"38757b31",
          9009 => x"90160c84",
          9010 => x"15338107",
          9011 => x"54738416",
          9012 => x"34775473",
          9013 => x"8287cc0c",
          9014 => x"903d0d04",
          9015 => x"e93d0d6b",
          9016 => x"6d028805",
          9017 => x"80eb0533",
          9018 => x"9d3d545a",
          9019 => x"5c59c5be",
          9020 => x"3f8b5680",
          9021 => x"0b8287cc",
          9022 => x"08248bf8",
          9023 => x"388287cc",
          9024 => x"08842982",
          9025 => x"9ef00570",
          9026 => x"08515574",
          9027 => x"802e8438",
          9028 => x"80753482",
          9029 => x"87cc0881",
          9030 => x"ff065f81",
          9031 => x"527e51ff",
          9032 => x"a0d13f82",
          9033 => x"87cc0881",
          9034 => x"ff067081",
          9035 => x"06565783",
          9036 => x"56748bc0",
          9037 => x"3876822a",
          9038 => x"70810651",
          9039 => x"558a5674",
          9040 => x"8bb23899",
          9041 => x"3dfc0553",
          9042 => x"83527e51",
          9043 => x"ffa4f13f",
          9044 => x"8287cc08",
          9045 => x"99386755",
          9046 => x"74802e92",
          9047 => x"38748280",
          9048 => x"80268b38",
          9049 => x"ff157506",
          9050 => x"5574802e",
          9051 => x"83388148",
          9052 => x"78802e87",
          9053 => x"38848079",
          9054 => x"26923878",
          9055 => x"81800a26",
          9056 => x"8b38ff19",
          9057 => x"79065574",
          9058 => x"802e8638",
          9059 => x"93568ae4",
          9060 => x"3978892a",
          9061 => x"6e892a70",
          9062 => x"892b7759",
          9063 => x"4843597a",
          9064 => x"83388156",
          9065 => x"61307080",
          9066 => x"25770751",
          9067 => x"55915674",
          9068 => x"8ac23899",
          9069 => x"3df80553",
          9070 => x"81527e51",
          9071 => x"ffa4813f",
          9072 => x"81568287",
          9073 => x"cc088aac",
          9074 => x"3877832a",
          9075 => x"70770682",
          9076 => x"87cc0843",
          9077 => x"56457483",
          9078 => x"38bf4166",
          9079 => x"558e5660",
          9080 => x"75268a90",
          9081 => x"38746131",
          9082 => x"70485580",
          9083 => x"ff75278a",
          9084 => x"83389356",
          9085 => x"78818026",
          9086 => x"89fa3877",
          9087 => x"812a7081",
          9088 => x"06564374",
          9089 => x"802e9538",
          9090 => x"77870655",
          9091 => x"74822e83",
          9092 => x"8d387781",
          9093 => x"06557480",
          9094 => x"2e838338",
          9095 => x"77810655",
          9096 => x"9356825e",
          9097 => x"74802e89",
          9098 => x"cb38785a",
          9099 => x"7d832e09",
          9100 => x"810680e1",
          9101 => x"3878ae38",
          9102 => x"66912a57",
          9103 => x"810b8282",
          9104 => x"b822565a",
          9105 => x"74802e9d",
          9106 => x"38747726",
          9107 => x"98388282",
          9108 => x"b8567910",
          9109 => x"82177022",
          9110 => x"57575a74",
          9111 => x"802e8638",
          9112 => x"767527ee",
          9113 => x"38795266",
          9114 => x"51ff8eff",
          9115 => x"3f8287cc",
          9116 => x"08842984",
          9117 => x"87057089",
          9118 => x"2a5e55a0",
          9119 => x"5c800b82",
          9120 => x"87cc08fc",
          9121 => x"808a0556",
          9122 => x"44fdfff0",
          9123 => x"0a752780",
          9124 => x"ec3888d3",
          9125 => x"3978ae38",
          9126 => x"668c2a57",
          9127 => x"810b8282",
          9128 => x"a822565a",
          9129 => x"74802e9d",
          9130 => x"38747726",
          9131 => x"98388282",
          9132 => x"a8567910",
          9133 => x"82177022",
          9134 => x"57575a74",
          9135 => x"802e8638",
          9136 => x"767527ee",
          9137 => x"38795266",
          9138 => x"51ff8e9f",
          9139 => x"3f8287cc",
          9140 => x"08108405",
          9141 => x"578287cc",
          9142 => x"089ff526",
          9143 => x"9638810b",
          9144 => x"8287cc08",
          9145 => x"108287cc",
          9146 => x"08057111",
          9147 => x"722a8305",
          9148 => x"59565e83",
          9149 => x"ff17892a",
          9150 => x"5d815ca0",
          9151 => x"44601c7d",
          9152 => x"11650569",
          9153 => x"7012ff05",
          9154 => x"71307072",
          9155 => x"0674315c",
          9156 => x"52595759",
          9157 => x"407d832e",
          9158 => x"09810689",
          9159 => x"38761c60",
          9160 => x"18415c84",
          9161 => x"39761d5d",
          9162 => x"79902918",
          9163 => x"70623168",
          9164 => x"58515574",
          9165 => x"762687af",
          9166 => x"38757c31",
          9167 => x"7d317a53",
          9168 => x"70653152",
          9169 => x"55ff8da3",
          9170 => x"3f8287cc",
          9171 => x"08587d83",
          9172 => x"2e098106",
          9173 => x"9b388287",
          9174 => x"cc0883ff",
          9175 => x"f52680dd",
          9176 => x"38788783",
          9177 => x"3879812a",
          9178 => x"5978fdbe",
          9179 => x"3886f839",
          9180 => x"7d822e09",
          9181 => x"810680c5",
          9182 => x"3883fff5",
          9183 => x"0b8287cc",
          9184 => x"0827a038",
          9185 => x"788f3879",
          9186 => x"1a557480",
          9187 => x"c0268638",
          9188 => x"7459fd96",
          9189 => x"39628106",
          9190 => x"5574802e",
          9191 => x"8f38835e",
          9192 => x"fd883982",
          9193 => x"87cc089f",
          9194 => x"f5269238",
          9195 => x"7886b838",
          9196 => x"791a5981",
          9197 => x"807927fc",
          9198 => x"f13886ab",
          9199 => x"3980557d",
          9200 => x"812e0981",
          9201 => x"0683387d",
          9202 => x"559ff578",
          9203 => x"278b3874",
          9204 => x"8106558e",
          9205 => x"5674869c",
          9206 => x"38848053",
          9207 => x"80527a51",
          9208 => x"ffa2ba3f",
          9209 => x"8b538280",
          9210 => x"d0527a51",
          9211 => x"ffa28b3f",
          9212 => x"8480528b",
          9213 => x"1b51ffa1",
          9214 => x"b43f798d",
          9215 => x"1c347b83",
          9216 => x"ffff0652",
          9217 => x"8e1b51ff",
          9218 => x"a1a33f81",
          9219 => x"0b901c34",
          9220 => x"7d833270",
          9221 => x"3070962a",
          9222 => x"84800654",
          9223 => x"5155911b",
          9224 => x"51ffa189",
          9225 => x"3f665574",
          9226 => x"83ffff26",
          9227 => x"90387483",
          9228 => x"ffff0652",
          9229 => x"931b51ff",
          9230 => x"a0f33f8a",
          9231 => x"397452a0",
          9232 => x"1b51ffa1",
          9233 => x"863ff80b",
          9234 => x"951c34bf",
          9235 => x"52981b51",
          9236 => x"ffa0da3f",
          9237 => x"81ff529a",
          9238 => x"1b51ffa0",
          9239 => x"d03f6052",
          9240 => x"9c1b51ff",
          9241 => x"a0e53f7d",
          9242 => x"832e0981",
          9243 => x"0680cb38",
          9244 => x"8288b20a",
          9245 => x"5280c31b",
          9246 => x"51ffa0cf",
          9247 => x"3f7c52a4",
          9248 => x"1b51ffa0",
          9249 => x"c63f8252",
          9250 => x"ac1b51ff",
          9251 => x"a0bd3f81",
          9252 => x"52b01b51",
          9253 => x"ffa0963f",
          9254 => x"8652b21b",
          9255 => x"51ffa08d",
          9256 => x"3fff800b",
          9257 => x"80c01c34",
          9258 => x"a90b80c2",
          9259 => x"1c349353",
          9260 => x"8280dc52",
          9261 => x"80c71b51",
          9262 => x"ae398288",
          9263 => x"b20a52a7",
          9264 => x"1b51ffa0",
          9265 => x"863f7c83",
          9266 => x"ffff0652",
          9267 => x"961b51ff",
          9268 => x"9fdb3fff",
          9269 => x"800ba41c",
          9270 => x"34a90ba6",
          9271 => x"1c349353",
          9272 => x"8280f052",
          9273 => x"ab1b51ff",
          9274 => x"a0903f82",
          9275 => x"d4d55283",
          9276 => x"fe1b7052",
          9277 => x"59ff9fb5",
          9278 => x"3f815460",
          9279 => x"537a527e",
          9280 => x"51ff9bd8",
          9281 => x"3f815682",
          9282 => x"87cc0883",
          9283 => x"e7387d83",
          9284 => x"2e098106",
          9285 => x"80ee3875",
          9286 => x"54608605",
          9287 => x"537a527e",
          9288 => x"51ff9bb8",
          9289 => x"3f848053",
          9290 => x"80527a51",
          9291 => x"ff9fee3f",
          9292 => x"848b85a4",
          9293 => x"d2527a51",
          9294 => x"ff9f903f",
          9295 => x"868a85e4",
          9296 => x"f25283e4",
          9297 => x"1b51ff9f",
          9298 => x"823fff18",
          9299 => x"5283e81b",
          9300 => x"51ff9ef7",
          9301 => x"3f825283",
          9302 => x"ec1b51ff",
          9303 => x"9eed3f82",
          9304 => x"d4d55278",
          9305 => x"51ff9ec5",
          9306 => x"3f755460",
          9307 => x"8705537a",
          9308 => x"527e51ff",
          9309 => x"9ae63f75",
          9310 => x"54601653",
          9311 => x"7a527e51",
          9312 => x"ff9ad93f",
          9313 => x"65538052",
          9314 => x"7a51ff9f",
          9315 => x"903f7f56",
          9316 => x"80587d83",
          9317 => x"2e098106",
          9318 => x"9a38f852",
          9319 => x"7a51ff9e",
          9320 => x"aa3fff52",
          9321 => x"841b51ff",
          9322 => x"9ea13ff0",
          9323 => x"0a52881b",
          9324 => x"51913987",
          9325 => x"fffff855",
          9326 => x"7d812e83",
          9327 => x"38f85574",
          9328 => x"527a51ff",
          9329 => x"9e853f7c",
          9330 => x"55615774",
          9331 => x"62268338",
          9332 => x"74577654",
          9333 => x"75537a52",
          9334 => x"7e51ff99",
          9335 => x"ff3f8287",
          9336 => x"cc088287",
          9337 => x"38848053",
          9338 => x"8287cc08",
          9339 => x"527a51ff",
          9340 => x"9eab3f76",
          9341 => x"16757831",
          9342 => x"565674cd",
          9343 => x"38811858",
          9344 => x"77802eff",
          9345 => x"8d387955",
          9346 => x"7d832e83",
          9347 => x"38635561",
          9348 => x"57746226",
          9349 => x"83387457",
          9350 => x"76547553",
          9351 => x"7a527e51",
          9352 => x"ff99b93f",
          9353 => x"8287cc08",
          9354 => x"81c13876",
          9355 => x"16757831",
          9356 => x"565674db",
          9357 => x"388c567d",
          9358 => x"832e9338",
          9359 => x"86566683",
          9360 => x"ffff268a",
          9361 => x"3884567d",
          9362 => x"822e8338",
          9363 => x"81566481",
          9364 => x"06587780",
          9365 => x"fe388480",
          9366 => x"5377527a",
          9367 => x"51ff9dbd",
          9368 => x"3f82d4d5",
          9369 => x"527851ff",
          9370 => x"9cc33f83",
          9371 => x"be1b5577",
          9372 => x"7534810b",
          9373 => x"81163481",
          9374 => x"0b821634",
          9375 => x"77831634",
          9376 => x"75841634",
          9377 => x"60670556",
          9378 => x"80fdc152",
          9379 => x"7551ff86",
          9380 => x"da3ffe0b",
          9381 => x"85163482",
          9382 => x"87cc0882",
          9383 => x"2abf0756",
          9384 => x"75861634",
          9385 => x"8287cc08",
          9386 => x"87163460",
          9387 => x"5283c61b",
          9388 => x"51ff9c97",
          9389 => x"3f665283",
          9390 => x"ca1b51ff",
          9391 => x"9c8d3f81",
          9392 => x"5477537a",
          9393 => x"527e51ff",
          9394 => x"98923f81",
          9395 => x"568287cc",
          9396 => x"08a23880",
          9397 => x"5380527e",
          9398 => x"51ff99e4",
          9399 => x"3f815682",
          9400 => x"87cc0890",
          9401 => x"3889398e",
          9402 => x"568a3981",
          9403 => x"56863982",
          9404 => x"87cc0856",
          9405 => x"758287cc",
          9406 => x"0c993d0d",
          9407 => x"04f53d0d",
          9408 => x"7d605b59",
          9409 => x"807960ff",
          9410 => x"055a5757",
          9411 => x"767825b4",
          9412 => x"388d3df8",
          9413 => x"11555581",
          9414 => x"53fc1552",
          9415 => x"7951c9dc",
          9416 => x"3f7a812e",
          9417 => x"0981069c",
          9418 => x"388c3d33",
          9419 => x"55748d2e",
          9420 => x"db387476",
          9421 => x"70810558",
          9422 => x"34811757",
          9423 => x"748a2e09",
          9424 => x"8106c938",
          9425 => x"80763478",
          9426 => x"55768338",
          9427 => x"76557482",
          9428 => x"87cc0c8d",
          9429 => x"3d0d04f7",
          9430 => x"3d0d7b02",
          9431 => x"8405b305",
          9432 => x"33595777",
          9433 => x"8a2e0981",
          9434 => x"0687388d",
          9435 => x"527651e7",
          9436 => x"3f841708",
          9437 => x"56807624",
          9438 => x"be388817",
          9439 => x"0877178c",
          9440 => x"05565977",
          9441 => x"75348116",
          9442 => x"56bb7625",
          9443 => x"a1388b3d",
          9444 => x"fc055475",
          9445 => x"538c1752",
          9446 => x"760851cb",
          9447 => x"dc3f7976",
          9448 => x"32703070",
          9449 => x"72079f2a",
          9450 => x"70305351",
          9451 => x"56567584",
          9452 => x"180c8119",
          9453 => x"88180c8b",
          9454 => x"3d0d04f9",
          9455 => x"3d0d7984",
          9456 => x"11085656",
          9457 => x"807524a7",
          9458 => x"38893dfc",
          9459 => x"05547453",
          9460 => x"8c165275",
          9461 => x"0851cba1",
          9462 => x"3f8287cc",
          9463 => x"08913884",
          9464 => x"1608782e",
          9465 => x"09810687",
          9466 => x"38881608",
          9467 => x"558339ff",
          9468 => x"55748287",
          9469 => x"cc0c893d",
          9470 => x"0d04fd3d",
          9471 => x"0d755480",
          9472 => x"cc538052",
          9473 => x"7351ff9a",
          9474 => x"943f7674",
          9475 => x"0c853d0d",
          9476 => x"04ea3d0d",
          9477 => x"0280e305",
          9478 => x"336a5386",
          9479 => x"3d705354",
          9480 => x"54d83f73",
          9481 => x"527251fe",
          9482 => x"ae3f7251",
          9483 => x"ff8d3f98",
          9484 => x"3d0d0400",
          9485 => x"00ffffff",
          9486 => x"ff00ffff",
          9487 => x"ffff00ff",
          9488 => x"ffffff00",
          9489 => x"00000e06",
          9490 => x"00000d8a",
          9491 => x"00000d91",
          9492 => x"00000d98",
          9493 => x"00000d9f",
          9494 => x"00000da6",
          9495 => x"00000dad",
          9496 => x"00000db4",
          9497 => x"00000dbb",
          9498 => x"00000dc2",
          9499 => x"00000dc9",
          9500 => x"00000dd0",
          9501 => x"00000dd6",
          9502 => x"00000ddc",
          9503 => x"00000de2",
          9504 => x"00000de8",
          9505 => x"00000dee",
          9506 => x"00000df4",
          9507 => x"00000dfa",
          9508 => x"00000e00",
          9509 => x"00002542",
          9510 => x"00002548",
          9511 => x"0000254e",
          9512 => x"00002554",
          9513 => x"0000255a",
          9514 => x"0000317c",
          9515 => x"00003270",
          9516 => x"00003363",
          9517 => x"00003597",
          9518 => x"00003258",
          9519 => x"00003051",
          9520 => x"00003413",
          9521 => x"0000356e",
          9522 => x"00003450",
          9523 => x"000034e6",
          9524 => x"0000346c",
          9525 => x"00003313",
          9526 => x"00003051",
          9527 => x"00003363",
          9528 => x"00003386",
          9529 => x"00003413",
          9530 => x"00003051",
          9531 => x"00003051",
          9532 => x"0000346c",
          9533 => x"000034e6",
          9534 => x"0000356e",
          9535 => x"00003597",
          9536 => x"64696e69",
          9537 => x"74000000",
          9538 => x"64696f63",
          9539 => x"746c0000",
          9540 => x"66696e69",
          9541 => x"74000000",
          9542 => x"666c6f61",
          9543 => x"64000000",
          9544 => x"66657865",
          9545 => x"63000000",
          9546 => x"6d636c65",
          9547 => x"61720000",
          9548 => x"6d636f70",
          9549 => x"79000000",
          9550 => x"6d646966",
          9551 => x"66000000",
          9552 => x"6d64756d",
          9553 => x"70000000",
          9554 => x"6d656200",
          9555 => x"6d656800",
          9556 => x"6d657700",
          9557 => x"68696400",
          9558 => x"68696500",
          9559 => x"68666400",
          9560 => x"68666500",
          9561 => x"63616c6c",
          9562 => x"00000000",
          9563 => x"6a6d7000",
          9564 => x"72657374",
          9565 => x"61727400",
          9566 => x"72657365",
          9567 => x"74000000",
          9568 => x"696e666f",
          9569 => x"00000000",
          9570 => x"74657374",
          9571 => x"00000000",
          9572 => x"74626173",
          9573 => x"69630000",
          9574 => x"6d626173",
          9575 => x"69630000",
          9576 => x"6b696c6f",
          9577 => x"00000000",
          9578 => x"65640000",
          9579 => x"4469736b",
          9580 => x"20457272",
          9581 => x"6f720a00",
          9582 => x"496e7465",
          9583 => x"726e616c",
          9584 => x"20657272",
          9585 => x"6f722e0a",
          9586 => x"00000000",
          9587 => x"4469736b",
          9588 => x"206e6f74",
          9589 => x"20726561",
          9590 => x"64792e0a",
          9591 => x"00000000",
          9592 => x"4e6f2066",
          9593 => x"696c6520",
          9594 => x"666f756e",
          9595 => x"642e0a00",
          9596 => x"4e6f2070",
          9597 => x"61746820",
          9598 => x"666f756e",
          9599 => x"642e0a00",
          9600 => x"496e7661",
          9601 => x"6c696420",
          9602 => x"66696c65",
          9603 => x"6e616d65",
          9604 => x"2e0a0000",
          9605 => x"41636365",
          9606 => x"73732064",
          9607 => x"656e6965",
          9608 => x"642e0a00",
          9609 => x"46696c65",
          9610 => x"20616c72",
          9611 => x"65616479",
          9612 => x"20657869",
          9613 => x"7374732e",
          9614 => x"0a000000",
          9615 => x"46696c65",
          9616 => x"2068616e",
          9617 => x"646c6520",
          9618 => x"696e7661",
          9619 => x"6c69642e",
          9620 => x"0a000000",
          9621 => x"53442069",
          9622 => x"73207772",
          9623 => x"69746520",
          9624 => x"70726f74",
          9625 => x"65637465",
          9626 => x"642e0a00",
          9627 => x"44726976",
          9628 => x"65206e75",
          9629 => x"6d626572",
          9630 => x"20697320",
          9631 => x"696e7661",
          9632 => x"6c69642e",
          9633 => x"0a000000",
          9634 => x"4469736b",
          9635 => x"206e6f74",
          9636 => x"20656e61",
          9637 => x"626c6564",
          9638 => x"2e0a0000",
          9639 => x"4e6f2063",
          9640 => x"6f6d7061",
          9641 => x"7469626c",
          9642 => x"65206669",
          9643 => x"6c657379",
          9644 => x"7374656d",
          9645 => x"20666f75",
          9646 => x"6e64206f",
          9647 => x"6e206469",
          9648 => x"736b2e0a",
          9649 => x"00000000",
          9650 => x"466f726d",
          9651 => x"61742061",
          9652 => x"626f7274",
          9653 => x"65642e0a",
          9654 => x"00000000",
          9655 => x"54696d65",
          9656 => x"6f75742c",
          9657 => x"206f7065",
          9658 => x"72617469",
          9659 => x"6f6e2063",
          9660 => x"616e6365",
          9661 => x"6c6c6564",
          9662 => x"2e0a0000",
          9663 => x"46696c65",
          9664 => x"20697320",
          9665 => x"6c6f636b",
          9666 => x"65642e0a",
          9667 => x"00000000",
          9668 => x"496e7375",
          9669 => x"66666963",
          9670 => x"69656e74",
          9671 => x"206d656d",
          9672 => x"6f72792e",
          9673 => x"0a000000",
          9674 => x"546f6f20",
          9675 => x"6d616e79",
          9676 => x"206f7065",
          9677 => x"6e206669",
          9678 => x"6c65732e",
          9679 => x"0a000000",
          9680 => x"50617261",
          9681 => x"6d657465",
          9682 => x"72732069",
          9683 => x"6e636f72",
          9684 => x"72656374",
          9685 => x"2e0a0000",
          9686 => x"53756363",
          9687 => x"6573732e",
          9688 => x"0a000000",
          9689 => x"556e6b6e",
          9690 => x"6f776e20",
          9691 => x"6572726f",
          9692 => x"722e0a00",
          9693 => x"0a256c75",
          9694 => x"20627974",
          9695 => x"65732025",
          9696 => x"73206174",
          9697 => x"20256c75",
          9698 => x"20627974",
          9699 => x"65732f73",
          9700 => x"65632e0a",
          9701 => x"00000000",
          9702 => x"72656164",
          9703 => x"00000000",
          9704 => x"25303858",
          9705 => x"00000000",
          9706 => x"3a202000",
          9707 => x"25303458",
          9708 => x"00000000",
          9709 => x"20202020",
          9710 => x"20202020",
          9711 => x"00000000",
          9712 => x"25303258",
          9713 => x"00000000",
          9714 => x"20200000",
          9715 => x"207c0000",
          9716 => x"7c0d0a00",
          9717 => x"5a505554",
          9718 => x"41000000",
          9719 => x"0a2a2a20",
          9720 => x"25732028",
          9721 => x"00000000",
          9722 => x"30322f30",
          9723 => x"352f3230",
          9724 => x"32300000",
          9725 => x"76312e35",
          9726 => x"32000000",
          9727 => x"205a5055",
          9728 => x"2c207265",
          9729 => x"76202530",
          9730 => x"32782920",
          9731 => x"25732025",
          9732 => x"73202a2a",
          9733 => x"0a0a0000",
          9734 => x"5a505554",
          9735 => x"4120496e",
          9736 => x"74657272",
          9737 => x"75707420",
          9738 => x"48616e64",
          9739 => x"6c65720a",
          9740 => x"00000000",
          9741 => x"54696d65",
          9742 => x"7220696e",
          9743 => x"74657272",
          9744 => x"7570740a",
          9745 => x"00000000",
          9746 => x"50533220",
          9747 => x"696e7465",
          9748 => x"72727570",
          9749 => x"740a0000",
          9750 => x"494f4354",
          9751 => x"4c205244",
          9752 => x"20696e74",
          9753 => x"65727275",
          9754 => x"70740a00",
          9755 => x"494f4354",
          9756 => x"4c205752",
          9757 => x"20696e74",
          9758 => x"65727275",
          9759 => x"70740a00",
          9760 => x"55415254",
          9761 => x"30205258",
          9762 => x"20696e74",
          9763 => x"65727275",
          9764 => x"70740a00",
          9765 => x"55415254",
          9766 => x"30205458",
          9767 => x"20696e74",
          9768 => x"65727275",
          9769 => x"70740a00",
          9770 => x"55415254",
          9771 => x"31205258",
          9772 => x"20696e74",
          9773 => x"65727275",
          9774 => x"70740a00",
          9775 => x"55415254",
          9776 => x"31205458",
          9777 => x"20696e74",
          9778 => x"65727275",
          9779 => x"70740a00",
          9780 => x"53657474",
          9781 => x"696e6720",
          9782 => x"75702074",
          9783 => x"696d6572",
          9784 => x"2e2e2e0a",
          9785 => x"00000000",
          9786 => x"456e6162",
          9787 => x"6c696e67",
          9788 => x"2074696d",
          9789 => x"65722e2e",
          9790 => x"2e0a0000",
          9791 => x"6175746f",
          9792 => x"65786563",
          9793 => x"2e626174",
          9794 => x"00000000",
          9795 => x"7a707574",
          9796 => x"612e6873",
          9797 => x"74000000",
          9798 => x"303a0000",
          9799 => x"4661696c",
          9800 => x"65642074",
          9801 => x"6f20696e",
          9802 => x"69746961",
          9803 => x"6c697365",
          9804 => x"20736420",
          9805 => x"63617264",
          9806 => x"20302c20",
          9807 => x"706c6561",
          9808 => x"73652069",
          9809 => x"6e697420",
          9810 => x"6d616e75",
          9811 => x"616c6c79",
          9812 => x"2e0a0000",
          9813 => x"2a200000",
          9814 => x"42616420",
          9815 => x"6469736b",
          9816 => x"20696421",
          9817 => x"0a000000",
          9818 => x"496e6974",
          9819 => x"69616c69",
          9820 => x"7365642e",
          9821 => x"0a000000",
          9822 => x"4661696c",
          9823 => x"65642074",
          9824 => x"6f20696e",
          9825 => x"69746961",
          9826 => x"6c697365",
          9827 => x"2e0a0000",
          9828 => x"72633d25",
          9829 => x"640a0000",
          9830 => x"25753a00",
          9831 => x"436c6561",
          9832 => x"72696e67",
          9833 => x"2e2e2e2e",
          9834 => x"00000000",
          9835 => x"436f7079",
          9836 => x"696e672e",
          9837 => x"2e2e0000",
          9838 => x"436f6d70",
          9839 => x"6172696e",
          9840 => x"672e2e2e",
          9841 => x"00000000",
          9842 => x"2530386c",
          9843 => x"78282530",
          9844 => x"3878292d",
          9845 => x"3e253038",
          9846 => x"6c782825",
          9847 => x"30387829",
          9848 => x"0a000000",
          9849 => x"44756d70",
          9850 => x"204d656d",
          9851 => x"6f72790a",
          9852 => x"00000000",
          9853 => x"0a436f6d",
          9854 => x"706c6574",
          9855 => x"652e0a00",
          9856 => x"25303858",
          9857 => x"20253032",
          9858 => x"582d0000",
          9859 => x"3f3f3f0a",
          9860 => x"00000000",
          9861 => x"25303858",
          9862 => x"20253034",
          9863 => x"582d0000",
          9864 => x"25303858",
          9865 => x"20253038",
          9866 => x"582d0000",
          9867 => x"44697361",
          9868 => x"626c696e",
          9869 => x"6720696e",
          9870 => x"74657272",
          9871 => x"75707473",
          9872 => x"0a000000",
          9873 => x"456e6162",
          9874 => x"6c696e67",
          9875 => x"20696e74",
          9876 => x"65727275",
          9877 => x"7074730a",
          9878 => x"00000000",
          9879 => x"44697361",
          9880 => x"626c6564",
          9881 => x"20756172",
          9882 => x"74206669",
          9883 => x"666f0a00",
          9884 => x"456e6162",
          9885 => x"6c696e67",
          9886 => x"20756172",
          9887 => x"74206669",
          9888 => x"666f0a00",
          9889 => x"45786563",
          9890 => x"7574696e",
          9891 => x"6720636f",
          9892 => x"64652040",
          9893 => x"20253038",
          9894 => x"78202e2e",
          9895 => x"2e0a0000",
          9896 => x"43616c6c",
          9897 => x"696e6720",
          9898 => x"636f6465",
          9899 => x"20402025",
          9900 => x"30387820",
          9901 => x"2e2e2e0a",
          9902 => x"00000000",
          9903 => x"43616c6c",
          9904 => x"20726574",
          9905 => x"75726e65",
          9906 => x"6420636f",
          9907 => x"64652028",
          9908 => x"2564292e",
          9909 => x"0a000000",
          9910 => x"52657374",
          9911 => x"61727469",
          9912 => x"6e672061",
          9913 => x"70706c69",
          9914 => x"63617469",
          9915 => x"6f6e2e2e",
          9916 => x"2e0a0000",
          9917 => x"436f6c64",
          9918 => x"20726562",
          9919 => x"6f6f7469",
          9920 => x"6e672e2e",
          9921 => x"2e0a0000",
          9922 => x"5a505500",
          9923 => x"62696e00",
          9924 => x"25643a5c",
          9925 => x"25735c25",
          9926 => x"732e2573",
          9927 => x"00000000",
          9928 => x"25643a5c",
          9929 => x"25735c25",
          9930 => x"73000000",
          9931 => x"25643a5c",
          9932 => x"25730000",
          9933 => x"42616420",
          9934 => x"636f6d6d",
          9935 => x"616e642e",
          9936 => x"0a000000",
          9937 => x"52756e6e",
          9938 => x"696e672e",
          9939 => x"2e2e0a00",
          9940 => x"456e6162",
          9941 => x"6c696e67",
          9942 => x"20696e74",
          9943 => x"65727275",
          9944 => x"7074732e",
          9945 => x"2e2e0a00",
          9946 => x"25642f25",
          9947 => x"642f2564",
          9948 => x"2025643a",
          9949 => x"25643a25",
          9950 => x"642e2564",
          9951 => x"25640a00",
          9952 => x"536f4320",
          9953 => x"436f6e66",
          9954 => x"69677572",
          9955 => x"6174696f",
          9956 => x"6e000000",
          9957 => x"20286672",
          9958 => x"6f6d2053",
          9959 => x"6f432063",
          9960 => x"6f6e6669",
          9961 => x"67290000",
          9962 => x"3a0a4465",
          9963 => x"76696365",
          9964 => x"7320696d",
          9965 => x"706c656d",
          9966 => x"656e7465",
          9967 => x"643a0a00",
          9968 => x"20202020",
          9969 => x"57422053",
          9970 => x"4452414d",
          9971 => x"20202825",
          9972 => x"3038583a",
          9973 => x"25303858",
          9974 => x"292e0a00",
          9975 => x"20202020",
          9976 => x"53445241",
          9977 => x"4d202020",
          9978 => x"20202825",
          9979 => x"3038583a",
          9980 => x"25303858",
          9981 => x"292e0a00",
          9982 => x"20202020",
          9983 => x"494e534e",
          9984 => x"20425241",
          9985 => x"4d202825",
          9986 => x"3038583a",
          9987 => x"25303858",
          9988 => x"292e0a00",
          9989 => x"20202020",
          9990 => x"4252414d",
          9991 => x"20202020",
          9992 => x"20202825",
          9993 => x"3038583a",
          9994 => x"25303858",
          9995 => x"292e0a00",
          9996 => x"20202020",
          9997 => x"52414d20",
          9998 => x"20202020",
          9999 => x"20202825",
         10000 => x"3038583a",
         10001 => x"25303858",
         10002 => x"292e0a00",
         10003 => x"20202020",
         10004 => x"53442043",
         10005 => x"41524420",
         10006 => x"20202844",
         10007 => x"65766963",
         10008 => x"6573203d",
         10009 => x"25303264",
         10010 => x"292e0a00",
         10011 => x"20202020",
         10012 => x"54494d45",
         10013 => x"52312020",
         10014 => x"20202854",
         10015 => x"696d6572",
         10016 => x"7320203d",
         10017 => x"25303264",
         10018 => x"292e0a00",
         10019 => x"20202020",
         10020 => x"494e5452",
         10021 => x"20435452",
         10022 => x"4c202843",
         10023 => x"68616e6e",
         10024 => x"656c733d",
         10025 => x"25303264",
         10026 => x"292e0a00",
         10027 => x"20202020",
         10028 => x"57495348",
         10029 => x"424f4e45",
         10030 => x"20425553",
         10031 => x"0a000000",
         10032 => x"20202020",
         10033 => x"57422049",
         10034 => x"32430a00",
         10035 => x"20202020",
         10036 => x"494f4354",
         10037 => x"4c0a0000",
         10038 => x"20202020",
         10039 => x"5053320a",
         10040 => x"00000000",
         10041 => x"20202020",
         10042 => x"5350490a",
         10043 => x"00000000",
         10044 => x"41646472",
         10045 => x"65737365",
         10046 => x"733a0a00",
         10047 => x"20202020",
         10048 => x"43505520",
         10049 => x"52657365",
         10050 => x"74205665",
         10051 => x"63746f72",
         10052 => x"20416464",
         10053 => x"72657373",
         10054 => x"203d2025",
         10055 => x"3038580a",
         10056 => x"00000000",
         10057 => x"20202020",
         10058 => x"43505520",
         10059 => x"4d656d6f",
         10060 => x"72792053",
         10061 => x"74617274",
         10062 => x"20416464",
         10063 => x"72657373",
         10064 => x"203d2025",
         10065 => x"3038580a",
         10066 => x"00000000",
         10067 => x"20202020",
         10068 => x"53746163",
         10069 => x"6b205374",
         10070 => x"61727420",
         10071 => x"41646472",
         10072 => x"65737320",
         10073 => x"20202020",
         10074 => x"203d2025",
         10075 => x"3038580a",
         10076 => x"00000000",
         10077 => x"4d697363",
         10078 => x"3a0a0000",
         10079 => x"20202020",
         10080 => x"5a505520",
         10081 => x"49642020",
         10082 => x"20202020",
         10083 => x"20202020",
         10084 => x"20202020",
         10085 => x"20202020",
         10086 => x"203d2025",
         10087 => x"3034580a",
         10088 => x"00000000",
         10089 => x"20202020",
         10090 => x"53797374",
         10091 => x"656d2043",
         10092 => x"6c6f636b",
         10093 => x"20467265",
         10094 => x"71202020",
         10095 => x"20202020",
         10096 => x"203d2025",
         10097 => x"642e2530",
         10098 => x"34644d48",
         10099 => x"7a0a0000",
         10100 => x"20202020",
         10101 => x"53445241",
         10102 => x"4d20436c",
         10103 => x"6f636b20",
         10104 => x"46726571",
         10105 => x"20202020",
         10106 => x"20202020",
         10107 => x"203d2025",
         10108 => x"642e2530",
         10109 => x"34644d48",
         10110 => x"7a0a0000",
         10111 => x"20202020",
         10112 => x"57697368",
         10113 => x"626f6e65",
         10114 => x"20534452",
         10115 => x"414d2043",
         10116 => x"6c6f636b",
         10117 => x"20467265",
         10118 => x"713d2025",
         10119 => x"642e2530",
         10120 => x"34644d48",
         10121 => x"7a0a0000",
         10122 => x"536d616c",
         10123 => x"6c000000",
         10124 => x"4d656469",
         10125 => x"756d0000",
         10126 => x"466c6578",
         10127 => x"00000000",
         10128 => x"45564f00",
         10129 => x"45564f6d",
         10130 => x"696e0000",
         10131 => x"556e6b6e",
         10132 => x"6f776e00",
         10133 => x"00007fb0",
         10134 => x"01000000",
         10135 => x"00000002",
         10136 => x"00007fac",
         10137 => x"01000000",
         10138 => x"00000003",
         10139 => x"00007fa8",
         10140 => x"01000000",
         10141 => x"00000004",
         10142 => x"00007fa4",
         10143 => x"01000000",
         10144 => x"00000005",
         10145 => x"00007fa0",
         10146 => x"01000000",
         10147 => x"00000006",
         10148 => x"00007f9c",
         10149 => x"01000000",
         10150 => x"00000007",
         10151 => x"00007f98",
         10152 => x"01000000",
         10153 => x"00000001",
         10154 => x"00007f94",
         10155 => x"01000000",
         10156 => x"00000008",
         10157 => x"00007f90",
         10158 => x"01000000",
         10159 => x"0000000b",
         10160 => x"00007f8c",
         10161 => x"01000000",
         10162 => x"00000009",
         10163 => x"00007f88",
         10164 => x"01000000",
         10165 => x"0000000a",
         10166 => x"00007f84",
         10167 => x"04000000",
         10168 => x"0000000d",
         10169 => x"00007f80",
         10170 => x"04000000",
         10171 => x"0000000c",
         10172 => x"00007f7c",
         10173 => x"04000000",
         10174 => x"0000000e",
         10175 => x"00007f78",
         10176 => x"03000000",
         10177 => x"0000000f",
         10178 => x"00007f74",
         10179 => x"04000000",
         10180 => x"0000000f",
         10181 => x"00007f70",
         10182 => x"04000000",
         10183 => x"00000010",
         10184 => x"00007f6c",
         10185 => x"04000000",
         10186 => x"00000011",
         10187 => x"00007f68",
         10188 => x"03000000",
         10189 => x"00000012",
         10190 => x"00007f64",
         10191 => x"03000000",
         10192 => x"00000013",
         10193 => x"00007f60",
         10194 => x"03000000",
         10195 => x"00000014",
         10196 => x"00007f5c",
         10197 => x"03000000",
         10198 => x"00000015",
         10199 => x"1b5b4400",
         10200 => x"1b5b4300",
         10201 => x"1b5b4200",
         10202 => x"1b5b4100",
         10203 => x"1b5b367e",
         10204 => x"1b5b357e",
         10205 => x"1b5b347e",
         10206 => x"1b304600",
         10207 => x"1b5b337e",
         10208 => x"1b5b327e",
         10209 => x"1b5b317e",
         10210 => x"10000000",
         10211 => x"0e000000",
         10212 => x"0d000000",
         10213 => x"0b000000",
         10214 => x"08000000",
         10215 => x"06000000",
         10216 => x"05000000",
         10217 => x"04000000",
         10218 => x"03000000",
         10219 => x"02000000",
         10220 => x"01000000",
         10221 => x"68697374",
         10222 => x"6f727900",
         10223 => x"68697374",
         10224 => x"00000000",
         10225 => x"21000000",
         10226 => x"25303464",
         10227 => x"20202573",
         10228 => x"0a000000",
         10229 => x"4661696c",
         10230 => x"65642074",
         10231 => x"6f207265",
         10232 => x"73657420",
         10233 => x"74686520",
         10234 => x"68697374",
         10235 => x"6f727920",
         10236 => x"66696c65",
         10237 => x"20746f20",
         10238 => x"454f462e",
         10239 => x"0a000000",
         10240 => x"43616e6e",
         10241 => x"6f74206f",
         10242 => x"70656e2f",
         10243 => x"63726561",
         10244 => x"74652068",
         10245 => x"6973746f",
         10246 => x"72792066",
         10247 => x"696c652c",
         10248 => x"20646973",
         10249 => x"61626c69",
         10250 => x"6e672e0a",
         10251 => x"00000000",
         10252 => x"53440000",
         10253 => x"222a2b2c",
         10254 => x"3a3b3c3d",
         10255 => x"3e3f5b5d",
         10256 => x"7c7f0000",
         10257 => x"46415400",
         10258 => x"46415433",
         10259 => x"32000000",
         10260 => x"ebfe904d",
         10261 => x"53444f53",
         10262 => x"352e3000",
         10263 => x"4e4f204e",
         10264 => x"414d4520",
         10265 => x"20202046",
         10266 => x"41543332",
         10267 => x"20202000",
         10268 => x"4e4f204e",
         10269 => x"414d4520",
         10270 => x"20202046",
         10271 => x"41542020",
         10272 => x"20202000",
         10273 => x"00008030",
         10274 => x"00000000",
         10275 => x"00000000",
         10276 => x"00000000",
         10277 => x"809a4541",
         10278 => x"8e418f80",
         10279 => x"45454549",
         10280 => x"49498e8f",
         10281 => x"9092924f",
         10282 => x"994f5555",
         10283 => x"59999a9b",
         10284 => x"9c9d9e9f",
         10285 => x"41494f55",
         10286 => x"a5a5a6a7",
         10287 => x"a8a9aaab",
         10288 => x"acadaeaf",
         10289 => x"b0b1b2b3",
         10290 => x"b4b5b6b7",
         10291 => x"b8b9babb",
         10292 => x"bcbdbebf",
         10293 => x"c0c1c2c3",
         10294 => x"c4c5c6c7",
         10295 => x"c8c9cacb",
         10296 => x"cccdcecf",
         10297 => x"d0d1d2d3",
         10298 => x"d4d5d6d7",
         10299 => x"d8d9dadb",
         10300 => x"dcdddedf",
         10301 => x"e0e1e2e3",
         10302 => x"e4e5e6e7",
         10303 => x"e8e9eaeb",
         10304 => x"ecedeeef",
         10305 => x"f0f1f2f3",
         10306 => x"f4f5f6f7",
         10307 => x"f8f9fafb",
         10308 => x"fcfdfeff",
         10309 => x"2b2e2c3b",
         10310 => x"3d5b5d2f",
         10311 => x"5c222a3a",
         10312 => x"3c3e3f7c",
         10313 => x"7f000000",
         10314 => x"00010004",
         10315 => x"00100040",
         10316 => x"01000200",
         10317 => x"00000000",
         10318 => x"00010002",
         10319 => x"00040008",
         10320 => x"00100020",
         10321 => x"00000000",
         10322 => x"00000000",
         10323 => x"00007500",
         10324 => x"01020100",
         10325 => x"00000000",
         10326 => x"00000000",
         10327 => x"00007508",
         10328 => x"01040100",
         10329 => x"00000000",
         10330 => x"00000000",
         10331 => x"00007510",
         10332 => x"01140300",
         10333 => x"00000000",
         10334 => x"00000000",
         10335 => x"00007518",
         10336 => x"012b0300",
         10337 => x"00000000",
         10338 => x"00000000",
         10339 => x"00007520",
         10340 => x"01300300",
         10341 => x"00000000",
         10342 => x"00000000",
         10343 => x"00007528",
         10344 => x"013c0400",
         10345 => x"00000000",
         10346 => x"00000000",
         10347 => x"00007530",
         10348 => x"013d0400",
         10349 => x"00000000",
         10350 => x"00000000",
         10351 => x"00007538",
         10352 => x"013f0400",
         10353 => x"00000000",
         10354 => x"00000000",
         10355 => x"00007540",
         10356 => x"01400400",
         10357 => x"00000000",
         10358 => x"00000000",
         10359 => x"00007548",
         10360 => x"01410400",
         10361 => x"00000000",
         10362 => x"00000000",
         10363 => x"0000754c",
         10364 => x"01420400",
         10365 => x"00000000",
         10366 => x"00000000",
         10367 => x"00007550",
         10368 => x"01430400",
         10369 => x"00000000",
         10370 => x"00000000",
         10371 => x"00007554",
         10372 => x"01500500",
         10373 => x"00000000",
         10374 => x"00000000",
         10375 => x"00007558",
         10376 => x"01510500",
         10377 => x"00000000",
         10378 => x"00000000",
         10379 => x"0000755c",
         10380 => x"01540500",
         10381 => x"00000000",
         10382 => x"00000000",
         10383 => x"00007560",
         10384 => x"01550500",
         10385 => x"00000000",
         10386 => x"00000000",
         10387 => x"00007564",
         10388 => x"01790700",
         10389 => x"00000000",
         10390 => x"00000000",
         10391 => x"0000756c",
         10392 => x"01780700",
         10393 => x"00000000",
         10394 => x"00000000",
         10395 => x"00007570",
         10396 => x"01820800",
         10397 => x"00000000",
         10398 => x"00000000",
         10399 => x"00007578",
         10400 => x"01830800",
         10401 => x"00000000",
         10402 => x"00000000",
         10403 => x"00007580",
         10404 => x"01850800",
         10405 => x"00000000",
         10406 => x"00000000",
         10407 => x"00007588",
         10408 => x"01870800",
         10409 => x"00000000",
         10410 => x"00000000",
         10411 => x"00007590",
         10412 => x"018c0900",
         10413 => x"00000000",
         10414 => x"00000000",
         10415 => x"00007598",
         10416 => x"018d0900",
         10417 => x"00000000",
         10418 => x"00000000",
         10419 => x"000075a0",
         10420 => x"018e0900",
         10421 => x"00000000",
         10422 => x"00000000",
         10423 => x"000075a8",
         10424 => x"018f0900",
         10425 => x"00000000",
         10426 => x"00000000",
         10427 => x"00000000",
         10428 => x"00000000",
         10429 => x"00007fff",
         10430 => x"00000000",
         10431 => x"00007fff",
         10432 => x"00010000",
         10433 => x"00007fff",
         10434 => x"00010000",
         10435 => x"00810000",
         10436 => x"01000000",
         10437 => x"017fffff",
         10438 => x"00000000",
         10439 => x"00000000",
         10440 => x"00007800",
         10441 => x"00000000",
         10442 => x"05f5e100",
         10443 => x"05f5e100",
         10444 => x"05f5e100",
         10445 => x"00000000",
         10446 => x"01010101",
         10447 => x"01010101",
         10448 => x"01011001",
         10449 => x"01000000",
         10450 => x"00000000",
         10451 => x"00000000",
         10452 => x"00000000",
         10453 => x"00000000",
         10454 => x"00000000",
         10455 => x"00000000",
         10456 => x"00000000",
         10457 => x"00000000",
         10458 => x"00000000",
         10459 => x"00000000",
         10460 => x"00000000",
         10461 => x"00000000",
         10462 => x"00000000",
         10463 => x"00000000",
         10464 => x"00000000",
         10465 => x"00000000",
         10466 => x"00000000",
         10467 => x"00000000",
         10468 => x"00000000",
         10469 => x"00000000",
         10470 => x"00000000",
         10471 => x"00000000",
         10472 => x"00000000",
         10473 => x"00000000",
         10474 => x"00007fb4",
         10475 => x"01000000",
         10476 => x"00007fbc",
         10477 => x"01000000",
         10478 => x"00007fc4",
         10479 => x"02000000",
         10480 => x"00000000",
         10481 => x"00000000",
         10482 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

