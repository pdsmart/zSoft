-- Byte Addressed 32bit/64bit BRAM module for the ZPU Evo implementation.
--
-- This template provides a 32bit wide bus on port A and a 64bit bus
-- on port B. This is typically used for the ZPU Boot BRAM where port B
-- is used exclusively for instruction storage.
--
-- Copyright 2018-2021 - Philip Smart for the ZPU Evo implementation.
-- History:
--   20190618  - Initial 32 bit dual port BRAM described by inference rather than
--               using an IP Megacore. This was to make it more portable but also
--               to allow 8/16/32 bit writes to the memory.
--   20210108  - Updated to 64bit on Port B to allow for the 64bit decoder on the ZPU.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPort3264BootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 3);
        memBWrite            : in  std_logic_vector(WORD_64BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_64BIT_RANGE)
    );
end DualPort3264BootBRAM;

architecture arch of DualPort3264BootBRAM is

    -- Declare 8 byte wide arrays for byte level addressing.
    type ramArray is array(natural range 0 to (2**(addrbits-3))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"fa",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"05",
            10 => x"52",
            11 => x"00",
            12 => x"08",
            13 => x"81",
            14 => x"06",
            15 => x"0b",
            16 => x"05",
            17 => x"06",
            18 => x"06",
            19 => x"00",
            20 => x"73",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"09",
            25 => x"72",
            26 => x"31",
            27 => x"51",
            28 => x"73",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"93",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"2b",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"06",
            45 => x"b0",
            46 => x"00",
            47 => x"00",
            48 => x"ff",
            49 => x"0a",
            50 => x"51",
            51 => x"00",
            52 => x"51",
            53 => x"05",
            54 => x"72",
            55 => x"00",
            56 => x"05",
            57 => x"06",
            58 => x"00",
            59 => x"00",
            60 => x"05",
            61 => x"06",
            62 => x"00",
            63 => x"00",
            64 => x"05",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"81",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"06",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"08",
            77 => x"05",
            78 => x"52",
            79 => x"00",
            80 => x"08",
            81 => x"06",
            82 => x"0b",
            83 => x"00",
            84 => x"08",
            85 => x"ac",
            86 => x"90",
            87 => x"00",
            88 => x"08",
            89 => x"ab",
            90 => x"90",
            91 => x"00",
            92 => x"81",
            93 => x"05",
            94 => x"74",
            95 => x"51",
            96 => x"81",
            97 => x"ff",
            98 => x"72",
            99 => x"51",
           100 => x"04",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"52",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"72",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"ff",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"8c",
           133 => x"04",
           134 => x"0b",
           135 => x"8c",
           136 => x"04",
           137 => x"0b",
           138 => x"8c",
           139 => x"04",
           140 => x"0b",
           141 => x"8d",
           142 => x"04",
           143 => x"0b",
           144 => x"8d",
           145 => x"04",
           146 => x"0b",
           147 => x"8e",
           148 => x"04",
           149 => x"0b",
           150 => x"8f",
           151 => x"04",
           152 => x"0b",
           153 => x"8f",
           154 => x"04",
           155 => x"0b",
           156 => x"90",
           157 => x"04",
           158 => x"0b",
           159 => x"90",
           160 => x"04",
           161 => x"0b",
           162 => x"91",
           163 => x"04",
           164 => x"0b",
           165 => x"91",
           166 => x"04",
           167 => x"0b",
           168 => x"92",
           169 => x"04",
           170 => x"0b",
           171 => x"92",
           172 => x"04",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"81",
           193 => x"97",
           194 => x"80",
           195 => x"ee",
           196 => x"80",
           197 => x"f3",
           198 => x"80",
           199 => x"e0",
           200 => x"80",
           201 => x"a3",
           202 => x"80",
           203 => x"f6",
           204 => x"80",
           205 => x"86",
           206 => x"80",
           207 => x"82",
           208 => x"80",
           209 => x"88",
           210 => x"80",
           211 => x"a8",
           212 => x"80",
           213 => x"d1",
           214 => x"80",
           215 => x"8a",
           216 => x"80",
           217 => x"d4",
           218 => x"c0",
           219 => x"80",
           220 => x"80",
           221 => x"0c",
           222 => x"08",
           223 => x"90",
           224 => x"90",
           225 => x"bb",
           226 => x"bb",
           227 => x"84",
           228 => x"84",
           229 => x"04",
           230 => x"2d",
           231 => x"90",
           232 => x"a5",
           233 => x"80",
           234 => x"ed",
           235 => x"c0",
           236 => x"82",
           237 => x"80",
           238 => x"0c",
           239 => x"08",
           240 => x"90",
           241 => x"90",
           242 => x"bb",
           243 => x"bb",
           244 => x"84",
           245 => x"84",
           246 => x"04",
           247 => x"2d",
           248 => x"90",
           249 => x"f6",
           250 => x"80",
           251 => x"8c",
           252 => x"c0",
           253 => x"82",
           254 => x"80",
           255 => x"0c",
           256 => x"08",
           257 => x"90",
           258 => x"90",
           259 => x"bb",
           260 => x"bb",
           261 => x"84",
           262 => x"84",
           263 => x"04",
           264 => x"2d",
           265 => x"90",
           266 => x"fe",
           267 => x"80",
           268 => x"97",
           269 => x"c0",
           270 => x"83",
           271 => x"80",
           272 => x"0c",
           273 => x"08",
           274 => x"90",
           275 => x"90",
           276 => x"bb",
           277 => x"bb",
           278 => x"84",
           279 => x"84",
           280 => x"04",
           281 => x"2d",
           282 => x"90",
           283 => x"ab",
           284 => x"80",
           285 => x"f6",
           286 => x"c0",
           287 => x"81",
           288 => x"80",
           289 => x"0c",
           290 => x"08",
           291 => x"90",
           292 => x"90",
           293 => x"bb",
           294 => x"bb",
           295 => x"84",
           296 => x"bb",
           297 => x"84",
           298 => x"84",
           299 => x"04",
           300 => x"2d",
           301 => x"90",
           302 => x"85",
           303 => x"80",
           304 => x"d6",
           305 => x"c0",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"00",
           311 => x"06",
           312 => x"10",
           313 => x"51",
           314 => x"ff",
           315 => x"52",
           316 => x"38",
           317 => x"84",
           318 => x"80",
           319 => x"0b",
           320 => x"80",
           321 => x"87",
           322 => x"56",
           323 => x"51",
           324 => x"fa",
           325 => x"33",
           326 => x"07",
           327 => x"72",
           328 => x"ff",
           329 => x"70",
           330 => x"56",
           331 => x"80",
           332 => x"3f",
           333 => x"84",
           334 => x"84",
           335 => x"ff",
           336 => x"72",
           337 => x"73",
           338 => x"76",
           339 => x"3d",
           340 => x"0c",
           341 => x"7d",
           342 => x"34",
           343 => x"88",
           344 => x"05",
           345 => x"74",
           346 => x"0d",
           347 => x"75",
           348 => x"f1",
           349 => x"5d",
           350 => x"33",
           351 => x"55",
           352 => x"09",
           353 => x"57",
           354 => x"1c",
           355 => x"2e",
           356 => x"89",
           357 => x"70",
           358 => x"78",
           359 => x"7a",
           360 => x"40",
           361 => x"82",
           362 => x"ff",
           363 => x"84",
           364 => x"7a",
           365 => x"79",
           366 => x"2c",
           367 => x"0a",
           368 => x"56",
           369 => x"73",
           370 => x"78",
           371 => x"38",
           372 => x"81",
           373 => x"5a",
           374 => x"fe",
           375 => x"76",
           376 => x"76",
           377 => x"83",
           378 => x"8a",
           379 => x"7e",
           380 => x"d8",
           381 => x"cb",
           382 => x"e0",
           383 => x"eb",
           384 => x"3f",
           385 => x"86",
           386 => x"fe",
           387 => x"05",
           388 => x"5e",
           389 => x"79",
           390 => x"bb",
           391 => x"84",
           392 => x"89",
           393 => x"b0",
           394 => x"40",
           395 => x"3f",
           396 => x"84",
           397 => x"31",
           398 => x"7e",
           399 => x"80",
           400 => x"2c",
           401 => x"06",
           402 => x"77",
           403 => x"05",
           404 => x"84",
           405 => x"53",
           406 => x"70",
           407 => x"9e",
           408 => x"06",
           409 => x"38",
           410 => x"2a",
           411 => x"81",
           412 => x"38",
           413 => x"2c",
           414 => x"73",
           415 => x"2a",
           416 => x"7a",
           417 => x"98",
           418 => x"73",
           419 => x"73",
           420 => x"06",
           421 => x"78",
           422 => x"05",
           423 => x"74",
           424 => x"88",
           425 => x"29",
           426 => x"5a",
           427 => x"74",
           428 => x"38",
           429 => x"ff",
           430 => x"55",
           431 => x"b0",
           432 => x"80",
           433 => x"98",
           434 => x"e5",
           435 => x"5c",
           436 => x"76",
           437 => x"80",
           438 => x"d3",
           439 => x"94",
           440 => x"70",
           441 => x"84",
           442 => x"38",
           443 => x"fc",
           444 => x"29",
           445 => x"5a",
           446 => x"38",
           447 => x"e2",
           448 => x"07",
           449 => x"38",
           450 => x"5b",
           451 => x"05",
           452 => x"5f",
           453 => x"7f",
           454 => x"06",
           455 => x"07",
           456 => x"80",
           457 => x"56",
           458 => x"81",
           459 => x"77",
           460 => x"80",
           461 => x"80",
           462 => x"a0",
           463 => x"1a",
           464 => x"79",
           465 => x"7c",
           466 => x"51",
           467 => x"70",
           468 => x"83",
           469 => x"52",
           470 => x"85",
           471 => x"06",
           472 => x"80",
           473 => x"2c",
           474 => x"2a",
           475 => x"fd",
           476 => x"84",
           477 => x"56",
           478 => x"83",
           479 => x"5e",
           480 => x"33",
           481 => x"ca",
           482 => x"33",
           483 => x"ba",
           484 => x"77",
           485 => x"82",
           486 => x"84",
           487 => x"78",
           488 => x"90",
           489 => x"c0",
           490 => x"be",
           491 => x"05",
           492 => x"41",
           493 => x"87",
           494 => x"ff",
           495 => x"54",
           496 => x"7c",
           497 => x"f7",
           498 => x"29",
           499 => x"5a",
           500 => x"38",
           501 => x"e2",
           502 => x"3f",
           503 => x"e3",
           504 => x"3f",
           505 => x"80",
           506 => x"75",
           507 => x"70",
           508 => x"5a",
           509 => x"a2",
           510 => x"3f",
           511 => x"fa",
           512 => x"75",
           513 => x"81",
           514 => x"38",
           515 => x"2b",
           516 => x"39",
           517 => x"c8",
           518 => x"3f",
           519 => x"88",
           520 => x"ff",
           521 => x"54",
           522 => x"7e",
           523 => x"57",
           524 => x"84",
           525 => x"51",
           526 => x"fa",
           527 => x"e6",
           528 => x"2a",
           529 => x"58",
           530 => x"09",
           531 => x"81",
           532 => x"b0",
           533 => x"51",
           534 => x"bb",
           535 => x"57",
           536 => x"72",
           537 => x"08",
           538 => x"54",
           539 => x"90",
           540 => x"84",
           541 => x"76",
           542 => x"3d",
           543 => x"56",
           544 => x"81",
           545 => x"55",
           546 => x"09",
           547 => x"05",
           548 => x"81",
           549 => x"bb",
           550 => x"70",
           551 => x"2e",
           552 => x"15",
           553 => x"08",
           554 => x"81",
           555 => x"38",
           556 => x"e8",
           557 => x"3d",
           558 => x"85",
           559 => x"81",
           560 => x"72",
           561 => x"54",
           562 => x"08",
           563 => x"38",
           564 => x"08",
           565 => x"53",
           566 => x"75",
           567 => x"04",
           568 => x"90",
           569 => x"84",
           570 => x"08",
           571 => x"d7",
           572 => x"33",
           573 => x"81",
           574 => x"71",
           575 => x"52",
           576 => x"06",
           577 => x"75",
           578 => x"2e",
           579 => x"8c",
           580 => x"71",
           581 => x"84",
           582 => x"bf",
           583 => x"16",
           584 => x"16",
           585 => x"0d",
           586 => x"74",
           587 => x"bb",
           588 => x"85",
           589 => x"84",
           590 => x"71",
           591 => x"ff",
           592 => x"3d",
           593 => x"85",
           594 => x"3d",
           595 => x"71",
           596 => x"f7",
           597 => x"05",
           598 => x"05",
           599 => x"bb",
           600 => x"3d",
           601 => x"52",
           602 => x"72",
           603 => x"38",
           604 => x"70",
           605 => x"70",
           606 => x"86",
           607 => x"75",
           608 => x"53",
           609 => x"33",
           610 => x"2e",
           611 => x"53",
           612 => x"70",
           613 => x"74",
           614 => x"53",
           615 => x"70",
           616 => x"84",
           617 => x"77",
           618 => x"05",
           619 => x"05",
           620 => x"bb",
           621 => x"3d",
           622 => x"52",
           623 => x"70",
           624 => x"05",
           625 => x"38",
           626 => x"0d",
           627 => x"55",
           628 => x"73",
           629 => x"52",
           630 => x"9a",
           631 => x"b7",
           632 => x"80",
           633 => x"3d",
           634 => x"73",
           635 => x"e9",
           636 => x"71",
           637 => x"84",
           638 => x"71",
           639 => x"04",
           640 => x"52",
           641 => x"08",
           642 => x"55",
           643 => x"08",
           644 => x"9b",
           645 => x"80",
           646 => x"bb",
           647 => x"bb",
           648 => x"0c",
           649 => x"75",
           650 => x"71",
           651 => x"05",
           652 => x"38",
           653 => x"81",
           654 => x"31",
           655 => x"85",
           656 => x"77",
           657 => x"80",
           658 => x"05",
           659 => x"38",
           660 => x"0d",
           661 => x"54",
           662 => x"76",
           663 => x"08",
           664 => x"8d",
           665 => x"84",
           666 => x"72",
           667 => x"72",
           668 => x"74",
           669 => x"2b",
           670 => x"76",
           671 => x"2a",
           672 => x"31",
           673 => x"7b",
           674 => x"5c",
           675 => x"74",
           676 => x"71",
           677 => x"04",
           678 => x"80",
           679 => x"25",
           680 => x"71",
           681 => x"30",
           682 => x"31",
           683 => x"70",
           684 => x"71",
           685 => x"1b",
           686 => x"80",
           687 => x"2a",
           688 => x"06",
           689 => x"19",
           690 => x"54",
           691 => x"55",
           692 => x"58",
           693 => x"fd",
           694 => x"53",
           695 => x"84",
           696 => x"bb",
           697 => x"fa",
           698 => x"53",
           699 => x"fe",
           700 => x"e0",
           701 => x"73",
           702 => x"84",
           703 => x"26",
           704 => x"2e",
           705 => x"a0",
           706 => x"54",
           707 => x"38",
           708 => x"10",
           709 => x"9f",
           710 => x"75",
           711 => x"52",
           712 => x"72",
           713 => x"04",
           714 => x"9f",
           715 => x"9f",
           716 => x"74",
           717 => x"56",
           718 => x"bb",
           719 => x"bb",
           720 => x"3d",
           721 => x"7b",
           722 => x"59",
           723 => x"38",
           724 => x"55",
           725 => x"ad",
           726 => x"81",
           727 => x"77",
           728 => x"80",
           729 => x"80",
           730 => x"70",
           731 => x"70",
           732 => x"27",
           733 => x"06",
           734 => x"38",
           735 => x"76",
           736 => x"70",
           737 => x"ff",
           738 => x"75",
           739 => x"75",
           740 => x"04",
           741 => x"33",
           742 => x"81",
           743 => x"78",
           744 => x"e2",
           745 => x"f8",
           746 => x"27",
           747 => x"88",
           748 => x"75",
           749 => x"04",
           750 => x"70",
           751 => x"39",
           752 => x"3d",
           753 => x"5b",
           754 => x"70",
           755 => x"09",
           756 => x"78",
           757 => x"2e",
           758 => x"38",
           759 => x"14",
           760 => x"db",
           761 => x"27",
           762 => x"89",
           763 => x"55",
           764 => x"51",
           765 => x"13",
           766 => x"73",
           767 => x"81",
           768 => x"16",
           769 => x"56",
           770 => x"80",
           771 => x"7a",
           772 => x"0c",
           773 => x"70",
           774 => x"73",
           775 => x"38",
           776 => x"55",
           777 => x"90",
           778 => x"81",
           779 => x"14",
           780 => x"27",
           781 => x"0c",
           782 => x"15",
           783 => x"80",
           784 => x"bb",
           785 => x"d8",
           786 => x"ff",
           787 => x"3d",
           788 => x"38",
           789 => x"52",
           790 => x"ef",
           791 => x"cf",
           792 => x"0d",
           793 => x"3f",
           794 => x"51",
           795 => x"83",
           796 => x"3d",
           797 => x"87",
           798 => x"b4",
           799 => x"04",
           800 => x"83",
           801 => x"ee",
           802 => x"d1",
           803 => x"0d",
           804 => x"3f",
           805 => x"51",
           806 => x"83",
           807 => x"3d",
           808 => x"af",
           809 => x"f4",
           810 => x"04",
           811 => x"83",
           812 => x"ee",
           813 => x"d2",
           814 => x"0d",
           815 => x"3f",
           816 => x"51",
           817 => x"83",
           818 => x"3d",
           819 => x"97",
           820 => x"05",
           821 => x"3d",
           822 => x"25",
           823 => x"87",
           824 => x"77",
           825 => x"93",
           826 => x"77",
           827 => x"97",
           828 => x"84",
           829 => x"38",
           830 => x"30",
           831 => x"70",
           832 => x"58",
           833 => x"98",
           834 => x"80",
           835 => x"29",
           836 => x"08",
           837 => x"83",
           838 => x"84",
           839 => x"04",
           840 => x"88",
           841 => x"96",
           842 => x"53",
           843 => x"3f",
           844 => x"84",
           845 => x"80",
           846 => x"17",
           847 => x"74",
           848 => x"08",
           849 => x"bb",
           850 => x"78",
           851 => x"3f",
           852 => x"02",
           853 => x"ff",
           854 => x"fd",
           855 => x"38",
           856 => x"2e",
           857 => x"8a",
           858 => x"e4",
           859 => x"84",
           860 => x"84",
           861 => x"8a",
           862 => x"61",
           863 => x"33",
           864 => x"5c",
           865 => x"82",
           866 => x"dd",
           867 => x"ec",
           868 => x"38",
           869 => x"a0",
           870 => x"72",
           871 => x"52",
           872 => x"81",
           873 => x"a0",
           874 => x"dc",
           875 => x"3f",
           876 => x"38",
           877 => x"55",
           878 => x"80",
           879 => x"53",
           880 => x"56",
           881 => x"fe",
           882 => x"e8",
           883 => x"81",
           884 => x"83",
           885 => x"18",
           886 => x"c8",
           887 => x"70",
           888 => x"81",
           889 => x"38",
           890 => x"b9",
           891 => x"8f",
           892 => x"dc",
           893 => x"08",
           894 => x"78",
           895 => x"39",
           896 => x"82",
           897 => x"a0",
           898 => x"fe",
           899 => x"27",
           900 => x"ac",
           901 => x"e6",
           902 => x"ba",
           903 => x"99",
           904 => x"3f",
           905 => x"54",
           906 => x"27",
           907 => x"7a",
           908 => x"d3",
           909 => x"84",
           910 => x"e9",
           911 => x"fd",
           912 => x"73",
           913 => x"fe",
           914 => x"bb",
           915 => x"59",
           916 => x"59",
           917 => x"fc",
           918 => x"80",
           919 => x"08",
           920 => x"32",
           921 => x"70",
           922 => x"55",
           923 => x"25",
           924 => x"3f",
           925 => x"98",
           926 => x"9b",
           927 => x"75",
           928 => x"58",
           929 => x"fd",
           930 => x"0c",
           931 => x"87",
           932 => x"3f",
           933 => x"d0",
           934 => x"81",
           935 => x"51",
           936 => x"2a",
           937 => x"89",
           938 => x"51",
           939 => x"2a",
           940 => x"ad",
           941 => x"51",
           942 => x"2a",
           943 => x"d2",
           944 => x"51",
           945 => x"81",
           946 => x"3f",
           947 => x"99",
           948 => x"3f",
           949 => x"3f",
           950 => x"81",
           951 => x"3f",
           952 => x"2a",
           953 => x"38",
           954 => x"83",
           955 => x"51",
           956 => x"81",
           957 => x"9c",
           958 => x"3f",
           959 => x"80",
           960 => x"70",
           961 => x"fe",
           962 => x"9b",
           963 => x"b1",
           964 => x"85",
           965 => x"80",
           966 => x"81",
           967 => x"51",
           968 => x"3f",
           969 => x"52",
           970 => x"bd",
           971 => x"d5",
           972 => x"9a",
           973 => x"06",
           974 => x"38",
           975 => x"3f",
           976 => x"80",
           977 => x"70",
           978 => x"fd",
           979 => x"0d",
           980 => x"de",
           981 => x"81",
           982 => x"81",
           983 => x"61",
           984 => x"51",
           985 => x"d6",
           986 => x"80",
           987 => x"a3",
           988 => x"70",
           989 => x"2e",
           990 => x"88",
           991 => x"82",
           992 => x"5a",
           993 => x"33",
           994 => x"8c",
           995 => x"7b",
           996 => x"9b",
           997 => x"ef",
           998 => x"f4",
           999 => x"84",
          1000 => x"5d",
          1001 => x"8b",
          1002 => x"2e",
          1003 => x"ff",
          1004 => x"38",
          1005 => x"fe",
          1006 => x"e9",
          1007 => x"84",
          1008 => x"38",
          1009 => x"ff",
          1010 => x"bb",
          1011 => x"7a",
          1012 => x"84",
          1013 => x"84",
          1014 => x"0b",
          1015 => x"8d",
          1016 => x"38",
          1017 => x"54",
          1018 => x"51",
          1019 => x"84",
          1020 => x"80",
          1021 => x"0a",
          1022 => x"bb",
          1023 => x"70",
          1024 => x"5b",
          1025 => x"83",
          1026 => x"78",
          1027 => x"81",
          1028 => x"38",
          1029 => x"5d",
          1030 => x"81",
          1031 => x"3f",
          1032 => x"7e",
          1033 => x"51",
          1034 => x"f8",
          1035 => x"79",
          1036 => x"a8",
          1037 => x"8a",
          1038 => x"38",
          1039 => x"34",
          1040 => x"7e",
          1041 => x"84",
          1042 => x"84",
          1043 => x"83",
          1044 => x"5f",
          1045 => x"fc",
          1046 => x"51",
          1047 => x"0b",
          1048 => x"d6",
          1049 => x"7e",
          1050 => x"5a",
          1051 => x"1a",
          1052 => x"81",
          1053 => x"10",
          1054 => x"04",
          1055 => x"51",
          1056 => x"84",
          1057 => x"84",
          1058 => x"06",
          1059 => x"45",
          1060 => x"8c",
          1061 => x"94",
          1062 => x"9c",
          1063 => x"80",
          1064 => x"d2",
          1065 => x"e4",
          1066 => x"fa",
          1067 => x"c0",
          1068 => x"8e",
          1069 => x"51",
          1070 => x"83",
          1071 => x"ed",
          1072 => x"84",
          1073 => x"fa",
          1074 => x"fa",
          1075 => x"51",
          1076 => x"84",
          1077 => x"38",
          1078 => x"80",
          1079 => x"b8",
          1080 => x"05",
          1081 => x"08",
          1082 => x"83",
          1083 => x"59",
          1084 => x"53",
          1085 => x"84",
          1086 => x"38",
          1087 => x"80",
          1088 => x"84",
          1089 => x"08",
          1090 => x"cf",
          1091 => x"80",
          1092 => x"7e",
          1093 => x"f9",
          1094 => x"38",
          1095 => x"39",
          1096 => x"80",
          1097 => x"84",
          1098 => x"3d",
          1099 => x"51",
          1100 => x"86",
          1101 => x"78",
          1102 => x"3f",
          1103 => x"52",
          1104 => x"7e",
          1105 => x"38",
          1106 => x"82",
          1107 => x"3d",
          1108 => x"51",
          1109 => x"80",
          1110 => x"fc",
          1111 => x"ca",
          1112 => x"f8",
          1113 => x"53",
          1114 => x"84",
          1115 => x"38",
          1116 => x"68",
          1117 => x"8d",
          1118 => x"5c",
          1119 => x"55",
          1120 => x"83",
          1121 => x"66",
          1122 => x"59",
          1123 => x"53",
          1124 => x"84",
          1125 => x"38",
          1126 => x"80",
          1127 => x"84",
          1128 => x"3d",
          1129 => x"51",
          1130 => x"80",
          1131 => x"51",
          1132 => x"27",
          1133 => x"81",
          1134 => x"05",
          1135 => x"11",
          1136 => x"3f",
          1137 => x"be",
          1138 => x"ff",
          1139 => x"bb",
          1140 => x"54",
          1141 => x"3f",
          1142 => x"52",
          1143 => x"7e",
          1144 => x"38",
          1145 => x"81",
          1146 => x"80",
          1147 => x"05",
          1148 => x"ff",
          1149 => x"bb",
          1150 => x"68",
          1151 => x"34",
          1152 => x"fc",
          1153 => x"fa",
          1154 => x"38",
          1155 => x"11",
          1156 => x"3f",
          1157 => x"9e",
          1158 => x"ff",
          1159 => x"bb",
          1160 => x"b8",
          1161 => x"05",
          1162 => x"08",
          1163 => x"83",
          1164 => x"67",
          1165 => x"65",
          1166 => x"0c",
          1167 => x"d9",
          1168 => x"ff",
          1169 => x"bb",
          1170 => x"52",
          1171 => x"bb",
          1172 => x"3f",
          1173 => x"9e",
          1174 => x"e6",
          1175 => x"84",
          1176 => x"c2",
          1177 => x"83",
          1178 => x"83",
          1179 => x"b8",
          1180 => x"05",
          1181 => x"08",
          1182 => x"79",
          1183 => x"c4",
          1184 => x"53",
          1185 => x"84",
          1186 => x"80",
          1187 => x"38",
          1188 => x"70",
          1189 => x"5f",
          1190 => x"a0",
          1191 => x"a8",
          1192 => x"54",
          1193 => x"a3",
          1194 => x"3f",
          1195 => x"59",
          1196 => x"f0",
          1197 => x"96",
          1198 => x"f2",
          1199 => x"64",
          1200 => x"11",
          1201 => x"3f",
          1202 => x"b6",
          1203 => x"22",
          1204 => x"45",
          1205 => x"80",
          1206 => x"84",
          1207 => x"5e",
          1208 => x"82",
          1209 => x"fe",
          1210 => x"e1",
          1211 => x"b9",
          1212 => x"fc",
          1213 => x"9a",
          1214 => x"81",
          1215 => x"05",
          1216 => x"fb",
          1217 => x"53",
          1218 => x"84",
          1219 => x"38",
          1220 => x"05",
          1221 => x"83",
          1222 => x"7b",
          1223 => x"83",
          1224 => x"3f",
          1225 => x"d9",
          1226 => x"cc",
          1227 => x"b8",
          1228 => x"05",
          1229 => x"08",
          1230 => x"80",
          1231 => x"5b",
          1232 => x"f4",
          1233 => x"cf",
          1234 => x"ea",
          1235 => x"80",
          1236 => x"49",
          1237 => x"d3",
          1238 => x"83",
          1239 => x"59",
          1240 => x"59",
          1241 => x"d0",
          1242 => x"f8",
          1243 => x"83",
          1244 => x"9b",
          1245 => x"92",
          1246 => x"80",
          1247 => x"49",
          1248 => x"5e",
          1249 => x"dc",
          1250 => x"86",
          1251 => x"83",
          1252 => x"83",
          1253 => x"94",
          1254 => x"ca",
          1255 => x"05",
          1256 => x"08",
          1257 => x"3d",
          1258 => x"87",
          1259 => x"87",
          1260 => x"3f",
          1261 => x"08",
          1262 => x"51",
          1263 => x"08",
          1264 => x"70",
          1265 => x"74",
          1266 => x"08",
          1267 => x"84",
          1268 => x"74",
          1269 => x"8c",
          1270 => x"0c",
          1271 => x"94",
          1272 => x"b9",
          1273 => x"34",
          1274 => x"3d",
          1275 => x"84",
          1276 => x"89",
          1277 => x"51",
          1278 => x"83",
          1279 => x"f3",
          1280 => x"3f",
          1281 => x"53",
          1282 => x"51",
          1283 => x"d3",
          1284 => x"83",
          1285 => x"80",
          1286 => x"d4",
          1287 => x"3d",
          1288 => x"75",
          1289 => x"38",
          1290 => x"52",
          1291 => x"38",
          1292 => x"06",
          1293 => x"38",
          1294 => x"2e",
          1295 => x"2e",
          1296 => x"81",
          1297 => x"2e",
          1298 => x"8b",
          1299 => x"12",
          1300 => x"06",
          1301 => x"06",
          1302 => x"70",
          1303 => x"52",
          1304 => x"72",
          1305 => x"0c",
          1306 => x"87",
          1307 => x"38",
          1308 => x"12",
          1309 => x"06",
          1310 => x"38",
          1311 => x"81",
          1312 => x"81",
          1313 => x"3d",
          1314 => x"80",
          1315 => x"0d",
          1316 => x"51",
          1317 => x"80",
          1318 => x"0c",
          1319 => x"76",
          1320 => x"81",
          1321 => x"83",
          1322 => x"73",
          1323 => x"33",
          1324 => x"fe",
          1325 => x"73",
          1326 => x"33",
          1327 => x"e6",
          1328 => x"74",
          1329 => x"13",
          1330 => x"26",
          1331 => x"98",
          1332 => x"bc",
          1333 => x"b8",
          1334 => x"b4",
          1335 => x"b0",
          1336 => x"ac",
          1337 => x"a8",
          1338 => x"73",
          1339 => x"87",
          1340 => x"84",
          1341 => x"f3",
          1342 => x"9c",
          1343 => x"bc",
          1344 => x"98",
          1345 => x"87",
          1346 => x"1c",
          1347 => x"7b",
          1348 => x"08",
          1349 => x"98",
          1350 => x"87",
          1351 => x"1c",
          1352 => x"79",
          1353 => x"83",
          1354 => x"ff",
          1355 => x"1b",
          1356 => x"1b",
          1357 => x"83",
          1358 => x"51",
          1359 => x"04",
          1360 => x"53",
          1361 => x"80",
          1362 => x"98",
          1363 => x"ff",
          1364 => x"83",
          1365 => x"0c",
          1366 => x"e9",
          1367 => x"2b",
          1368 => x"2e",
          1369 => x"80",
          1370 => x"98",
          1371 => x"ff",
          1372 => x"0d",
          1373 => x"54",
          1374 => x"bb",
          1375 => x"51",
          1376 => x"72",
          1377 => x"25",
          1378 => x"85",
          1379 => x"9b",
          1380 => x"81",
          1381 => x"2e",
          1382 => x"08",
          1383 => x"54",
          1384 => x"91",
          1385 => x"e3",
          1386 => x"72",
          1387 => x"81",
          1388 => x"ff",
          1389 => x"70",
          1390 => x"90",
          1391 => x"84",
          1392 => x"2a",
          1393 => x"38",
          1394 => x"80",
          1395 => x"06",
          1396 => x"c0",
          1397 => x"81",
          1398 => x"d8",
          1399 => x"33",
          1400 => x"52",
          1401 => x"0d",
          1402 => x"75",
          1403 => x"2e",
          1404 => x"bc",
          1405 => x"55",
          1406 => x"c0",
          1407 => x"81",
          1408 => x"8c",
          1409 => x"51",
          1410 => x"81",
          1411 => x"71",
          1412 => x"38",
          1413 => x"94",
          1414 => x"87",
          1415 => x"81",
          1416 => x"9b",
          1417 => x"3d",
          1418 => x"06",
          1419 => x"32",
          1420 => x"38",
          1421 => x"80",
          1422 => x"84",
          1423 => x"53",
          1424 => x"ff",
          1425 => x"70",
          1426 => x"80",
          1427 => x"a4",
          1428 => x"9e",
          1429 => x"c0",
          1430 => x"87",
          1431 => x"0c",
          1432 => x"d0",
          1433 => x"f3",
          1434 => x"83",
          1435 => x"08",
          1436 => x"b4",
          1437 => x"9e",
          1438 => x"c0",
          1439 => x"87",
          1440 => x"0c",
          1441 => x"f0",
          1442 => x"71",
          1443 => x"84",
          1444 => x"9e",
          1445 => x"c0",
          1446 => x"81",
          1447 => x"87",
          1448 => x"0a",
          1449 => x"38",
          1450 => x"87",
          1451 => x"0a",
          1452 => x"83",
          1453 => x"34",
          1454 => x"70",
          1455 => x"70",
          1456 => x"83",
          1457 => x"9e",
          1458 => x"51",
          1459 => x"81",
          1460 => x"0b",
          1461 => x"80",
          1462 => x"2e",
          1463 => x"89",
          1464 => x"08",
          1465 => x"52",
          1466 => x"71",
          1467 => x"c0",
          1468 => x"06",
          1469 => x"38",
          1470 => x"80",
          1471 => x"82",
          1472 => x"80",
          1473 => x"f4",
          1474 => x"90",
          1475 => x"52",
          1476 => x"52",
          1477 => x"87",
          1478 => x"80",
          1479 => x"83",
          1480 => x"34",
          1481 => x"70",
          1482 => x"80",
          1483 => x"f4",
          1484 => x"98",
          1485 => x"71",
          1486 => x"c0",
          1487 => x"51",
          1488 => x"81",
          1489 => x"c0",
          1490 => x"84",
          1491 => x"34",
          1492 => x"70",
          1493 => x"2e",
          1494 => x"93",
          1495 => x"06",
          1496 => x"3d",
          1497 => x"fb",
          1498 => x"b6",
          1499 => x"73",
          1500 => x"c3",
          1501 => x"74",
          1502 => x"54",
          1503 => x"33",
          1504 => x"89",
          1505 => x"f4",
          1506 => x"83",
          1507 => x"38",
          1508 => x"86",
          1509 => x"83",
          1510 => x"75",
          1511 => x"54",
          1512 => x"33",
          1513 => x"8d",
          1514 => x"f4",
          1515 => x"83",
          1516 => x"f3",
          1517 => x"ff",
          1518 => x"52",
          1519 => x"3f",
          1520 => x"9c",
          1521 => x"c4",
          1522 => x"22",
          1523 => x"ec",
          1524 => x"84",
          1525 => x"84",
          1526 => x"76",
          1527 => x"08",
          1528 => x"c4",
          1529 => x"b9",
          1530 => x"85",
          1531 => x"80",
          1532 => x"51",
          1533 => x"bd",
          1534 => x"54",
          1535 => x"a0",
          1536 => x"0d",
          1537 => x"84",
          1538 => x"84",
          1539 => x"76",
          1540 => x"08",
          1541 => x"dc",
          1542 => x"80",
          1543 => x"83",
          1544 => x"da",
          1545 => x"e8",
          1546 => x"b3",
          1547 => x"83",
          1548 => x"83",
          1549 => x"51",
          1550 => x"51",
          1551 => x"22",
          1552 => x"84",
          1553 => x"84",
          1554 => x"84",
          1555 => x"76",
          1556 => x"08",
          1557 => x"dc",
          1558 => x"80",
          1559 => x"83",
          1560 => x"83",
          1561 => x"fd",
          1562 => x"88",
          1563 => x"8d",
          1564 => x"38",
          1565 => x"bf",
          1566 => x"74",
          1567 => x"83",
          1568 => x"83",
          1569 => x"fc",
          1570 => x"33",
          1571 => x"ec",
          1572 => x"80",
          1573 => x"f4",
          1574 => x"ff",
          1575 => x"55",
          1576 => x"39",
          1577 => x"f4",
          1578 => x"93",
          1579 => x"38",
          1580 => x"f3",
          1581 => x"94",
          1582 => x"8f",
          1583 => x"38",
          1584 => x"f3",
          1585 => x"b0",
          1586 => x"8a",
          1587 => x"38",
          1588 => x"f3",
          1589 => x"cc",
          1590 => x"89",
          1591 => x"38",
          1592 => x"f3",
          1593 => x"e8",
          1594 => x"88",
          1595 => x"38",
          1596 => x"f3",
          1597 => x"84",
          1598 => x"8b",
          1599 => x"38",
          1600 => x"b0",
          1601 => x"bc",
          1602 => x"74",
          1603 => x"ff",
          1604 => x"71",
          1605 => x"83",
          1606 => x"83",
          1607 => x"83",
          1608 => x"ff",
          1609 => x"83",
          1610 => x"83",
          1611 => x"ff",
          1612 => x"83",
          1613 => x"83",
          1614 => x"ff",
          1615 => x"71",
          1616 => x"c0",
          1617 => x"08",
          1618 => x"3d",
          1619 => x"5a",
          1620 => x"83",
          1621 => x"3f",
          1622 => x"8b",
          1623 => x"08",
          1624 => x"82",
          1625 => x"80",
          1626 => x"3f",
          1627 => x"55",
          1628 => x"8e",
          1629 => x"70",
          1630 => x"09",
          1631 => x"51",
          1632 => x"73",
          1633 => x"8c",
          1634 => x"3f",
          1635 => x"76",
          1636 => x"0c",
          1637 => x"51",
          1638 => x"09",
          1639 => x"51",
          1640 => x"e4",
          1641 => x"84",
          1642 => x"e4",
          1643 => x"84",
          1644 => x"d8",
          1645 => x"08",
          1646 => x"5a",
          1647 => x"80",
          1648 => x"10",
          1649 => x"52",
          1650 => x"84",
          1651 => x"ff",
          1652 => x"90",
          1653 => x"2e",
          1654 => x"38",
          1655 => x"54",
          1656 => x"73",
          1657 => x"04",
          1658 => x"11",
          1659 => x"3f",
          1660 => x"38",
          1661 => x"fd",
          1662 => x"ff",
          1663 => x"81",
          1664 => x"82",
          1665 => x"39",
          1666 => x"27",
          1667 => x"70",
          1668 => x"81",
          1669 => x"eb",
          1670 => x"fe",
          1671 => x"53",
          1672 => x"84",
          1673 => x"d0",
          1674 => x"f8",
          1675 => x"84",
          1676 => x"77",
          1677 => x"84",
          1678 => x"08",
          1679 => x"ff",
          1680 => x"34",
          1681 => x"e3",
          1682 => x"74",
          1683 => x"38",
          1684 => x"3d",
          1685 => x"08",
          1686 => x"3d",
          1687 => x"42",
          1688 => x"f4",
          1689 => x"34",
          1690 => x"38",
          1691 => x"74",
          1692 => x"2e",
          1693 => x"5a",
          1694 => x"2e",
          1695 => x"40",
          1696 => x"bb",
          1697 => x"5b",
          1698 => x"79",
          1699 => x"70",
          1700 => x"bc",
          1701 => x"71",
          1702 => x"df",
          1703 => x"51",
          1704 => x"5c",
          1705 => x"cd",
          1706 => x"75",
          1707 => x"05",
          1708 => x"24",
          1709 => x"82",
          1710 => x"e4",
          1711 => x"91",
          1712 => x"70",
          1713 => x"b6",
          1714 => x"84",
          1715 => x"2e",
          1716 => x"2b",
          1717 => x"70",
          1718 => x"2c",
          1719 => x"11",
          1720 => x"57",
          1721 => x"76",
          1722 => x"a8",
          1723 => x"70",
          1724 => x"09",
          1725 => x"2e",
          1726 => x"39",
          1727 => x"81",
          1728 => x"70",
          1729 => x"57",
          1730 => x"75",
          1731 => x"80",
          1732 => x"57",
          1733 => x"e0",
          1734 => x"78",
          1735 => x"2e",
          1736 => x"57",
          1737 => x"c6",
          1738 => x"57",
          1739 => x"c0",
          1740 => x"7f",
          1741 => x"95",
          1742 => x"83",
          1743 => x"83",
          1744 => x"0b",
          1745 => x"e2",
          1746 => x"33",
          1747 => x"84",
          1748 => x"b5",
          1749 => x"05",
          1750 => x"c9",
          1751 => x"ff",
          1752 => x"55",
          1753 => x"e6",
          1754 => x"84",
          1755 => x"52",
          1756 => x"39",
          1757 => x"92",
          1758 => x"f4",
          1759 => x"8f",
          1760 => x"34",
          1761 => x"84",
          1762 => x"2e",
          1763 => x"88",
          1764 => x"e8",
          1765 => x"3f",
          1766 => x"ff",
          1767 => x"ff",
          1768 => x"78",
          1769 => x"7b",
          1770 => x"e2",
          1771 => x"38",
          1772 => x"f1",
          1773 => x"58",
          1774 => x"10",
          1775 => x"57",
          1776 => x"26",
          1777 => x"f4",
          1778 => x"80",
          1779 => x"b7",
          1780 => x"e2",
          1781 => x"ff",
          1782 => x"51",
          1783 => x"33",
          1784 => x"80",
          1785 => x"08",
          1786 => x"84",
          1787 => x"b3",
          1788 => x"88",
          1789 => x"c8",
          1790 => x"c8",
          1791 => x"39",
          1792 => x"06",
          1793 => x"75",
          1794 => x"e8",
          1795 => x"e2",
          1796 => x"55",
          1797 => x"33",
          1798 => x"33",
          1799 => x"c1",
          1800 => x"15",
          1801 => x"16",
          1802 => x"3f",
          1803 => x"06",
          1804 => x"77",
          1805 => x"39",
          1806 => x"33",
          1807 => x"38",
          1808 => x"34",
          1809 => x"81",
          1810 => x"24",
          1811 => x"52",
          1812 => x"e2",
          1813 => x"2c",
          1814 => x"56",
          1815 => x"e6",
          1816 => x"aa",
          1817 => x"80",
          1818 => x"c4",
          1819 => x"f8",
          1820 => x"88",
          1821 => x"80",
          1822 => x"98",
          1823 => x"59",
          1824 => x"f9",
          1825 => x"78",
          1826 => x"33",
          1827 => x"80",
          1828 => x"98",
          1829 => x"55",
          1830 => x"16",
          1831 => x"e6",
          1832 => x"b0",
          1833 => x"81",
          1834 => x"e2",
          1835 => x"24",
          1836 => x"e2",
          1837 => x"91",
          1838 => x"51",
          1839 => x"33",
          1840 => x"34",
          1841 => x"84",
          1842 => x"61",
          1843 => x"51",
          1844 => x"52",
          1845 => x"84",
          1846 => x"da",
          1847 => x"80",
          1848 => x"33",
          1849 => x"70",
          1850 => x"38",
          1851 => x"f4",
          1852 => x"59",
          1853 => x"08",
          1854 => x"10",
          1855 => x"54",
          1856 => x"a0",
          1857 => x"10",
          1858 => x"57",
          1859 => x"f4",
          1860 => x"38",
          1861 => x"2e",
          1862 => x"c8",
          1863 => x"7b",
          1864 => x"04",
          1865 => x"2e",
          1866 => x"88",
          1867 => x"e8",
          1868 => x"3f",
          1869 => x"ff",
          1870 => x"ff",
          1871 => x"61",
          1872 => x"83",
          1873 => x"80",
          1874 => x"84",
          1875 => x"e2",
          1876 => x"56",
          1877 => x"e2",
          1878 => x"e2",
          1879 => x"e2",
          1880 => x"88",
          1881 => x"c8",
          1882 => x"84",
          1883 => x"76",
          1884 => x"e8",
          1885 => x"3f",
          1886 => x"70",
          1887 => x"57",
          1888 => x"38",
          1889 => x"ff",
          1890 => x"29",
          1891 => x"84",
          1892 => x"7a",
          1893 => x"08",
          1894 => x"74",
          1895 => x"05",
          1896 => x"5c",
          1897 => x"38",
          1898 => x"17",
          1899 => x"52",
          1900 => x"75",
          1901 => x"05",
          1902 => x"44",
          1903 => x"38",
          1904 => x"34",
          1905 => x"51",
          1906 => x"0a",
          1907 => x"2c",
          1908 => x"61",
          1909 => x"39",
          1910 => x"34",
          1911 => x"2e",
          1912 => x"88",
          1913 => x"e8",
          1914 => x"3f",
          1915 => x"ff",
          1916 => x"ff",
          1917 => x"7c",
          1918 => x"83",
          1919 => x"80",
          1920 => x"84",
          1921 => x"0c",
          1922 => x"33",
          1923 => x"61",
          1924 => x"33",
          1925 => x"98",
          1926 => x"76",
          1927 => x"33",
          1928 => x"29",
          1929 => x"84",
          1930 => x"78",
          1931 => x"84",
          1932 => x"7c",
          1933 => x"84",
          1934 => x"8b",
          1935 => x"c4",
          1936 => x"70",
          1937 => x"05",
          1938 => x"45",
          1939 => x"90",
          1940 => x"78",
          1941 => x"79",
          1942 => x"08",
          1943 => x"75",
          1944 => x"05",
          1945 => x"57",
          1946 => x"38",
          1947 => x"ff",
          1948 => x"29",
          1949 => x"84",
          1950 => x"76",
          1951 => x"84",
          1952 => x"bb",
          1953 => x"bb",
          1954 => x"ff",
          1955 => x"55",
          1956 => x"f0",
          1957 => x"39",
          1958 => x"70",
          1959 => x"75",
          1960 => x"05",
          1961 => x"52",
          1962 => x"84",
          1963 => x"98",
          1964 => x"5b",
          1965 => x"fe",
          1966 => x"2e",
          1967 => x"93",
          1968 => x"ff",
          1969 => x"25",
          1970 => x"34",
          1971 => x"2e",
          1972 => x"e5",
          1973 => x"db",
          1974 => x"0c",
          1975 => x"c1",
          1976 => x"80",
          1977 => x"56",
          1978 => x"ba",
          1979 => x"84",
          1980 => x"84",
          1981 => x"05",
          1982 => x"f6",
          1983 => x"84",
          1984 => x"80",
          1985 => x"08",
          1986 => x"84",
          1987 => x"a6",
          1988 => x"88",
          1989 => x"c8",
          1990 => x"c8",
          1991 => x"39",
          1992 => x"bb",
          1993 => x"bb",
          1994 => x"53",
          1995 => x"3f",
          1996 => x"c8",
          1997 => x"f1",
          1998 => x"88",
          1999 => x"e8",
          2000 => x"3f",
          2001 => x"ff",
          2002 => x"ff",
          2003 => x"76",
          2004 => x"51",
          2005 => x"08",
          2006 => x"08",
          2007 => x"52",
          2008 => x"1d",
          2009 => x"33",
          2010 => x"56",
          2011 => x"e6",
          2012 => x"8a",
          2013 => x"51",
          2014 => x"08",
          2015 => x"84",
          2016 => x"84",
          2017 => x"55",
          2018 => x"84",
          2019 => x"c4",
          2020 => x"3d",
          2021 => x"75",
          2022 => x"ff",
          2023 => x"84",
          2024 => x"81",
          2025 => x"7b",
          2026 => x"c4",
          2027 => x"74",
          2028 => x"e8",
          2029 => x"3f",
          2030 => x"ff",
          2031 => x"52",
          2032 => x"e2",
          2033 => x"e2",
          2034 => x"c7",
          2035 => x"83",
          2036 => x"fc",
          2037 => x"70",
          2038 => x"3f",
          2039 => x"f4",
          2040 => x"9c",
          2041 => x"94",
          2042 => x"f4",
          2043 => x"9c",
          2044 => x"80",
          2045 => x"52",
          2046 => x"f4",
          2047 => x"06",
          2048 => x"38",
          2049 => x"39",
          2050 => x"53",
          2051 => x"3f",
          2052 => x"82",
          2053 => x"51",
          2054 => x"e2",
          2055 => x"34",
          2056 => x"0d",
          2057 => x"81",
          2058 => x"82",
          2059 => x"3d",
          2060 => x"80",
          2061 => x"3f",
          2062 => x"84",
          2063 => x"f5",
          2064 => x"a5",
          2065 => x"80",
          2066 => x"fb",
          2067 => x"70",
          2068 => x"81",
          2069 => x"10",
          2070 => x"58",
          2071 => x"75",
          2072 => x"9c",
          2073 => x"80",
          2074 => x"7f",
          2075 => x"10",
          2076 => x"56",
          2077 => x"9c",
          2078 => x"10",
          2079 => x"41",
          2080 => x"81",
          2081 => x"83",
          2082 => x"81",
          2083 => x"38",
          2084 => x"74",
          2085 => x"f4",
          2086 => x"5b",
          2087 => x"80",
          2088 => x"39",
          2089 => x"f4",
          2090 => x"06",
          2091 => x"54",
          2092 => x"84",
          2093 => x"f4",
          2094 => x"05",
          2095 => x"52",
          2096 => x"f4",
          2097 => x"05",
          2098 => x"2e",
          2099 => x"83",
          2100 => x"83",
          2101 => x"e2",
          2102 => x"e6",
          2103 => x"0d",
          2104 => x"05",
          2105 => x"83",
          2106 => x"81",
          2107 => x"38",
          2108 => x"c7",
          2109 => x"70",
          2110 => x"79",
          2111 => x"b4",
          2112 => x"83",
          2113 => x"70",
          2114 => x"88",
          2115 => x"56",
          2116 => x"80",
          2117 => x"73",
          2118 => x"26",
          2119 => x"83",
          2120 => x"79",
          2121 => x"e0",
          2122 => x"05",
          2123 => x"38",
          2124 => x"80",
          2125 => x"10",
          2126 => x"29",
          2127 => x"59",
          2128 => x"f8",
          2129 => x"f7",
          2130 => x"b2",
          2131 => x"75",
          2132 => x"5b",
          2133 => x"74",
          2134 => x"06",
          2135 => x"06",
          2136 => x"ff",
          2137 => x"57",
          2138 => x"38",
          2139 => x"05",
          2140 => x"83",
          2141 => x"38",
          2142 => x"fe",
          2143 => x"55",
          2144 => x"81",
          2145 => x"a0",
          2146 => x"84",
          2147 => x"84",
          2148 => x"83",
          2149 => x"5b",
          2150 => x"78",
          2151 => x"06",
          2152 => x"18",
          2153 => x"bb",
          2154 => x"80",
          2155 => x"b0",
          2156 => x"07",
          2157 => x"7f",
          2158 => x"fd",
          2159 => x"e6",
          2160 => x"ff",
          2161 => x"b5",
          2162 => x"a0",
          2163 => x"5f",
          2164 => x"b8",
          2165 => x"b8",
          2166 => x"fa",
          2167 => x"7c",
          2168 => x"5f",
          2169 => x"26",
          2170 => x"7d",
          2171 => x"06",
          2172 => x"7d",
          2173 => x"06",
          2174 => x"5d",
          2175 => x"75",
          2176 => x"83",
          2177 => x"76",
          2178 => x"fb",
          2179 => x"56",
          2180 => x"8e",
          2181 => x"87",
          2182 => x"34",
          2183 => x"75",
          2184 => x"80",
          2185 => x"34",
          2186 => x"34",
          2187 => x"81",
          2188 => x"c0",
          2189 => x"f8",
          2190 => x"06",
          2191 => x"73",
          2192 => x"07",
          2193 => x"87",
          2194 => x"51",
          2195 => x"73",
          2196 => x"72",
          2197 => x"f8",
          2198 => x"87",
          2199 => x"84",
          2200 => x"02",
          2201 => x"05",
          2202 => x"56",
          2203 => x"38",
          2204 => x"33",
          2205 => x"12",
          2206 => x"b2",
          2207 => x"29",
          2208 => x"f9",
          2209 => x"81",
          2210 => x"22",
          2211 => x"23",
          2212 => x"81",
          2213 => x"5b",
          2214 => x"ff",
          2215 => x"83",
          2216 => x"06",
          2217 => x"79",
          2218 => x"f8",
          2219 => x"54",
          2220 => x"99",
          2221 => x"13",
          2222 => x"81",
          2223 => x"57",
          2224 => x"73",
          2225 => x"a1",
          2226 => x"d6",
          2227 => x"14",
          2228 => x"34",
          2229 => x"eb",
          2230 => x"56",
          2231 => x"78",
          2232 => x"06",
          2233 => x"38",
          2234 => x"f8",
          2235 => x"75",
          2236 => x"c7",
          2237 => x"81",
          2238 => x"5c",
          2239 => x"84",
          2240 => x"33",
          2241 => x"70",
          2242 => x"05",
          2243 => x"34",
          2244 => x"b8",
          2245 => x"5c",
          2246 => x"80",
          2247 => x"3d",
          2248 => x"83",
          2249 => x"06",
          2250 => x"73",
          2251 => x"2e",
          2252 => x"ff",
          2253 => x"72",
          2254 => x"38",
          2255 => x"f8",
          2256 => x"11",
          2257 => x"fe",
          2258 => x"99",
          2259 => x"56",
          2260 => x"75",
          2261 => x"53",
          2262 => x"0b",
          2263 => x"81",
          2264 => x"d8",
          2265 => x"b8",
          2266 => x"83",
          2267 => x"80",
          2268 => x"33",
          2269 => x"76",
          2270 => x"51",
          2271 => x"10",
          2272 => x"04",
          2273 => x"27",
          2274 => x"80",
          2275 => x"0d",
          2276 => x"83",
          2277 => x"54",
          2278 => x"12",
          2279 => x"0b",
          2280 => x"04",
          2281 => x"70",
          2282 => x"55",
          2283 => x"de",
          2284 => x"84",
          2285 => x"51",
          2286 => x"72",
          2287 => x"bb",
          2288 => x"fa",
          2289 => x"70",
          2290 => x"55",
          2291 => x"84",
          2292 => x"83",
          2293 => x"f8",
          2294 => x"74",
          2295 => x"fa",
          2296 => x"0c",
          2297 => x"fa",
          2298 => x"b8",
          2299 => x"75",
          2300 => x"70",
          2301 => x"ff",
          2302 => x"70",
          2303 => x"83",
          2304 => x"83",
          2305 => x"71",
          2306 => x"84",
          2307 => x"80",
          2308 => x"80",
          2309 => x"0b",
          2310 => x"04",
          2311 => x"90",
          2312 => x"80",
          2313 => x"0d",
          2314 => x"07",
          2315 => x"39",
          2316 => x"86",
          2317 => x"d7",
          2318 => x"34",
          2319 => x"3d",
          2320 => x"fc",
          2321 => x"b0",
          2322 => x"33",
          2323 => x"34",
          2324 => x"81",
          2325 => x"fa",
          2326 => x"b0",
          2327 => x"70",
          2328 => x"83",
          2329 => x"07",
          2330 => x"ef",
          2331 => x"06",
          2332 => x"df",
          2333 => x"06",
          2334 => x"b0",
          2335 => x"33",
          2336 => x"83",
          2337 => x"fa",
          2338 => x"07",
          2339 => x"a7",
          2340 => x"06",
          2341 => x"b0",
          2342 => x"33",
          2343 => x"83",
          2344 => x"fa",
          2345 => x"83",
          2346 => x"fa",
          2347 => x"51",
          2348 => x"39",
          2349 => x"02",
          2350 => x"fa",
          2351 => x"fa",
          2352 => x"41",
          2353 => x"82",
          2354 => x"78",
          2355 => x"b8",
          2356 => x"34",
          2357 => x"fa",
          2358 => x"8f",
          2359 => x"81",
          2360 => x"fa",
          2361 => x"82",
          2362 => x"83",
          2363 => x"b2",
          2364 => x"57",
          2365 => x"f6",
          2366 => x"52",
          2367 => x"3f",
          2368 => x"84",
          2369 => x"34",
          2370 => x"fa",
          2371 => x"0b",
          2372 => x"b8",
          2373 => x"34",
          2374 => x"0b",
          2375 => x"33",
          2376 => x"ba",
          2377 => x"7c",
          2378 => x"fe",
          2379 => x"85",
          2380 => x"38",
          2381 => x"22",
          2382 => x"ff",
          2383 => x"06",
          2384 => x"78",
          2385 => x"51",
          2386 => x"fa",
          2387 => x"7a",
          2388 => x"b2",
          2389 => x"3d",
          2390 => x"34",
          2391 => x"0b",
          2392 => x"fa",
          2393 => x"23",
          2394 => x"3f",
          2395 => x"b0",
          2396 => x"83",
          2397 => x"78",
          2398 => x"38",
          2399 => x"e5",
          2400 => x"19",
          2401 => x"39",
          2402 => x"a7",
          2403 => x"fa",
          2404 => x"71",
          2405 => x"83",
          2406 => x"71",
          2407 => x"06",
          2408 => x"55",
          2409 => x"38",
          2410 => x"89",
          2411 => x"83",
          2412 => x"38",
          2413 => x"33",
          2414 => x"05",
          2415 => x"33",
          2416 => x"b8",
          2417 => x"fa",
          2418 => x"5a",
          2419 => x"34",
          2420 => x"16",
          2421 => x"c7",
          2422 => x"33",
          2423 => x"22",
          2424 => x"11",
          2425 => x"b0",
          2426 => x"18",
          2427 => x"78",
          2428 => x"33",
          2429 => x"53",
          2430 => x"fb",
          2431 => x"84",
          2432 => x"80",
          2433 => x"0c",
          2434 => x"97",
          2435 => x"75",
          2436 => x"38",
          2437 => x"80",
          2438 => x"39",
          2439 => x"b9",
          2440 => x"2e",
          2441 => x"53",
          2442 => x"81",
          2443 => x"72",
          2444 => x"a0",
          2445 => x"81",
          2446 => x"d8",
          2447 => x"b5",
          2448 => x"51",
          2449 => x"84",
          2450 => x"ff",
          2451 => x"83",
          2452 => x"55",
          2453 => x"53",
          2454 => x"a0",
          2455 => x"33",
          2456 => x"53",
          2457 => x"83",
          2458 => x"0b",
          2459 => x"51",
          2460 => x"52",
          2461 => x"39",
          2462 => x"33",
          2463 => x"81",
          2464 => x"83",
          2465 => x"38",
          2466 => x"88",
          2467 => x"88",
          2468 => x"fa",
          2469 => x"72",
          2470 => x"80",
          2471 => x"34",
          2472 => x"33",
          2473 => x"12",
          2474 => x"b6",
          2475 => x"71",
          2476 => x"b0",
          2477 => x"34",
          2478 => x"06",
          2479 => x"33",
          2480 => x"58",
          2481 => x"d6",
          2482 => x"06",
          2483 => x"38",
          2484 => x"f1",
          2485 => x"b5",
          2486 => x"9c",
          2487 => x"8a",
          2488 => x"78",
          2489 => x"db",
          2490 => x"ba",
          2491 => x"fa",
          2492 => x"72",
          2493 => x"80",
          2494 => x"34",
          2495 => x"33",
          2496 => x"12",
          2497 => x"b6",
          2498 => x"71",
          2499 => x"33",
          2500 => x"b8",
          2501 => x"fa",
          2502 => x"72",
          2503 => x"83",
          2504 => x"05",
          2505 => x"06",
          2506 => x"77",
          2507 => x"bb",
          2508 => x"9b",
          2509 => x"83",
          2510 => x"06",
          2511 => x"b5",
          2512 => x"9c",
          2513 => x"aa",
          2514 => x"84",
          2515 => x"11",
          2516 => x"78",
          2517 => x"ff",
          2518 => x"1a",
          2519 => x"9c",
          2520 => x"e9",
          2521 => x"84",
          2522 => x"83",
          2523 => x"5e",
          2524 => x"86",
          2525 => x"f8",
          2526 => x"b2",
          2527 => x"59",
          2528 => x"83",
          2529 => x"5b",
          2530 => x"b0",
          2531 => x"70",
          2532 => x"83",
          2533 => x"44",
          2534 => x"33",
          2535 => x"1f",
          2536 => x"51",
          2537 => x"b5",
          2538 => x"33",
          2539 => x"06",
          2540 => x"12",
          2541 => x"b2",
          2542 => x"05",
          2543 => x"8a",
          2544 => x"81",
          2545 => x"06",
          2546 => x"38",
          2547 => x"fc",
          2548 => x"34",
          2549 => x"0b",
          2550 => x"ba",
          2551 => x"0c",
          2552 => x"3d",
          2553 => x"ba",
          2554 => x"ba",
          2555 => x"ba",
          2556 => x"0c",
          2557 => x"3d",
          2558 => x"81",
          2559 => x"33",
          2560 => x"06",
          2561 => x"06",
          2562 => x"80",
          2563 => x"72",
          2564 => x"06",
          2565 => x"5c",
          2566 => x"fe",
          2567 => x"58",
          2568 => x"83",
          2569 => x"7a",
          2570 => x"72",
          2571 => x"b9",
          2572 => x"34",
          2573 => x"33",
          2574 => x"12",
          2575 => x"fa",
          2576 => x"60",
          2577 => x"fa",
          2578 => x"34",
          2579 => x"06",
          2580 => x"33",
          2581 => x"5e",
          2582 => x"99",
          2583 => x"ff",
          2584 => x"ea",
          2585 => x"96",
          2586 => x"fa",
          2587 => x"81",
          2588 => x"ac",
          2589 => x"78",
          2590 => x"2e",
          2591 => x"5f",
          2592 => x"56",
          2593 => x"10",
          2594 => x"08",
          2595 => x"80",
          2596 => x"0b",
          2597 => x"04",
          2598 => x"33",
          2599 => x"33",
          2600 => x"11",
          2601 => x"b2",
          2602 => x"70",
          2603 => x"33",
          2604 => x"7f",
          2605 => x"7a",
          2606 => x"7a",
          2607 => x"5c",
          2608 => x"c7",
          2609 => x"33",
          2610 => x"22",
          2611 => x"56",
          2612 => x"83",
          2613 => x"5a",
          2614 => x"b0",
          2615 => x"70",
          2616 => x"83",
          2617 => x"5b",
          2618 => x"33",
          2619 => x"05",
          2620 => x"7a",
          2621 => x"33",
          2622 => x"56",
          2623 => x"70",
          2624 => x"26",
          2625 => x"84",
          2626 => x"72",
          2627 => x"72",
          2628 => x"54",
          2629 => x"a0",
          2630 => x"84",
          2631 => x"83",
          2632 => x"5e",
          2633 => x"b6",
          2634 => x"71",
          2635 => x"33",
          2636 => x"b8",
          2637 => x"fa",
          2638 => x"72",
          2639 => x"83",
          2640 => x"34",
          2641 => x"5b",
          2642 => x"77",
          2643 => x"82",
          2644 => x"84",
          2645 => x"83",
          2646 => x"80",
          2647 => x"33",
          2648 => x"56",
          2649 => x"86",
          2650 => x"9c",
          2651 => x"33",
          2652 => x"34",
          2653 => x"33",
          2654 => x"80",
          2655 => x"42",
          2656 => x"51",
          2657 => x"08",
          2658 => x"85",
          2659 => x"ba",
          2660 => x"41",
          2661 => x"ba",
          2662 => x"fa",
          2663 => x"1c",
          2664 => x"84",
          2665 => x"5b",
          2666 => x"f8",
          2667 => x"b5",
          2668 => x"5b",
          2669 => x"c7",
          2670 => x"33",
          2671 => x"22",
          2672 => x"56",
          2673 => x"fa",
          2674 => x"5e",
          2675 => x"b0",
          2676 => x"70",
          2677 => x"83",
          2678 => x"41",
          2679 => x"33",
          2680 => x"70",
          2681 => x"26",
          2682 => x"58",
          2683 => x"75",
          2684 => x"ba",
          2685 => x"7f",
          2686 => x"fc",
          2687 => x"52",
          2688 => x"84",
          2689 => x"84",
          2690 => x"84",
          2691 => x"84",
          2692 => x"b2",
          2693 => x"33",
          2694 => x"33",
          2695 => x"33",
          2696 => x"84",
          2697 => x"ff",
          2698 => x"7c",
          2699 => x"38",
          2700 => x"83",
          2701 => x"53",
          2702 => x"52",
          2703 => x"fe",
          2704 => x"81",
          2705 => x"76",
          2706 => x"38",
          2707 => x"fb",
          2708 => x"84",
          2709 => x"ff",
          2710 => x"38",
          2711 => x"11",
          2712 => x"a5",
          2713 => x"05",
          2714 => x"33",
          2715 => x"83",
          2716 => x"71",
          2717 => x"72",
          2718 => x"83",
          2719 => x"ba",
          2720 => x"e7",
          2721 => x"70",
          2722 => x"5d",
          2723 => x"38",
          2724 => x"39",
          2725 => x"fa",
          2726 => x"57",
          2727 => x"17",
          2728 => x"9c",
          2729 => x"83",
          2730 => x"ff",
          2731 => x"84",
          2732 => x"b4",
          2733 => x"33",
          2734 => x"83",
          2735 => x"71",
          2736 => x"72",
          2737 => x"83",
          2738 => x"ba",
          2739 => x"c4",
          2740 => x"99",
          2741 => x"84",
          2742 => x"83",
          2743 => x"86",
          2744 => x"22",
          2745 => x"05",
          2746 => x"88",
          2747 => x"5a",
          2748 => x"92",
          2749 => x"34",
          2750 => x"5a",
          2751 => x"ba",
          2752 => x"81",
          2753 => x"f9",
          2754 => x"85",
          2755 => x"38",
          2756 => x"33",
          2757 => x"ff",
          2758 => x"83",
          2759 => x"34",
          2760 => x"57",
          2761 => x"ba",
          2762 => x"61",
          2763 => x"59",
          2764 => x"75",
          2765 => x"f4",
          2766 => x"94",
          2767 => x"57",
          2768 => x"76",
          2769 => x"53",
          2770 => x"f4",
          2771 => x"84",
          2772 => x"39",
          2773 => x"57",
          2774 => x"d8",
          2775 => x"75",
          2776 => x"51",
          2777 => x"ba",
          2778 => x"b7",
          2779 => x"70",
          2780 => x"ff",
          2781 => x"f7",
          2782 => x"40",
          2783 => x"7e",
          2784 => x"fa",
          2785 => x"18",
          2786 => x"77",
          2787 => x"b8",
          2788 => x"60",
          2789 => x"83",
          2790 => x"ba",
          2791 => x"ef",
          2792 => x"f7",
          2793 => x"94",
          2794 => x"f8",
          2795 => x"b5",
          2796 => x"a0",
          2797 => x"40",
          2798 => x"ff",
          2799 => x"59",
          2800 => x"f0",
          2801 => x"7c",
          2802 => x"fe",
          2803 => x"76",
          2804 => x"75",
          2805 => x"06",
          2806 => x"24",
          2807 => x"56",
          2808 => x"16",
          2809 => x"81",
          2810 => x"57",
          2811 => x"75",
          2812 => x"06",
          2813 => x"58",
          2814 => x"b0",
          2815 => x"ff",
          2816 => x"42",
          2817 => x"84",
          2818 => x"33",
          2819 => x"70",
          2820 => x"05",
          2821 => x"34",
          2822 => x"b8",
          2823 => x"40",
          2824 => x"38",
          2825 => x"80",
          2826 => x"34",
          2827 => x"70",
          2828 => x"b8",
          2829 => x"71",
          2830 => x"78",
          2831 => x"84",
          2832 => x"87",
          2833 => x"33",
          2834 => x"80",
          2835 => x"84",
          2836 => x"79",
          2837 => x"22",
          2838 => x"8b",
          2839 => x"76",
          2840 => x"79",
          2841 => x"ed",
          2842 => x"60",
          2843 => x"06",
          2844 => x"7b",
          2845 => x"76",
          2846 => x"70",
          2847 => x"80",
          2848 => x"b0",
          2849 => x"5d",
          2850 => x"57",
          2851 => x"33",
          2852 => x"71",
          2853 => x"59",
          2854 => x"38",
          2855 => x"7d",
          2856 => x"77",
          2857 => x"84",
          2858 => x"ff",
          2859 => x"b2",
          2860 => x"59",
          2861 => x"76",
          2862 => x"05",
          2863 => x"76",
          2864 => x"b0",
          2865 => x"a0",
          2866 => x"70",
          2867 => x"76",
          2868 => x"e0",
          2869 => x"05",
          2870 => x"27",
          2871 => x"70",
          2872 => x"39",
          2873 => x"06",
          2874 => x"84",
          2875 => x"f0",
          2876 => x"f2",
          2877 => x"70",
          2878 => x"39",
          2879 => x"b9",
          2880 => x"b4",
          2881 => x"b2",
          2882 => x"5f",
          2883 => x"33",
          2884 => x"34",
          2885 => x"56",
          2886 => x"81",
          2887 => x"fa",
          2888 => x"33",
          2889 => x"83",
          2890 => x"b0",
          2891 => x"75",
          2892 => x"fa",
          2893 => x"56",
          2894 => x"39",
          2895 => x"81",
          2896 => x"f4",
          2897 => x"8f",
          2898 => x"ff",
          2899 => x"9f",
          2900 => x"b0",
          2901 => x"33",
          2902 => x"75",
          2903 => x"83",
          2904 => x"c0",
          2905 => x"fe",
          2906 => x"af",
          2907 => x"b0",
          2908 => x"33",
          2909 => x"83",
          2910 => x"fa",
          2911 => x"56",
          2912 => x"39",
          2913 => x"82",
          2914 => x"fe",
          2915 => x"f8",
          2916 => x"fd",
          2917 => x"f0",
          2918 => x"fd",
          2919 => x"f0",
          2920 => x"fd",
          2921 => x"df",
          2922 => x"fa",
          2923 => x"b0",
          2924 => x"75",
          2925 => x"80",
          2926 => x"81",
          2927 => x"84",
          2928 => x"84",
          2929 => x"84",
          2930 => x"b2",
          2931 => x"e8",
          2932 => x"34",
          2933 => x"3d",
          2934 => x"83",
          2935 => x"58",
          2936 => x"ba",
          2937 => x"d8",
          2938 => x"bb",
          2939 => x"08",
          2940 => x"ba",
          2941 => x"0c",
          2942 => x"b5",
          2943 => x"33",
          2944 => x"85",
          2945 => x"02",
          2946 => x"1e",
          2947 => x"ca",
          2948 => x"80",
          2949 => x"fa",
          2950 => x"ff",
          2951 => x"83",
          2952 => x"d0",
          2953 => x"fe",
          2954 => x"fa",
          2955 => x"9f",
          2956 => x"a6",
          2957 => x"84",
          2958 => x"ee",
          2959 => x"ee",
          2960 => x"05",
          2961 => x"58",
          2962 => x"b4",
          2963 => x"ff",
          2964 => x"f3",
          2965 => x"84",
          2966 => x"58",
          2967 => x"83",
          2968 => x"70",
          2969 => x"71",
          2970 => x"05",
          2971 => x"7e",
          2972 => x"83",
          2973 => x"5f",
          2974 => x"79",
          2975 => x"57",
          2976 => x"b8",
          2977 => x"98",
          2978 => x"b2",
          2979 => x"57",
          2980 => x"84",
          2981 => x"82",
          2982 => x"fa",
          2983 => x"fa",
          2984 => x"76",
          2985 => x"05",
          2986 => x"5c",
          2987 => x"80",
          2988 => x"ff",
          2989 => x"29",
          2990 => x"27",
          2991 => x"57",
          2992 => x"80",
          2993 => x"34",
          2994 => x"70",
          2995 => x"b8",
          2996 => x"71",
          2997 => x"76",
          2998 => x"33",
          2999 => x"70",
          3000 => x"05",
          3001 => x"34",
          3002 => x"b8",
          3003 => x"41",
          3004 => x"38",
          3005 => x"33",
          3006 => x"34",
          3007 => x"33",
          3008 => x"33",
          3009 => x"76",
          3010 => x"70",
          3011 => x"58",
          3012 => x"79",
          3013 => x"06",
          3014 => x"83",
          3015 => x"34",
          3016 => x"06",
          3017 => x"27",
          3018 => x"fa",
          3019 => x"b5",
          3020 => x"ff",
          3021 => x"ef",
          3022 => x"75",
          3023 => x"38",
          3024 => x"06",
          3025 => x"5d",
          3026 => x"f4",
          3027 => x"56",
          3028 => x"39",
          3029 => x"23",
          3030 => x"75",
          3031 => x"77",
          3032 => x"8d",
          3033 => x"34",
          3034 => x"05",
          3035 => x"38",
          3036 => x"83",
          3037 => x"59",
          3038 => x"d3",
          3039 => x"fa",
          3040 => x"83",
          3041 => x"83",
          3042 => x"0b",
          3043 => x"80",
          3044 => x"39",
          3045 => x"b9",
          3046 => x"83",
          3047 => x"3d",
          3048 => x"fa",
          3049 => x"38",
          3050 => x"84",
          3051 => x"76",
          3052 => x"0b",
          3053 => x"04",
          3054 => x"5c",
          3055 => x"81",
          3056 => x"58",
          3057 => x"d6",
          3058 => x"88",
          3059 => x"0c",
          3060 => x"08",
          3061 => x"38",
          3062 => x"70",
          3063 => x"58",
          3064 => x"80",
          3065 => x"83",
          3066 => x"30",
          3067 => x"5d",
          3068 => x"b8",
          3069 => x"fa",
          3070 => x"c7",
          3071 => x"5b",
          3072 => x"83",
          3073 => x"58",
          3074 => x"8c",
          3075 => x"80",
          3076 => x"88",
          3077 => x"75",
          3078 => x"84",
          3079 => x"34",
          3080 => x"55",
          3081 => x"54",
          3082 => x"ff",
          3083 => x"54",
          3084 => x"72",
          3085 => x"83",
          3086 => x"06",
          3087 => x"38",
          3088 => x"f8",
          3089 => x"34",
          3090 => x"5e",
          3091 => x"f8",
          3092 => x"25",
          3093 => x"34",
          3094 => x"81",
          3095 => x"72",
          3096 => x"83",
          3097 => x"53",
          3098 => x"0b",
          3099 => x"f8",
          3100 => x"f8",
          3101 => x"83",
          3102 => x"5c",
          3103 => x"55",
          3104 => x"f8",
          3105 => x"82",
          3106 => x"53",
          3107 => x"f8",
          3108 => x"38",
          3109 => x"ff",
          3110 => x"33",
          3111 => x"74",
          3112 => x"2e",
          3113 => x"33",
          3114 => x"83",
          3115 => x"c0",
          3116 => x"27",
          3117 => x"98",
          3118 => x"81",
          3119 => x"89",
          3120 => x"f8",
          3121 => x"fe",
          3122 => x"8b",
          3123 => x"05",
          3124 => x"08",
          3125 => x"f4",
          3126 => x"5e",
          3127 => x"0b",
          3128 => x"81",
          3129 => x"f9",
          3130 => x"83",
          3131 => x"58",
          3132 => x"b6",
          3133 => x"33",
          3134 => x"39",
          3135 => x"2e",
          3136 => x"f4",
          3137 => x"54",
          3138 => x"39",
          3139 => x"81",
          3140 => x"81",
          3141 => x"80",
          3142 => x"38",
          3143 => x"27",
          3144 => x"25",
          3145 => x"81",
          3146 => x"81",
          3147 => x"2b",
          3148 => x"24",
          3149 => x"10",
          3150 => x"83",
          3151 => x"54",
          3152 => x"f8",
          3153 => x"59",
          3154 => x"81",
          3155 => x"59",
          3156 => x"9f",
          3157 => x"54",
          3158 => x"7b",
          3159 => x"76",
          3160 => x"7b",
          3161 => x"38",
          3162 => x"53",
          3163 => x"05",
          3164 => x"83",
          3165 => x"06",
          3166 => x"84",
          3167 => x"f9",
          3168 => x"74",
          3169 => x"52",
          3170 => x"bb",
          3171 => x"76",
          3172 => x"72",
          3173 => x"cc",
          3174 => x"f8",
          3175 => x"0b",
          3176 => x"83",
          3177 => x"f8",
          3178 => x"81",
          3179 => x"fc",
          3180 => x"55",
          3181 => x"81",
          3182 => x"81",
          3183 => x"08",
          3184 => x"08",
          3185 => x"38",
          3186 => x"d8",
          3187 => x"d7",
          3188 => x"34",
          3189 => x"34",
          3190 => x"9e",
          3191 => x"0b",
          3192 => x"08",
          3193 => x"e0",
          3194 => x"42",
          3195 => x"79",
          3196 => x"38",
          3197 => x"38",
          3198 => x"c0",
          3199 => x"81",
          3200 => x"84",
          3201 => x"38",
          3202 => x"ff",
          3203 => x"b8",
          3204 => x"81",
          3205 => x"59",
          3206 => x"e4",
          3207 => x"0b",
          3208 => x"84",
          3209 => x"ff",
          3210 => x"83",
          3211 => x"23",
          3212 => x"53",
          3213 => x"73",
          3214 => x"33",
          3215 => x"53",
          3216 => x"72",
          3217 => x"b7",
          3218 => x"a5",
          3219 => x"54",
          3220 => x"83",
          3221 => x"81",
          3222 => x"e8",
          3223 => x"0d",
          3224 => x"0d",
          3225 => x"f5",
          3226 => x"33",
          3227 => x"51",
          3228 => x"f5",
          3229 => x"15",
          3230 => x"34",
          3231 => x"90",
          3232 => x"87",
          3233 => x"98",
          3234 => x"38",
          3235 => x"08",
          3236 => x"71",
          3237 => x"98",
          3238 => x"27",
          3239 => x"2e",
          3240 => x"08",
          3241 => x"98",
          3242 => x"08",
          3243 => x"14",
          3244 => x"52",
          3245 => x"ff",
          3246 => x"08",
          3247 => x"52",
          3248 => x"06",
          3249 => x"74",
          3250 => x"38",
          3251 => x"bb",
          3252 => x"0b",
          3253 => x"04",
          3254 => x"a3",
          3255 => x"f5",
          3256 => x"80",
          3257 => x"51",
          3258 => x"72",
          3259 => x"71",
          3260 => x"72",
          3261 => x"52",
          3262 => x"08",
          3263 => x"83",
          3264 => x"81",
          3265 => x"e8",
          3266 => x"f5",
          3267 => x"53",
          3268 => x"c0",
          3269 => x"f6",
          3270 => x"9c",
          3271 => x"38",
          3272 => x"c0",
          3273 => x"73",
          3274 => x"ff",
          3275 => x"9c",
          3276 => x"c0",
          3277 => x"9c",
          3278 => x"81",
          3279 => x"52",
          3280 => x"81",
          3281 => x"a4",
          3282 => x"ff",
          3283 => x"ff",
          3284 => x"c7",
          3285 => x"fe",
          3286 => x"06",
          3287 => x"7b",
          3288 => x"73",
          3289 => x"53",
          3290 => x"72",
          3291 => x"84",
          3292 => x"84",
          3293 => x"ff",
          3294 => x"02",
          3295 => x"80",
          3296 => x"2b",
          3297 => x"98",
          3298 => x"83",
          3299 => x"84",
          3300 => x"85",
          3301 => x"83",
          3302 => x"80",
          3303 => x"27",
          3304 => x"33",
          3305 => x"71",
          3306 => x"54",
          3307 => x"08",
          3308 => x"83",
          3309 => x"81",
          3310 => x"e8",
          3311 => x"f5",
          3312 => x"53",
          3313 => x"c0",
          3314 => x"f6",
          3315 => x"9c",
          3316 => x"38",
          3317 => x"c0",
          3318 => x"73",
          3319 => x"ff",
          3320 => x"9c",
          3321 => x"c0",
          3322 => x"9c",
          3323 => x"81",
          3324 => x"52",
          3325 => x"81",
          3326 => x"a4",
          3327 => x"ff",
          3328 => x"ff",
          3329 => x"38",
          3330 => x"d5",
          3331 => x"54",
          3332 => x"76",
          3333 => x"04",
          3334 => x"83",
          3335 => x"34",
          3336 => x"56",
          3337 => x"87",
          3338 => x"9c",
          3339 => x"ce",
          3340 => x"08",
          3341 => x"72",
          3342 => x"87",
          3343 => x"74",
          3344 => x"db",
          3345 => x"ff",
          3346 => x"71",
          3347 => x"87",
          3348 => x"05",
          3349 => x"87",
          3350 => x"2e",
          3351 => x"98",
          3352 => x"87",
          3353 => x"87",
          3354 => x"26",
          3355 => x"16",
          3356 => x"80",
          3357 => x"54",
          3358 => x"3d",
          3359 => x"f7",
          3360 => x"0d",
          3361 => x"83",
          3362 => x"83",
          3363 => x"33",
          3364 => x"77",
          3365 => x"98",
          3366 => x"41",
          3367 => x"57",
          3368 => x"72",
          3369 => x"71",
          3370 => x"05",
          3371 => x"2b",
          3372 => x"52",
          3373 => x"9e",
          3374 => x"71",
          3375 => x"05",
          3376 => x"74",
          3377 => x"54",
          3378 => x"08",
          3379 => x"33",
          3380 => x"5c",
          3381 => x"34",
          3382 => x"08",
          3383 => x"80",
          3384 => x"08",
          3385 => x"14",
          3386 => x"33",
          3387 => x"82",
          3388 => x"58",
          3389 => x"13",
          3390 => x"33",
          3391 => x"83",
          3392 => x"85",
          3393 => x"88",
          3394 => x"58",
          3395 => x"34",
          3396 => x"11",
          3397 => x"71",
          3398 => x"72",
          3399 => x"71",
          3400 => x"55",
          3401 => x"87",
          3402 => x"70",
          3403 => x"07",
          3404 => x"5a",
          3405 => x"81",
          3406 => x"17",
          3407 => x"2b",
          3408 => x"33",
          3409 => x"70",
          3410 => x"05",
          3411 => x"5c",
          3412 => x"34",
          3413 => x"08",
          3414 => x"71",
          3415 => x"05",
          3416 => x"2b",
          3417 => x"2a",
          3418 => x"52",
          3419 => x"84",
          3420 => x"33",
          3421 => x"83",
          3422 => x"12",
          3423 => x"07",
          3424 => x"53",
          3425 => x"33",
          3426 => x"82",
          3427 => x"59",
          3428 => x"34",
          3429 => x"33",
          3430 => x"83",
          3431 => x"83",
          3432 => x"88",
          3433 => x"52",
          3434 => x"15",
          3435 => x"0d",
          3436 => x"76",
          3437 => x"86",
          3438 => x"3d",
          3439 => x"ba",
          3440 => x"f0",
          3441 => x"84",
          3442 => x"84",
          3443 => x"81",
          3444 => x"08",
          3445 => x"85",
          3446 => x"76",
          3447 => x"34",
          3448 => x"22",
          3449 => x"83",
          3450 => x"51",
          3451 => x"89",
          3452 => x"10",
          3453 => x"f8",
          3454 => x"81",
          3455 => x"f7",
          3456 => x"51",
          3457 => x"83",
          3458 => x"06",
          3459 => x"84",
          3460 => x"12",
          3461 => x"59",
          3462 => x"75",
          3463 => x"10",
          3464 => x"71",
          3465 => x"06",
          3466 => x"70",
          3467 => x"52",
          3468 => x"2e",
          3469 => x"12",
          3470 => x"07",
          3471 => x"ff",
          3472 => x"56",
          3473 => x"33",
          3474 => x"70",
          3475 => x"56",
          3476 => x"81",
          3477 => x"8d",
          3478 => x"85",
          3479 => x"74",
          3480 => x"82",
          3481 => x"5c",
          3482 => x"81",
          3483 => x"76",
          3484 => x"34",
          3485 => x"08",
          3486 => x"71",
          3487 => x"ff",
          3488 => x"ff",
          3489 => x"57",
          3490 => x"72",
          3491 => x"34",
          3492 => x"74",
          3493 => x"f4",
          3494 => x"12",
          3495 => x"07",
          3496 => x"75",
          3497 => x"84",
          3498 => x"05",
          3499 => x"88",
          3500 => x"58",
          3501 => x"15",
          3502 => x"84",
          3503 => x"2b",
          3504 => x"5a",
          3505 => x"72",
          3506 => x"70",
          3507 => x"85",
          3508 => x"88",
          3509 => x"15",
          3510 => x"f4",
          3511 => x"bb",
          3512 => x"14",
          3513 => x"71",
          3514 => x"33",
          3515 => x"70",
          3516 => x"52",
          3517 => x"34",
          3518 => x"11",
          3519 => x"71",
          3520 => x"33",
          3521 => x"70",
          3522 => x"5b",
          3523 => x"87",
          3524 => x"70",
          3525 => x"07",
          3526 => x"59",
          3527 => x"81",
          3528 => x"84",
          3529 => x"0d",
          3530 => x"76",
          3531 => x"8a",
          3532 => x"3d",
          3533 => x"84",
          3534 => x"89",
          3535 => x"84",
          3536 => x"ba",
          3537 => x"52",
          3538 => x"3f",
          3539 => x"34",
          3540 => x"f4",
          3541 => x"0b",
          3542 => x"56",
          3543 => x"17",
          3544 => x"f0",
          3545 => x"70",
          3546 => x"58",
          3547 => x"73",
          3548 => x"70",
          3549 => x"05",
          3550 => x"34",
          3551 => x"77",
          3552 => x"39",
          3553 => x"80",
          3554 => x"41",
          3555 => x"80",
          3556 => x"88",
          3557 => x"8f",
          3558 => x"05",
          3559 => x"73",
          3560 => x"83",
          3561 => x"83",
          3562 => x"33",
          3563 => x"70",
          3564 => x"10",
          3565 => x"70",
          3566 => x"07",
          3567 => x"42",
          3568 => x"5c",
          3569 => x"7a",
          3570 => x"83",
          3571 => x"10",
          3572 => x"33",
          3573 => x"53",
          3574 => x"24",
          3575 => x"f6",
          3576 => x"87",
          3577 => x"38",
          3578 => x"be",
          3579 => x"92",
          3580 => x"12",
          3581 => x"07",
          3582 => x"71",
          3583 => x"43",
          3584 => x"60",
          3585 => x"11",
          3586 => x"71",
          3587 => x"33",
          3588 => x"83",
          3589 => x"85",
          3590 => x"88",
          3591 => x"58",
          3592 => x"34",
          3593 => x"08",
          3594 => x"33",
          3595 => x"74",
          3596 => x"71",
          3597 => x"42",
          3598 => x"86",
          3599 => x"ba",
          3600 => x"33",
          3601 => x"06",
          3602 => x"76",
          3603 => x"ba",
          3604 => x"83",
          3605 => x"2b",
          3606 => x"33",
          3607 => x"41",
          3608 => x"79",
          3609 => x"ba",
          3610 => x"12",
          3611 => x"07",
          3612 => x"33",
          3613 => x"41",
          3614 => x"79",
          3615 => x"84",
          3616 => x"33",
          3617 => x"66",
          3618 => x"52",
          3619 => x"fe",
          3620 => x"1e",
          3621 => x"83",
          3622 => x"62",
          3623 => x"84",
          3624 => x"84",
          3625 => x"a0",
          3626 => x"80",
          3627 => x"51",
          3628 => x"08",
          3629 => x"1f",
          3630 => x"84",
          3631 => x"84",
          3632 => x"34",
          3633 => x"f4",
          3634 => x"fe",
          3635 => x"06",
          3636 => x"78",
          3637 => x"84",
          3638 => x"84",
          3639 => x"56",
          3640 => x"15",
          3641 => x"fa",
          3642 => x"38",
          3643 => x"38",
          3644 => x"84",
          3645 => x"0d",
          3646 => x"71",
          3647 => x"05",
          3648 => x"2b",
          3649 => x"2a",
          3650 => x"34",
          3651 => x"f4",
          3652 => x"75",
          3653 => x"84",
          3654 => x"81",
          3655 => x"83",
          3656 => x"64",
          3657 => x"4a",
          3658 => x"63",
          3659 => x"41",
          3660 => x"f4",
          3661 => x"81",
          3662 => x"05",
          3663 => x"54",
          3664 => x"83",
          3665 => x"39",
          3666 => x"70",
          3667 => x"83",
          3668 => x"10",
          3669 => x"33",
          3670 => x"53",
          3671 => x"73",
          3672 => x"39",
          3673 => x"7a",
          3674 => x"ff",
          3675 => x"38",
          3676 => x"84",
          3677 => x"ba",
          3678 => x"52",
          3679 => x"3f",
          3680 => x"34",
          3681 => x"f4",
          3682 => x"0b",
          3683 => x"58",
          3684 => x"19",
          3685 => x"f0",
          3686 => x"70",
          3687 => x"58",
          3688 => x"34",
          3689 => x"f0",
          3690 => x"f4",
          3691 => x"61",
          3692 => x"34",
          3693 => x"de",
          3694 => x"61",
          3695 => x"39",
          3696 => x"51",
          3697 => x"bb",
          3698 => x"1e",
          3699 => x"8b",
          3700 => x"86",
          3701 => x"2b",
          3702 => x"14",
          3703 => x"07",
          3704 => x"5b",
          3705 => x"64",
          3706 => x"34",
          3707 => x"11",
          3708 => x"71",
          3709 => x"33",
          3710 => x"70",
          3711 => x"59",
          3712 => x"7a",
          3713 => x"08",
          3714 => x"88",
          3715 => x"88",
          3716 => x"34",
          3717 => x"08",
          3718 => x"33",
          3719 => x"74",
          3720 => x"88",
          3721 => x"5e",
          3722 => x"34",
          3723 => x"08",
          3724 => x"71",
          3725 => x"05",
          3726 => x"88",
          3727 => x"40",
          3728 => x"18",
          3729 => x"f4",
          3730 => x"12",
          3731 => x"62",
          3732 => x"5d",
          3733 => x"96",
          3734 => x"05",
          3735 => x"fc",
          3736 => x"ba",
          3737 => x"f0",
          3738 => x"84",
          3739 => x"84",
          3740 => x"81",
          3741 => x"08",
          3742 => x"85",
          3743 => x"7f",
          3744 => x"34",
          3745 => x"22",
          3746 => x"83",
          3747 => x"43",
          3748 => x"89",
          3749 => x"10",
          3750 => x"f8",
          3751 => x"81",
          3752 => x"bd",
          3753 => x"19",
          3754 => x"71",
          3755 => x"33",
          3756 => x"70",
          3757 => x"55",
          3758 => x"85",
          3759 => x"1e",
          3760 => x"8b",
          3761 => x"86",
          3762 => x"2b",
          3763 => x"48",
          3764 => x"05",
          3765 => x"ba",
          3766 => x"33",
          3767 => x"06",
          3768 => x"75",
          3769 => x"ba",
          3770 => x"12",
          3771 => x"07",
          3772 => x"71",
          3773 => x"ff",
          3774 => x"48",
          3775 => x"41",
          3776 => x"34",
          3777 => x"33",
          3778 => x"83",
          3779 => x"12",
          3780 => x"ff",
          3781 => x"5e",
          3782 => x"76",
          3783 => x"ff",
          3784 => x"33",
          3785 => x"83",
          3786 => x"85",
          3787 => x"88",
          3788 => x"78",
          3789 => x"84",
          3790 => x"33",
          3791 => x"83",
          3792 => x"87",
          3793 => x"88",
          3794 => x"55",
          3795 => x"60",
          3796 => x"18",
          3797 => x"2b",
          3798 => x"2a",
          3799 => x"78",
          3800 => x"70",
          3801 => x"8b",
          3802 => x"70",
          3803 => x"07",
          3804 => x"77",
          3805 => x"5f",
          3806 => x"17",
          3807 => x"f4",
          3808 => x"33",
          3809 => x"74",
          3810 => x"88",
          3811 => x"88",
          3812 => x"5d",
          3813 => x"34",
          3814 => x"11",
          3815 => x"71",
          3816 => x"33",
          3817 => x"83",
          3818 => x"85",
          3819 => x"88",
          3820 => x"59",
          3821 => x"1d",
          3822 => x"f4",
          3823 => x"12",
          3824 => x"07",
          3825 => x"33",
          3826 => x"5f",
          3827 => x"77",
          3828 => x"84",
          3829 => x"12",
          3830 => x"ff",
          3831 => x"59",
          3832 => x"84",
          3833 => x"33",
          3834 => x"83",
          3835 => x"15",
          3836 => x"2a",
          3837 => x"55",
          3838 => x"84",
          3839 => x"81",
          3840 => x"2b",
          3841 => x"15",
          3842 => x"2a",
          3843 => x"55",
          3844 => x"34",
          3845 => x"11",
          3846 => x"07",
          3847 => x"42",
          3848 => x"51",
          3849 => x"08",
          3850 => x"70",
          3851 => x"f1",
          3852 => x"33",
          3853 => x"79",
          3854 => x"71",
          3855 => x"48",
          3856 => x"05",
          3857 => x"ba",
          3858 => x"85",
          3859 => x"2b",
          3860 => x"15",
          3861 => x"2a",
          3862 => x"56",
          3863 => x"87",
          3864 => x"70",
          3865 => x"07",
          3866 => x"5c",
          3867 => x"81",
          3868 => x"1f",
          3869 => x"2b",
          3870 => x"33",
          3871 => x"70",
          3872 => x"05",
          3873 => x"58",
          3874 => x"34",
          3875 => x"08",
          3876 => x"71",
          3877 => x"05",
          3878 => x"2b",
          3879 => x"2a",
          3880 => x"5b",
          3881 => x"77",
          3882 => x"39",
          3883 => x"84",
          3884 => x"08",
          3885 => x"52",
          3886 => x"f6",
          3887 => x"5b",
          3888 => x"e9",
          3889 => x"84",
          3890 => x"2e",
          3891 => x"73",
          3892 => x"04",
          3893 => x"84",
          3894 => x"2e",
          3895 => x"bb",
          3896 => x"73",
          3897 => x"04",
          3898 => x"0c",
          3899 => x"82",
          3900 => x"f4",
          3901 => x"f4",
          3902 => x"81",
          3903 => x"76",
          3904 => x"34",
          3905 => x"17",
          3906 => x"ba",
          3907 => x"05",
          3908 => x"ff",
          3909 => x"56",
          3910 => x"34",
          3911 => x"10",
          3912 => x"55",
          3913 => x"83",
          3914 => x"fe",
          3915 => x"0d",
          3916 => x"70",
          3917 => x"11",
          3918 => x"83",
          3919 => x"93",
          3920 => x"26",
          3921 => x"84",
          3922 => x"72",
          3923 => x"34",
          3924 => x"84",
          3925 => x"f7",
          3926 => x"05",
          3927 => x"81",
          3928 => x"bb",
          3929 => x"54",
          3930 => x"85",
          3931 => x"53",
          3932 => x"84",
          3933 => x"74",
          3934 => x"8c",
          3935 => x"26",
          3936 => x"54",
          3937 => x"73",
          3938 => x"3d",
          3939 => x"70",
          3940 => x"78",
          3941 => x"3d",
          3942 => x"af",
          3943 => x"54",
          3944 => x"80",
          3945 => x"83",
          3946 => x"0b",
          3947 => x"75",
          3948 => x"bb",
          3949 => x"80",
          3950 => x"08",
          3951 => x"d6",
          3952 => x"73",
          3953 => x"55",
          3954 => x"0d",
          3955 => x"81",
          3956 => x"26",
          3957 => x"0d",
          3958 => x"02",
          3959 => x"55",
          3960 => x"84",
          3961 => x"06",
          3962 => x"0b",
          3963 => x"70",
          3964 => x"ad",
          3965 => x"53",
          3966 => x"0d",
          3967 => x"84",
          3968 => x"81",
          3969 => x"84",
          3970 => x"2b",
          3971 => x"70",
          3972 => x"81",
          3973 => x"38",
          3974 => x"ea",
          3975 => x"70",
          3976 => x"92",
          3977 => x"54",
          3978 => x"08",
          3979 => x"90",
          3980 => x"0b",
          3981 => x"74",
          3982 => x"77",
          3983 => x"38",
          3984 => x"51",
          3985 => x"80",
          3986 => x"bb",
          3987 => x"54",
          3988 => x"53",
          3989 => x"3f",
          3990 => x"2e",
          3991 => x"84",
          3992 => x"70",
          3993 => x"84",
          3994 => x"74",
          3995 => x"33",
          3996 => x"ff",
          3997 => x"79",
          3998 => x"3f",
          3999 => x"2e",
          4000 => x"18",
          4001 => x"06",
          4002 => x"80",
          4003 => x"05",
          4004 => x"38",
          4005 => x"ff",
          4006 => x"d2",
          4007 => x"34",
          4008 => x"c1",
          4009 => x"84",
          4010 => x"9d",
          4011 => x"19",
          4012 => x"34",
          4013 => x"19",
          4014 => x"a1",
          4015 => x"84",
          4016 => x"7a",
          4017 => x"5b",
          4018 => x"2a",
          4019 => x"90",
          4020 => x"7a",
          4021 => x"34",
          4022 => x"1a",
          4023 => x"52",
          4024 => x"76",
          4025 => x"81",
          4026 => x"bb",
          4027 => x"fd",
          4028 => x"70",
          4029 => x"88",
          4030 => x"38",
          4031 => x"8f",
          4032 => x"58",
          4033 => x"82",
          4034 => x"09",
          4035 => x"16",
          4036 => x"5a",
          4037 => x"2e",
          4038 => x"7b",
          4039 => x"81",
          4040 => x"17",
          4041 => x"84",
          4042 => x"81",
          4043 => x"9a",
          4044 => x"11",
          4045 => x"1b",
          4046 => x"17",
          4047 => x"83",
          4048 => x"7d",
          4049 => x"81",
          4050 => x"17",
          4051 => x"84",
          4052 => x"81",
          4053 => x"ca",
          4054 => x"11",
          4055 => x"81",
          4056 => x"59",
          4057 => x"ff",
          4058 => x"0d",
          4059 => x"05",
          4060 => x"38",
          4061 => x"5d",
          4062 => x"81",
          4063 => x"17",
          4064 => x"3f",
          4065 => x"38",
          4066 => x"0c",
          4067 => x"fe",
          4068 => x"33",
          4069 => x"bb",
          4070 => x"04",
          4071 => x"b8",
          4072 => x"05",
          4073 => x"38",
          4074 => x"5e",
          4075 => x"82",
          4076 => x"17",
          4077 => x"3f",
          4078 => x"38",
          4079 => x"0c",
          4080 => x"83",
          4081 => x"11",
          4082 => x"71",
          4083 => x"72",
          4084 => x"ff",
          4085 => x"84",
          4086 => x"8f",
          4087 => x"08",
          4088 => x"33",
          4089 => x"84",
          4090 => x"06",
          4091 => x"83",
          4092 => x"08",
          4093 => x"7d",
          4094 => x"82",
          4095 => x"81",
          4096 => x"17",
          4097 => x"52",
          4098 => x"7a",
          4099 => x"17",
          4100 => x"18",
          4101 => x"bb",
          4102 => x"82",
          4103 => x"18",
          4104 => x"31",
          4105 => x"38",
          4106 => x"81",
          4107 => x"fb",
          4108 => x"53",
          4109 => x"52",
          4110 => x"bb",
          4111 => x"fd",
          4112 => x"18",
          4113 => x"31",
          4114 => x"a0",
          4115 => x"17",
          4116 => x"06",
          4117 => x"08",
          4118 => x"81",
          4119 => x"5a",
          4120 => x"08",
          4121 => x"33",
          4122 => x"84",
          4123 => x"06",
          4124 => x"83",
          4125 => x"08",
          4126 => x"74",
          4127 => x"82",
          4128 => x"81",
          4129 => x"17",
          4130 => x"52",
          4131 => x"7c",
          4132 => x"17",
          4133 => x"52",
          4134 => x"fa",
          4135 => x"38",
          4136 => x"62",
          4137 => x"76",
          4138 => x"27",
          4139 => x"2e",
          4140 => x"38",
          4141 => x"84",
          4142 => x"75",
          4143 => x"80",
          4144 => x"78",
          4145 => x"7c",
          4146 => x"06",
          4147 => x"b8",
          4148 => x"87",
          4149 => x"85",
          4150 => x"1a",
          4151 => x"75",
          4152 => x"83",
          4153 => x"1f",
          4154 => x"1f",
          4155 => x"84",
          4156 => x"74",
          4157 => x"38",
          4158 => x"58",
          4159 => x"76",
          4160 => x"33",
          4161 => x"81",
          4162 => x"53",
          4163 => x"f1",
          4164 => x"2e",
          4165 => x"b4",
          4166 => x"38",
          4167 => x"05",
          4168 => x"2b",
          4169 => x"07",
          4170 => x"7d",
          4171 => x"7d",
          4172 => x"7d",
          4173 => x"81",
          4174 => x"75",
          4175 => x"1b",
          4176 => x"5a",
          4177 => x"83",
          4178 => x"7d",
          4179 => x"81",
          4180 => x"19",
          4181 => x"84",
          4182 => x"81",
          4183 => x"7b",
          4184 => x"19",
          4185 => x"5f",
          4186 => x"8f",
          4187 => x"77",
          4188 => x"74",
          4189 => x"7d",
          4190 => x"80",
          4191 => x"76",
          4192 => x"53",
          4193 => x"52",
          4194 => x"bb",
          4195 => x"80",
          4196 => x"1a",
          4197 => x"08",
          4198 => x"08",
          4199 => x"8b",
          4200 => x"2e",
          4201 => x"76",
          4202 => x"3f",
          4203 => x"38",
          4204 => x"0c",
          4205 => x"06",
          4206 => x"56",
          4207 => x"33",
          4208 => x"56",
          4209 => x"1a",
          4210 => x"53",
          4211 => x"52",
          4212 => x"bb",
          4213 => x"fc",
          4214 => x"1a",
          4215 => x"08",
          4216 => x"08",
          4217 => x"fb",
          4218 => x"82",
          4219 => x"81",
          4220 => x"19",
          4221 => x"fb",
          4222 => x"19",
          4223 => x"ee",
          4224 => x"08",
          4225 => x"38",
          4226 => x"b4",
          4227 => x"a0",
          4228 => x"40",
          4229 => x"38",
          4230 => x"09",
          4231 => x"7d",
          4232 => x"51",
          4233 => x"39",
          4234 => x"53",
          4235 => x"3f",
          4236 => x"2e",
          4237 => x"bb",
          4238 => x"08",
          4239 => x"08",
          4240 => x"5e",
          4241 => x"19",
          4242 => x"06",
          4243 => x"53",
          4244 => x"86",
          4245 => x"54",
          4246 => x"33",
          4247 => x"8b",
          4248 => x"7a",
          4249 => x"5f",
          4250 => x"2a",
          4251 => x"39",
          4252 => x"82",
          4253 => x"11",
          4254 => x"0a",
          4255 => x"58",
          4256 => x"88",
          4257 => x"90",
          4258 => x"98",
          4259 => x"cf",
          4260 => x"08",
          4261 => x"90",
          4262 => x"f4",
          4263 => x"ec",
          4264 => x"73",
          4265 => x"2e",
          4266 => x"56",
          4267 => x"82",
          4268 => x"75",
          4269 => x"bb",
          4270 => x"80",
          4271 => x"b1",
          4272 => x"30",
          4273 => x"07",
          4274 => x"38",
          4275 => x"b5",
          4276 => x"0c",
          4277 => x"91",
          4278 => x"39",
          4279 => x"81",
          4280 => x"db",
          4281 => x"bb",
          4282 => x"19",
          4283 => x"38",
          4284 => x"56",
          4285 => x"82",
          4286 => x"3f",
          4287 => x"2e",
          4288 => x"09",
          4289 => x"70",
          4290 => x"51",
          4291 => x"84",
          4292 => x"90",
          4293 => x"a3",
          4294 => x"9b",
          4295 => x"39",
          4296 => x"53",
          4297 => x"84",
          4298 => x"30",
          4299 => x"25",
          4300 => x"74",
          4301 => x"9c",
          4302 => x"56",
          4303 => x"15",
          4304 => x"07",
          4305 => x"74",
          4306 => x"04",
          4307 => x"3d",
          4308 => x"fe",
          4309 => x"38",
          4310 => x"8b",
          4311 => x"a7",
          4312 => x"84",
          4313 => x"74",
          4314 => x"ff",
          4315 => x"71",
          4316 => x"0a",
          4317 => x"53",
          4318 => x"0c",
          4319 => x"38",
          4320 => x"cc",
          4321 => x"88",
          4322 => x"a9",
          4323 => x"74",
          4324 => x"82",
          4325 => x"89",
          4326 => x"ff",
          4327 => x"80",
          4328 => x"3d",
          4329 => x"0c",
          4330 => x"55",
          4331 => x"17",
          4332 => x"76",
          4333 => x"fe",
          4334 => x"75",
          4335 => x"76",
          4336 => x"53",
          4337 => x"74",
          4338 => x"bb",
          4339 => x"ff",
          4340 => x"84",
          4341 => x"08",
          4342 => x"ff",
          4343 => x"76",
          4344 => x"0b",
          4345 => x"04",
          4346 => x"12",
          4347 => x"80",
          4348 => x"98",
          4349 => x"56",
          4350 => x"ff",
          4351 => x"94",
          4352 => x"79",
          4353 => x"74",
          4354 => x"18",
          4355 => x"b8",
          4356 => x"84",
          4357 => x"77",
          4358 => x"05",
          4359 => x"38",
          4360 => x"84",
          4361 => x"0b",
          4362 => x"81",
          4363 => x"c6",
          4364 => x"08",
          4365 => x"81",
          4366 => x"51",
          4367 => x"5d",
          4368 => x"2e",
          4369 => x"84",
          4370 => x"56",
          4371 => x"86",
          4372 => x"33",
          4373 => x"18",
          4374 => x"80",
          4375 => x"19",
          4376 => x"05",
          4377 => x"19",
          4378 => x"76",
          4379 => x"55",
          4380 => x"22",
          4381 => x"81",
          4382 => x"19",
          4383 => x"84",
          4384 => x"dd",
          4385 => x"84",
          4386 => x"75",
          4387 => x"70",
          4388 => x"86",
          4389 => x"38",
          4390 => x"b4",
          4391 => x"74",
          4392 => x"82",
          4393 => x"81",
          4394 => x"19",
          4395 => x"52",
          4396 => x"fe",
          4397 => x"83",
          4398 => x"09",
          4399 => x"0c",
          4400 => x"5e",
          4401 => x"85",
          4402 => x"b0",
          4403 => x"fc",
          4404 => x"0c",
          4405 => x"64",
          4406 => x"5b",
          4407 => x"5e",
          4408 => x"b8",
          4409 => x"19",
          4410 => x"19",
          4411 => x"09",
          4412 => x"75",
          4413 => x"51",
          4414 => x"80",
          4415 => x"79",
          4416 => x"90",
          4417 => x"58",
          4418 => x"18",
          4419 => x"5b",
          4420 => x"e5",
          4421 => x"30",
          4422 => x"54",
          4423 => x"74",
          4424 => x"2e",
          4425 => x"86",
          4426 => x"51",
          4427 => x"5b",
          4428 => x"98",
          4429 => x"7a",
          4430 => x"04",
          4431 => x"52",
          4432 => x"81",
          4433 => x"09",
          4434 => x"84",
          4435 => x"a8",
          4436 => x"58",
          4437 => x"b5",
          4438 => x"2e",
          4439 => x"54",
          4440 => x"53",
          4441 => x"de",
          4442 => x"8f",
          4443 => x"76",
          4444 => x"2e",
          4445 => x"bf",
          4446 => x"05",
          4447 => x"ab",
          4448 => x"cc",
          4449 => x"81",
          4450 => x"5b",
          4451 => x"bb",
          4452 => x"5b",
          4453 => x"7d",
          4454 => x"8c",
          4455 => x"33",
          4456 => x"75",
          4457 => x"bf",
          4458 => x"81",
          4459 => x"33",
          4460 => x"71",
          4461 => x"80",
          4462 => x"26",
          4463 => x"76",
          4464 => x"5a",
          4465 => x"38",
          4466 => x"59",
          4467 => x"81",
          4468 => x"61",
          4469 => x"70",
          4470 => x"39",
          4471 => x"81",
          4472 => x"38",
          4473 => x"75",
          4474 => x"05",
          4475 => x"ff",
          4476 => x"e4",
          4477 => x"ff",
          4478 => x"84",
          4479 => x"0d",
          4480 => x"7b",
          4481 => x"08",
          4482 => x"38",
          4483 => x"ac",
          4484 => x"08",
          4485 => x"2e",
          4486 => x"58",
          4487 => x"81",
          4488 => x"1b",
          4489 => x"3f",
          4490 => x"38",
          4491 => x"0c",
          4492 => x"1c",
          4493 => x"2e",
          4494 => x"06",
          4495 => x"86",
          4496 => x"f2",
          4497 => x"75",
          4498 => x"e2",
          4499 => x"7c",
          4500 => x"57",
          4501 => x"05",
          4502 => x"76",
          4503 => x"59",
          4504 => x"2e",
          4505 => x"06",
          4506 => x"1d",
          4507 => x"33",
          4508 => x"71",
          4509 => x"76",
          4510 => x"2e",
          4511 => x"ac",
          4512 => x"c8",
          4513 => x"bb",
          4514 => x"79",
          4515 => x"04",
          4516 => x"52",
          4517 => x"81",
          4518 => x"09",
          4519 => x"84",
          4520 => x"a8",
          4521 => x"58",
          4522 => x"ea",
          4523 => x"2e",
          4524 => x"54",
          4525 => x"53",
          4526 => x"b6",
          4527 => x"5a",
          4528 => x"86",
          4529 => x"f2",
          4530 => x"79",
          4531 => x"77",
          4532 => x"7f",
          4533 => x"7d",
          4534 => x"5d",
          4535 => x"84",
          4536 => x"08",
          4537 => x"39",
          4538 => x"ff",
          4539 => x"a2",
          4540 => x"2e",
          4541 => x"08",
          4542 => x"88",
          4543 => x"b3",
          4544 => x"29",
          4545 => x"56",
          4546 => x"81",
          4547 => x"07",
          4548 => x"ed",
          4549 => x"38",
          4550 => x"bb",
          4551 => x"22",
          4552 => x"a0",
          4553 => x"2e",
          4554 => x"56",
          4555 => x"b0",
          4556 => x"06",
          4557 => x"74",
          4558 => x"05",
          4559 => x"38",
          4560 => x"5a",
          4561 => x"84",
          4562 => x"ff",
          4563 => x"55",
          4564 => x"70",
          4565 => x"06",
          4566 => x"85",
          4567 => x"22",
          4568 => x"38",
          4569 => x"51",
          4570 => x"a0",
          4571 => x"58",
          4572 => x"77",
          4573 => x"55",
          4574 => x"33",
          4575 => x"2e",
          4576 => x"1f",
          4577 => x"8c",
          4578 => x"61",
          4579 => x"59",
          4580 => x"ff",
          4581 => x"27",
          4582 => x"57",
          4583 => x"1a",
          4584 => x"77",
          4585 => x"ff",
          4586 => x"44",
          4587 => x"38",
          4588 => x"18",
          4589 => x"22",
          4590 => x"05",
          4591 => x"07",
          4592 => x"38",
          4593 => x"16",
          4594 => x"56",
          4595 => x"fe",
          4596 => x"78",
          4597 => x"a0",
          4598 => x"78",
          4599 => x"33",
          4600 => x"06",
          4601 => x"77",
          4602 => x"05",
          4603 => x"59",
          4604 => x"87",
          4605 => x"84",
          4606 => x"5b",
          4607 => x"87",
          4608 => x"38",
          4609 => x"84",
          4610 => x"d6",
          4611 => x"1f",
          4612 => x"db",
          4613 => x"81",
          4614 => x"90",
          4615 => x"88",
          4616 => x"5b",
          4617 => x"84",
          4618 => x"08",
          4619 => x"b8",
          4620 => x"80",
          4621 => x"f3",
          4622 => x"2e",
          4623 => x"54",
          4624 => x"33",
          4625 => x"08",
          4626 => x"57",
          4627 => x"bc",
          4628 => x"42",
          4629 => x"74",
          4630 => x"5f",
          4631 => x"19",
          4632 => x"81",
          4633 => x"bb",
          4634 => x"80",
          4635 => x"84",
          4636 => x"81",
          4637 => x"f3",
          4638 => x"08",
          4639 => x"78",
          4640 => x"54",
          4641 => x"33",
          4642 => x"08",
          4643 => x"56",
          4644 => x"80",
          4645 => x"57",
          4646 => x"34",
          4647 => x"0b",
          4648 => x"75",
          4649 => x"81",
          4650 => x"ef",
          4651 => x"98",
          4652 => x"81",
          4653 => x"84",
          4654 => x"81",
          4655 => x"57",
          4656 => x"59",
          4657 => x"84",
          4658 => x"08",
          4659 => x"39",
          4660 => x"52",
          4661 => x"84",
          4662 => x"06",
          4663 => x"83",
          4664 => x"08",
          4665 => x"8b",
          4666 => x"2e",
          4667 => x"57",
          4668 => x"1f",
          4669 => x"e9",
          4670 => x"84",
          4671 => x"84",
          4672 => x"74",
          4673 => x"78",
          4674 => x"05",
          4675 => x"56",
          4676 => x"06",
          4677 => x"57",
          4678 => x"b2",
          4679 => x"2e",
          4680 => x"54",
          4681 => x"33",
          4682 => x"08",
          4683 => x"56",
          4684 => x"fe",
          4685 => x"08",
          4686 => x"60",
          4687 => x"34",
          4688 => x"34",
          4689 => x"f3",
          4690 => x"83",
          4691 => x"1f",
          4692 => x"83",
          4693 => x"76",
          4694 => x"88",
          4695 => x"38",
          4696 => x"8c",
          4697 => x"ff",
          4698 => x"70",
          4699 => x"a6",
          4700 => x"1d",
          4701 => x"3f",
          4702 => x"84",
          4703 => x"40",
          4704 => x"81",
          4705 => x"70",
          4706 => x"96",
          4707 => x"fc",
          4708 => x"1d",
          4709 => x"31",
          4710 => x"a0",
          4711 => x"1c",
          4712 => x"06",
          4713 => x"08",
          4714 => x"81",
          4715 => x"56",
          4716 => x"70",
          4717 => x"2e",
          4718 => x"ff",
          4719 => x"2e",
          4720 => x"80",
          4721 => x"54",
          4722 => x"1c",
          4723 => x"84",
          4724 => x"38",
          4725 => x"b4",
          4726 => x"74",
          4727 => x"1c",
          4728 => x"84",
          4729 => x"75",
          4730 => x"fa",
          4731 => x"57",
          4732 => x"75",
          4733 => x"39",
          4734 => x"08",
          4735 => x"51",
          4736 => x"54",
          4737 => x"53",
          4738 => x"96",
          4739 => x"7f",
          4740 => x"0b",
          4741 => x"2e",
          4742 => x"2e",
          4743 => x"8c",
          4744 => x"5c",
          4745 => x"54",
          4746 => x"55",
          4747 => x"80",
          4748 => x"5a",
          4749 => x"73",
          4750 => x"58",
          4751 => x"70",
          4752 => x"5c",
          4753 => x"0b",
          4754 => x"59",
          4755 => x"33",
          4756 => x"2e",
          4757 => x"38",
          4758 => x"07",
          4759 => x"26",
          4760 => x"ae",
          4761 => x"18",
          4762 => x"34",
          4763 => x"ba",
          4764 => x"0b",
          4765 => x"72",
          4766 => x"0b",
          4767 => x"94",
          4768 => x"9c",
          4769 => x"73",
          4770 => x"1c",
          4771 => x"34",
          4772 => x"33",
          4773 => x"88",
          4774 => x"07",
          4775 => x"0c",
          4776 => x"71",
          4777 => x"5a",
          4778 => x"99",
          4779 => x"2b",
          4780 => x"8f",
          4781 => x"c0",
          4782 => x"7a",
          4783 => x"7a",
          4784 => x"d0",
          4785 => x"ff",
          4786 => x"38",
          4787 => x"88",
          4788 => x"18",
          4789 => x"8c",
          4790 => x"11",
          4791 => x"90",
          4792 => x"30",
          4793 => x"25",
          4794 => x"38",
          4795 => x"80",
          4796 => x"39",
          4797 => x"57",
          4798 => x"96",
          4799 => x"33",
          4800 => x"26",
          4801 => x"33",
          4802 => x"72",
          4803 => x"7d",
          4804 => x"83",
          4805 => x"70",
          4806 => x"16",
          4807 => x"57",
          4808 => x"fd",
          4809 => x"39",
          4810 => x"30",
          4811 => x"a9",
          4812 => x"70",
          4813 => x"57",
          4814 => x"81",
          4815 => x"38",
          4816 => x"16",
          4817 => x"3d",
          4818 => x"27",
          4819 => x"08",
          4820 => x"05",
          4821 => x"38",
          4822 => x"ec",
          4823 => x"38",
          4824 => x"81",
          4825 => x"70",
          4826 => x"71",
          4827 => x"73",
          4828 => x"82",
          4829 => x"38",
          4830 => x"33",
          4831 => x"73",
          4832 => x"2e",
          4833 => x"81",
          4834 => x"38",
          4835 => x"84",
          4836 => x"38",
          4837 => x"81",
          4838 => x"33",
          4839 => x"f0",
          4840 => x"dc",
          4841 => x"07",
          4842 => x"a1",
          4843 => x"74",
          4844 => x"38",
          4845 => x"80",
          4846 => x"e1",
          4847 => x"96",
          4848 => x"9f",
          4849 => x"b5",
          4850 => x"84",
          4851 => x"54",
          4852 => x"84",
          4853 => x"83",
          4854 => x"5c",
          4855 => x"e4",
          4856 => x"80",
          4857 => x"bb",
          4858 => x"3d",
          4859 => x"70",
          4860 => x"55",
          4861 => x"81",
          4862 => x"55",
          4863 => x"80",
          4864 => x"78",
          4865 => x"73",
          4866 => x"5a",
          4867 => x"82",
          4868 => x"76",
          4869 => x"11",
          4870 => x"70",
          4871 => x"5f",
          4872 => x"72",
          4873 => x"38",
          4874 => x"23",
          4875 => x"78",
          4876 => x"58",
          4877 => x"e6",
          4878 => x"72",
          4879 => x"2e",
          4880 => x"22",
          4881 => x"76",
          4882 => x"57",
          4883 => x"70",
          4884 => x"81",
          4885 => x"55",
          4886 => x"34",
          4887 => x"73",
          4888 => x"81",
          4889 => x"2e",
          4890 => x"d0",
          4891 => x"80",
          4892 => x"85",
          4893 => x"59",
          4894 => x"75",
          4895 => x"80",
          4896 => x"54",
          4897 => x"8b",
          4898 => x"8a",
          4899 => x"26",
          4900 => x"7e",
          4901 => x"57",
          4902 => x"18",
          4903 => x"a0",
          4904 => x"83",
          4905 => x"38",
          4906 => x"82",
          4907 => x"83",
          4908 => x"81",
          4909 => x"06",
          4910 => x"90",
          4911 => x"5e",
          4912 => x"07",
          4913 => x"e4",
          4914 => x"1d",
          4915 => x"80",
          4916 => x"08",
          4917 => x"38",
          4918 => x"80",
          4919 => x"81",
          4920 => x"08",
          4921 => x"08",
          4922 => x"16",
          4923 => x"40",
          4924 => x"75",
          4925 => x"07",
          4926 => x"56",
          4927 => x"ac",
          4928 => x"09",
          4929 => x"18",
          4930 => x"1d",
          4931 => x"83",
          4932 => x"05",
          4933 => x"27",
          4934 => x"ab",
          4935 => x"84",
          4936 => x"54",
          4937 => x"74",
          4938 => x"ce",
          4939 => x"81",
          4940 => x"cd",
          4941 => x"60",
          4942 => x"12",
          4943 => x"41",
          4944 => x"d8",
          4945 => x"65",
          4946 => x"55",
          4947 => x"17",
          4948 => x"39",
          4949 => x"fd",
          4950 => x"06",
          4951 => x"2e",
          4952 => x"82",
          4953 => x"a0",
          4954 => x"06",
          4955 => x"0b",
          4956 => x"84",
          4957 => x"ff",
          4958 => x"80",
          4959 => x"26",
          4960 => x"77",
          4961 => x"79",
          4962 => x"51",
          4963 => x"08",
          4964 => x"81",
          4965 => x"38",
          4966 => x"11",
          4967 => x"ff",
          4968 => x"38",
          4969 => x"33",
          4970 => x"73",
          4971 => x"2e",
          4972 => x"81",
          4973 => x"38",
          4974 => x"d4",
          4975 => x"26",
          4976 => x"ff",
          4977 => x"78",
          4978 => x"70",
          4979 => x"ff",
          4980 => x"1b",
          4981 => x"1b",
          4982 => x"80",
          4983 => x"33",
          4984 => x"80",
          4985 => x"83",
          4986 => x"55",
          4987 => x"39",
          4988 => x"33",
          4989 => x"77",
          4990 => x"95",
          4991 => x"2a",
          4992 => x"7c",
          4993 => x"34",
          4994 => x"83",
          4995 => x"81",
          4996 => x"38",
          4997 => x"06",
          4998 => x"84",
          4999 => x"eb",
          5000 => x"80",
          5001 => x"61",
          5002 => x"42",
          5003 => x"70",
          5004 => x"56",
          5005 => x"74",
          5006 => x"38",
          5007 => x"24",
          5008 => x"e2",
          5009 => x"58",
          5010 => x"61",
          5011 => x"5d",
          5012 => x"17",
          5013 => x"bb",
          5014 => x"06",
          5015 => x"38",
          5016 => x"ba",
          5017 => x"52",
          5018 => x"3f",
          5019 => x"70",
          5020 => x"84",
          5021 => x"75",
          5022 => x"60",
          5023 => x"18",
          5024 => x"7b",
          5025 => x"17",
          5026 => x"ff",
          5027 => x"7b",
          5028 => x"74",
          5029 => x"38",
          5030 => x"33",
          5031 => x"56",
          5032 => x"38",
          5033 => x"f9",
          5034 => x"81",
          5035 => x"8d",
          5036 => x"80",
          5037 => x"71",
          5038 => x"80",
          5039 => x"80",
          5040 => x"71",
          5041 => x"38",
          5042 => x"12",
          5043 => x"07",
          5044 => x"2b",
          5045 => x"43",
          5046 => x"80",
          5047 => x"c8",
          5048 => x"06",
          5049 => x"26",
          5050 => x"76",
          5051 => x"5f",
          5052 => x"77",
          5053 => x"78",
          5054 => x"ca",
          5055 => x"88",
          5056 => x"23",
          5057 => x"58",
          5058 => x"33",
          5059 => x"07",
          5060 => x"17",
          5061 => x"90",
          5062 => x"33",
          5063 => x"71",
          5064 => x"42",
          5065 => x"33",
          5066 => x"58",
          5067 => x"1c",
          5068 => x"26",
          5069 => x"31",
          5070 => x"84",
          5071 => x"2e",
          5072 => x"80",
          5073 => x"83",
          5074 => x"38",
          5075 => x"eb",
          5076 => x"19",
          5077 => x"70",
          5078 => x"0c",
          5079 => x"38",
          5080 => x"80",
          5081 => x"18",
          5082 => x"8d",
          5083 => x"7a",
          5084 => x"15",
          5085 => x"18",
          5086 => x"18",
          5087 => x"80",
          5088 => x"86",
          5089 => x"dc",
          5090 => x"dc",
          5091 => x"e4",
          5092 => x"18",
          5093 => x"0c",
          5094 => x"bb",
          5095 => x"33",
          5096 => x"57",
          5097 => x"17",
          5098 => x"59",
          5099 => x"7e",
          5100 => x"7c",
          5101 => x"05",
          5102 => x"33",
          5103 => x"99",
          5104 => x"ff",
          5105 => x"77",
          5106 => x"81",
          5107 => x"9f",
          5108 => x"81",
          5109 => x"78",
          5110 => x"9f",
          5111 => x"80",
          5112 => x"1e",
          5113 => x"38",
          5114 => x"2e",
          5115 => x"06",
          5116 => x"80",
          5117 => x"57",
          5118 => x"06",
          5119 => x"32",
          5120 => x"5a",
          5121 => x"81",
          5122 => x"77",
          5123 => x"33",
          5124 => x"38",
          5125 => x"33",
          5126 => x"83",
          5127 => x"2b",
          5128 => x"59",
          5129 => x"84",
          5130 => x"57",
          5131 => x"84",
          5132 => x"9f",
          5133 => x"10",
          5134 => x"44",
          5135 => x"5b",
          5136 => x"38",
          5137 => x"b4",
          5138 => x"ff",
          5139 => x"b8",
          5140 => x"b4",
          5141 => x"2e",
          5142 => x"b4",
          5143 => x"81",
          5144 => x"07",
          5145 => x"d5",
          5146 => x"0b",
          5147 => x"e9",
          5148 => x"32",
          5149 => x"42",
          5150 => x"e8",
          5151 => x"ff",
          5152 => x"1e",
          5153 => x"81",
          5154 => x"27",
          5155 => x"b7",
          5156 => x"83",
          5157 => x"39",
          5158 => x"b4",
          5159 => x"5d",
          5160 => x"71",
          5161 => x"56",
          5162 => x"80",
          5163 => x"18",
          5164 => x"70",
          5165 => x"05",
          5166 => x"5b",
          5167 => x"8e",
          5168 => x"58",
          5169 => x"93",
          5170 => x"3d",
          5171 => x"fe",
          5172 => x"83",
          5173 => x"39",
          5174 => x"3d",
          5175 => x"83",
          5176 => x"81",
          5177 => x"5c",
          5178 => x"57",
          5179 => x"38",
          5180 => x"81",
          5181 => x"58",
          5182 => x"70",
          5183 => x"ff",
          5184 => x"2e",
          5185 => x"38",
          5186 => x"fc",
          5187 => x"80",
          5188 => x"71",
          5189 => x"2e",
          5190 => x"1b",
          5191 => x"2e",
          5192 => x"7a",
          5193 => x"81",
          5194 => x"17",
          5195 => x"bb",
          5196 => x"58",
          5197 => x"f9",
          5198 => x"b7",
          5199 => x"88",
          5200 => x"d5",
          5201 => x"b8",
          5202 => x"71",
          5203 => x"14",
          5204 => x"33",
          5205 => x"5c",
          5206 => x"2e",
          5207 => x"9c",
          5208 => x"71",
          5209 => x"14",
          5210 => x"33",
          5211 => x"5a",
          5212 => x"2e",
          5213 => x"a0",
          5214 => x"71",
          5215 => x"14",
          5216 => x"33",
          5217 => x"a4",
          5218 => x"71",
          5219 => x"14",
          5220 => x"33",
          5221 => x"44",
          5222 => x"56",
          5223 => x"22",
          5224 => x"23",
          5225 => x"0b",
          5226 => x"0c",
          5227 => x"f0",
          5228 => x"95",
          5229 => x"b8",
          5230 => x"59",
          5231 => x"08",
          5232 => x"38",
          5233 => x"b4",
          5234 => x"7f",
          5235 => x"17",
          5236 => x"38",
          5237 => x"39",
          5238 => x"38",
          5239 => x"b8",
          5240 => x"e3",
          5241 => x"88",
          5242 => x"f6",
          5243 => x"f6",
          5244 => x"33",
          5245 => x"88",
          5246 => x"07",
          5247 => x"1e",
          5248 => x"44",
          5249 => x"58",
          5250 => x"58",
          5251 => x"a8",
          5252 => x"59",
          5253 => x"da",
          5254 => x"17",
          5255 => x"52",
          5256 => x"3f",
          5257 => x"80",
          5258 => x"3d",
          5259 => x"75",
          5260 => x"81",
          5261 => x"55",
          5262 => x"ed",
          5263 => x"84",
          5264 => x"80",
          5265 => x"cc",
          5266 => x"2e",
          5267 => x"73",
          5268 => x"62",
          5269 => x"80",
          5270 => x"70",
          5271 => x"84",
          5272 => x"84",
          5273 => x"84",
          5274 => x"75",
          5275 => x"56",
          5276 => x"82",
          5277 => x"5c",
          5278 => x"80",
          5279 => x"5b",
          5280 => x"81",
          5281 => x"5a",
          5282 => x"76",
          5283 => x"81",
          5284 => x"57",
          5285 => x"70",
          5286 => x"70",
          5287 => x"09",
          5288 => x"38",
          5289 => x"07",
          5290 => x"79",
          5291 => x"1d",
          5292 => x"38",
          5293 => x"24",
          5294 => x"fe",
          5295 => x"84",
          5296 => x"89",
          5297 => x"bf",
          5298 => x"53",
          5299 => x"9f",
          5300 => x"bb",
          5301 => x"7a",
          5302 => x"0c",
          5303 => x"52",
          5304 => x"3f",
          5305 => x"84",
          5306 => x"9c",
          5307 => x"38",
          5308 => x"84",
          5309 => x"59",
          5310 => x"81",
          5311 => x"38",
          5312 => x"71",
          5313 => x"58",
          5314 => x"97",
          5315 => x"0b",
          5316 => x"34",
          5317 => x"56",
          5318 => x"57",
          5319 => x"0b",
          5320 => x"83",
          5321 => x"0b",
          5322 => x"34",
          5323 => x"9f",
          5324 => x"16",
          5325 => x"7e",
          5326 => x"57",
          5327 => x"9c",
          5328 => x"82",
          5329 => x"02",
          5330 => x"5c",
          5331 => x"86",
          5332 => x"b8",
          5333 => x"c2",
          5334 => x"5d",
          5335 => x"2a",
          5336 => x"38",
          5337 => x"38",
          5338 => x"80",
          5339 => x"59",
          5340 => x"67",
          5341 => x"9a",
          5342 => x"33",
          5343 => x"2e",
          5344 => x"9c",
          5345 => x"71",
          5346 => x"14",
          5347 => x"33",
          5348 => x"7f",
          5349 => x"86",
          5350 => x"1b",
          5351 => x"0b",
          5352 => x"0c",
          5353 => x"55",
          5354 => x"ff",
          5355 => x"2a",
          5356 => x"c9",
          5357 => x"2e",
          5358 => x"8a",
          5359 => x"08",
          5360 => x"70",
          5361 => x"76",
          5362 => x"06",
          5363 => x"38",
          5364 => x"3f",
          5365 => x"84",
          5366 => x"84",
          5367 => x"75",
          5368 => x"c2",
          5369 => x"38",
          5370 => x"80",
          5371 => x"7a",
          5372 => x"7a",
          5373 => x"7a",
          5374 => x"31",
          5375 => x"33",
          5376 => x"90",
          5377 => x"9c",
          5378 => x"71",
          5379 => x"14",
          5380 => x"33",
          5381 => x"61",
          5382 => x"5e",
          5383 => x"78",
          5384 => x"34",
          5385 => x"94",
          5386 => x"7c",
          5387 => x"cc",
          5388 => x"88",
          5389 => x"fb",
          5390 => x"aa",
          5391 => x"84",
          5392 => x"38",
          5393 => x"f7",
          5394 => x"82",
          5395 => x"51",
          5396 => x"08",
          5397 => x"11",
          5398 => x"75",
          5399 => x"0c",
          5400 => x"84",
          5401 => x"ff",
          5402 => x"59",
          5403 => x"af",
          5404 => x"2e",
          5405 => x"54",
          5406 => x"33",
          5407 => x"84",
          5408 => x"81",
          5409 => x"7b",
          5410 => x"80",
          5411 => x"f9",
          5412 => x"80",
          5413 => x"95",
          5414 => x"2b",
          5415 => x"56",
          5416 => x"0b",
          5417 => x"34",
          5418 => x"56",
          5419 => x"57",
          5420 => x"0b",
          5421 => x"83",
          5422 => x"ff",
          5423 => x"f8",
          5424 => x"78",
          5425 => x"19",
          5426 => x"59",
          5427 => x"19",
          5428 => x"05",
          5429 => x"38",
          5430 => x"0c",
          5431 => x"81",
          5432 => x"84",
          5433 => x"38",
          5434 => x"39",
          5435 => x"16",
          5436 => x"ff",
          5437 => x"7d",
          5438 => x"84",
          5439 => x"16",
          5440 => x"84",
          5441 => x"27",
          5442 => x"74",
          5443 => x"38",
          5444 => x"08",
          5445 => x"51",
          5446 => x"b6",
          5447 => x"7a",
          5448 => x"c5",
          5449 => x"64",
          5450 => x"89",
          5451 => x"08",
          5452 => x"33",
          5453 => x"16",
          5454 => x"78",
          5455 => x"5f",
          5456 => x"19",
          5457 => x"19",
          5458 => x"80",
          5459 => x"8c",
          5460 => x"75",
          5461 => x"81",
          5462 => x"7b",
          5463 => x"ff",
          5464 => x"7b",
          5465 => x"19",
          5466 => x"38",
          5467 => x"98",
          5468 => x"fe",
          5469 => x"57",
          5470 => x"18",
          5471 => x"05",
          5472 => x"38",
          5473 => x"7a",
          5474 => x"55",
          5475 => x"31",
          5476 => x"81",
          5477 => x"84",
          5478 => x"19",
          5479 => x"78",
          5480 => x"57",
          5481 => x"0c",
          5482 => x"59",
          5483 => x"d2",
          5484 => x"0c",
          5485 => x"84",
          5486 => x"fe",
          5487 => x"77",
          5488 => x"70",
          5489 => x"7b",
          5490 => x"53",
          5491 => x"9f",
          5492 => x"e3",
          5493 => x"55",
          5494 => x"54",
          5495 => x"51",
          5496 => x"08",
          5497 => x"94",
          5498 => x"84",
          5499 => x"27",
          5500 => x"17",
          5501 => x"2e",
          5502 => x"56",
          5503 => x"ff",
          5504 => x"38",
          5505 => x"70",
          5506 => x"75",
          5507 => x"08",
          5508 => x"84",
          5509 => x"81",
          5510 => x"84",
          5511 => x"fc",
          5512 => x"fc",
          5513 => x"56",
          5514 => x"80",
          5515 => x"58",
          5516 => x"77",
          5517 => x"55",
          5518 => x"70",
          5519 => x"05",
          5520 => x"38",
          5521 => x"34",
          5522 => x"3d",
          5523 => x"82",
          5524 => x"0d",
          5525 => x"65",
          5526 => x"89",
          5527 => x"08",
          5528 => x"33",
          5529 => x"16",
          5530 => x"78",
          5531 => x"40",
          5532 => x"19",
          5533 => x"19",
          5534 => x"58",
          5535 => x"38",
          5536 => x"7b",
          5537 => x"7a",
          5538 => x"ff",
          5539 => x"8a",
          5540 => x"06",
          5541 => x"f9",
          5542 => x"2e",
          5543 => x"ed",
          5544 => x"74",
          5545 => x"38",
          5546 => x"19",
          5547 => x"7a",
          5548 => x"fe",
          5549 => x"57",
          5550 => x"18",
          5551 => x"05",
          5552 => x"38",
          5553 => x"79",
          5554 => x"55",
          5555 => x"31",
          5556 => x"81",
          5557 => x"84",
          5558 => x"19",
          5559 => x"ab",
          5560 => x"72",
          5561 => x"70",
          5562 => x"05",
          5563 => x"38",
          5564 => x"7c",
          5565 => x"7a",
          5566 => x"78",
          5567 => x"94",
          5568 => x"58",
          5569 => x"75",
          5570 => x"fd",
          5571 => x"c0",
          5572 => x"56",
          5573 => x"0d",
          5574 => x"3d",
          5575 => x"a2",
          5576 => x"1a",
          5577 => x"53",
          5578 => x"ff",
          5579 => x"81",
          5580 => x"9c",
          5581 => x"80",
          5582 => x"83",
          5583 => x"05",
          5584 => x"93",
          5585 => x"75",
          5586 => x"56",
          5587 => x"80",
          5588 => x"c7",
          5589 => x"ff",
          5590 => x"55",
          5591 => x"90",
          5592 => x"52",
          5593 => x"bb",
          5594 => x"fc",
          5595 => x"19",
          5596 => x"33",
          5597 => x"84",
          5598 => x"ff",
          5599 => x"58",
          5600 => x"ff",
          5601 => x"81",
          5602 => x"79",
          5603 => x"0b",
          5604 => x"84",
          5605 => x"91",
          5606 => x"0c",
          5607 => x"7d",
          5608 => x"38",
          5609 => x"38",
          5610 => x"38",
          5611 => x"5a",
          5612 => x"55",
          5613 => x"38",
          5614 => x"06",
          5615 => x"38",
          5616 => x"83",
          5617 => x"56",
          5618 => x"80",
          5619 => x"5a",
          5620 => x"c0",
          5621 => x"52",
          5622 => x"3f",
          5623 => x"38",
          5624 => x"0c",
          5625 => x"18",
          5626 => x"57",
          5627 => x"19",
          5628 => x"5a",
          5629 => x"2a",
          5630 => x"76",
          5631 => x"83",
          5632 => x"55",
          5633 => x"7a",
          5634 => x"75",
          5635 => x"78",
          5636 => x"0b",
          5637 => x"34",
          5638 => x"0b",
          5639 => x"34",
          5640 => x"7b",
          5641 => x"84",
          5642 => x"5b",
          5643 => x"74",
          5644 => x"04",
          5645 => x"16",
          5646 => x"ff",
          5647 => x"84",
          5648 => x"c0",
          5649 => x"34",
          5650 => x"84",
          5651 => x"17",
          5652 => x"33",
          5653 => x"fd",
          5654 => x"a0",
          5655 => x"16",
          5656 => x"59",
          5657 => x"74",
          5658 => x"75",
          5659 => x"74",
          5660 => x"9d",
          5661 => x"9e",
          5662 => x"9f",
          5663 => x"97",
          5664 => x"80",
          5665 => x"92",
          5666 => x"7b",
          5667 => x"51",
          5668 => x"08",
          5669 => x"56",
          5670 => x"81",
          5671 => x"84",
          5672 => x"fc",
          5673 => x"fc",
          5674 => x"53",
          5675 => x"52",
          5676 => x"84",
          5677 => x"18",
          5678 => x"19",
          5679 => x"b4",
          5680 => x"fc",
          5681 => x"0d",
          5682 => x"84",
          5683 => x"08",
          5684 => x"9e",
          5685 => x"96",
          5686 => x"8e",
          5687 => x"58",
          5688 => x"52",
          5689 => x"75",
          5690 => x"89",
          5691 => x"ff",
          5692 => x"81",
          5693 => x"08",
          5694 => x"ff",
          5695 => x"2e",
          5696 => x"33",
          5697 => x"2e",
          5698 => x"2e",
          5699 => x"80",
          5700 => x"e0",
          5701 => x"8c",
          5702 => x"84",
          5703 => x"d0",
          5704 => x"53",
          5705 => x"73",
          5706 => x"73",
          5707 => x"83",
          5708 => x"56",
          5709 => x"75",
          5710 => x"12",
          5711 => x"38",
          5712 => x"54",
          5713 => x"89",
          5714 => x"54",
          5715 => x"51",
          5716 => x"38",
          5717 => x"70",
          5718 => x"07",
          5719 => x"38",
          5720 => x"78",
          5721 => x"cf",
          5722 => x"76",
          5723 => x"0d",
          5724 => x"99",
          5725 => x"84",
          5726 => x"2e",
          5727 => x"98",
          5728 => x"98",
          5729 => x"84",
          5730 => x"08",
          5731 => x"33",
          5732 => x"24",
          5733 => x"70",
          5734 => x"80",
          5735 => x"33",
          5736 => x"73",
          5737 => x"83",
          5738 => x"74",
          5739 => x"04",
          5740 => x"81",
          5741 => x"bb",
          5742 => x"16",
          5743 => x"71",
          5744 => x"0c",
          5745 => x"12",
          5746 => x"98",
          5747 => x"80",
          5748 => x"5d",
          5749 => x"e4",
          5750 => x"3d",
          5751 => x"08",
          5752 => x"38",
          5753 => x"98",
          5754 => x"80",
          5755 => x"2e",
          5756 => x"3d",
          5757 => x"a5",
          5758 => x"84",
          5759 => x"80",
          5760 => x"08",
          5761 => x"08",
          5762 => x"c7",
          5763 => x"52",
          5764 => x"3f",
          5765 => x"38",
          5766 => x"0c",
          5767 => x"08",
          5768 => x"88",
          5769 => x"59",
          5770 => x"38",
          5771 => x"7a",
          5772 => x"84",
          5773 => x"9f",
          5774 => x"b4",
          5775 => x"bb",
          5776 => x"08",
          5777 => x"88",
          5778 => x"59",
          5779 => x"38",
          5780 => x"84",
          5781 => x"3f",
          5782 => x"84",
          5783 => x"84",
          5784 => x"38",
          5785 => x"7a",
          5786 => x"82",
          5787 => x"90",
          5788 => x"17",
          5789 => x"38",
          5790 => x"95",
          5791 => x"17",
          5792 => x"3d",
          5793 => x"59",
          5794 => x"eb",
          5795 => x"11",
          5796 => x"3d",
          5797 => x"60",
          5798 => x"e2",
          5799 => x"f4",
          5800 => x"59",
          5801 => x"81",
          5802 => x"5a",
          5803 => x"78",
          5804 => x"27",
          5805 => x"7c",
          5806 => x"57",
          5807 => x"70",
          5808 => x"09",
          5809 => x"80",
          5810 => x"80",
          5811 => x"94",
          5812 => x"2b",
          5813 => x"f0",
          5814 => x"71",
          5815 => x"07",
          5816 => x"52",
          5817 => x"bb",
          5818 => x"80",
          5819 => x"81",
          5820 => x"70",
          5821 => x"8a",
          5822 => x"08",
          5823 => x"83",
          5824 => x"08",
          5825 => x"74",
          5826 => x"82",
          5827 => x"81",
          5828 => x"16",
          5829 => x"52",
          5830 => x"3f",
          5831 => x"80",
          5832 => x"7b",
          5833 => x"70",
          5834 => x"08",
          5835 => x"7e",
          5836 => x"38",
          5837 => x"18",
          5838 => x"70",
          5839 => x"fe",
          5840 => x"81",
          5841 => x"81",
          5842 => x"38",
          5843 => x"34",
          5844 => x"3d",
          5845 => x"5a",
          5846 => x"38",
          5847 => x"38",
          5848 => x"38",
          5849 => x"5b",
          5850 => x"55",
          5851 => x"38",
          5852 => x"38",
          5853 => x"82",
          5854 => x"5a",
          5855 => x"8a",
          5856 => x"58",
          5857 => x"52",
          5858 => x"84",
          5859 => x"70",
          5860 => x"84",
          5861 => x"38",
          5862 => x"0c",
          5863 => x"5a",
          5864 => x"77",
          5865 => x"31",
          5866 => x"90",
          5867 => x"51",
          5868 => x"38",
          5869 => x"3f",
          5870 => x"84",
          5871 => x"2e",
          5872 => x"82",
          5873 => x"27",
          5874 => x"ff",
          5875 => x"94",
          5876 => x"83",
          5877 => x"38",
          5878 => x"05",
          5879 => x"ca",
          5880 => x"b0",
          5881 => x"5c",
          5882 => x"38",
          5883 => x"56",
          5884 => x"18",
          5885 => x"59",
          5886 => x"06",
          5887 => x"9c",
          5888 => x"a1",
          5889 => x"a8",
          5890 => x"a2",
          5891 => x"7b",
          5892 => x"86",
          5893 => x"90",
          5894 => x"90",
          5895 => x"52",
          5896 => x"84",
          5897 => x"2e",
          5898 => x"34",
          5899 => x"8d",
          5900 => x"81",
          5901 => x"82",
          5902 => x"80",
          5903 => x"fc",
          5904 => x"d4",
          5905 => x"17",
          5906 => x"38",
          5907 => x"fe",
          5908 => x"18",
          5909 => x"8d",
          5910 => x"ff",
          5911 => x"56",
          5912 => x"ff",
          5913 => x"81",
          5914 => x"77",
          5915 => x"52",
          5916 => x"bb",
          5917 => x"81",
          5918 => x"ff",
          5919 => x"08",
          5920 => x"ff",
          5921 => x"82",
          5922 => x"0d",
          5923 => x"54",
          5924 => x"8c",
          5925 => x"05",
          5926 => x"08",
          5927 => x"8f",
          5928 => x"84",
          5929 => x"7a",
          5930 => x"ba",
          5931 => x"84",
          5932 => x"16",
          5933 => x"78",
          5934 => x"84",
          5935 => x"2e",
          5936 => x"11",
          5937 => x"07",
          5938 => x"57",
          5939 => x"17",
          5940 => x"17",
          5941 => x"aa",
          5942 => x"84",
          5943 => x"84",
          5944 => x"85",
          5945 => x"95",
          5946 => x"2b",
          5947 => x"19",
          5948 => x"3d",
          5949 => x"2e",
          5950 => x"2e",
          5951 => x"2e",
          5952 => x"22",
          5953 => x"80",
          5954 => x"75",
          5955 => x"3d",
          5956 => x"80",
          5957 => x"06",
          5958 => x"53",
          5959 => x"7c",
          5960 => x"9f",
          5961 => x"97",
          5962 => x"8f",
          5963 => x"59",
          5964 => x"80",
          5965 => x"c7",
          5966 => x"75",
          5967 => x"84",
          5968 => x"08",
          5969 => x"08",
          5970 => x"b3",
          5971 => x"9a",
          5972 => x"32",
          5973 => x"84",
          5974 => x"72",
          5975 => x"04",
          5976 => x"b2",
          5977 => x"99",
          5978 => x"32",
          5979 => x"84",
          5980 => x"cf",
          5981 => x"ea",
          5982 => x"84",
          5983 => x"33",
          5984 => x"84",
          5985 => x"38",
          5986 => x"39",
          5987 => x"89",
          5988 => x"c2",
          5989 => x"84",
          5990 => x"74",
          5991 => x"04",
          5992 => x"3f",
          5993 => x"84",
          5994 => x"33",
          5995 => x"24",
          5996 => x"76",
          5997 => x"74",
          5998 => x"04",
          5999 => x"3d",
          6000 => x"56",
          6001 => x"52",
          6002 => x"bb",
          6003 => x"9a",
          6004 => x"11",
          6005 => x"57",
          6006 => x"75",
          6007 => x"95",
          6008 => x"77",
          6009 => x"93",
          6010 => x"84",
          6011 => x"38",
          6012 => x"b4",
          6013 => x"83",
          6014 => x"8d",
          6015 => x"52",
          6016 => x"3f",
          6017 => x"38",
          6018 => x"0c",
          6019 => x"38",
          6020 => x"8d",
          6021 => x"33",
          6022 => x"88",
          6023 => x"07",
          6024 => x"ff",
          6025 => x"80",
          6026 => x"ff",
          6027 => x"53",
          6028 => x"78",
          6029 => x"94",
          6030 => x"58",
          6031 => x"84",
          6032 => x"b4",
          6033 => x"81",
          6034 => x"3f",
          6035 => x"f8",
          6036 => x"34",
          6037 => x"84",
          6038 => x"18",
          6039 => x"33",
          6040 => x"fe",
          6041 => x"a0",
          6042 => x"17",
          6043 => x"5e",
          6044 => x"3d",
          6045 => x"81",
          6046 => x"2e",
          6047 => x"81",
          6048 => x"08",
          6049 => x"80",
          6050 => x"58",
          6051 => x"ca",
          6052 => x"0c",
          6053 => x"84",
          6054 => x"b8",
          6055 => x"88",
          6056 => x"1f",
          6057 => x"5f",
          6058 => x"fd",
          6059 => x"fd",
          6060 => x"7f",
          6061 => x"33",
          6062 => x"fe",
          6063 => x"39",
          6064 => x"77",
          6065 => x"75",
          6066 => x"74",
          6067 => x"84",
          6068 => x"82",
          6069 => x"81",
          6070 => x"80",
          6071 => x"2a",
          6072 => x"80",
          6073 => x"55",
          6074 => x"38",
          6075 => x"78",
          6076 => x"38",
          6077 => x"38",
          6078 => x"94",
          6079 => x"c0",
          6080 => x"a8",
          6081 => x"25",
          6082 => x"53",
          6083 => x"52",
          6084 => x"84",
          6085 => x"57",
          6086 => x"84",
          6087 => x"79",
          6088 => x"74",
          6089 => x"84",
          6090 => x"08",
          6091 => x"84",
          6092 => x"bb",
          6093 => x"80",
          6094 => x"cb",
          6095 => x"38",
          6096 => x"08",
          6097 => x"af",
          6098 => x"17",
          6099 => x"34",
          6100 => x"38",
          6101 => x"f7",
          6102 => x"06",
          6103 => x"08",
          6104 => x"90",
          6105 => x"0b",
          6106 => x"18",
          6107 => x"3f",
          6108 => x"c2",
          6109 => x"81",
          6110 => x"59",
          6111 => x"27",
          6112 => x"98",
          6113 => x"81",
          6114 => x"a1",
          6115 => x"08",
          6116 => x"97",
          6117 => x"ff",
          6118 => x"56",
          6119 => x"74",
          6120 => x"84",
          6121 => x"08",
          6122 => x"84",
          6123 => x"bb",
          6124 => x"80",
          6125 => x"d3",
          6126 => x"38",
          6127 => x"08",
          6128 => x"38",
          6129 => x"33",
          6130 => x"79",
          6131 => x"80",
          6132 => x"fc",
          6133 => x"82",
          6134 => x"bf",
          6135 => x"33",
          6136 => x"34",
          6137 => x"90",
          6138 => x"84",
          6139 => x"55",
          6140 => x"33",
          6141 => x"84",
          6142 => x"ff",
          6143 => x"a7",
          6144 => x"51",
          6145 => x"08",
          6146 => x"8a",
          6147 => x"3d",
          6148 => x"52",
          6149 => x"b1",
          6150 => x"bb",
          6151 => x"05",
          6152 => x"57",
          6153 => x"2b",
          6154 => x"80",
          6155 => x"57",
          6156 => x"a3",
          6157 => x"33",
          6158 => x"5e",
          6159 => x"d5",
          6160 => x"76",
          6161 => x"98",
          6162 => x"77",
          6163 => x"52",
          6164 => x"b2",
          6165 => x"bb",
          6166 => x"84",
          6167 => x"3f",
          6168 => x"84",
          6169 => x"84",
          6170 => x"33",
          6171 => x"90",
          6172 => x"ff",
          6173 => x"2e",
          6174 => x"a1",
          6175 => x"57",
          6176 => x"38",
          6177 => x"3f",
          6178 => x"84",
          6179 => x"70",
          6180 => x"80",
          6181 => x"38",
          6182 => x"27",
          6183 => x"81",
          6184 => x"38",
          6185 => x"bb",
          6186 => x"3d",
          6187 => x"08",
          6188 => x"2e",
          6189 => x"59",
          6190 => x"80",
          6191 => x"17",
          6192 => x"a7",
          6193 => x"85",
          6194 => x"18",
          6195 => x"19",
          6196 => x"83",
          6197 => x"fe",
          6198 => x"8c",
          6199 => x"84",
          6200 => x"38",
          6201 => x"cd",
          6202 => x"54",
          6203 => x"17",
          6204 => x"58",
          6205 => x"81",
          6206 => x"08",
          6207 => x"18",
          6208 => x"55",
          6209 => x"38",
          6210 => x"09",
          6211 => x"b4",
          6212 => x"7c",
          6213 => x"fe",
          6214 => x"55",
          6215 => x"52",
          6216 => x"bb",
          6217 => x"80",
          6218 => x"08",
          6219 => x"84",
          6220 => x"53",
          6221 => x"3f",
          6222 => x"17",
          6223 => x"5c",
          6224 => x"81",
          6225 => x"81",
          6226 => x"55",
          6227 => x"56",
          6228 => x"39",
          6229 => x"39",
          6230 => x"0d",
          6231 => x"52",
          6232 => x"84",
          6233 => x"08",
          6234 => x"84",
          6235 => x"6f",
          6236 => x"a6",
          6237 => x"84",
          6238 => x"84",
          6239 => x"84",
          6240 => x"06",
          6241 => x"70",
          6242 => x"56",
          6243 => x"52",
          6244 => x"f9",
          6245 => x"5c",
          6246 => x"56",
          6247 => x"f9",
          6248 => x"81",
          6249 => x"84",
          6250 => x"5a",
          6251 => x"9c",
          6252 => x"5b",
          6253 => x"22",
          6254 => x"5c",
          6255 => x"59",
          6256 => x"70",
          6257 => x"74",
          6258 => x"55",
          6259 => x"54",
          6260 => x"33",
          6261 => x"84",
          6262 => x"dc",
          6263 => x"54",
          6264 => x"53",
          6265 => x"de",
          6266 => x"be",
          6267 => x"34",
          6268 => x"55",
          6269 => x"38",
          6270 => x"09",
          6271 => x"b4",
          6272 => x"77",
          6273 => x"9e",
          6274 => x"7d",
          6275 => x"b4",
          6276 => x"ac",
          6277 => x"b2",
          6278 => x"bb",
          6279 => x"84",
          6280 => x"38",
          6281 => x"84",
          6282 => x"fe",
          6283 => x"fc",
          6284 => x"94",
          6285 => x"27",
          6286 => x"84",
          6287 => x"18",
          6288 => x"a1",
          6289 => x"3d",
          6290 => x"83",
          6291 => x"78",
          6292 => x"8b",
          6293 => x"70",
          6294 => x"75",
          6295 => x"18",
          6296 => x"19",
          6297 => x"34",
          6298 => x"80",
          6299 => x"d1",
          6300 => x"06",
          6301 => x"77",
          6302 => x"34",
          6303 => x"cc",
          6304 => x"1a",
          6305 => x"81",
          6306 => x"59",
          6307 => x"7d",
          6308 => x"64",
          6309 => x"57",
          6310 => x"88",
          6311 => x"75",
          6312 => x"38",
          6313 => x"79",
          6314 => x"84",
          6315 => x"b6",
          6316 => x"96",
          6317 => x"17",
          6318 => x"cc",
          6319 => x"5d",
          6320 => x"59",
          6321 => x"79",
          6322 => x"90",
          6323 => x"0b",
          6324 => x"b9",
          6325 => x"84",
          6326 => x"76",
          6327 => x"34",
          6328 => x"17",
          6329 => x"5b",
          6330 => x"2a",
          6331 => x"59",
          6332 => x"57",
          6333 => x"2a",
          6334 => x"2a",
          6335 => x"90",
          6336 => x"0b",
          6337 => x"d1",
          6338 => x"96",
          6339 => x"3d",
          6340 => x"2e",
          6341 => x"33",
          6342 => x"2e",
          6343 => x"ba",
          6344 => x"3d",
          6345 => x"ff",
          6346 => x"56",
          6347 => x"38",
          6348 => x"0d",
          6349 => x"08",
          6350 => x"9f",
          6351 => x"84",
          6352 => x"bb",
          6353 => x"56",
          6354 => x"ae",
          6355 => x"81",
          6356 => x"59",
          6357 => x"99",
          6358 => x"55",
          6359 => x"70",
          6360 => x"74",
          6361 => x"51",
          6362 => x"08",
          6363 => x"38",
          6364 => x"38",
          6365 => x"3d",
          6366 => x"81",
          6367 => x"26",
          6368 => x"06",
          6369 => x"80",
          6370 => x"f4",
          6371 => x"5c",
          6372 => x"70",
          6373 => x"5a",
          6374 => x"e0",
          6375 => x"ff",
          6376 => x"38",
          6377 => x"55",
          6378 => x"75",
          6379 => x"77",
          6380 => x"30",
          6381 => x"5d",
          6382 => x"81",
          6383 => x"24",
          6384 => x"5b",
          6385 => x"b4",
          6386 => x"3d",
          6387 => x"ff",
          6388 => x"56",
          6389 => x"fd",
          6390 => x"09",
          6391 => x"ff",
          6392 => x"56",
          6393 => x"6f",
          6394 => x"05",
          6395 => x"70",
          6396 => x"05",
          6397 => x"38",
          6398 => x"34",
          6399 => x"06",
          6400 => x"07",
          6401 => x"81",
          6402 => x"70",
          6403 => x"80",
          6404 => x"6b",
          6405 => x"33",
          6406 => x"72",
          6407 => x"2e",
          6408 => x"08",
          6409 => x"82",
          6410 => x"29",
          6411 => x"80",
          6412 => x"58",
          6413 => x"83",
          6414 => x"81",
          6415 => x"17",
          6416 => x"bb",
          6417 => x"58",
          6418 => x"57",
          6419 => x"fb",
          6420 => x"ae",
          6421 => x"70",
          6422 => x"80",
          6423 => x"77",
          6424 => x"7a",
          6425 => x"75",
          6426 => x"34",
          6427 => x"18",
          6428 => x"34",
          6429 => x"08",
          6430 => x"38",
          6431 => x"3f",
          6432 => x"84",
          6433 => x"98",
          6434 => x"08",
          6435 => x"7a",
          6436 => x"06",
          6437 => x"b8",
          6438 => x"e2",
          6439 => x"2e",
          6440 => x"b4",
          6441 => x"9c",
          6442 => x"0b",
          6443 => x"27",
          6444 => x"fc",
          6445 => x"84",
          6446 => x"38",
          6447 => x"38",
          6448 => x"51",
          6449 => x"08",
          6450 => x"04",
          6451 => x"3d",
          6452 => x"33",
          6453 => x"78",
          6454 => x"84",
          6455 => x"38",
          6456 => x"a0",
          6457 => x"3d",
          6458 => x"53",
          6459 => x"e2",
          6460 => x"08",
          6461 => x"38",
          6462 => x"b4",
          6463 => x"bb",
          6464 => x"08",
          6465 => x"5d",
          6466 => x"93",
          6467 => x"17",
          6468 => x"33",
          6469 => x"fd",
          6470 => x"53",
          6471 => x"52",
          6472 => x"84",
          6473 => x"bb",
          6474 => x"08",
          6475 => x"08",
          6476 => x"fc",
          6477 => x"82",
          6478 => x"81",
          6479 => x"05",
          6480 => x"fe",
          6481 => x"39",
          6482 => x"33",
          6483 => x"56",
          6484 => x"52",
          6485 => x"84",
          6486 => x"08",
          6487 => x"84",
          6488 => x"66",
          6489 => x"97",
          6490 => x"84",
          6491 => x"cf",
          6492 => x"56",
          6493 => x"71",
          6494 => x"74",
          6495 => x"8b",
          6496 => x"16",
          6497 => x"84",
          6498 => x"96",
          6499 => x"57",
          6500 => x"97",
          6501 => x"bb",
          6502 => x"80",
          6503 => x"0c",
          6504 => x"52",
          6505 => x"91",
          6506 => x"bb",
          6507 => x"05",
          6508 => x"75",
          6509 => x"19",
          6510 => x"56",
          6511 => x"55",
          6512 => x"58",
          6513 => x"54",
          6514 => x"0b",
          6515 => x"c1",
          6516 => x"84",
          6517 => x"0d",
          6518 => x"3d",
          6519 => x"a0",
          6520 => x"bb",
          6521 => x"08",
          6522 => x"80",
          6523 => x"5a",
          6524 => x"70",
          6525 => x"80",
          6526 => x"06",
          6527 => x"38",
          6528 => x"5a",
          6529 => x"38",
          6530 => x"7a",
          6531 => x"81",
          6532 => x"16",
          6533 => x"bb",
          6534 => x"57",
          6535 => x"57",
          6536 => x"58",
          6537 => x"38",
          6538 => x"38",
          6539 => x"11",
          6540 => x"71",
          6541 => x"72",
          6542 => x"62",
          6543 => x"76",
          6544 => x"04",
          6545 => x"3d",
          6546 => x"84",
          6547 => x"08",
          6548 => x"2e",
          6549 => x"7b",
          6550 => x"54",
          6551 => x"53",
          6552 => x"e6",
          6553 => x"7a",
          6554 => x"84",
          6555 => x"16",
          6556 => x"84",
          6557 => x"27",
          6558 => x"74",
          6559 => x"38",
          6560 => x"08",
          6561 => x"51",
          6562 => x"54",
          6563 => x"33",
          6564 => x"84",
          6565 => x"86",
          6566 => x"f4",
          6567 => x"bb",
          6568 => x"84",
          6569 => x"59",
          6570 => x"57",
          6571 => x"19",
          6572 => x"70",
          6573 => x"80",
          6574 => x"11",
          6575 => x"2e",
          6576 => x"fd",
          6577 => x"a1",
          6578 => x"51",
          6579 => x"08",
          6580 => x"38",
          6581 => x"a0",
          6582 => x"15",
          6583 => x"08",
          6584 => x"58",
          6585 => x"38",
          6586 => x"81",
          6587 => x"81",
          6588 => x"ff",
          6589 => x"a1",
          6590 => x"84",
          6591 => x"84",
          6592 => x"80",
          6593 => x"0b",
          6594 => x"06",
          6595 => x"d6",
          6596 => x"38",
          6597 => x"06",
          6598 => x"38",
          6599 => x"38",
          6600 => x"a3",
          6601 => x"38",
          6602 => x"ff",
          6603 => x"55",
          6604 => x"81",
          6605 => x"5d",
          6606 => x"33",
          6607 => x"5a",
          6608 => x"3d",
          6609 => x"2e",
          6610 => x"02",
          6611 => x"5c",
          6612 => x"87",
          6613 => x"7d",
          6614 => x"70",
          6615 => x"bb",
          6616 => x"80",
          6617 => x"bb",
          6618 => x"b5",
          6619 => x"bb",
          6620 => x"74",
          6621 => x"bb",
          6622 => x"e8",
          6623 => x"52",
          6624 => x"bb",
          6625 => x"80",
          6626 => x"38",
          6627 => x"70",
          6628 => x"05",
          6629 => x"38",
          6630 => x"7d",
          6631 => x"84",
          6632 => x"8a",
          6633 => x"ff",
          6634 => x"2e",
          6635 => x"55",
          6636 => x"08",
          6637 => x"ea",
          6638 => x"bb",
          6639 => x"81",
          6640 => x"19",
          6641 => x"59",
          6642 => x"83",
          6643 => x"81",
          6644 => x"53",
          6645 => x"fe",
          6646 => x"80",
          6647 => x"76",
          6648 => x"38",
          6649 => x"5a",
          6650 => x"38",
          6651 => x"56",
          6652 => x"81",
          6653 => x"81",
          6654 => x"84",
          6655 => x"08",
          6656 => x"76",
          6657 => x"76",
          6658 => x"80",
          6659 => x"15",
          6660 => x"0b",
          6661 => x"57",
          6662 => x"76",
          6663 => x"55",
          6664 => x"70",
          6665 => x"05",
          6666 => x"38",
          6667 => x"34",
          6668 => x"7d",
          6669 => x"84",
          6670 => x"fe",
          6671 => x"53",
          6672 => x"d5",
          6673 => x"2e",
          6674 => x"bb",
          6675 => x"08",
          6676 => x"19",
          6677 => x"55",
          6678 => x"84",
          6679 => x"81",
          6680 => x"84",
          6681 => x"08",
          6682 => x"39",
          6683 => x"fd",
          6684 => x"b4",
          6685 => x"7a",
          6686 => x"b6",
          6687 => x"60",
          6688 => x"33",
          6689 => x"2e",
          6690 => x"2e",
          6691 => x"2e",
          6692 => x"22",
          6693 => x"38",
          6694 => x"38",
          6695 => x"38",
          6696 => x"17",
          6697 => x"70",
          6698 => x"80",
          6699 => x"22",
          6700 => x"57",
          6701 => x"15",
          6702 => x"9f",
          6703 => x"1c",
          6704 => x"81",
          6705 => x"78",
          6706 => x"56",
          6707 => x"fe",
          6708 => x"55",
          6709 => x"82",
          6710 => x"81",
          6711 => x"2e",
          6712 => x"81",
          6713 => x"2e",
          6714 => x"06",
          6715 => x"84",
          6716 => x"87",
          6717 => x"0d",
          6718 => x"e5",
          6719 => x"54",
          6720 => x"55",
          6721 => x"81",
          6722 => x"80",
          6723 => x"81",
          6724 => x"52",
          6725 => x"bb",
          6726 => x"ff",
          6727 => x"57",
          6728 => x"90",
          6729 => x"8c",
          6730 => x"18",
          6731 => x"5c",
          6732 => x"fe",
          6733 => x"7a",
          6734 => x"94",
          6735 => x"5d",
          6736 => x"d6",
          6737 => x"5b",
          6738 => x"fe",
          6739 => x"ff",
          6740 => x"90",
          6741 => x"a5",
          6742 => x"05",
          6743 => x"3d",
          6744 => x"2e",
          6745 => x"5b",
          6746 => x"ba",
          6747 => x"75",
          6748 => x"e0",
          6749 => x"38",
          6750 => x"70",
          6751 => x"38",
          6752 => x"f8",
          6753 => x"40",
          6754 => x"ce",
          6755 => x"ff",
          6756 => x"57",
          6757 => x"81",
          6758 => x"38",
          6759 => x"79",
          6760 => x"84",
          6761 => x"80",
          6762 => x"80",
          6763 => x"06",
          6764 => x"2e",
          6765 => x"f8",
          6766 => x"f0",
          6767 => x"83",
          6768 => x"08",
          6769 => x"4c",
          6770 => x"38",
          6771 => x"56",
          6772 => x"7d",
          6773 => x"74",
          6774 => x"f7",
          6775 => x"83",
          6776 => x"61",
          6777 => x"07",
          6778 => x"d5",
          6779 => x"7d",
          6780 => x"33",
          6781 => x"38",
          6782 => x"12",
          6783 => x"07",
          6784 => x"2b",
          6785 => x"83",
          6786 => x"2b",
          6787 => x"70",
          6788 => x"07",
          6789 => x"0c",
          6790 => x"59",
          6791 => x"57",
          6792 => x"93",
          6793 => x"38",
          6794 => x"49",
          6795 => x"87",
          6796 => x"61",
          6797 => x"83",
          6798 => x"58",
          6799 => x"ae",
          6800 => x"83",
          6801 => x"2e",
          6802 => x"83",
          6803 => x"70",
          6804 => x"86",
          6805 => x"52",
          6806 => x"bb",
          6807 => x"bb",
          6808 => x"81",
          6809 => x"bb",
          6810 => x"83",
          6811 => x"89",
          6812 => x"1f",
          6813 => x"05",
          6814 => x"57",
          6815 => x"74",
          6816 => x"60",
          6817 => x"f2",
          6818 => x"53",
          6819 => x"89",
          6820 => x"83",
          6821 => x"09",
          6822 => x"f5",
          6823 => x"ac",
          6824 => x"55",
          6825 => x"74",
          6826 => x"84",
          6827 => x"bb",
          6828 => x"39",
          6829 => x"3d",
          6830 => x"33",
          6831 => x"57",
          6832 => x"1d",
          6833 => x"58",
          6834 => x"0b",
          6835 => x"7d",
          6836 => x"33",
          6837 => x"9f",
          6838 => x"89",
          6839 => x"58",
          6840 => x"26",
          6841 => x"06",
          6842 => x"5a",
          6843 => x"85",
          6844 => x"32",
          6845 => x"7b",
          6846 => x"80",
          6847 => x"5c",
          6848 => x"56",
          6849 => x"53",
          6850 => x"3f",
          6851 => x"b6",
          6852 => x"bb",
          6853 => x"bf",
          6854 => x"26",
          6855 => x"fb",
          6856 => x"7b",
          6857 => x"a3",
          6858 => x"81",
          6859 => x"fd",
          6860 => x"46",
          6861 => x"08",
          6862 => x"38",
          6863 => x"fb",
          6864 => x"84",
          6865 => x"0c",
          6866 => x"99",
          6867 => x"74",
          6868 => x"ae",
          6869 => x"76",
          6870 => x"55",
          6871 => x"c0",
          6872 => x"58",
          6873 => x"ff",
          6874 => x"05",
          6875 => x"05",
          6876 => x"83",
          6877 => x"05",
          6878 => x"8f",
          6879 => x"62",
          6880 => x"61",
          6881 => x"06",
          6882 => x"56",
          6883 => x"38",
          6884 => x"61",
          6885 => x"6b",
          6886 => x"05",
          6887 => x"61",
          6888 => x"34",
          6889 => x"9c",
          6890 => x"61",
          6891 => x"6b",
          6892 => x"84",
          6893 => x"61",
          6894 => x"f7",
          6895 => x"61",
          6896 => x"34",
          6897 => x"83",
          6898 => x"05",
          6899 => x"97",
          6900 => x"34",
          6901 => x"ab",
          6902 => x"76",
          6903 => x"81",
          6904 => x"ef",
          6905 => x"d5",
          6906 => x"ff",
          6907 => x"60",
          6908 => x"81",
          6909 => x"38",
          6910 => x"9c",
          6911 => x"70",
          6912 => x"74",
          6913 => x"83",
          6914 => x"f8",
          6915 => x"57",
          6916 => x"45",
          6917 => x"34",
          6918 => x"81",
          6919 => x"75",
          6920 => x"66",
          6921 => x"7a",
          6922 => x"d6",
          6923 => x"38",
          6924 => x"70",
          6925 => x"74",
          6926 => x"58",
          6927 => x"40",
          6928 => x"56",
          6929 => x"65",
          6930 => x"55",
          6931 => x"51",
          6932 => x"08",
          6933 => x"31",
          6934 => x"62",
          6935 => x"83",
          6936 => x"62",
          6937 => x"84",
          6938 => x"5e",
          6939 => x"56",
          6940 => x"34",
          6941 => x"d5",
          6942 => x"83",
          6943 => x"67",
          6944 => x"34",
          6945 => x"84",
          6946 => x"52",
          6947 => x"fe",
          6948 => x"08",
          6949 => x"86",
          6950 => x"87",
          6951 => x"34",
          6952 => x"61",
          6953 => x"08",
          6954 => x"83",
          6955 => x"64",
          6956 => x"2a",
          6957 => x"62",
          6958 => x"05",
          6959 => x"79",
          6960 => x"84",
          6961 => x"53",
          6962 => x"3f",
          6963 => x"b6",
          6964 => x"84",
          6965 => x"0c",
          6966 => x"1c",
          6967 => x"7a",
          6968 => x"0b",
          6969 => x"80",
          6970 => x"38",
          6971 => x"17",
          6972 => x"2e",
          6973 => x"77",
          6974 => x"84",
          6975 => x"05",
          6976 => x"80",
          6977 => x"8a",
          6978 => x"77",
          6979 => x"e4",
          6980 => x"f5",
          6981 => x"38",
          6982 => x"38",
          6983 => x"06",
          6984 => x"83",
          6985 => x"05",
          6986 => x"a1",
          6987 => x"61",
          6988 => x"76",
          6989 => x"80",
          6990 => x"80",
          6991 => x"05",
          6992 => x"34",
          6993 => x"2a",
          6994 => x"90",
          6995 => x"7c",
          6996 => x"34",
          6997 => x"ad",
          6998 => x"80",
          6999 => x"05",
          7000 => x"61",
          7001 => x"34",
          7002 => x"a9",
          7003 => x"80",
          7004 => x"55",
          7005 => x"70",
          7006 => x"74",
          7007 => x"81",
          7008 => x"58",
          7009 => x"f9",
          7010 => x"52",
          7011 => x"57",
          7012 => x"7d",
          7013 => x"83",
          7014 => x"84",
          7015 => x"bf",
          7016 => x"84",
          7017 => x"bb",
          7018 => x"4a",
          7019 => x"ff",
          7020 => x"6a",
          7021 => x"61",
          7022 => x"34",
          7023 => x"88",
          7024 => x"ff",
          7025 => x"7c",
          7026 => x"1f",
          7027 => x"8e",
          7028 => x"75",
          7029 => x"57",
          7030 => x"7c",
          7031 => x"80",
          7032 => x"80",
          7033 => x"80",
          7034 => x"e4",
          7035 => x"05",
          7036 => x"34",
          7037 => x"7f",
          7038 => x"05",
          7039 => x"83",
          7040 => x"75",
          7041 => x"2a",
          7042 => x"82",
          7043 => x"83",
          7044 => x"05",
          7045 => x"80",
          7046 => x"81",
          7047 => x"51",
          7048 => x"1f",
          7049 => x"de",
          7050 => x"39",
          7051 => x"80",
          7052 => x"76",
          7053 => x"8e",
          7054 => x"52",
          7055 => x"81",
          7056 => x"3d",
          7057 => x"74",
          7058 => x"17",
          7059 => x"77",
          7060 => x"55",
          7061 => x"bb",
          7062 => x"3d",
          7063 => x"33",
          7064 => x"38",
          7065 => x"9e",
          7066 => x"05",
          7067 => x"55",
          7068 => x"18",
          7069 => x"3d",
          7070 => x"74",
          7071 => x"ff",
          7072 => x"30",
          7073 => x"84",
          7074 => x"5a",
          7075 => x"51",
          7076 => x"3d",
          7077 => x"3d",
          7078 => x"80",
          7079 => x"15",
          7080 => x"77",
          7081 => x"7c",
          7082 => x"7d",
          7083 => x"75",
          7084 => x"b8",
          7085 => x"88",
          7086 => x"9e",
          7087 => x"75",
          7088 => x"ff",
          7089 => x"86",
          7090 => x"0b",
          7091 => x"04",
          7092 => x"54",
          7093 => x"9d",
          7094 => x"70",
          7095 => x"5a",
          7096 => x"76",
          7097 => x"7d",
          7098 => x"04",
          7099 => x"9a",
          7100 => x"80",
          7101 => x"ff",
          7102 => x"85",
          7103 => x"27",
          7104 => x"06",
          7105 => x"83",
          7106 => x"9c",
          7107 => x"06",
          7108 => x"38",
          7109 => x"22",
          7110 => x"70",
          7111 => x"53",
          7112 => x"02",
          7113 => x"05",
          7114 => x"ff",
          7115 => x"bb",
          7116 => x"83",
          7117 => x"70",
          7118 => x"83",
          7119 => x"84",
          7120 => x"3d",
          7121 => x"26",
          7122 => x"06",
          7123 => x"ff",
          7124 => x"05",
          7125 => x"25",
          7126 => x"53",
          7127 => x"53",
          7128 => x"81",
          7129 => x"76",
          7130 => x"10",
          7131 => x"54",
          7132 => x"26",
          7133 => x"cb",
          7134 => x"0c",
          7135 => x"55",
          7136 => x"38",
          7137 => x"54",
          7138 => x"83",
          7139 => x"d3",
          7140 => x"ff",
          7141 => x"70",
          7142 => x"39",
          7143 => x"57",
          7144 => x"ff",
          7145 => x"16",
          7146 => x"c5",
          7147 => x"06",
          7148 => x"31",
          7149 => x"ff",
          7150 => x"39",
          7151 => x"22",
          7152 => x"00",
          7153 => x"ff",
          7154 => x"00",
          7155 => x"80",
          7156 => x"6a",
          7157 => x"54",
          7158 => x"3e",
          7159 => x"28",
          7160 => x"12",
          7161 => x"fc",
          7162 => x"e6",
          7163 => x"d0",
          7164 => x"ba",
          7165 => x"64",
          7166 => x"64",
          7167 => x"64",
          7168 => x"64",
          7169 => x"64",
          7170 => x"64",
          7171 => x"64",
          7172 => x"64",
          7173 => x"64",
          7174 => x"64",
          7175 => x"64",
          7176 => x"64",
          7177 => x"64",
          7178 => x"64",
          7179 => x"64",
          7180 => x"64",
          7181 => x"64",
          7182 => x"64",
          7183 => x"64",
          7184 => x"64",
          7185 => x"64",
          7186 => x"81",
          7187 => x"64",
          7188 => x"64",
          7189 => x"64",
          7190 => x"64",
          7191 => x"64",
          7192 => x"64",
          7193 => x"64",
          7194 => x"64",
          7195 => x"16",
          7196 => x"9a",
          7197 => x"77",
          7198 => x"de",
          7199 => x"64",
          7200 => x"64",
          7201 => x"64",
          7202 => x"64",
          7203 => x"64",
          7204 => x"64",
          7205 => x"64",
          7206 => x"64",
          7207 => x"64",
          7208 => x"64",
          7209 => x"64",
          7210 => x"64",
          7211 => x"64",
          7212 => x"64",
          7213 => x"64",
          7214 => x"64",
          7215 => x"64",
          7216 => x"64",
          7217 => x"64",
          7218 => x"64",
          7219 => x"64",
          7220 => x"64",
          7221 => x"64",
          7222 => x"64",
          7223 => x"64",
          7224 => x"64",
          7225 => x"80",
          7226 => x"64",
          7227 => x"64",
          7228 => x"64",
          7229 => x"64",
          7230 => x"68",
          7231 => x"50",
          7232 => x"61",
          7233 => x"49",
          7234 => x"4b",
          7235 => x"63",
          7236 => x"3f",
          7237 => x"9a",
          7238 => x"90",
          7239 => x"fd",
          7240 => x"b5",
          7241 => x"e4",
          7242 => x"8b",
          7243 => x"62",
          7244 => x"fc",
          7245 => x"fd",
          7246 => x"e4",
          7247 => x"90",
          7248 => x"5d",
          7249 => x"a3",
          7250 => x"c8",
          7251 => x"6d",
          7252 => x"2a",
          7253 => x"2a",
          7254 => x"2a",
          7255 => x"2a",
          7256 => x"2a",
          7257 => x"2a",
          7258 => x"2a",
          7259 => x"2a",
          7260 => x"2a",
          7261 => x"2a",
          7262 => x"2a",
          7263 => x"2a",
          7264 => x"2a",
          7265 => x"2a",
          7266 => x"42",
          7267 => x"1d",
          7268 => x"34",
          7269 => x"e5",
          7270 => x"2a",
          7271 => x"d5",
          7272 => x"7e",
          7273 => x"c3",
          7274 => x"9f",
          7275 => x"2a",
          7276 => x"d0",
          7277 => x"11",
          7278 => x"45",
          7279 => x"fa",
          7280 => x"51",
          7281 => x"93",
          7282 => x"51",
          7283 => x"51",
          7284 => x"51",
          7285 => x"7b",
          7286 => x"51",
          7287 => x"51",
          7288 => x"51",
          7289 => x"51",
          7290 => x"51",
          7291 => x"51",
          7292 => x"51",
          7293 => x"51",
          7294 => x"51",
          7295 => x"51",
          7296 => x"51",
          7297 => x"51",
          7298 => x"a1",
          7299 => x"51",
          7300 => x"51",
          7301 => x"28",
          7302 => x"0b",
          7303 => x"e9",
          7304 => x"e9",
          7305 => x"e9",
          7306 => x"c4",
          7307 => x"e9",
          7308 => x"e9",
          7309 => x"e9",
          7310 => x"e9",
          7311 => x"e9",
          7312 => x"e9",
          7313 => x"e9",
          7314 => x"e9",
          7315 => x"e9",
          7316 => x"e9",
          7317 => x"e9",
          7318 => x"ce",
          7319 => x"a8",
          7320 => x"59",
          7321 => x"36",
          7322 => x"26",
          7323 => x"04",
          7324 => x"e0",
          7325 => x"40",
          7326 => x"18",
          7327 => x"62",
          7328 => x"9f",
          7329 => x"9f",
          7330 => x"9f",
          7331 => x"9f",
          7332 => x"9f",
          7333 => x"9f",
          7334 => x"9f",
          7335 => x"9f",
          7336 => x"9f",
          7337 => x"9f",
          7338 => x"8d",
          7339 => x"9f",
          7340 => x"9f",
          7341 => x"a0",
          7342 => x"74",
          7343 => x"55",
          7344 => x"3f",
          7345 => x"29",
          7346 => x"0f",
          7347 => x"fd",
          7348 => x"49",
          7349 => x"fd",
          7350 => x"fd",
          7351 => x"fd",
          7352 => x"fd",
          7353 => x"7f",
          7354 => x"fd",
          7355 => x"fd",
          7356 => x"fd",
          7357 => x"fd",
          7358 => x"fd",
          7359 => x"fd",
          7360 => x"fd",
          7361 => x"fd",
          7362 => x"fd",
          7363 => x"fd",
          7364 => x"fd",
          7365 => x"fd",
          7366 => x"fd",
          7367 => x"fd",
          7368 => x"fd",
          7369 => x"fd",
          7370 => x"fd",
          7371 => x"fd",
          7372 => x"1d",
          7373 => x"fd",
          7374 => x"fd",
          7375 => x"fd",
          7376 => x"fd",
          7377 => x"fd",
          7378 => x"fd",
          7379 => x"fd",
          7380 => x"2b",
          7381 => x"b8",
          7382 => x"b8",
          7383 => x"e1",
          7384 => x"fd",
          7385 => x"fd",
          7386 => x"16",
          7387 => x"fd",
          7388 => x"58",
          7389 => x"18",
          7390 => x"fd",
          7391 => x"69",
          7392 => x"63",
          7393 => x"69",
          7394 => x"61",
          7395 => x"65",
          7396 => x"65",
          7397 => x"70",
          7398 => x"66",
          7399 => x"6d",
          7400 => x"00",
          7401 => x"00",
          7402 => x"00",
          7403 => x"00",
          7404 => x"00",
          7405 => x"74",
          7406 => x"65",
          7407 => x"6f",
          7408 => x"74",
          7409 => x"00",
          7410 => x"73",
          7411 => x"73",
          7412 => x"6f",
          7413 => x"00",
          7414 => x"20",
          7415 => x"00",
          7416 => x"65",
          7417 => x"72",
          7418 => x"00",
          7419 => x"79",
          7420 => x"69",
          7421 => x"00",
          7422 => x"63",
          7423 => x"6d",
          7424 => x"00",
          7425 => x"20",
          7426 => x"00",
          7427 => x"2c",
          7428 => x"69",
          7429 => x"65",
          7430 => x"00",
          7431 => x"61",
          7432 => x"00",
          7433 => x"61",
          7434 => x"69",
          7435 => x"6d",
          7436 => x"6f",
          7437 => x"00",
          7438 => x"74",
          7439 => x"64",
          7440 => x"76",
          7441 => x"72",
          7442 => x"61",
          7443 => x"00",
          7444 => x"72",
          7445 => x"74",
          7446 => x"00",
          7447 => x"6e",
          7448 => x"61",
          7449 => x"00",
          7450 => x"72",
          7451 => x"69",
          7452 => x"00",
          7453 => x"64",
          7454 => x"00",
          7455 => x"20",
          7456 => x"65",
          7457 => x"70",
          7458 => x"6e",
          7459 => x"66",
          7460 => x"6e",
          7461 => x"6b",
          7462 => x"61",
          7463 => x"65",
          7464 => x"72",
          7465 => x"6b",
          7466 => x"00",
          7467 => x"2e",
          7468 => x"75",
          7469 => x"25",
          7470 => x"75",
          7471 => x"73",
          7472 => x"00",
          7473 => x"00",
          7474 => x"00",
          7475 => x"58",
          7476 => x"00",
          7477 => x"00",
          7478 => x"00",
          7479 => x"20",
          7480 => x"00",
          7481 => x"00",
          7482 => x"30",
          7483 => x"33",
          7484 => x"55",
          7485 => x"30",
          7486 => x"25",
          7487 => x"00",
          7488 => x"20",
          7489 => x"64",
          7490 => x"20",
          7491 => x"20",
          7492 => x"78",
          7493 => x"20",
          7494 => x"72",
          7495 => x"20",
          7496 => x"20",
          7497 => x"78",
          7498 => x"20",
          7499 => x"70",
          7500 => x"65",
          7501 => x"54",
          7502 => x"74",
          7503 => x"00",
          7504 => x"58",
          7505 => x"75",
          7506 => x"54",
          7507 => x"74",
          7508 => x"00",
          7509 => x"58",
          7510 => x"75",
          7511 => x"54",
          7512 => x"74",
          7513 => x"00",
          7514 => x"44",
          7515 => x"75",
          7516 => x"20",
          7517 => x"70",
          7518 => x"65",
          7519 => x"72",
          7520 => x"74",
          7521 => x"74",
          7522 => x"00",
          7523 => x"67",
          7524 => x"2e",
          7525 => x"6f",
          7526 => x"74",
          7527 => x"5f",
          7528 => x"00",
          7529 => x"74",
          7530 => x"61",
          7531 => x"20",
          7532 => x"20",
          7533 => x"69",
          7534 => x"75",
          7535 => x"00",
          7536 => x"5c",
          7537 => x"00",
          7538 => x"6d",
          7539 => x"00",
          7540 => x"00",
          7541 => x"25",
          7542 => x"00",
          7543 => x"62",
          7544 => x"2e",
          7545 => x"74",
          7546 => x"61",
          7547 => x"69",
          7548 => x"00",
          7549 => x"20",
          7550 => x"25",
          7551 => x"2e",
          7552 => x"6c",
          7553 => x"65",
          7554 => x"28",
          7555 => x"00",
          7556 => x"6e",
          7557 => x"40",
          7558 => x"2e",
          7559 => x"6c",
          7560 => x"2d",
          7561 => x"6c",
          7562 => x"00",
          7563 => x"6e",
          7564 => x"00",
          7565 => x"30",
          7566 => x"38",
          7567 => x"29",
          7568 => x"79",
          7569 => x"00",
          7570 => x"30",
          7571 => x"61",
          7572 => x"2e",
          7573 => x"70",
          7574 => x"00",
          7575 => x"74",
          7576 => x"5c",
          7577 => x"00",
          7578 => x"65",
          7579 => x"64",
          7580 => x"74",
          7581 => x"73",
          7582 => x"64",
          7583 => x"00",
          7584 => x"64",
          7585 => x"25",
          7586 => x"00",
          7587 => x"66",
          7588 => x"6f",
          7589 => x"65",
          7590 => x"6d",
          7591 => x"65",
          7592 => x"72",
          7593 => x"00",
          7594 => x"20",
          7595 => x"65",
          7596 => x"64",
          7597 => x"25",
          7598 => x"00",
          7599 => x"20",
          7600 => x"53",
          7601 => x"64",
          7602 => x"25",
          7603 => x"00",
          7604 => x"63",
          7605 => x"20",
          7606 => x"20",
          7607 => x"25",
          7608 => x"00",
          7609 => x"00",
          7610 => x"20",
          7611 => x"20",
          7612 => x"20",
          7613 => x"25",
          7614 => x"00",
          7615 => x"74",
          7616 => x"6b",
          7617 => x"20",
          7618 => x"25",
          7619 => x"48",
          7620 => x"20",
          7621 => x"65",
          7622 => x"43",
          7623 => x"65",
          7624 => x"30",
          7625 => x"00",
          7626 => x"41",
          7627 => x"20",
          7628 => x"20",
          7629 => x"25",
          7630 => x"48",
          7631 => x"20",
          7632 => x"20",
          7633 => x"20",
          7634 => x"00",
          7635 => x"49",
          7636 => x"20",
          7637 => x"45",
          7638 => x"00",
          7639 => x"52",
          7640 => x"43",
          7641 => x"3d",
          7642 => x"00",
          7643 => x"45",
          7644 => x"54",
          7645 => x"3d",
          7646 => x"00",
          7647 => x"43",
          7648 => x"44",
          7649 => x"3d",
          7650 => x"00",
          7651 => x"20",
          7652 => x"25",
          7653 => x"58",
          7654 => x"20",
          7655 => x"20",
          7656 => x"3a",
          7657 => x"00",
          7658 => x"4e",
          7659 => x"25",
          7660 => x"58",
          7661 => x"20",
          7662 => x"20",
          7663 => x"3a",
          7664 => x"00",
          7665 => x"53",
          7666 => x"25",
          7667 => x"58",
          7668 => x"72",
          7669 => x"63",
          7670 => x"00",
          7671 => x"00",
          7672 => x"00",
          7673 => x"00",
          7674 => x"00",
          7675 => x"00",
          7676 => x"3c",
          7677 => x"02",
          7678 => x"00",
          7679 => x"34",
          7680 => x"04",
          7681 => x"00",
          7682 => x"2c",
          7683 => x"06",
          7684 => x"00",
          7685 => x"24",
          7686 => x"01",
          7687 => x"00",
          7688 => x"1c",
          7689 => x"0b",
          7690 => x"00",
          7691 => x"14",
          7692 => x"0a",
          7693 => x"00",
          7694 => x"0c",
          7695 => x"0c",
          7696 => x"00",
          7697 => x"04",
          7698 => x"0f",
          7699 => x"00",
          7700 => x"fc",
          7701 => x"10",
          7702 => x"00",
          7703 => x"f4",
          7704 => x"12",
          7705 => x"00",
          7706 => x"ec",
          7707 => x"14",
          7708 => x"00",
          7709 => x"00",
          7710 => x"00",
          7711 => x"7e",
          7712 => x"7e",
          7713 => x"7e",
          7714 => x"7e",
          7715 => x"00",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"74",
          7721 => x"70",
          7722 => x"00",
          7723 => x"6f",
          7724 => x"61",
          7725 => x"6f",
          7726 => x"2c",
          7727 => x"69",
          7728 => x"74",
          7729 => x"74",
          7730 => x"00",
          7731 => x"20",
          7732 => x"25",
          7733 => x"00",
          7734 => x"25",
          7735 => x"6c",
          7736 => x"65",
          7737 => x"20",
          7738 => x"20",
          7739 => x"20",
          7740 => x"00",
          7741 => x"00",
          7742 => x"00",
          7743 => x"00",
          7744 => x"00",
          7745 => x"00",
          7746 => x"00",
          7747 => x"00",
          7748 => x"00",
          7749 => x"00",
          7750 => x"00",
          7751 => x"00",
          7752 => x"00",
          7753 => x"00",
          7754 => x"00",
          7755 => x"00",
          7756 => x"00",
          7757 => x"7e",
          7758 => x"7e",
          7759 => x"64",
          7760 => x"25",
          7761 => x"3a",
          7762 => x"00",
          7763 => x"2d",
          7764 => x"64",
          7765 => x"00",
          7766 => x"64",
          7767 => x"78",
          7768 => x"25",
          7769 => x"00",
          7770 => x"43",
          7771 => x"00",
          7772 => x"20",
          7773 => x"00",
          7774 => x"20",
          7775 => x"00",
          7776 => x"20",
          7777 => x"74",
          7778 => x"69",
          7779 => x"00",
          7780 => x"3c",
          7781 => x"00",
          7782 => x"00",
          7783 => x"33",
          7784 => x"4d",
          7785 => x"00",
          7786 => x"20",
          7787 => x"20",
          7788 => x"4e",
          7789 => x"46",
          7790 => x"00",
          7791 => x"00",
          7792 => x"00",
          7793 => x"12",
          7794 => x"00",
          7795 => x"80",
          7796 => x"8f",
          7797 => x"55",
          7798 => x"9f",
          7799 => x"a7",
          7800 => x"af",
          7801 => x"b7",
          7802 => x"bf",
          7803 => x"c7",
          7804 => x"cf",
          7805 => x"d7",
          7806 => x"df",
          7807 => x"e7",
          7808 => x"ef",
          7809 => x"f7",
          7810 => x"ff",
          7811 => x"2f",
          7812 => x"7c",
          7813 => x"04",
          7814 => x"00",
          7815 => x"02",
          7816 => x"20",
          7817 => x"fc",
          7818 => x"e0",
          7819 => x"eb",
          7820 => x"ec",
          7821 => x"e6",
          7822 => x"f2",
          7823 => x"d6",
          7824 => x"a5",
          7825 => x"ed",
          7826 => x"d1",
          7827 => x"10",
          7828 => x"a1",
          7829 => x"92",
          7830 => x"61",
          7831 => x"63",
          7832 => x"5c",
          7833 => x"34",
          7834 => x"3c",
          7835 => x"54",
          7836 => x"50",
          7837 => x"64",
          7838 => x"52",
          7839 => x"18",
          7840 => x"8c",
          7841 => x"df",
          7842 => x"c3",
          7843 => x"98",
          7844 => x"c6",
          7845 => x"b1",
          7846 => x"21",
          7847 => x"19",
          7848 => x"b2",
          7849 => x"1a",
          7850 => x"07",
          7851 => x"00",
          7852 => x"39",
          7853 => x"79",
          7854 => x"43",
          7855 => x"84",
          7856 => x"87",
          7857 => x"8b",
          7858 => x"90",
          7859 => x"94",
          7860 => x"98",
          7861 => x"9c",
          7862 => x"a0",
          7863 => x"a4",
          7864 => x"a7",
          7865 => x"ac",
          7866 => x"af",
          7867 => x"b3",
          7868 => x"b8",
          7869 => x"bc",
          7870 => x"c0",
          7871 => x"c4",
          7872 => x"c8",
          7873 => x"ca",
          7874 => x"01",
          7875 => x"f3",
          7876 => x"f4",
          7877 => x"12",
          7878 => x"3b",
          7879 => x"3f",
          7880 => x"46",
          7881 => x"81",
          7882 => x"8a",
          7883 => x"90",
          7884 => x"5f",
          7885 => x"94",
          7886 => x"67",
          7887 => x"62",
          7888 => x"9c",
          7889 => x"73",
          7890 => x"77",
          7891 => x"7b",
          7892 => x"7f",
          7893 => x"a9",
          7894 => x"87",
          7895 => x"b2",
          7896 => x"8f",
          7897 => x"7b",
          7898 => x"ff",
          7899 => x"88",
          7900 => x"11",
          7901 => x"a3",
          7902 => x"03",
          7903 => x"d8",
          7904 => x"f9",
          7905 => x"f6",
          7906 => x"fa",
          7907 => x"50",
          7908 => x"8a",
          7909 => x"cf",
          7910 => x"44",
          7911 => x"00",
          7912 => x"00",
          7913 => x"00",
          7914 => x"20",
          7915 => x"40",
          7916 => x"59",
          7917 => x"5d",
          7918 => x"08",
          7919 => x"bb",
          7920 => x"cb",
          7921 => x"f9",
          7922 => x"fb",
          7923 => x"08",
          7924 => x"04",
          7925 => x"bc",
          7926 => x"d0",
          7927 => x"e5",
          7928 => x"01",
          7929 => x"32",
          7930 => x"01",
          7931 => x"30",
          7932 => x"67",
          7933 => x"80",
          7934 => x"41",
          7935 => x"00",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"00",
          7940 => x"00",
          7941 => x"00",
          7942 => x"00",
          7943 => x"00",
          7944 => x"00",
          7945 => x"00",
          7946 => x"00",
          7947 => x"00",
          7948 => x"00",
          7949 => x"00",
          7950 => x"00",
          7951 => x"00",
          7952 => x"00",
          7953 => x"00",
          7954 => x"00",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"00",
          7959 => x"00",
          7960 => x"00",
          7961 => x"00",
          7962 => x"00",
          7963 => x"00",
          7964 => x"00",
          7965 => x"00",
          7966 => x"00",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"00",
          7983 => x"00",
          7984 => x"00",
          7985 => x"00",
          7986 => x"00",
          7987 => x"00",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"00",
          7996 => x"00",
          7997 => x"00",
          7998 => x"00",
          7999 => x"00",
          8000 => x"00",
          8001 => x"01",
          8002 => x"01",
          8003 => x"00",
          8004 => x"00",
          8005 => x"00",
          8006 => x"00",
          8007 => x"00",
          8008 => x"00",
          8009 => x"00",
          8010 => x"00",
          8011 => x"00",
          8012 => x"00",
          8013 => x"00",
          8014 => x"00",
          8015 => x"80",
          8016 => x"88",
          8017 => x"90",
          8018 => x"80",
          8019 => x"0d",
          8020 => x"f0",
          8021 => x"78",
          8022 => x"70",
          8023 => x"68",
          8024 => x"38",
          8025 => x"2e",
          8026 => x"2f",
          8027 => x"f0",
          8028 => x"f0",
          8029 => x"0d",
          8030 => x"f0",
          8031 => x"58",
          8032 => x"50",
          8033 => x"48",
          8034 => x"38",
          8035 => x"2e",
          8036 => x"2f",
          8037 => x"f0",
          8038 => x"f0",
          8039 => x"0d",
          8040 => x"f0",
          8041 => x"58",
          8042 => x"50",
          8043 => x"48",
          8044 => x"28",
          8045 => x"3e",
          8046 => x"2f",
          8047 => x"f0",
          8048 => x"f0",
          8049 => x"f0",
          8050 => x"f0",
          8051 => x"18",
          8052 => x"10",
          8053 => x"08",
          8054 => x"f0",
          8055 => x"f0",
          8056 => x"1c",
          8057 => x"f0",
          8058 => x"f0",
          8059 => x"cd",
          8060 => x"f0",
          8061 => x"dd",
          8062 => x"b1",
          8063 => x"73",
          8064 => x"a2",
          8065 => x"b9",
          8066 => x"be",
          8067 => x"f0",
          8068 => x"f0",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"f3",
          9105 => x"fb",
          9106 => x"c3",
          9107 => x"e6",
          9108 => x"63",
          9109 => x"6a",
          9110 => x"23",
          9111 => x"2c",
          9112 => x"03",
          9113 => x"0b",
          9114 => x"13",
          9115 => x"52",
          9116 => x"83",
          9117 => x"8b",
          9118 => x"93",
          9119 => x"bc",
          9120 => x"00",
          9121 => x"00",
          9122 => x"00",
          9123 => x"00",
          9124 => x"00",
          9125 => x"00",
          9126 => x"00",
          9127 => x"00",
          9128 => x"00",
          9129 => x"00",
          9130 => x"00",
          9131 => x"00",
          9132 => x"00",
          9133 => x"00",
          9134 => x"00",
          9135 => x"03",
          9136 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"87",
             1 => x"e9",
             2 => x"00",
             3 => x"00",
             4 => x"8c",
             5 => x"90",
             6 => x"00",
             7 => x"00",
             8 => x"06",
             9 => x"82",
            10 => x"06",
            11 => x"00",
            12 => x"06",
            13 => x"09",
            14 => x"09",
            15 => x"0b",
            16 => x"81",
            17 => x"09",
            18 => x"81",
            19 => x"00",
            20 => x"24",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"05",
            26 => x"0a",
            27 => x"53",
            28 => x"26",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"9f",
            45 => x"93",
            46 => x"00",
            47 => x"00",
            48 => x"2a",
            49 => x"09",
            50 => x"53",
            51 => x"00",
            52 => x"53",
            53 => x"81",
            54 => x"07",
            55 => x"00",
            56 => x"81",
            57 => x"09",
            58 => x"00",
            59 => x"00",
            60 => x"81",
            61 => x"09",
            62 => x"04",
            63 => x"00",
            64 => x"81",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"09",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"72",
            73 => x"51",
            74 => x"00",
            75 => x"00",
            76 => x"06",
            77 => x"83",
            78 => x"06",
            79 => x"00",
            80 => x"06",
            81 => x"83",
            82 => x"0b",
            83 => x"00",
            84 => x"8c",
            85 => x"0b",
            86 => x"56",
            87 => x"04",
            88 => x"8c",
            89 => x"0b",
            90 => x"56",
            91 => x"04",
            92 => x"70",
            93 => x"ff",
            94 => x"72",
            95 => x"51",
            96 => x"70",
            97 => x"06",
            98 => x"09",
            99 => x"51",
           100 => x"05",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"05",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"05",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"05",
           125 => x"04",
           126 => x"ff",
           127 => x"ff",
           128 => x"06",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"85",
           134 => x"0b",
           135 => x"0b",
           136 => x"c6",
           137 => x"0b",
           138 => x"0b",
           139 => x"86",
           140 => x"0b",
           141 => x"0b",
           142 => x"c6",
           143 => x"0b",
           144 => x"0b",
           145 => x"8a",
           146 => x"0b",
           147 => x"0b",
           148 => x"ce",
           149 => x"0b",
           150 => x"0b",
           151 => x"92",
           152 => x"0b",
           153 => x"0b",
           154 => x"d6",
           155 => x"0b",
           156 => x"0b",
           157 => x"9a",
           158 => x"0b",
           159 => x"0b",
           160 => x"de",
           161 => x"0b",
           162 => x"0b",
           163 => x"a2",
           164 => x"0b",
           165 => x"0b",
           166 => x"e6",
           167 => x"0b",
           168 => x"0b",
           169 => x"aa",
           170 => x"0b",
           171 => x"0b",
           172 => x"ed",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"8c",
           193 => x"d6",
           194 => x"c0",
           195 => x"a2",
           196 => x"c0",
           197 => x"a0",
           198 => x"c0",
           199 => x"a0",
           200 => x"c0",
           201 => x"94",
           202 => x"c0",
           203 => x"a1",
           204 => x"c0",
           205 => x"af",
           206 => x"c0",
           207 => x"ad",
           208 => x"c0",
           209 => x"94",
           210 => x"c0",
           211 => x"95",
           212 => x"c0",
           213 => x"95",
           214 => x"c0",
           215 => x"b1",
           216 => x"c0",
           217 => x"80",
           218 => x"80",
           219 => x"0c",
           220 => x"08",
           221 => x"90",
           222 => x"90",
           223 => x"bb",
           224 => x"bb",
           225 => x"84",
           226 => x"84",
           227 => x"04",
           228 => x"2d",
           229 => x"90",
           230 => x"c5",
           231 => x"80",
           232 => x"d9",
           233 => x"c0",
           234 => x"82",
           235 => x"80",
           236 => x"0c",
           237 => x"08",
           238 => x"90",
           239 => x"90",
           240 => x"bb",
           241 => x"bb",
           242 => x"84",
           243 => x"84",
           244 => x"04",
           245 => x"2d",
           246 => x"90",
           247 => x"b1",
           248 => x"80",
           249 => x"ff",
           250 => x"c0",
           251 => x"83",
           252 => x"80",
           253 => x"0c",
           254 => x"08",
           255 => x"90",
           256 => x"90",
           257 => x"bb",
           258 => x"bb",
           259 => x"84",
           260 => x"84",
           261 => x"04",
           262 => x"2d",
           263 => x"90",
           264 => x"97",
           265 => x"80",
           266 => x"f6",
           267 => x"c0",
           268 => x"83",
           269 => x"80",
           270 => x"0c",
           271 => x"08",
           272 => x"90",
           273 => x"90",
           274 => x"bb",
           275 => x"bb",
           276 => x"84",
           277 => x"84",
           278 => x"04",
           279 => x"2d",
           280 => x"90",
           281 => x"d4",
           282 => x"80",
           283 => x"f5",
           284 => x"c0",
           285 => x"81",
           286 => x"80",
           287 => x"0c",
           288 => x"08",
           289 => x"90",
           290 => x"90",
           291 => x"bb",
           292 => x"bb",
           293 => x"84",
           294 => x"84",
           295 => x"04",
           296 => x"84",
           297 => x"04",
           298 => x"2d",
           299 => x"90",
           300 => x"84",
           301 => x"80",
           302 => x"f3",
           303 => x"c0",
           304 => x"81",
           305 => x"80",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"04",
           311 => x"83",
           312 => x"10",
           313 => x"51",
           314 => x"06",
           315 => x"10",
           316 => x"ed",
           317 => x"bb",
           318 => x"38",
           319 => x"0b",
           320 => x"51",
           321 => x"0d",
           322 => x"08",
           323 => x"08",
           324 => x"04",
           325 => x"11",
           326 => x"25",
           327 => x"72",
           328 => x"38",
           329 => x"30",
           330 => x"55",
           331 => x"71",
           332 => x"fa",
           333 => x"bb",
           334 => x"bb",
           335 => x"34",
           336 => x"70",
           337 => x"54",
           338 => x"34",
           339 => x"88",
           340 => x"84",
           341 => x"0d",
           342 => x"05",
           343 => x"3d",
           344 => x"e4",
           345 => x"80",
           346 => x"3d",
           347 => x"52",
           348 => x"04",
           349 => x"5d",
           350 => x"1e",
           351 => x"06",
           352 => x"2e",
           353 => x"33",
           354 => x"81",
           355 => x"80",
           356 => x"7e",
           357 => x"32",
           358 => x"55",
           359 => x"38",
           360 => x"06",
           361 => x"7a",
           362 => x"76",
           363 => x"73",
           364 => x"04",
           365 => x"10",
           366 => x"98",
           367 => x"8b",
           368 => x"5b",
           369 => x"38",
           370 => x"38",
           371 => x"f7",
           372 => x"09",
           373 => x"5a",
           374 => x"76",
           375 => x"52",
           376 => x"57",
           377 => x"7a",
           378 => x"78",
           379 => x"54",
           380 => x"80",
           381 => x"83",
           382 => x"73",
           383 => x"27",
           384 => x"eb",
           385 => x"fe",
           386 => x"59",
           387 => x"84",
           388 => x"06",
           389 => x"5e",
           390 => x"84",
           391 => x"bb",
           392 => x"72",
           393 => x"08",
           394 => x"05",
           395 => x"ca",
           396 => x"bb",
           397 => x"94",
           398 => x"56",
           399 => x"80",
           400 => x"90",
           401 => x"81",
           402 => x"38",
           403 => x"80",
           404 => x"77",
           405 => x"05",
           406 => x"2a",
           407 => x"2e",
           408 => x"ff",
           409 => x"cc",
           410 => x"83",
           411 => x"74",
           412 => x"f0",
           413 => x"90",
           414 => x"53",
           415 => x"81",
           416 => x"38",
           417 => x"86",
           418 => x"54",
           419 => x"54",
           420 => x"81",
           421 => x"77",
           422 => x"80",
           423 => x"80",
           424 => x"51",
           425 => x"80",
           426 => x"2c",
           427 => x"38",
           428 => x"b2",
           429 => x"81",
           430 => x"55",
           431 => x"52",
           432 => x"81",
           433 => x"70",
           434 => x"24",
           435 => x"06",
           436 => x"38",
           437 => x"76",
           438 => x"80",
           439 => x"bb",
           440 => x"1e",
           441 => x"7d",
           442 => x"ec",
           443 => x"2e",
           444 => x"80",
           445 => x"2c",
           446 => x"91",
           447 => x"3f",
           448 => x"a0",
           449 => x"87",
           450 => x"07",
           451 => x"84",
           452 => x"06",
           453 => x"39",
           454 => x"0a",
           455 => x"72",
           456 => x"80",
           457 => x"5a",
           458 => x"70",
           459 => x"38",
           460 => x"80",
           461 => x"5f",
           462 => x"52",
           463 => x"ff",
           464 => x"57",
           465 => x"38",
           466 => x"33",
           467 => x"1a",
           468 => x"79",
           469 => x"7c",
           470 => x"51",
           471 => x"0a",
           472 => x"80",
           473 => x"90",
           474 => x"87",
           475 => x"7a",
           476 => x"60",
           477 => x"41",
           478 => x"7a",
           479 => x"94",
           480 => x"7c",
           481 => x"f8",
           482 => x"7c",
           483 => x"f8",
           484 => x"08",
           485 => x"72",
           486 => x"3f",
           487 => x"06",
           488 => x"72",
           489 => x"80",
           490 => x"f7",
           491 => x"84",
           492 => x"58",
           493 => x"51",
           494 => x"83",
           495 => x"2b",
           496 => x"07",
           497 => x"38",
           498 => x"80",
           499 => x"2c",
           500 => x"d6",
           501 => x"3f",
           502 => x"bb",
           503 => x"fa",
           504 => x"ab",
           505 => x"7e",
           506 => x"39",
           507 => x"2b",
           508 => x"57",
           509 => x"ff",
           510 => x"fb",
           511 => x"2e",
           512 => x"52",
           513 => x"74",
           514 => x"f1",
           515 => x"98",
           516 => x"b7",
           517 => x"3f",
           518 => x"bb",
           519 => x"51",
           520 => x"83",
           521 => x"2b",
           522 => x"07",
           523 => x"52",
           524 => x"0d",
           525 => x"74",
           526 => x"04",
           527 => x"84",
           528 => x"81",
           529 => x"56",
           530 => x"2e",
           531 => x"70",
           532 => x"2e",
           533 => x"72",
           534 => x"84",
           535 => x"ff",
           536 => x"53",
           537 => x"e8",
           538 => x"08",
           539 => x"51",
           540 => x"bb",
           541 => x"57",
           542 => x"88",
           543 => x"7a",
           544 => x"70",
           545 => x"51",
           546 => x"2e",
           547 => x"81",
           548 => x"09",
           549 => x"84",
           550 => x"73",
           551 => x"80",
           552 => x"90",
           553 => x"84",
           554 => x"70",
           555 => x"e3",
           556 => x"e6",
           557 => x"83",
           558 => x"7a",
           559 => x"32",
           560 => x"56",
           561 => x"06",
           562 => x"15",
           563 => x"91",
           564 => x"74",
           565 => x"08",
           566 => x"56",
           567 => x"0d",
           568 => x"51",
           569 => x"56",
           570 => x"15",
           571 => x"56",
           572 => x"11",
           573 => x"32",
           574 => x"54",
           575 => x"06",
           576 => x"81",
           577 => x"38",
           578 => x"80",
           579 => x"0c",
           580 => x"0c",
           581 => x"bb",
           582 => x"ff",
           583 => x"8c",
           584 => x"84",
           585 => x"3d",
           586 => x"55",
           587 => x"84",
           588 => x"38",
           589 => x"52",
           590 => x"38",
           591 => x"34",
           592 => x"87",
           593 => x"72",
           594 => x"fd",
           595 => x"54",
           596 => x"70",
           597 => x"81",
           598 => x"81",
           599 => x"84",
           600 => x"fc",
           601 => x"55",
           602 => x"73",
           603 => x"93",
           604 => x"73",
           605 => x"51",
           606 => x"0c",
           607 => x"73",
           608 => x"53",
           609 => x"71",
           610 => x"80",
           611 => x"53",
           612 => x"51",
           613 => x"0d",
           614 => x"05",
           615 => x"12",
           616 => x"51",
           617 => x"75",
           618 => x"81",
           619 => x"81",
           620 => x"84",
           621 => x"fd",
           622 => x"55",
           623 => x"71",
           624 => x"81",
           625 => x"ef",
           626 => x"3d",
           627 => x"7a",
           628 => x"38",
           629 => x"33",
           630 => x"06",
           631 => x"2e",
           632 => x"38",
           633 => x"86",
           634 => x"38",
           635 => x"2e",
           636 => x"51",
           637 => x"31",
           638 => x"04",
           639 => x"0d",
           640 => x"70",
           641 => x"84",
           642 => x"52",
           643 => x"84",
           644 => x"2e",
           645 => x"54",
           646 => x"84",
           647 => x"84",
           648 => x"84",
           649 => x"0d",
           650 => x"54",
           651 => x"81",
           652 => x"8c",
           653 => x"09",
           654 => x"75",
           655 => x"0c",
           656 => x"75",
           657 => x"70",
           658 => x"81",
           659 => x"f4",
           660 => x"3d",
           661 => x"58",
           662 => x"38",
           663 => x"84",
           664 => x"2e",
           665 => x"71",
           666 => x"52",
           667 => x"52",
           668 => x"13",
           669 => x"71",
           670 => x"74",
           671 => x"9f",
           672 => x"72",
           673 => x"06",
           674 => x"1c",
           675 => x"53",
           676 => x"52",
           677 => x"0d",
           678 => x"80",
           679 => x"80",
           680 => x"75",
           681 => x"70",
           682 => x"71",
           683 => x"06",
           684 => x"84",
           685 => x"75",
           686 => x"70",
           687 => x"71",
           688 => x"81",
           689 => x"75",
           690 => x"52",
           691 => x"55",
           692 => x"51",
           693 => x"04",
           694 => x"71",
           695 => x"bb",
           696 => x"84",
           697 => x"04",
           698 => x"a0",
           699 => x"51",
           700 => x"53",
           701 => x"38",
           702 => x"bb",
           703 => x"9f",
           704 => x"9f",
           705 => x"2a",
           706 => x"54",
           707 => x"a8",
           708 => x"74",
           709 => x"11",
           710 => x"06",
           711 => x"52",
           712 => x"38",
           713 => x"0d",
           714 => x"7a",
           715 => x"7c",
           716 => x"71",
           717 => x"59",
           718 => x"84",
           719 => x"84",
           720 => x"f7",
           721 => x"70",
           722 => x"56",
           723 => x"8f",
           724 => x"33",
           725 => x"73",
           726 => x"2e",
           727 => x"56",
           728 => x"58",
           729 => x"38",
           730 => x"14",
           731 => x"14",
           732 => x"73",
           733 => x"ff",
           734 => x"89",
           735 => x"77",
           736 => x"0c",
           737 => x"26",
           738 => x"38",
           739 => x"56",
           740 => x"0d",
           741 => x"70",
           742 => x"09",
           743 => x"70",
           744 => x"80",
           745 => x"80",
           746 => x"74",
           747 => x"56",
           748 => x"38",
           749 => x"0d",
           750 => x"0c",
           751 => x"ca",
           752 => x"8b",
           753 => x"7d",
           754 => x"08",
           755 => x"2e",
           756 => x"70",
           757 => x"a0",
           758 => x"f5",
           759 => x"d0",
           760 => x"80",
           761 => x"74",
           762 => x"27",
           763 => x"06",
           764 => x"06",
           765 => x"f9",
           766 => x"89",
           767 => x"27",
           768 => x"81",
           769 => x"56",
           770 => x"78",
           771 => x"75",
           772 => x"84",
           773 => x"16",
           774 => x"59",
           775 => x"ff",
           776 => x"33",
           777 => x"38",
           778 => x"38",
           779 => x"d0",
           780 => x"73",
           781 => x"84",
           782 => x"81",
           783 => x"55",
           784 => x"84",
           785 => x"80",
           786 => x"81",
           787 => x"ff",
           788 => x"8c",
           789 => x"05",
           790 => x"51",
           791 => x"83",
           792 => x"3d",
           793 => x"a8",
           794 => x"ec",
           795 => x"04",
           796 => x"83",
           797 => x"ef",
           798 => x"d0",
           799 => x"0d",
           800 => x"3f",
           801 => x"51",
           802 => x"83",
           803 => x"3d",
           804 => x"d0",
           805 => x"b4",
           806 => x"04",
           807 => x"83",
           808 => x"ee",
           809 => x"d1",
           810 => x"0d",
           811 => x"3f",
           812 => x"51",
           813 => x"83",
           814 => x"3d",
           815 => x"f8",
           816 => x"c8",
           817 => x"04",
           818 => x"83",
           819 => x"81",
           820 => x"e3",
           821 => x"99",
           822 => x"73",
           823 => x"75",
           824 => x"74",
           825 => x"55",
           826 => x"53",
           827 => x"82",
           828 => x"57",
           829 => x"d1",
           830 => x"76",
           831 => x"30",
           832 => x"57",
           833 => x"c0",
           834 => x"26",
           835 => x"e8",
           836 => x"84",
           837 => x"52",
           838 => x"76",
           839 => x"0d",
           840 => x"98",
           841 => x"81",
           842 => x"80",
           843 => x"ea",
           844 => x"bb",
           845 => x"74",
           846 => x"75",
           847 => x"52",
           848 => x"84",
           849 => x"84",
           850 => x"53",
           851 => x"ed",
           852 => x"7c",
           853 => x"59",
           854 => x"51",
           855 => x"8b",
           856 => x"81",
           857 => x"0c",
           858 => x"e6",
           859 => x"bb",
           860 => x"2d",
           861 => x"0c",
           862 => x"7f",
           863 => x"05",
           864 => x"5c",
           865 => x"83",
           866 => x"51",
           867 => x"dd",
           868 => x"b2",
           869 => x"7c",
           870 => x"53",
           871 => x"33",
           872 => x"3f",
           873 => x"54",
           874 => x"26",
           875 => x"ad",
           876 => x"c0",
           877 => x"80",
           878 => x"55",
           879 => x"81",
           880 => x"06",
           881 => x"80",
           882 => x"e6",
           883 => x"3f",
           884 => x"38",
           885 => x"78",
           886 => x"9d",
           887 => x"2b",
           888 => x"2e",
           889 => x"c3",
           890 => x"fe",
           891 => x"0c",
           892 => x"51",
           893 => x"e8",
           894 => x"3f",
           895 => x"da",
           896 => x"3f",
           897 => x"54",
           898 => x"27",
           899 => x"7a",
           900 => x"d3",
           901 => x"84",
           902 => x"ea",
           903 => x"fe",
           904 => x"c5",
           905 => x"53",
           906 => x"79",
           907 => x"72",
           908 => x"83",
           909 => x"14",
           910 => x"51",
           911 => x"38",
           912 => x"52",
           913 => x"56",
           914 => x"84",
           915 => x"88",
           916 => x"a0",
           917 => x"06",
           918 => x"39",
           919 => x"84",
           920 => x"a0",
           921 => x"30",
           922 => x"51",
           923 => x"80",
           924 => x"99",
           925 => x"70",
           926 => x"72",
           927 => x"73",
           928 => x"57",
           929 => x"38",
           930 => x"84",
           931 => x"0d",
           932 => x"dd",
           933 => x"d4",
           934 => x"9d",
           935 => x"06",
           936 => x"82",
           937 => x"82",
           938 => x"06",
           939 => x"84",
           940 => x"81",
           941 => x"06",
           942 => x"86",
           943 => x"80",
           944 => x"06",
           945 => x"2a",
           946 => x"f5",
           947 => x"9c",
           948 => x"aa",
           949 => x"dd",
           950 => x"9c",
           951 => x"92",
           952 => x"88",
           953 => x"c6",
           954 => x"3f",
           955 => x"80",
           956 => x"70",
           957 => x"ff",
           958 => x"c2",
           959 => x"3f",
           960 => x"2a",
           961 => x"2e",
           962 => x"51",
           963 => x"9b",
           964 => x"72",
           965 => x"71",
           966 => x"39",
           967 => x"cc",
           968 => x"f2",
           969 => x"51",
           970 => x"ff",
           971 => x"83",
           972 => x"51",
           973 => x"81",
           974 => x"e6",
           975 => x"ba",
           976 => x"3f",
           977 => x"2a",
           978 => x"2e",
           979 => x"3d",
           980 => x"84",
           981 => x"51",
           982 => x"08",
           983 => x"78",
           984 => x"c4",
           985 => x"83",
           986 => x"48",
           987 => x"eb",
           988 => x"33",
           989 => x"80",
           990 => x"83",
           991 => x"7d",
           992 => x"5a",
           993 => x"79",
           994 => x"06",
           995 => x"5a",
           996 => x"7b",
           997 => x"83",
           998 => x"e7",
           999 => x"bb",
          1000 => x"52",
          1001 => x"08",
          1002 => x"81",
          1003 => x"81",
          1004 => x"c4",
          1005 => x"2e",
          1006 => x"51",
          1007 => x"5e",
          1008 => x"ce",
          1009 => x"3d",
          1010 => x"84",
          1011 => x"5c",
          1012 => x"bb",
          1013 => x"bb",
          1014 => x"81",
          1015 => x"2e",
          1016 => x"e7",
          1017 => x"7b",
          1018 => x"7c",
          1019 => x"58",
          1020 => x"55",
          1021 => x"80",
          1022 => x"84",
          1023 => x"09",
          1024 => x"51",
          1025 => x"26",
          1026 => x"59",
          1027 => x"70",
          1028 => x"95",
          1029 => x"07",
          1030 => x"2e",
          1031 => x"9e",
          1032 => x"3f",
          1033 => x"7e",
          1034 => x"ef",
          1035 => x"59",
          1036 => x"d6",
          1037 => x"8a",
          1038 => x"c5",
          1039 => x"f8",
          1040 => x"52",
          1041 => x"bb",
          1042 => x"bb",
          1043 => x"0b",
          1044 => x"06",
          1045 => x"06",
          1046 => x"94",
          1047 => x"0b",
          1048 => x"83",
          1049 => x"52",
          1050 => x"5a",
          1051 => x"7c",
          1052 => x"78",
          1053 => x"10",
          1054 => x"08",
          1055 => x"7e",
          1056 => x"52",
          1057 => x"3f",
          1058 => x"81",
          1059 => x"3d",
          1060 => x"d7",
          1061 => x"81",
          1062 => x"d7",
          1063 => x"54",
          1064 => x"51",
          1065 => x"8d",
          1066 => x"3f",
          1067 => x"80",
          1068 => x"8f",
          1069 => x"b4",
          1070 => x"04",
          1071 => x"d0",
          1072 => x"ff",
          1073 => x"eb",
          1074 => x"2e",
          1075 => x"e4",
          1076 => x"2d",
          1077 => x"9f",
          1078 => x"d8",
          1079 => x"39",
          1080 => x"80",
          1081 => x"84",
          1082 => x"52",
          1083 => x"68",
          1084 => x"11",
          1085 => x"3f",
          1086 => x"d7",
          1087 => x"ff",
          1088 => x"bb",
          1089 => x"78",
          1090 => x"51",
          1091 => x"53",
          1092 => x"3f",
          1093 => x"2e",
          1094 => x"d3",
          1095 => x"cf",
          1096 => x"ff",
          1097 => x"bb",
          1098 => x"b8",
          1099 => x"05",
          1100 => x"08",
          1101 => x"53",
          1102 => x"95",
          1103 => x"f8",
          1104 => x"48",
          1105 => x"bf",
          1106 => x"64",
          1107 => x"b8",
          1108 => x"05",
          1109 => x"08",
          1110 => x"fe",
          1111 => x"e9",
          1112 => x"2e",
          1113 => x"11",
          1114 => x"3f",
          1115 => x"ef",
          1116 => x"3f",
          1117 => x"83",
          1118 => x"5f",
          1119 => x"7a",
          1120 => x"52",
          1121 => x"66",
          1122 => x"47",
          1123 => x"11",
          1124 => x"3f",
          1125 => x"9f",
          1126 => x"ff",
          1127 => x"bb",
          1128 => x"b8",
          1129 => x"05",
          1130 => x"08",
          1131 => x"80",
          1132 => x"67",
          1133 => x"70",
          1134 => x"81",
          1135 => x"84",
          1136 => x"83",
          1137 => x"f6",
          1138 => x"53",
          1139 => x"84",
          1140 => x"33",
          1141 => x"dd",
          1142 => x"f8",
          1143 => x"48",
          1144 => x"87",
          1145 => x"68",
          1146 => x"02",
          1147 => x"81",
          1148 => x"53",
          1149 => x"84",
          1150 => x"38",
          1151 => x"79",
          1152 => x"fe",
          1153 => x"e6",
          1154 => x"bd",
          1155 => x"84",
          1156 => x"e3",
          1157 => x"f5",
          1158 => x"53",
          1159 => x"84",
          1160 => x"38",
          1161 => x"80",
          1162 => x"84",
          1163 => x"46",
          1164 => x"68",
          1165 => x"38",
          1166 => x"5b",
          1167 => x"51",
          1168 => x"3d",
          1169 => x"84",
          1170 => x"05",
          1171 => x"84",
          1172 => x"f3",
          1173 => x"f4",
          1174 => x"e7",
          1175 => x"ff",
          1176 => x"e5",
          1177 => x"38",
          1178 => x"2e",
          1179 => x"49",
          1180 => x"80",
          1181 => x"84",
          1182 => x"5a",
          1183 => x"f3",
          1184 => x"11",
          1185 => x"3f",
          1186 => x"38",
          1187 => x"83",
          1188 => x"30",
          1189 => x"5c",
          1190 => x"7a",
          1191 => x"d9",
          1192 => x"68",
          1193 => x"eb",
          1194 => x"a0",
          1195 => x"0c",
          1196 => x"fe",
          1197 => x"e2",
          1198 => x"2e",
          1199 => x"59",
          1200 => x"f0",
          1201 => x"f7",
          1202 => x"f2",
          1203 => x"05",
          1204 => x"7d",
          1205 => x"ff",
          1206 => x"bb",
          1207 => x"64",
          1208 => x"70",
          1209 => x"3d",
          1210 => x"51",
          1211 => x"ff",
          1212 => x"fe",
          1213 => x"e3",
          1214 => x"2e",
          1215 => x"db",
          1216 => x"49",
          1217 => x"11",
          1218 => x"3f",
          1219 => x"98",
          1220 => x"84",
          1221 => x"7a",
          1222 => x"38",
          1223 => x"53",
          1224 => x"e5",
          1225 => x"51",
          1226 => x"d9",
          1227 => x"39",
          1228 => x"80",
          1229 => x"84",
          1230 => x"02",
          1231 => x"05",
          1232 => x"83",
          1233 => x"80",
          1234 => x"fc",
          1235 => x"7b",
          1236 => x"08",
          1237 => x"51",
          1238 => x"39",
          1239 => x"64",
          1240 => x"33",
          1241 => x"f3",
          1242 => x"d9",
          1243 => x"39",
          1244 => x"2e",
          1245 => x"fc",
          1246 => x"7d",
          1247 => x"08",
          1248 => x"33",
          1249 => x"f3",
          1250 => x"f4",
          1251 => x"38",
          1252 => x"39",
          1253 => x"2e",
          1254 => x"fb",
          1255 => x"80",
          1256 => x"f0",
          1257 => x"f3",
          1258 => x"34",
          1259 => x"57",
          1260 => x"c2",
          1261 => x"77",
          1262 => x"75",
          1263 => x"84",
          1264 => x"9c",
          1265 => x"52",
          1266 => x"84",
          1267 => x"87",
          1268 => x"3f",
          1269 => x"0c",
          1270 => x"84",
          1271 => x"94",
          1272 => x"c9",
          1273 => x"05",
          1274 => x"89",
          1275 => x"0c",
          1276 => x"3f",
          1277 => x"98",
          1278 => x"52",
          1279 => x"83",
          1280 => x"98",
          1281 => x"d8",
          1282 => x"e0",
          1283 => x"83",
          1284 => x"52",
          1285 => x"90",
          1286 => x"c3",
          1287 => x"fb",
          1288 => x"80",
          1289 => x"83",
          1290 => x"52",
          1291 => x"91",
          1292 => x"ff",
          1293 => x"f1",
          1294 => x"a2",
          1295 => x"81",
          1296 => x"70",
          1297 => x"a0",
          1298 => x"2e",
          1299 => x"81",
          1300 => x"ff",
          1301 => x"81",
          1302 => x"32",
          1303 => x"52",
          1304 => x"80",
          1305 => x"76",
          1306 => x"0c",
          1307 => x"c4",
          1308 => x"81",
          1309 => x"ff",
          1310 => x"e4",
          1311 => x"55",
          1312 => x"09",
          1313 => x"fc",
          1314 => x"38",
          1315 => x"3d",
          1316 => x"72",
          1317 => x"08",
          1318 => x"84",
          1319 => x"0d",
          1320 => x"53",
          1321 => x"38",
          1322 => x"52",
          1323 => x"13",
          1324 => x"80",
          1325 => x"52",
          1326 => x"13",
          1327 => x"80",
          1328 => x"52",
          1329 => x"8a",
          1330 => x"e7",
          1331 => x"c0",
          1332 => x"98",
          1333 => x"98",
          1334 => x"98",
          1335 => x"98",
          1336 => x"98",
          1337 => x"98",
          1338 => x"0c",
          1339 => x"0b",
          1340 => x"71",
          1341 => x"04",
          1342 => x"98",
          1343 => x"98",
          1344 => x"c0",
          1345 => x"34",
          1346 => x"83",
          1347 => x"5c",
          1348 => x"ac",
          1349 => x"c0",
          1350 => x"34",
          1351 => x"88",
          1352 => x"5a",
          1353 => x"79",
          1354 => x"ff",
          1355 => x"85",
          1356 => x"83",
          1357 => x"7d",
          1358 => x"fc",
          1359 => x"0d",
          1360 => x"33",
          1361 => x"51",
          1362 => x"08",
          1363 => x"71",
          1364 => x"72",
          1365 => x"84",
          1366 => x"80",
          1367 => x"98",
          1368 => x"ff",
          1369 => x"51",
          1370 => x"08",
          1371 => x"71",
          1372 => x"3d",
          1373 => x"2b",
          1374 => x"84",
          1375 => x"2c",
          1376 => x"73",
          1377 => x"73",
          1378 => x"0c",
          1379 => x"02",
          1380 => x"70",
          1381 => x"80",
          1382 => x"94",
          1383 => x"53",
          1384 => x"71",
          1385 => x"70",
          1386 => x"53",
          1387 => x"2a",
          1388 => x"81",
          1389 => x"52",
          1390 => x"94",
          1391 => x"bb",
          1392 => x"91",
          1393 => x"97",
          1394 => x"72",
          1395 => x"81",
          1396 => x"87",
          1397 => x"70",
          1398 => x"38",
          1399 => x"05",
          1400 => x"52",
          1401 => x"3d",
          1402 => x"80",
          1403 => x"77",
          1404 => x"f3",
          1405 => x"57",
          1406 => x"87",
          1407 => x"70",
          1408 => x"2e",
          1409 => x"06",
          1410 => x"32",
          1411 => x"38",
          1412 => x"cf",
          1413 => x"c0",
          1414 => x"38",
          1415 => x"0c",
          1416 => x"ff",
          1417 => x"88",
          1418 => x"81",
          1419 => x"81",
          1420 => x"c1",
          1421 => x"71",
          1422 => x"94",
          1423 => x"06",
          1424 => x"39",
          1425 => x"08",
          1426 => x"70",
          1427 => x"9e",
          1428 => x"c0",
          1429 => x"87",
          1430 => x"0c",
          1431 => x"cc",
          1432 => x"f3",
          1433 => x"83",
          1434 => x"08",
          1435 => x"b0",
          1436 => x"9e",
          1437 => x"c0",
          1438 => x"87",
          1439 => x"0c",
          1440 => x"ec",
          1441 => x"f3",
          1442 => x"52",
          1443 => x"9e",
          1444 => x"c0",
          1445 => x"87",
          1446 => x"0c",
          1447 => x"0b",
          1448 => x"80",
          1449 => x"fb",
          1450 => x"0b",
          1451 => x"80",
          1452 => x"2e",
          1453 => x"86",
          1454 => x"08",
          1455 => x"52",
          1456 => x"71",
          1457 => x"c0",
          1458 => x"06",
          1459 => x"38",
          1460 => x"80",
          1461 => x"a0",
          1462 => x"80",
          1463 => x"f4",
          1464 => x"90",
          1465 => x"52",
          1466 => x"52",
          1467 => x"87",
          1468 => x"80",
          1469 => x"83",
          1470 => x"34",
          1471 => x"70",
          1472 => x"70",
          1473 => x"83",
          1474 => x"9e",
          1475 => x"51",
          1476 => x"81",
          1477 => x"0b",
          1478 => x"c0",
          1479 => x"2e",
          1480 => x"8e",
          1481 => x"08",
          1482 => x"70",
          1483 => x"83",
          1484 => x"08",
          1485 => x"51",
          1486 => x"87",
          1487 => x"06",
          1488 => x"38",
          1489 => x"87",
          1490 => x"70",
          1491 => x"92",
          1492 => x"08",
          1493 => x"80",
          1494 => x"f4",
          1495 => x"87",
          1496 => x"83",
          1497 => x"39",
          1498 => x"ff",
          1499 => x"54",
          1500 => x"51",
          1501 => x"55",
          1502 => x"33",
          1503 => x"88",
          1504 => x"f4",
          1505 => x"83",
          1506 => x"38",
          1507 => x"a9",
          1508 => x"84",
          1509 => x"74",
          1510 => x"56",
          1511 => x"33",
          1512 => x"8c",
          1513 => x"f4",
          1514 => x"83",
          1515 => x"38",
          1516 => x"83",
          1517 => x"51",
          1518 => x"08",
          1519 => x"8d",
          1520 => x"db",
          1521 => x"db",
          1522 => x"f4",
          1523 => x"b4",
          1524 => x"bd",
          1525 => x"3f",
          1526 => x"29",
          1527 => x"84",
          1528 => x"b4",
          1529 => x"74",
          1530 => x"74",
          1531 => x"f4",
          1532 => x"75",
          1533 => x"08",
          1534 => x"54",
          1535 => x"dc",
          1536 => x"3d",
          1537 => x"bd",
          1538 => x"3f",
          1539 => x"29",
          1540 => x"84",
          1541 => x"b3",
          1542 => x"74",
          1543 => x"39",
          1544 => x"83",
          1545 => x"f3",
          1546 => x"ff",
          1547 => x"52",
          1548 => x"3f",
          1549 => x"9c",
          1550 => x"c4",
          1551 => x"f4",
          1552 => x"b3",
          1553 => x"bd",
          1554 => x"3f",
          1555 => x"29",
          1556 => x"84",
          1557 => x"b2",
          1558 => x"74",
          1559 => x"39",
          1560 => x"3f",
          1561 => x"2e",
          1562 => x"dd",
          1563 => x"f4",
          1564 => x"ef",
          1565 => x"ff",
          1566 => x"55",
          1567 => x"39",
          1568 => x"3f",
          1569 => x"2e",
          1570 => x"92",
          1571 => x"b1",
          1572 => x"75",
          1573 => x"83",
          1574 => x"51",
          1575 => x"33",
          1576 => x"cd",
          1577 => x"dd",
          1578 => x"f4",
          1579 => x"ca",
          1580 => x"83",
          1581 => x"de",
          1582 => x"f4",
          1583 => x"a1",
          1584 => x"83",
          1585 => x"de",
          1586 => x"f4",
          1587 => x"f8",
          1588 => x"83",
          1589 => x"de",
          1590 => x"f4",
          1591 => x"cf",
          1592 => x"83",
          1593 => x"de",
          1594 => x"f4",
          1595 => x"a6",
          1596 => x"83",
          1597 => x"df",
          1598 => x"f4",
          1599 => x"fd",
          1600 => x"ff",
          1601 => x"ff",
          1602 => x"55",
          1603 => x"39",
          1604 => x"52",
          1605 => x"10",
          1606 => x"04",
          1607 => x"3f",
          1608 => x"51",
          1609 => x"04",
          1610 => x"3f",
          1611 => x"51",
          1612 => x"04",
          1613 => x"3f",
          1614 => x"51",
          1615 => x"04",
          1616 => x"87",
          1617 => x"98",
          1618 => x"d9",
          1619 => x"08",
          1620 => x"52",
          1621 => x"fb",
          1622 => x"38",
          1623 => x"ec",
          1624 => x"51",
          1625 => x"08",
          1626 => x"d5",
          1627 => x"57",
          1628 => x"25",
          1629 => x"05",
          1630 => x"74",
          1631 => x"2a",
          1632 => x"38",
          1633 => x"08",
          1634 => x"93",
          1635 => x"78",
          1636 => x"84",
          1637 => x"b8",
          1638 => x"2e",
          1639 => x"79",
          1640 => x"bf",
          1641 => x"bb",
          1642 => x"e3",
          1643 => x"0b",
          1644 => x"04",
          1645 => x"3d",
          1646 => x"57",
          1647 => x"38",
          1648 => x"10",
          1649 => x"08",
          1650 => x"bb",
          1651 => x"51",
          1652 => x"08",
          1653 => x"81",
          1654 => x"99",
          1655 => x"57",
          1656 => x"54",
          1657 => x"0d",
          1658 => x"84",
          1659 => x"ab",
          1660 => x"d1",
          1661 => x"51",
          1662 => x"81",
          1663 => x"38",
          1664 => x"54",
          1665 => x"b6",
          1666 => x"76",
          1667 => x"5b",
          1668 => x"09",
          1669 => x"26",
          1670 => x"56",
          1671 => x"08",
          1672 => x"82",
          1673 => x"80",
          1674 => x"80",
          1675 => x"3f",
          1676 => x"38",
          1677 => x"bb",
          1678 => x"84",
          1679 => x"08",
          1680 => x"77",
          1681 => x"83",
          1682 => x"3f",
          1683 => x"b2",
          1684 => x"aa",
          1685 => x"3d",
          1686 => x"bc",
          1687 => x"58",
          1688 => x"83",
          1689 => x"f0",
          1690 => x"9e",
          1691 => x"57",
          1692 => x"80",
          1693 => x"06",
          1694 => x"80",
          1695 => x"3d",
          1696 => x"84",
          1697 => x"2c",
          1698 => x"38",
          1699 => x"33",
          1700 => x"e2",
          1701 => x"2c",
          1702 => x"83",
          1703 => x"33",
          1704 => x"58",
          1705 => x"80",
          1706 => x"38",
          1707 => x"0a",
          1708 => x"76",
          1709 => x"70",
          1710 => x"df",
          1711 => x"25",
          1712 => x"18",
          1713 => x"81",
          1714 => x"75",
          1715 => x"80",
          1716 => x"98",
          1717 => x"33",
          1718 => x"98",
          1719 => x"e4",
          1720 => x"5d",
          1721 => x"38",
          1722 => x"e9",
          1723 => x"2b",
          1724 => x"2e",
          1725 => x"80",
          1726 => x"8a",
          1727 => x"75",
          1728 => x"05",
          1729 => x"59",
          1730 => x"38",
          1731 => x"55",
          1732 => x"43",
          1733 => x"df",
          1734 => x"55",
          1735 => x"80",
          1736 => x"81",
          1737 => x"fe",
          1738 => x"80",
          1739 => x"e2",
          1740 => x"79",
          1741 => x"74",
          1742 => x"10",
          1743 => x"04",
          1744 => x"80",
          1745 => x"84",
          1746 => x"c8",
          1747 => x"38",
          1748 => x"ff",
          1749 => x"ff",
          1750 => x"fc",
          1751 => x"81",
          1752 => x"57",
          1753 => x"84",
          1754 => x"61",
          1755 => x"33",
          1756 => x"9a",
          1757 => x"7c",
          1758 => x"83",
          1759 => x"75",
          1760 => x"c4",
          1761 => x"33",
          1762 => x"80",
          1763 => x"52",
          1764 => x"e6",
          1765 => x"c3",
          1766 => x"51",
          1767 => x"33",
          1768 => x"34",
          1769 => x"38",
          1770 => x"84",
          1771 => x"8a",
          1772 => x"8c",
          1773 => x"06",
          1774 => x"7c",
          1775 => x"08",
          1776 => x"93",
          1777 => x"83",
          1778 => x"75",
          1779 => x"ff",
          1780 => x"84",
          1781 => x"81",
          1782 => x"7b",
          1783 => x"c4",
          1784 => x"74",
          1785 => x"e8",
          1786 => x"3f",
          1787 => x"ff",
          1788 => x"52",
          1789 => x"e2",
          1790 => x"e2",
          1791 => x"c7",
          1792 => x"ff",
          1793 => x"55",
          1794 => x"e6",
          1795 => x"84",
          1796 => x"52",
          1797 => x"c8",
          1798 => x"c4",
          1799 => x"f9",
          1800 => x"81",
          1801 => x"7b",
          1802 => x"9b",
          1803 => x"ff",
          1804 => x"55",
          1805 => x"92",
          1806 => x"c4",
          1807 => x"82",
          1808 => x"c4",
          1809 => x"7c",
          1810 => x"76",
          1811 => x"08",
          1812 => x"84",
          1813 => x"98",
          1814 => x"43",
          1815 => x"84",
          1816 => x"b1",
          1817 => x"81",
          1818 => x"e2",
          1819 => x"24",
          1820 => x"52",
          1821 => x"81",
          1822 => x"70",
          1823 => x"56",
          1824 => x"f7",
          1825 => x"33",
          1826 => x"77",
          1827 => x"81",
          1828 => x"70",
          1829 => x"57",
          1830 => x"7b",
          1831 => x"84",
          1832 => x"ff",
          1833 => x"29",
          1834 => x"84",
          1835 => x"76",
          1836 => x"84",
          1837 => x"f7",
          1838 => x"88",
          1839 => x"c8",
          1840 => x"c8",
          1841 => x"39",
          1842 => x"80",
          1843 => x"8a",
          1844 => x"c4",
          1845 => x"bb",
          1846 => x"8a",
          1847 => x"76",
          1848 => x"f4",
          1849 => x"05",
          1850 => x"c2",
          1851 => x"83",
          1852 => x"57",
          1853 => x"84",
          1854 => x"70",
          1855 => x"08",
          1856 => x"ff",
          1857 => x"70",
          1858 => x"08",
          1859 => x"83",
          1860 => x"8c",
          1861 => x"80",
          1862 => x"e2",
          1863 => x"34",
          1864 => x"0d",
          1865 => x"80",
          1866 => x"52",
          1867 => x"e6",
          1868 => x"8b",
          1869 => x"51",
          1870 => x"33",
          1871 => x"34",
          1872 => x"38",
          1873 => x"3f",
          1874 => x"0b",
          1875 => x"84",
          1876 => x"5c",
          1877 => x"84",
          1878 => x"84",
          1879 => x"84",
          1880 => x"52",
          1881 => x"e2",
          1882 => x"2c",
          1883 => x"56",
          1884 => x"e6",
          1885 => x"83",
          1886 => x"2b",
          1887 => x"5c",
          1888 => x"fa",
          1889 => x"51",
          1890 => x"0a",
          1891 => x"2c",
          1892 => x"74",
          1893 => x"e8",
          1894 => x"3f",
          1895 => x"0a",
          1896 => x"33",
          1897 => x"b9",
          1898 => x"81",
          1899 => x"08",
          1900 => x"3f",
          1901 => x"0a",
          1902 => x"33",
          1903 => x"e6",
          1904 => x"77",
          1905 => x"33",
          1906 => x"80",
          1907 => x"98",
          1908 => x"5b",
          1909 => x"b6",
          1910 => x"1d",
          1911 => x"80",
          1912 => x"52",
          1913 => x"e6",
          1914 => x"9b",
          1915 => x"51",
          1916 => x"33",
          1917 => x"34",
          1918 => x"38",
          1919 => x"3f",
          1920 => x"0b",
          1921 => x"84",
          1922 => x"c8",
          1923 => x"76",
          1924 => x"c4",
          1925 => x"74",
          1926 => x"76",
          1927 => x"7a",
          1928 => x"0a",
          1929 => x"2c",
          1930 => x"75",
          1931 => x"74",
          1932 => x"06",
          1933 => x"34",
          1934 => x"25",
          1935 => x"e2",
          1936 => x"33",
          1937 => x"0a",
          1938 => x"06",
          1939 => x"81",
          1940 => x"2c",
          1941 => x"75",
          1942 => x"e8",
          1943 => x"3f",
          1944 => x"0a",
          1945 => x"33",
          1946 => x"aa",
          1947 => x"51",
          1948 => x"0a",
          1949 => x"2c",
          1950 => x"74",
          1951 => x"39",
          1952 => x"84",
          1953 => x"84",
          1954 => x"51",
          1955 => x"08",
          1956 => x"f4",
          1957 => x"c3",
          1958 => x"16",
          1959 => x"3f",
          1960 => x"0a",
          1961 => x"33",
          1962 => x"38",
          1963 => x"70",
          1964 => x"58",
          1965 => x"38",
          1966 => x"80",
          1967 => x"57",
          1968 => x"38",
          1969 => x"80",
          1970 => x"f4",
          1971 => x"80",
          1972 => x"e7",
          1973 => x"80",
          1974 => x"ec",
          1975 => x"ee",
          1976 => x"3f",
          1977 => x"58",
          1978 => x"ff",
          1979 => x"3f",
          1980 => x"34",
          1981 => x"81",
          1982 => x"aa",
          1983 => x"33",
          1984 => x"74",
          1985 => x"e8",
          1986 => x"3f",
          1987 => x"ff",
          1988 => x"52",
          1989 => x"e2",
          1990 => x"e2",
          1991 => x"c7",
          1992 => x"84",
          1993 => x"84",
          1994 => x"05",
          1995 => x"8f",
          1996 => x"e2",
          1997 => x"2e",
          1998 => x"52",
          1999 => x"e6",
          2000 => x"eb",
          2001 => x"51",
          2002 => x"33",
          2003 => x"34",
          2004 => x"75",
          2005 => x"84",
          2006 => x"84",
          2007 => x"75",
          2008 => x"81",
          2009 => x"c4",
          2010 => x"5e",
          2011 => x"84",
          2012 => x"a5",
          2013 => x"a0",
          2014 => x"e8",
          2015 => x"3f",
          2016 => x"7a",
          2017 => x"06",
          2018 => x"0b",
          2019 => x"e2",
          2020 => x"b5",
          2021 => x"56",
          2022 => x"51",
          2023 => x"08",
          2024 => x"08",
          2025 => x"52",
          2026 => x"e2",
          2027 => x"56",
          2028 => x"e6",
          2029 => x"83",
          2030 => x"51",
          2031 => x"08",
          2032 => x"84",
          2033 => x"84",
          2034 => x"55",
          2035 => x"3f",
          2036 => x"87",
          2037 => x"19",
          2038 => x"96",
          2039 => x"83",
          2040 => x"f4",
          2041 => x"e3",
          2042 => x"83",
          2043 => x"f4",
          2044 => x"74",
          2045 => x"7b",
          2046 => x"83",
          2047 => x"ff",
          2048 => x"9f",
          2049 => x"8f",
          2050 => x"76",
          2051 => x"8a",
          2052 => x"51",
          2053 => x"08",
          2054 => x"84",
          2055 => x"c4",
          2056 => x"3d",
          2057 => x"51",
          2058 => x"08",
          2059 => x"97",
          2060 => x"53",
          2061 => x"e9",
          2062 => x"bb",
          2063 => x"e8",
          2064 => x"ff",
          2065 => x"57",
          2066 => x"80",
          2067 => x"05",
          2068 => x"76",
          2069 => x"70",
          2070 => x"08",
          2071 => x"38",
          2072 => x"f4",
          2073 => x"5f",
          2074 => x"08",
          2075 => x"10",
          2076 => x"54",
          2077 => x"92",
          2078 => x"10",
          2079 => x"57",
          2080 => x"70",
          2081 => x"27",
          2082 => x"09",
          2083 => x"dc",
          2084 => x"52",
          2085 => x"f4",
          2086 => x"06",
          2087 => x"38",
          2088 => x"bd",
          2089 => x"83",
          2090 => x"fc",
          2091 => x"70",
          2092 => x"3f",
          2093 => x"f4",
          2094 => x"9c",
          2095 => x"94",
          2096 => x"f4",
          2097 => x"9c",
          2098 => x"80",
          2099 => x"75",
          2100 => x"75",
          2101 => x"83",
          2102 => x"77",
          2103 => x"3d",
          2104 => x"84",
          2105 => x"72",
          2106 => x"2e",
          2107 => x"9e",
          2108 => x"86",
          2109 => x"80",
          2110 => x"58",
          2111 => x"fa",
          2112 => x"75",
          2113 => x"33",
          2114 => x"71",
          2115 => x"56",
          2116 => x"38",
          2117 => x"74",
          2118 => x"74",
          2119 => x"38",
          2120 => x"17",
          2121 => x"0b",
          2122 => x"81",
          2123 => x"ee",
          2124 => x"a0",
          2125 => x"10",
          2126 => x"90",
          2127 => x"40",
          2128 => x"b8",
          2129 => x"b8",
          2130 => x"fa",
          2131 => x"70",
          2132 => x"57",
          2133 => x"72",
          2134 => x"ff",
          2135 => x"ff",
          2136 => x"81",
          2137 => x"42",
          2138 => x"8f",
          2139 => x"31",
          2140 => x"76",
          2141 => x"9c",
          2142 => x"26",
          2143 => x"05",
          2144 => x"70",
          2145 => x"c7",
          2146 => x"70",
          2147 => x"06",
          2148 => x"06",
          2149 => x"5d",
          2150 => x"74",
          2151 => x"ff",
          2152 => x"29",
          2153 => x"fd",
          2154 => x"34",
          2155 => x"fa",
          2156 => x"2b",
          2157 => x"7a",
          2158 => x"26",
          2159 => x"fc",
          2160 => x"81",
          2161 => x"fa",
          2162 => x"c7",
          2163 => x"56",
          2164 => x"84",
          2165 => x"84",
          2166 => x"83",
          2167 => x"06",
          2168 => x"41",
          2169 => x"73",
          2170 => x"70",
          2171 => x"ff",
          2172 => x"29",
          2173 => x"ff",
          2174 => x"5c",
          2175 => x"77",
          2176 => x"79",
          2177 => x"38",
          2178 => x"38",
          2179 => x"29",
          2180 => x"87",
          2181 => x"34",
          2182 => x"73",
          2183 => x"f4",
          2184 => x"8e",
          2185 => x"76",
          2186 => x"74",
          2187 => x"34",
          2188 => x"86",
          2189 => x"81",
          2190 => x"77",
          2191 => x"34",
          2192 => x"c0",
          2193 => x"c0",
          2194 => x"07",
          2195 => x"34",
          2196 => x"53",
          2197 => x"b8",
          2198 => x"0c",
          2199 => x"33",
          2200 => x"0d",
          2201 => x"b3",
          2202 => x"59",
          2203 => x"da",
          2204 => x"b5",
          2205 => x"29",
          2206 => x"fa",
          2207 => x"7c",
          2208 => x"83",
          2209 => x"72",
          2210 => x"b2",
          2211 => x"b2",
          2212 => x"70",
          2213 => x"55",
          2214 => x"38",
          2215 => x"34",
          2216 => x"ff",
          2217 => x"57",
          2218 => x"b8",
          2219 => x"80",
          2220 => x"84",
          2221 => x"e0",
          2222 => x"70",
          2223 => x"05",
          2224 => x"f5",
          2225 => x"26",
          2226 => x"99",
          2227 => x"e0",
          2228 => x"55",
          2229 => x"27",
          2230 => x"05",
          2231 => x"57",
          2232 => x"ff",
          2233 => x"fd",
          2234 => x"b8",
          2235 => x"57",
          2236 => x"86",
          2237 => x"75",
          2238 => x"5c",
          2239 => x"38",
          2240 => x"14",
          2241 => x"78",
          2242 => x"81",
          2243 => x"59",
          2244 => x"84",
          2245 => x"56",
          2246 => x"38",
          2247 => x"8b",
          2248 => x"34",
          2249 => x"ff",
          2250 => x"57",
          2251 => x"80",
          2252 => x"06",
          2253 => x"53",
          2254 => x"c8",
          2255 => x"b8",
          2256 => x"29",
          2257 => x"27",
          2258 => x"84",
          2259 => x"56",
          2260 => x"75",
          2261 => x"13",
          2262 => x"a0",
          2263 => x"70",
          2264 => x"72",
          2265 => x"84",
          2266 => x"39",
          2267 => x"b9",
          2268 => x"f7",
          2269 => x"0d",
          2270 => x"53",
          2271 => x"10",
          2272 => x"08",
          2273 => x"71",
          2274 => x"34",
          2275 => x"3d",
          2276 => x"34",
          2277 => x"06",
          2278 => x"ff",
          2279 => x"80",
          2280 => x"0d",
          2281 => x"31",
          2282 => x"54",
          2283 => x"34",
          2284 => x"05",
          2285 => x"56",
          2286 => x"53",
          2287 => x"84",
          2288 => x"83",
          2289 => x"09",
          2290 => x"53",
          2291 => x"0b",
          2292 => x"04",
          2293 => x"b8",
          2294 => x"70",
          2295 => x"83",
          2296 => x"84",
          2297 => x"83",
          2298 => x"84",
          2299 => x"71",
          2300 => x"51",
          2301 => x"39",
          2302 => x"51",
          2303 => x"10",
          2304 => x"04",
          2305 => x"06",
          2306 => x"72",
          2307 => x"71",
          2308 => x"38",
          2309 => x"80",
          2310 => x"0d",
          2311 => x"06",
          2312 => x"34",
          2313 => x"3d",
          2314 => x"f0",
          2315 => x"e8",
          2316 => x"06",
          2317 => x"34",
          2318 => x"b0",
          2319 => x"83",
          2320 => x"81",
          2321 => x"fa",
          2322 => x"b0",
          2323 => x"b0",
          2324 => x"33",
          2325 => x"83",
          2326 => x"fa",
          2327 => x"51",
          2328 => x"39",
          2329 => x"81",
          2330 => x"fe",
          2331 => x"f8",
          2332 => x"fe",
          2333 => x"df",
          2334 => x"fa",
          2335 => x"b0",
          2336 => x"70",
          2337 => x"83",
          2338 => x"e0",
          2339 => x"fe",
          2340 => x"cf",
          2341 => x"fa",
          2342 => x"b0",
          2343 => x"70",
          2344 => x"83",
          2345 => x"70",
          2346 => x"83",
          2347 => x"07",
          2348 => x"e0",
          2349 => x"33",
          2350 => x"83",
          2351 => x"83",
          2352 => x"43",
          2353 => x"2e",
          2354 => x"38",
          2355 => x"84",
          2356 => x"fc",
          2357 => x"83",
          2358 => x"34",
          2359 => x"09",
          2360 => x"b8",
          2361 => x"34",
          2362 => x"0b",
          2363 => x"fa",
          2364 => x"33",
          2365 => x"b8",
          2366 => x"7a",
          2367 => x"8d",
          2368 => x"0b",
          2369 => x"b4",
          2370 => x"83",
          2371 => x"80",
          2372 => x"84",
          2373 => x"b4",
          2374 => x"80",
          2375 => x"87",
          2376 => x"84",
          2377 => x"54",
          2378 => x"51",
          2379 => x"ba",
          2380 => x"a5",
          2381 => x"70",
          2382 => x"fe",
          2383 => x"ff",
          2384 => x"59",
          2385 => x"b4",
          2386 => x"b8",
          2387 => x"34",
          2388 => x"fa",
          2389 => x"8f",
          2390 => x"fa",
          2391 => x"81",
          2392 => x"83",
          2393 => x"b2",
          2394 => x"d5",
          2395 => x"e5",
          2396 => x"59",
          2397 => x"3f",
          2398 => x"a6",
          2399 => x"83",
          2400 => x"81",
          2401 => x"d8",
          2402 => x"05",
          2403 => x"83",
          2404 => x"72",
          2405 => x"11",
          2406 => x"5c",
          2407 => x"ff",
          2408 => x"51",
          2409 => x"e9",
          2410 => x"75",
          2411 => x"2e",
          2412 => x"d5",
          2413 => x"b4",
          2414 => x"29",
          2415 => x"16",
          2416 => x"84",
          2417 => x"83",
          2418 => x"5a",
          2419 => x"18",
          2420 => x"29",
          2421 => x"86",
          2422 => x"f8",
          2423 => x"b2",
          2424 => x"29",
          2425 => x"fa",
          2426 => x"81",
          2427 => x"73",
          2428 => x"f9",
          2429 => x"17",
          2430 => x"b8",
          2431 => x"38",
          2432 => x"2e",
          2433 => x"84",
          2434 => x"2e",
          2435 => x"38",
          2436 => x"c1",
          2437 => x"3f",
          2438 => x"be",
          2439 => x"84",
          2440 => x"89",
          2441 => x"80",
          2442 => x"3f",
          2443 => x"54",
          2444 => x"52",
          2445 => x"70",
          2446 => x"27",
          2447 => x"fa",
          2448 => x"83",
          2449 => x"bb",
          2450 => x"80",
          2451 => x"38",
          2452 => x"06",
          2453 => x"73",
          2454 => x"52",
          2455 => x"b5",
          2456 => x"05",
          2457 => x"72",
          2458 => x"80",
          2459 => x"81",
          2460 => x"80",
          2461 => x"86",
          2462 => x"05",
          2463 => x"75",
          2464 => x"2e",
          2465 => x"b5",
          2466 => x"78",
          2467 => x"2e",
          2468 => x"83",
          2469 => x"72",
          2470 => x"b9",
          2471 => x"17",
          2472 => x"b5",
          2473 => x"29",
          2474 => x"fa",
          2475 => x"60",
          2476 => x"fa",
          2477 => x"05",
          2478 => x"ff",
          2479 => x"b5",
          2480 => x"5d",
          2481 => x"99",
          2482 => x"ff",
          2483 => x"b8",
          2484 => x"86",
          2485 => x"fa",
          2486 => x"0c",
          2487 => x"84",
          2488 => x"38",
          2489 => x"80",
          2490 => x"84",
          2491 => x"83",
          2492 => x"72",
          2493 => x"b9",
          2494 => x"1d",
          2495 => x"b5",
          2496 => x"29",
          2497 => x"fa",
          2498 => x"76",
          2499 => x"b0",
          2500 => x"84",
          2501 => x"83",
          2502 => x"72",
          2503 => x"59",
          2504 => x"d6",
          2505 => x"ff",
          2506 => x"38",
          2507 => x"84",
          2508 => x"78",
          2509 => x"24",
          2510 => x"81",
          2511 => x"fa",
          2512 => x"0c",
          2513 => x"82",
          2514 => x"26",
          2515 => x"81",
          2516 => x"34",
          2517 => x"81",
          2518 => x"88",
          2519 => x"0c",
          2520 => x"fd",
          2521 => x"0c",
          2522 => x"33",
          2523 => x"05",
          2524 => x"33",
          2525 => x"b8",
          2526 => x"fa",
          2527 => x"5f",
          2528 => x"34",
          2529 => x"19",
          2530 => x"c7",
          2531 => x"33",
          2532 => x"22",
          2533 => x"11",
          2534 => x"b0",
          2535 => x"81",
          2536 => x"81",
          2537 => x"fa",
          2538 => x"f8",
          2539 => x"ff",
          2540 => x"29",
          2541 => x"fa",
          2542 => x"29",
          2543 => x"f9",
          2544 => x"75",
          2545 => x"ff",
          2546 => x"95",
          2547 => x"34",
          2548 => x"84",
          2549 => x"80",
          2550 => x"84",
          2551 => x"80",
          2552 => x"9c",
          2553 => x"84",
          2554 => x"84",
          2555 => x"84",
          2556 => x"80",
          2557 => x"9c",
          2558 => x"09",
          2559 => x"b4",
          2560 => x"ff",
          2561 => x"ff",
          2562 => x"a0",
          2563 => x"40",
          2564 => x"ff",
          2565 => x"43",
          2566 => x"85",
          2567 => x"1a",
          2568 => x"76",
          2569 => x"06",
          2570 => x"06",
          2571 => x"84",
          2572 => x"1e",
          2573 => x"b5",
          2574 => x"29",
          2575 => x"83",
          2576 => x"33",
          2577 => x"83",
          2578 => x"1a",
          2579 => x"ff",
          2580 => x"b5",
          2581 => x"5a",
          2582 => x"84",
          2583 => x"81",
          2584 => x"95",
          2585 => x"79",
          2586 => x"83",
          2587 => x"70",
          2588 => x"fd",
          2589 => x"38",
          2590 => x"bf",
          2591 => x"33",
          2592 => x"19",
          2593 => x"75",
          2594 => x"77",
          2595 => x"34",
          2596 => x"80",
          2597 => x"0d",
          2598 => x"f8",
          2599 => x"b5",
          2600 => x"29",
          2601 => x"fa",
          2602 => x"05",
          2603 => x"8a",
          2604 => x"5b",
          2605 => x"5c",
          2606 => x"06",
          2607 => x"05",
          2608 => x"86",
          2609 => x"f8",
          2610 => x"b2",
          2611 => x"5e",
          2612 => x"34",
          2613 => x"1e",
          2614 => x"c7",
          2615 => x"33",
          2616 => x"22",
          2617 => x"11",
          2618 => x"b0",
          2619 => x"81",
          2620 => x"7e",
          2621 => x"f9",
          2622 => x"19",
          2623 => x"1c",
          2624 => x"83",
          2625 => x"33",
          2626 => x"33",
          2627 => x"06",
          2628 => x"05",
          2629 => x"b9",
          2630 => x"34",
          2631 => x"33",
          2632 => x"12",
          2633 => x"fa",
          2634 => x"76",
          2635 => x"b0",
          2636 => x"84",
          2637 => x"83",
          2638 => x"72",
          2639 => x"59",
          2640 => x"18",
          2641 => x"06",
          2642 => x"38",
          2643 => x"39",
          2644 => x"0b",
          2645 => x"04",
          2646 => x"b9",
          2647 => x"b5",
          2648 => x"05",
          2649 => x"ba",
          2650 => x"0c",
          2651 => x"17",
          2652 => x"7c",
          2653 => x"f8",
          2654 => x"5b",
          2655 => x"88",
          2656 => x"05",
          2657 => x"84",
          2658 => x"ba",
          2659 => x"84",
          2660 => x"06",
          2661 => x"84",
          2662 => x"83",
          2663 => x"80",
          2664 => x"33",
          2665 => x"33",
          2666 => x"b8",
          2667 => x"fa",
          2668 => x"5d",
          2669 => x"86",
          2670 => x"f8",
          2671 => x"b2",
          2672 => x"5b",
          2673 => x"83",
          2674 => x"41",
          2675 => x"c7",
          2676 => x"33",
          2677 => x"22",
          2678 => x"11",
          2679 => x"b0",
          2680 => x"1c",
          2681 => x"7b",
          2682 => x"33",
          2683 => x"56",
          2684 => x"84",
          2685 => x"40",
          2686 => x"b8",
          2687 => x"78",
          2688 => x"0b",
          2689 => x"04",
          2690 => x"34",
          2691 => x"34",
          2692 => x"fa",
          2693 => x"b4",
          2694 => x"b5",
          2695 => x"b3",
          2696 => x"39",
          2697 => x"2e",
          2698 => x"5d",
          2699 => x"85",
          2700 => x"55",
          2701 => x"9b",
          2702 => x"70",
          2703 => x"51",
          2704 => x"08",
          2705 => x"57",
          2706 => x"cd",
          2707 => x"fe",
          2708 => x"0b",
          2709 => x"81",
          2710 => x"ad",
          2711 => x"81",
          2712 => x"8a",
          2713 => x"b4",
          2714 => x"85",
          2715 => x"38",
          2716 => x"33",
          2717 => x"2c",
          2718 => x"75",
          2719 => x"84",
          2720 => x"8e",
          2721 => x"05",
          2722 => x"33",
          2723 => x"c5",
          2724 => x"bd",
          2725 => x"83",
          2726 => x"5d",
          2727 => x"ff",
          2728 => x"fd",
          2729 => x"34",
          2730 => x"33",
          2731 => x"fd",
          2732 => x"fa",
          2733 => x"85",
          2734 => x"38",
          2735 => x"33",
          2736 => x"2c",
          2737 => x"75",
          2738 => x"84",
          2739 => x"fc",
          2740 => x"60",
          2741 => x"38",
          2742 => x"33",
          2743 => x"12",
          2744 => x"b2",
          2745 => x"29",
          2746 => x"f9",
          2747 => x"42",
          2748 => x"2e",
          2749 => x"89",
          2750 => x"33",
          2751 => x"84",
          2752 => x"09",
          2753 => x"83",
          2754 => x"ba",
          2755 => x"be",
          2756 => x"b5",
          2757 => x"33",
          2758 => x"25",
          2759 => x"b5",
          2760 => x"33",
          2761 => x"84",
          2762 => x"42",
          2763 => x"11",
          2764 => x"38",
          2765 => x"fa",
          2766 => x"e7",
          2767 => x"33",
          2768 => x"38",
          2769 => x"22",
          2770 => x"e6",
          2771 => x"06",
          2772 => x"da",
          2773 => x"5f",
          2774 => x"ba",
          2775 => x"38",
          2776 => x"06",
          2777 => x"84",
          2778 => x"8e",
          2779 => x"05",
          2780 => x"33",
          2781 => x"b8",
          2782 => x"11",
          2783 => x"77",
          2784 => x"83",
          2785 => x"ff",
          2786 => x"38",
          2787 => x"84",
          2788 => x"7a",
          2789 => x"75",
          2790 => x"84",
          2791 => x"8a",
          2792 => x"b8",
          2793 => x"f9",
          2794 => x"b8",
          2795 => x"fa",
          2796 => x"c7",
          2797 => x"5f",
          2798 => x"ff",
          2799 => x"52",
          2800 => x"84",
          2801 => x"70",
          2802 => x"8e",
          2803 => x"76",
          2804 => x"56",
          2805 => x"ff",
          2806 => x"60",
          2807 => x"33",
          2808 => x"ff",
          2809 => x"7e",
          2810 => x"57",
          2811 => x"38",
          2812 => x"ff",
          2813 => x"79",
          2814 => x"c7",
          2815 => x"81",
          2816 => x"58",
          2817 => x"38",
          2818 => x"17",
          2819 => x"7b",
          2820 => x"81",
          2821 => x"5e",
          2822 => x"84",
          2823 => x"43",
          2824 => x"9d",
          2825 => x"b9",
          2826 => x"5d",
          2827 => x"7c",
          2828 => x"84",
          2829 => x"71",
          2830 => x"7f",
          2831 => x"39",
          2832 => x"2e",
          2833 => x"d9",
          2834 => x"39",
          2835 => x"11",
          2836 => x"58",
          2837 => x"d8",
          2838 => x"06",
          2839 => x"58",
          2840 => x"33",
          2841 => x"81",
          2842 => x"7a",
          2843 => x"ff",
          2844 => x"38",
          2845 => x"57",
          2846 => x"1b",
          2847 => x"a0",
          2848 => x"c7",
          2849 => x"51",
          2850 => x"06",
          2851 => x"b0",
          2852 => x"07",
          2853 => x"7f",
          2854 => x"9e",
          2855 => x"0c",
          2856 => x"79",
          2857 => x"33",
          2858 => x"81",
          2859 => x"fa",
          2860 => x"59",
          2861 => x"38",
          2862 => x"62",
          2863 => x"57",
          2864 => x"fa",
          2865 => x"5a",
          2866 => x"78",
          2867 => x"57",
          2868 => x"0b",
          2869 => x"81",
          2870 => x"77",
          2871 => x"1f",
          2872 => x"8a",
          2873 => x"f0",
          2874 => x"71",
          2875 => x"80",
          2876 => x"80",
          2877 => x"18",
          2878 => x"b6",
          2879 => x"84",
          2880 => x"fa",
          2881 => x"fa",
          2882 => x"5c",
          2883 => x"b0",
          2884 => x"b0",
          2885 => x"59",
          2886 => x"33",
          2887 => x"83",
          2888 => x"b0",
          2889 => x"75",
          2890 => x"fa",
          2891 => x"56",
          2892 => x"83",
          2893 => x"07",
          2894 => x"b1",
          2895 => x"34",
          2896 => x"56",
          2897 => x"81",
          2898 => x"34",
          2899 => x"81",
          2900 => x"fa",
          2901 => x"b0",
          2902 => x"56",
          2903 => x"39",
          2904 => x"80",
          2905 => x"34",
          2906 => x"81",
          2907 => x"fa",
          2908 => x"b0",
          2909 => x"75",
          2910 => x"83",
          2911 => x"07",
          2912 => x"a1",
          2913 => x"06",
          2914 => x"34",
          2915 => x"81",
          2916 => x"34",
          2917 => x"80",
          2918 => x"34",
          2919 => x"80",
          2920 => x"34",
          2921 => x"81",
          2922 => x"83",
          2923 => x"fa",
          2924 => x"56",
          2925 => x"39",
          2926 => x"52",
          2927 => x"39",
          2928 => x"34",
          2929 => x"34",
          2930 => x"fa",
          2931 => x"0c",
          2932 => x"87",
          2933 => x"9c",
          2934 => x"34",
          2935 => x"06",
          2936 => x"84",
          2937 => x"53",
          2938 => x"84",
          2939 => x"84",
          2940 => x"84",
          2941 => x"84",
          2942 => x"fa",
          2943 => x"85",
          2944 => x"ba",
          2945 => x"5d",
          2946 => x"d8",
          2947 => x"34",
          2948 => x"34",
          2949 => x"83",
          2950 => x"58",
          2951 => x"0b",
          2952 => x"51",
          2953 => x"51",
          2954 => x"83",
          2955 => x"70",
          2956 => x"f2",
          2957 => x"39",
          2958 => x"27",
          2959 => x"34",
          2960 => x"ff",
          2961 => x"06",
          2962 => x"fa",
          2963 => x"33",
          2964 => x"25",
          2965 => x"39",
          2966 => x"06",
          2967 => x"38",
          2968 => x"33",
          2969 => x"33",
          2970 => x"80",
          2971 => x"71",
          2972 => x"06",
          2973 => x"42",
          2974 => x"38",
          2975 => x"5c",
          2976 => x"84",
          2977 => x"83",
          2978 => x"fa",
          2979 => x"11",
          2980 => x"38",
          2981 => x"27",
          2982 => x"83",
          2983 => x"83",
          2984 => x"76",
          2985 => x"81",
          2986 => x"29",
          2987 => x"a0",
          2988 => x"81",
          2989 => x"71",
          2990 => x"7e",
          2991 => x"1a",
          2992 => x"b9",
          2993 => x"5d",
          2994 => x"7d",
          2995 => x"84",
          2996 => x"71",
          2997 => x"77",
          2998 => x"17",
          2999 => x"7b",
          3000 => x"81",
          3001 => x"5f",
          3002 => x"84",
          3003 => x"59",
          3004 => x"99",
          3005 => x"17",
          3006 => x"7b",
          3007 => x"f8",
          3008 => x"f7",
          3009 => x"39",
          3010 => x"33",
          3011 => x"42",
          3012 => x"5a",
          3013 => x"ff",
          3014 => x"27",
          3015 => x"b4",
          3016 => x"ff",
          3017 => x"78",
          3018 => x"83",
          3019 => x"fa",
          3020 => x"33",
          3021 => x"25",
          3022 => x"39",
          3023 => x"c0",
          3024 => x"ff",
          3025 => x"5d",
          3026 => x"06",
          3027 => x"1d",
          3028 => x"93",
          3029 => x"b2",
          3030 => x"56",
          3031 => x"39",
          3032 => x"f5",
          3033 => x"58",
          3034 => x"81",
          3035 => x"ec",
          3036 => x"34",
          3037 => x"05",
          3038 => x"f4",
          3039 => x"83",
          3040 => x"0b",
          3041 => x"7e",
          3042 => x"80",
          3043 => x"39",
          3044 => x"a7",
          3045 => x"84",
          3046 => x"0b",
          3047 => x"fd",
          3048 => x"b8",
          3049 => x"90",
          3050 => x"0b",
          3051 => x"04",
          3052 => x"80",
          3053 => x"0d",
          3054 => x"33",
          3055 => x"70",
          3056 => x"33",
          3057 => x"80",
          3058 => x"f9",
          3059 => x"84",
          3060 => x"e4",
          3061 => x"91",
          3062 => x"07",
          3063 => x"5e",
          3064 => x"59",
          3065 => x"06",
          3066 => x"70",
          3067 => x"5c",
          3068 => x"84",
          3069 => x"83",
          3070 => x"86",
          3071 => x"22",
          3072 => x"70",
          3073 => x"33",
          3074 => x"83",
          3075 => x"8e",
          3076 => x"98",
          3077 => x"56",
          3078 => x"80",
          3079 => x"15",
          3080 => x"55",
          3081 => x"80",
          3082 => x"81",
          3083 => x"58",
          3084 => x"38",
          3085 => x"74",
          3086 => x"ff",
          3087 => x"cd",
          3088 => x"83",
          3089 => x"15",
          3090 => x"55",
          3091 => x"83",
          3092 => x"80",
          3093 => x"dc",
          3094 => x"2a",
          3095 => x"58",
          3096 => x"0b",
          3097 => x"06",
          3098 => x"81",
          3099 => x"83",
          3100 => x"83",
          3101 => x"33",
          3102 => x"5e",
          3103 => x"33",
          3104 => x"83",
          3105 => x"2e",
          3106 => x"33",
          3107 => x"83",
          3108 => x"ec",
          3109 => x"81",
          3110 => x"16",
          3111 => x"38",
          3112 => x"ff",
          3113 => x"16",
          3114 => x"38",
          3115 => x"87",
          3116 => x"73",
          3117 => x"c0",
          3118 => x"58",
          3119 => x"54",
          3120 => x"83",
          3121 => x"34",
          3122 => x"82",
          3123 => x"fc",
          3124 => x"8c",
          3125 => x"83",
          3126 => x"5e",
          3127 => x"80",
          3128 => x"72",
          3129 => x"83",
          3130 => x"08",
          3131 => x"06",
          3132 => x"fa",
          3133 => x"14",
          3134 => x"a5",
          3135 => x"80",
          3136 => x"83",
          3137 => x"f0",
          3138 => x"e0",
          3139 => x"7c",
          3140 => x"09",
          3141 => x"2e",
          3142 => x"d7",
          3143 => x"77",
          3144 => x"80",
          3145 => x"38",
          3146 => x"10",
          3147 => x"98",
          3148 => x"73",
          3149 => x"79",
          3150 => x"05",
          3151 => x"56",
          3152 => x"83",
          3153 => x"80",
          3154 => x"79",
          3155 => x"82",
          3156 => x"fa",
          3157 => x"33",
          3158 => x"38",
          3159 => x"25",
          3160 => x"38",
          3161 => x"cc",
          3162 => x"80",
          3163 => x"90",
          3164 => x"2e",
          3165 => x"ff",
          3166 => x"38",
          3167 => x"2e",
          3168 => x"55",
          3169 => x"06",
          3170 => x"84",
          3171 => x"be",
          3172 => x"39",
          3173 => x"f8",
          3174 => x"83",
          3175 => x"80",
          3176 => x"0b",
          3177 => x"83",
          3178 => x"74",
          3179 => x"2e",
          3180 => x"33",
          3181 => x"77",
          3182 => x"09",
          3183 => x"d8",
          3184 => x"9c",
          3185 => x"e8",
          3186 => x"f8",
          3187 => x"fb",
          3188 => x"15",
          3189 => x"dd",
          3190 => x"fa",
          3191 => x"80",
          3192 => x"e4",
          3193 => x"f8",
          3194 => x"5d",
          3195 => x"39",
          3196 => x"cb",
          3197 => x"ce",
          3198 => x"fc",
          3199 => x"34",
          3200 => x"0b",
          3201 => x"83",
          3202 => x"34",
          3203 => x"84",
          3204 => x"38",
          3205 => x"ff",
          3206 => x"f8",
          3207 => x"84",
          3208 => x"39",
          3209 => x"06",
          3210 => x"27",
          3211 => x"b2",
          3212 => x"55",
          3213 => x"54",
          3214 => x"f8",
          3215 => x"05",
          3216 => x"53",
          3217 => x"f6",
          3218 => x"ba",
          3219 => x"72",
          3220 => x"52",
          3221 => x"3f",
          3222 => x"f8",
          3223 => x"3d",
          3224 => x"3d",
          3225 => x"83",
          3226 => x"05",
          3227 => x"08",
          3228 => x"83",
          3229 => x"81",
          3230 => x"e8",
          3231 => x"f5",
          3232 => x"53",
          3233 => x"c0",
          3234 => x"f6",
          3235 => x"9c",
          3236 => x"38",
          3237 => x"c0",
          3238 => x"73",
          3239 => x"ff",
          3240 => x"9c",
          3241 => x"c0",
          3242 => x"9c",
          3243 => x"81",
          3244 => x"52",
          3245 => x"81",
          3246 => x"a4",
          3247 => x"ff",
          3248 => x"ff",
          3249 => x"38",
          3250 => x"d5",
          3251 => x"84",
          3252 => x"81",
          3253 => x"0d",
          3254 => x"05",
          3255 => x"83",
          3256 => x"fc",
          3257 => x"07",
          3258 => x"34",
          3259 => x"34",
          3260 => x"34",
          3261 => x"08",
          3262 => x"90",
          3263 => x"0b",
          3264 => x"0b",
          3265 => x"80",
          3266 => x"83",
          3267 => x"05",
          3268 => x"87",
          3269 => x"2e",
          3270 => x"98",
          3271 => x"87",
          3272 => x"87",
          3273 => x"70",
          3274 => x"71",
          3275 => x"98",
          3276 => x"87",
          3277 => x"98",
          3278 => x"38",
          3279 => x"08",
          3280 => x"71",
          3281 => x"98",
          3282 => x"38",
          3283 => x"81",
          3284 => x"80",
          3285 => x"71",
          3286 => x"ff",
          3287 => x"14",
          3288 => x"70",
          3289 => x"05",
          3290 => x"34",
          3291 => x"bb",
          3292 => x"0b",
          3293 => x"04",
          3294 => x"79",
          3295 => x"56",
          3296 => x"88",
          3297 => x"79",
          3298 => x"75",
          3299 => x"70",
          3300 => x"71",
          3301 => x"7a",
          3302 => x"84",
          3303 => x"73",
          3304 => x"52",
          3305 => x"72",
          3306 => x"08",
          3307 => x"90",
          3308 => x"0b",
          3309 => x"0b",
          3310 => x"80",
          3311 => x"83",
          3312 => x"05",
          3313 => x"87",
          3314 => x"2e",
          3315 => x"98",
          3316 => x"87",
          3317 => x"87",
          3318 => x"70",
          3319 => x"71",
          3320 => x"98",
          3321 => x"87",
          3322 => x"98",
          3323 => x"38",
          3324 => x"08",
          3325 => x"71",
          3326 => x"98",
          3327 => x"38",
          3328 => x"81",
          3329 => x"a1",
          3330 => x"fe",
          3331 => x"06",
          3332 => x"57",
          3333 => x"0d",
          3334 => x"0d",
          3335 => x"71",
          3336 => x"56",
          3337 => x"0b",
          3338 => x"98",
          3339 => x"80",
          3340 => x"9c",
          3341 => x"53",
          3342 => x"33",
          3343 => x"70",
          3344 => x"2e",
          3345 => x"51",
          3346 => x"38",
          3347 => x"38",
          3348 => x"90",
          3349 => x"52",
          3350 => x"72",
          3351 => x"c0",
          3352 => x"27",
          3353 => x"38",
          3354 => x"71",
          3355 => x"ff",
          3356 => x"75",
          3357 => x"06",
          3358 => x"80",
          3359 => x"ce",
          3360 => x"3d",
          3361 => x"31",
          3362 => x"70",
          3363 => x"12",
          3364 => x"07",
          3365 => x"71",
          3366 => x"54",
          3367 => x"56",
          3368 => x"38",
          3369 => x"33",
          3370 => x"76",
          3371 => x"98",
          3372 => x"5c",
          3373 => x"83",
          3374 => x"33",
          3375 => x"75",
          3376 => x"57",
          3377 => x"06",
          3378 => x"f4",
          3379 => x"13",
          3380 => x"2a",
          3381 => x"14",
          3382 => x"f4",
          3383 => x"34",
          3384 => x"f4",
          3385 => x"85",
          3386 => x"70",
          3387 => x"07",
          3388 => x"58",
          3389 => x"81",
          3390 => x"12",
          3391 => x"71",
          3392 => x"33",
          3393 => x"70",
          3394 => x"58",
          3395 => x"12",
          3396 => x"84",
          3397 => x"2b",
          3398 => x"52",
          3399 => x"33",
          3400 => x"52",
          3401 => x"72",
          3402 => x"15",
          3403 => x"2b",
          3404 => x"2a",
          3405 => x"77",
          3406 => x"70",
          3407 => x"8b",
          3408 => x"70",
          3409 => x"07",
          3410 => x"77",
          3411 => x"54",
          3412 => x"14",
          3413 => x"f4",
          3414 => x"33",
          3415 => x"74",
          3416 => x"88",
          3417 => x"88",
          3418 => x"54",
          3419 => x"34",
          3420 => x"11",
          3421 => x"71",
          3422 => x"81",
          3423 => x"2b",
          3424 => x"53",
          3425 => x"71",
          3426 => x"07",
          3427 => x"59",
          3428 => x"16",
          3429 => x"70",
          3430 => x"71",
          3431 => x"33",
          3432 => x"70",
          3433 => x"56",
          3434 => x"83",
          3435 => x"3d",
          3436 => x"58",
          3437 => x"2e",
          3438 => x"89",
          3439 => x"84",
          3440 => x"ba",
          3441 => x"52",
          3442 => x"3f",
          3443 => x"34",
          3444 => x"f4",
          3445 => x"0b",
          3446 => x"56",
          3447 => x"17",
          3448 => x"f0",
          3449 => x"70",
          3450 => x"58",
          3451 => x"73",
          3452 => x"70",
          3453 => x"05",
          3454 => x"34",
          3455 => x"39",
          3456 => x"81",
          3457 => x"12",
          3458 => x"ff",
          3459 => x"06",
          3460 => x"85",
          3461 => x"52",
          3462 => x"54",
          3463 => x"10",
          3464 => x"33",
          3465 => x"ff",
          3466 => x"06",
          3467 => x"54",
          3468 => x"80",
          3469 => x"84",
          3470 => x"2b",
          3471 => x"81",
          3472 => x"54",
          3473 => x"70",
          3474 => x"07",
          3475 => x"5d",
          3476 => x"38",
          3477 => x"82",
          3478 => x"82",
          3479 => x"38",
          3480 => x"74",
          3481 => x"5b",
          3482 => x"78",
          3483 => x"15",
          3484 => x"14",
          3485 => x"f4",
          3486 => x"33",
          3487 => x"8f",
          3488 => x"ff",
          3489 => x"53",
          3490 => x"34",
          3491 => x"12",
          3492 => x"75",
          3493 => x"ba",
          3494 => x"87",
          3495 => x"2b",
          3496 => x"57",
          3497 => x"34",
          3498 => x"78",
          3499 => x"71",
          3500 => x"54",
          3501 => x"87",
          3502 => x"19",
          3503 => x"8b",
          3504 => x"58",
          3505 => x"34",
          3506 => x"08",
          3507 => x"33",
          3508 => x"70",
          3509 => x"84",
          3510 => x"ba",
          3511 => x"84",
          3512 => x"86",
          3513 => x"2b",
          3514 => x"17",
          3515 => x"07",
          3516 => x"54",
          3517 => x"12",
          3518 => x"84",
          3519 => x"2b",
          3520 => x"14",
          3521 => x"07",
          3522 => x"56",
          3523 => x"76",
          3524 => x"18",
          3525 => x"2b",
          3526 => x"2a",
          3527 => x"74",
          3528 => x"18",
          3529 => x"3d",
          3530 => x"58",
          3531 => x"77",
          3532 => x"89",
          3533 => x"3f",
          3534 => x"0c",
          3535 => x"0b",
          3536 => x"84",
          3537 => x"76",
          3538 => x"ec",
          3539 => x"75",
          3540 => x"ba",
          3541 => x"81",
          3542 => x"08",
          3543 => x"87",
          3544 => x"ba",
          3545 => x"07",
          3546 => x"2a",
          3547 => x"34",
          3548 => x"22",
          3549 => x"08",
          3550 => x"15",
          3551 => x"54",
          3552 => x"e3",
          3553 => x"5f",
          3554 => x"45",
          3555 => x"7e",
          3556 => x"2e",
          3557 => x"27",
          3558 => x"82",
          3559 => x"58",
          3560 => x"31",
          3561 => x"70",
          3562 => x"12",
          3563 => x"31",
          3564 => x"10",
          3565 => x"11",
          3566 => x"2b",
          3567 => x"53",
          3568 => x"44",
          3569 => x"80",
          3570 => x"33",
          3571 => x"70",
          3572 => x"12",
          3573 => x"07",
          3574 => x"74",
          3575 => x"82",
          3576 => x"2e",
          3577 => x"f9",
          3578 => x"87",
          3579 => x"24",
          3580 => x"81",
          3581 => x"2b",
          3582 => x"33",
          3583 => x"47",
          3584 => x"80",
          3585 => x"82",
          3586 => x"2b",
          3587 => x"11",
          3588 => x"71",
          3589 => x"33",
          3590 => x"70",
          3591 => x"41",
          3592 => x"1d",
          3593 => x"f4",
          3594 => x"12",
          3595 => x"07",
          3596 => x"33",
          3597 => x"5f",
          3598 => x"77",
          3599 => x"84",
          3600 => x"12",
          3601 => x"ff",
          3602 => x"59",
          3603 => x"84",
          3604 => x"33",
          3605 => x"83",
          3606 => x"15",
          3607 => x"2a",
          3608 => x"55",
          3609 => x"84",
          3610 => x"81",
          3611 => x"2b",
          3612 => x"15",
          3613 => x"2a",
          3614 => x"55",
          3615 => x"34",
          3616 => x"11",
          3617 => x"07",
          3618 => x"42",
          3619 => x"51",
          3620 => x"08",
          3621 => x"70",
          3622 => x"7a",
          3623 => x"73",
          3624 => x"04",
          3625 => x"0c",
          3626 => x"82",
          3627 => x"f4",
          3628 => x"f4",
          3629 => x"81",
          3630 => x"60",
          3631 => x"34",
          3632 => x"1d",
          3633 => x"ba",
          3634 => x"05",
          3635 => x"ff",
          3636 => x"57",
          3637 => x"34",
          3638 => x"10",
          3639 => x"55",
          3640 => x"83",
          3641 => x"7e",
          3642 => x"8c",
          3643 => x"df",
          3644 => x"bb",
          3645 => x"3d",
          3646 => x"08",
          3647 => x"7f",
          3648 => x"88",
          3649 => x"88",
          3650 => x"7b",
          3651 => x"ba",
          3652 => x"58",
          3653 => x"34",
          3654 => x"33",
          3655 => x"70",
          3656 => x"05",
          3657 => x"2a",
          3658 => x"63",
          3659 => x"06",
          3660 => x"ba",
          3661 => x"60",
          3662 => x"08",
          3663 => x"7e",
          3664 => x"70",
          3665 => x"ac",
          3666 => x"31",
          3667 => x"33",
          3668 => x"70",
          3669 => x"12",
          3670 => x"07",
          3671 => x"54",
          3672 => x"bc",
          3673 => x"80",
          3674 => x"ff",
          3675 => x"dd",
          3676 => x"0b",
          3677 => x"84",
          3678 => x"7e",
          3679 => x"84",
          3680 => x"7a",
          3681 => x"ba",
          3682 => x"81",
          3683 => x"08",
          3684 => x"87",
          3685 => x"ba",
          3686 => x"07",
          3687 => x"2a",
          3688 => x"05",
          3689 => x"ba",
          3690 => x"ba",
          3691 => x"7e",
          3692 => x"05",
          3693 => x"83",
          3694 => x"5b",
          3695 => x"f2",
          3696 => x"7e",
          3697 => x"84",
          3698 => x"76",
          3699 => x"71",
          3700 => x"11",
          3701 => x"8b",
          3702 => x"84",
          3703 => x"2b",
          3704 => x"56",
          3705 => x"78",
          3706 => x"05",
          3707 => x"84",
          3708 => x"2b",
          3709 => x"14",
          3710 => x"07",
          3711 => x"5d",
          3712 => x"34",
          3713 => x"f4",
          3714 => x"71",
          3715 => x"70",
          3716 => x"7d",
          3717 => x"f4",
          3718 => x"12",
          3719 => x"07",
          3720 => x"71",
          3721 => x"5c",
          3722 => x"7c",
          3723 => x"f4",
          3724 => x"33",
          3725 => x"74",
          3726 => x"71",
          3727 => x"47",
          3728 => x"82",
          3729 => x"ba",
          3730 => x"83",
          3731 => x"57",
          3732 => x"58",
          3733 => x"bc",
          3734 => x"84",
          3735 => x"5f",
          3736 => x"84",
          3737 => x"ba",
          3738 => x"52",
          3739 => x"3f",
          3740 => x"34",
          3741 => x"f4",
          3742 => x"0b",
          3743 => x"54",
          3744 => x"15",
          3745 => x"f0",
          3746 => x"70",
          3747 => x"45",
          3748 => x"60",
          3749 => x"70",
          3750 => x"05",
          3751 => x"34",
          3752 => x"e7",
          3753 => x"86",
          3754 => x"2b",
          3755 => x"1c",
          3756 => x"07",
          3757 => x"59",
          3758 => x"61",
          3759 => x"70",
          3760 => x"71",
          3761 => x"05",
          3762 => x"88",
          3763 => x"48",
          3764 => x"86",
          3765 => x"84",
          3766 => x"12",
          3767 => x"ff",
          3768 => x"58",
          3769 => x"84",
          3770 => x"81",
          3771 => x"2b",
          3772 => x"33",
          3773 => x"8f",
          3774 => x"2a",
          3775 => x"44",
          3776 => x"17",
          3777 => x"70",
          3778 => x"71",
          3779 => x"81",
          3780 => x"ff",
          3781 => x"5e",
          3782 => x"34",
          3783 => x"ff",
          3784 => x"15",
          3785 => x"71",
          3786 => x"33",
          3787 => x"70",
          3788 => x"5d",
          3789 => x"34",
          3790 => x"11",
          3791 => x"71",
          3792 => x"33",
          3793 => x"70",
          3794 => x"42",
          3795 => x"75",
          3796 => x"08",
          3797 => x"88",
          3798 => x"88",
          3799 => x"34",
          3800 => x"08",
          3801 => x"71",
          3802 => x"05",
          3803 => x"2b",
          3804 => x"06",
          3805 => x"5f",
          3806 => x"82",
          3807 => x"ba",
          3808 => x"12",
          3809 => x"07",
          3810 => x"71",
          3811 => x"70",
          3812 => x"59",
          3813 => x"1d",
          3814 => x"82",
          3815 => x"2b",
          3816 => x"11",
          3817 => x"71",
          3818 => x"33",
          3819 => x"70",
          3820 => x"42",
          3821 => x"84",
          3822 => x"ba",
          3823 => x"85",
          3824 => x"2b",
          3825 => x"15",
          3826 => x"2a",
          3827 => x"57",
          3828 => x"34",
          3829 => x"81",
          3830 => x"ff",
          3831 => x"5e",
          3832 => x"34",
          3833 => x"11",
          3834 => x"71",
          3835 => x"81",
          3836 => x"88",
          3837 => x"55",
          3838 => x"34",
          3839 => x"33",
          3840 => x"83",
          3841 => x"83",
          3842 => x"88",
          3843 => x"55",
          3844 => x"1a",
          3845 => x"82",
          3846 => x"2b",
          3847 => x"2b",
          3848 => x"05",
          3849 => x"f4",
          3850 => x"1c",
          3851 => x"5f",
          3852 => x"1a",
          3853 => x"07",
          3854 => x"33",
          3855 => x"40",
          3856 => x"84",
          3857 => x"84",
          3858 => x"33",
          3859 => x"83",
          3860 => x"87",
          3861 => x"88",
          3862 => x"41",
          3863 => x"64",
          3864 => x"1d",
          3865 => x"2b",
          3866 => x"2a",
          3867 => x"7c",
          3868 => x"70",
          3869 => x"8b",
          3870 => x"70",
          3871 => x"07",
          3872 => x"77",
          3873 => x"49",
          3874 => x"1e",
          3875 => x"f4",
          3876 => x"33",
          3877 => x"74",
          3878 => x"88",
          3879 => x"88",
          3880 => x"5e",
          3881 => x"34",
          3882 => x"83",
          3883 => x"3f",
          3884 => x"84",
          3885 => x"73",
          3886 => x"b3",
          3887 => x"61",
          3888 => x"f0",
          3889 => x"29",
          3890 => x"80",
          3891 => x"38",
          3892 => x"0d",
          3893 => x"bb",
          3894 => x"80",
          3895 => x"84",
          3896 => x"3f",
          3897 => x"0d",
          3898 => x"f4",
          3899 => x"23",
          3900 => x"ff",
          3901 => x"ba",
          3902 => x"0b",
          3903 => x"54",
          3904 => x"15",
          3905 => x"86",
          3906 => x"84",
          3907 => x"ff",
          3908 => x"ff",
          3909 => x"55",
          3910 => x"17",
          3911 => x"10",
          3912 => x"05",
          3913 => x"0b",
          3914 => x"2e",
          3915 => x"3d",
          3916 => x"52",
          3917 => x"80",
          3918 => x"0c",
          3919 => x"02",
          3920 => x"81",
          3921 => x"3f",
          3922 => x"53",
          3923 => x"13",
          3924 => x"72",
          3925 => x"04",
          3926 => x"8c",
          3927 => x"59",
          3928 => x"84",
          3929 => x"06",
          3930 => x"58",
          3931 => x"78",
          3932 => x"3f",
          3933 => x"55",
          3934 => x"98",
          3935 => x"78",
          3936 => x"06",
          3937 => x"54",
          3938 => x"8b",
          3939 => x"19",
          3940 => x"79",
          3941 => x"f7",
          3942 => x"05",
          3943 => x"81",
          3944 => x"bb",
          3945 => x"54",
          3946 => x"85",
          3947 => x"53",
          3948 => x"84",
          3949 => x"74",
          3950 => x"8c",
          3951 => x"26",
          3952 => x"54",
          3953 => x"73",
          3954 => x"3d",
          3955 => x"70",
          3956 => x"78",
          3957 => x"3d",
          3958 => x"33",
          3959 => x"53",
          3960 => x"38",
          3961 => x"81",
          3962 => x"85",
          3963 => x"53",
          3964 => x"25",
          3965 => x"84",
          3966 => x"3d",
          3967 => x"73",
          3968 => x"04",
          3969 => x"bb",
          3970 => x"84",
          3971 => x"54",
          3972 => x"2a",
          3973 => x"8a",
          3974 => x"74",
          3975 => x"51",
          3976 => x"c0",
          3977 => x"06",
          3978 => x"71",
          3979 => x"ff",
          3980 => x"80",
          3981 => x"57",
          3982 => x"38",
          3983 => x"87",
          3984 => x"33",
          3985 => x"08",
          3986 => x"84",
          3987 => x"81",
          3988 => x"70",
          3989 => x"ff",
          3990 => x"77",
          3991 => x"bb",
          3992 => x"08",
          3993 => x"08",
          3994 => x"5b",
          3995 => x"18",
          3996 => x"06",
          3997 => x"53",
          3998 => x"b7",
          3999 => x"83",
          4000 => x"84",
          4001 => x"81",
          4002 => x"84",
          4003 => x"81",
          4004 => x"f4",
          4005 => x"34",
          4006 => x"80",
          4007 => x"19",
          4008 => x"80",
          4009 => x"0b",
          4010 => x"84",
          4011 => x"9e",
          4012 => x"19",
          4013 => x"a0",
          4014 => x"84",
          4015 => x"75",
          4016 => x"5b",
          4017 => x"08",
          4018 => x"88",
          4019 => x"7a",
          4020 => x"34",
          4021 => x"19",
          4022 => x"b4",
          4023 => x"79",
          4024 => x"3f",
          4025 => x"52",
          4026 => x"84",
          4027 => x"38",
          4028 => x"60",
          4029 => x"27",
          4030 => x"8c",
          4031 => x"0c",
          4032 => x"56",
          4033 => x"74",
          4034 => x"2e",
          4035 => x"2a",
          4036 => x"05",
          4037 => x"79",
          4038 => x"7b",
          4039 => x"38",
          4040 => x"81",
          4041 => x"bb",
          4042 => x"59",
          4043 => x"ff",
          4044 => x"b8",
          4045 => x"a8",
          4046 => x"b4",
          4047 => x"0b",
          4048 => x"74",
          4049 => x"38",
          4050 => x"81",
          4051 => x"bb",
          4052 => x"59",
          4053 => x"fe",
          4054 => x"b8",
          4055 => x"78",
          4056 => x"59",
          4057 => x"9f",
          4058 => x"3d",
          4059 => x"08",
          4060 => x"b5",
          4061 => x"5c",
          4062 => x"06",
          4063 => x"b8",
          4064 => x"a8",
          4065 => x"85",
          4066 => x"18",
          4067 => x"83",
          4068 => x"11",
          4069 => x"84",
          4070 => x"0d",
          4071 => x"fd",
          4072 => x"08",
          4073 => x"b5",
          4074 => x"5c",
          4075 => x"06",
          4076 => x"b8",
          4077 => x"c0",
          4078 => x"85",
          4079 => x"18",
          4080 => x"2b",
          4081 => x"83",
          4082 => x"2b",
          4083 => x"70",
          4084 => x"80",
          4085 => x"bb",
          4086 => x"56",
          4087 => x"17",
          4088 => x"18",
          4089 => x"5a",
          4090 => x"81",
          4091 => x"08",
          4092 => x"18",
          4093 => x"5e",
          4094 => x"38",
          4095 => x"09",
          4096 => x"b4",
          4097 => x"7b",
          4098 => x"3f",
          4099 => x"b4",
          4100 => x"81",
          4101 => x"84",
          4102 => x"06",
          4103 => x"83",
          4104 => x"08",
          4105 => x"8b",
          4106 => x"2e",
          4107 => x"5b",
          4108 => x"08",
          4109 => x"33",
          4110 => x"84",
          4111 => x"06",
          4112 => x"83",
          4113 => x"08",
          4114 => x"7d",
          4115 => x"82",
          4116 => x"81",
          4117 => x"17",
          4118 => x"52",
          4119 => x"7a",
          4120 => x"17",
          4121 => x"18",
          4122 => x"5a",
          4123 => x"81",
          4124 => x"08",
          4125 => x"18",
          4126 => x"55",
          4127 => x"38",
          4128 => x"09",
          4129 => x"b4",
          4130 => x"7d",
          4131 => x"3f",
          4132 => x"b4",
          4133 => x"7b",
          4134 => x"3f",
          4135 => x"bb",
          4136 => x"60",
          4137 => x"81",
          4138 => x"08",
          4139 => x"78",
          4140 => x"80",
          4141 => x"77",
          4142 => x"04",
          4143 => x"58",
          4144 => x"76",
          4145 => x"33",
          4146 => x"81",
          4147 => x"53",
          4148 => x"f2",
          4149 => x"2e",
          4150 => x"b4",
          4151 => x"38",
          4152 => x"7b",
          4153 => x"b8",
          4154 => x"b9",
          4155 => x"77",
          4156 => x"04",
          4157 => x"ff",
          4158 => x"05",
          4159 => x"5c",
          4160 => x"19",
          4161 => x"09",
          4162 => x"77",
          4163 => x"51",
          4164 => x"80",
          4165 => x"77",
          4166 => x"b7",
          4167 => x"79",
          4168 => x"98",
          4169 => x"06",
          4170 => x"34",
          4171 => x"34",
          4172 => x"34",
          4173 => x"34",
          4174 => x"39",
          4175 => x"a8",
          4176 => x"59",
          4177 => x"0b",
          4178 => x"74",
          4179 => x"38",
          4180 => x"81",
          4181 => x"bb",
          4182 => x"58",
          4183 => x"58",
          4184 => x"06",
          4185 => x"06",
          4186 => x"2e",
          4187 => x"06",
          4188 => x"5a",
          4189 => x"34",
          4190 => x"56",
          4191 => x"74",
          4192 => x"74",
          4193 => x"33",
          4194 => x"84",
          4195 => x"06",
          4196 => x"83",
          4197 => x"1b",
          4198 => x"84",
          4199 => x"27",
          4200 => x"82",
          4201 => x"53",
          4202 => x"d8",
          4203 => x"85",
          4204 => x"1a",
          4205 => x"ff",
          4206 => x"56",
          4207 => x"76",
          4208 => x"07",
          4209 => x"83",
          4210 => x"76",
          4211 => x"33",
          4212 => x"84",
          4213 => x"06",
          4214 => x"83",
          4215 => x"1b",
          4216 => x"84",
          4217 => x"27",
          4218 => x"74",
          4219 => x"38",
          4220 => x"81",
          4221 => x"5a",
          4222 => x"b8",
          4223 => x"57",
          4224 => x"84",
          4225 => x"ae",
          4226 => x"34",
          4227 => x"31",
          4228 => x"5f",
          4229 => x"f0",
          4230 => x"2e",
          4231 => x"54",
          4232 => x"33",
          4233 => x"d0",
          4234 => x"70",
          4235 => x"cf",
          4236 => x"7c",
          4237 => x"84",
          4238 => x"19",
          4239 => x"1b",
          4240 => x"40",
          4241 => x"82",
          4242 => x"81",
          4243 => x"1e",
          4244 => x"ed",
          4245 => x"81",
          4246 => x"19",
          4247 => x"fd",
          4248 => x"06",
          4249 => x"59",
          4250 => x"88",
          4251 => x"fa",
          4252 => x"76",
          4253 => x"b8",
          4254 => x"8f",
          4255 => x"42",
          4256 => x"7d",
          4257 => x"7d",
          4258 => x"7d",
          4259 => x"fa",
          4260 => x"71",
          4261 => x"38",
          4262 => x"80",
          4263 => x"80",
          4264 => x"54",
          4265 => x"7b",
          4266 => x"16",
          4267 => x"38",
          4268 => x"38",
          4269 => x"84",
          4270 => x"38",
          4271 => x"2e",
          4272 => x"70",
          4273 => x"7b",
          4274 => x"aa",
          4275 => x"ff",
          4276 => x"84",
          4277 => x"ff",
          4278 => x"ca",
          4279 => x"3f",
          4280 => x"27",
          4281 => x"84",
          4282 => x"9c",
          4283 => x"c4",
          4284 => x"1b",
          4285 => x"38",
          4286 => x"eb",
          4287 => x"81",
          4288 => x"08",
          4289 => x"25",
          4290 => x"54",
          4291 => x"38",
          4292 => x"38",
          4293 => x"fe",
          4294 => x"fe",
          4295 => x"96",
          4296 => x"ff",
          4297 => x"3f",
          4298 => x"08",
          4299 => x"80",
          4300 => x"38",
          4301 => x"0c",
          4302 => x"08",
          4303 => x"ff",
          4304 => x"81",
          4305 => x"55",
          4306 => x"0d",
          4307 => x"8c",
          4308 => x"58",
          4309 => x"b8",
          4310 => x"f5",
          4311 => x"ff",
          4312 => x"bb",
          4313 => x"56",
          4314 => x"55",
          4315 => x"7c",
          4316 => x"80",
          4317 => x"06",
          4318 => x"19",
          4319 => x"df",
          4320 => x"80",
          4321 => x"0b",
          4322 => x"27",
          4323 => x"0c",
          4324 => x"53",
          4325 => x"73",
          4326 => x"83",
          4327 => x"0c",
          4328 => x"8a",
          4329 => x"84",
          4330 => x"08",
          4331 => x"8a",
          4332 => x"73",
          4333 => x"53",
          4334 => x"59",
          4335 => x"22",
          4336 => x"5a",
          4337 => x"39",
          4338 => x"84",
          4339 => x"08",
          4340 => x"bb",
          4341 => x"17",
          4342 => x"27",
          4343 => x"73",
          4344 => x"81",
          4345 => x"0d",
          4346 => x"90",
          4347 => x"f0",
          4348 => x"0b",
          4349 => x"84",
          4350 => x"83",
          4351 => x"15",
          4352 => x"38",
          4353 => x"55",
          4354 => x"98",
          4355 => x"1b",
          4356 => x"75",
          4357 => x"04",
          4358 => x"ff",
          4359 => x"da",
          4360 => x"3f",
          4361 => x"81",
          4362 => x"38",
          4363 => x"2e",
          4364 => x"84",
          4365 => x"2e",
          4366 => x"76",
          4367 => x"08",
          4368 => x"80",
          4369 => x"bb",
          4370 => x"81",
          4371 => x"ff",
          4372 => x"1a",
          4373 => x"fe",
          4374 => x"56",
          4375 => x"8a",
          4376 => x"08",
          4377 => x"b8",
          4378 => x"80",
          4379 => x"15",
          4380 => x"19",
          4381 => x"38",
          4382 => x"81",
          4383 => x"bb",
          4384 => x"56",
          4385 => x"0b",
          4386 => x"04",
          4387 => x"19",
          4388 => x"e4",
          4389 => x"f3",
          4390 => x"34",
          4391 => x"55",
          4392 => x"38",
          4393 => x"09",
          4394 => x"b4",
          4395 => x"75",
          4396 => x"3f",
          4397 => x"74",
          4398 => x"2e",
          4399 => x"18",
          4400 => x"05",
          4401 => x"fd",
          4402 => x"29",
          4403 => x"5c",
          4404 => x"84",
          4405 => x"0d",
          4406 => x"5a",
          4407 => x"58",
          4408 => x"38",
          4409 => x"b4",
          4410 => x"83",
          4411 => x"2e",
          4412 => x"54",
          4413 => x"33",
          4414 => x"08",
          4415 => x"57",
          4416 => x"82",
          4417 => x"58",
          4418 => x"8b",
          4419 => x"06",
          4420 => x"81",
          4421 => x"70",
          4422 => x"07",
          4423 => x"38",
          4424 => x"88",
          4425 => x"81",
          4426 => x"7b",
          4427 => x"08",
          4428 => x"38",
          4429 => x"38",
          4430 => x"0d",
          4431 => x"7e",
          4432 => x"3f",
          4433 => x"2e",
          4434 => x"bb",
          4435 => x"08",
          4436 => x"08",
          4437 => x"fe",
          4438 => x"82",
          4439 => x"81",
          4440 => x"05",
          4441 => x"e0",
          4442 => x"79",
          4443 => x"38",
          4444 => x"80",
          4445 => x"81",
          4446 => x"ac",
          4447 => x"2e",
          4448 => x"fe",
          4449 => x"09",
          4450 => x"84",
          4451 => x"84",
          4452 => x"77",
          4453 => x"57",
          4454 => x"38",
          4455 => x"1a",
          4456 => x"41",
          4457 => x"81",
          4458 => x"5a",
          4459 => x"17",
          4460 => x"33",
          4461 => x"7a",
          4462 => x"fe",
          4463 => x"05",
          4464 => x"1a",
          4465 => x"cc",
          4466 => x"06",
          4467 => x"79",
          4468 => x"10",
          4469 => x"1d",
          4470 => x"9d",
          4471 => x"38",
          4472 => x"a8",
          4473 => x"2a",
          4474 => x"81",
          4475 => x"81",
          4476 => x"76",
          4477 => x"38",
          4478 => x"bb",
          4479 => x"3d",
          4480 => x"52",
          4481 => x"84",
          4482 => x"80",
          4483 => x"0b",
          4484 => x"1c",
          4485 => x"76",
          4486 => x"78",
          4487 => x"06",
          4488 => x"b8",
          4489 => x"e0",
          4490 => x"85",
          4491 => x"1c",
          4492 => x"9c",
          4493 => x"80",
          4494 => x"bf",
          4495 => x"77",
          4496 => x"80",
          4497 => x"55",
          4498 => x"80",
          4499 => x"38",
          4500 => x"8b",
          4501 => x"29",
          4502 => x"57",
          4503 => x"19",
          4504 => x"7f",
          4505 => x"81",
          4506 => x"a0",
          4507 => x"5a",
          4508 => x"71",
          4509 => x"40",
          4510 => x"80",
          4511 => x"0b",
          4512 => x"f5",
          4513 => x"84",
          4514 => x"38",
          4515 => x"0d",
          4516 => x"7d",
          4517 => x"3f",
          4518 => x"2e",
          4519 => x"bb",
          4520 => x"08",
          4521 => x"08",
          4522 => x"fd",
          4523 => x"82",
          4524 => x"81",
          4525 => x"05",
          4526 => x"db",
          4527 => x"77",
          4528 => x"70",
          4529 => x"fe",
          4530 => x"5a",
          4531 => x"33",
          4532 => x"08",
          4533 => x"76",
          4534 => x"74",
          4535 => x"3f",
          4536 => x"84",
          4537 => x"c8",
          4538 => x"81",
          4539 => x"fe",
          4540 => x"77",
          4541 => x"1b",
          4542 => x"71",
          4543 => x"ff",
          4544 => x"8d",
          4545 => x"59",
          4546 => x"05",
          4547 => x"2b",
          4548 => x"80",
          4549 => x"84",
          4550 => x"84",
          4551 => x"70",
          4552 => x"81",
          4553 => x"08",
          4554 => x"76",
          4555 => x"ff",
          4556 => x"81",
          4557 => x"38",
          4558 => x"60",
          4559 => x"b4",
          4560 => x"5e",
          4561 => x"bb",
          4562 => x"83",
          4563 => x"ff",
          4564 => x"68",
          4565 => x"a0",
          4566 => x"74",
          4567 => x"70",
          4568 => x"8e",
          4569 => x"22",
          4570 => x"3d",
          4571 => x"58",
          4572 => x"33",
          4573 => x"15",
          4574 => x"05",
          4575 => x"80",
          4576 => x"ab",
          4577 => x"5b",
          4578 => x"7a",
          4579 => x"05",
          4580 => x"34",
          4581 => x"7b",
          4582 => x"56",
          4583 => x"82",
          4584 => x"06",
          4585 => x"83",
          4586 => x"06",
          4587 => x"87",
          4588 => x"ff",
          4589 => x"78",
          4590 => x"84",
          4591 => x"b0",
          4592 => x"84",
          4593 => x"ff",
          4594 => x"59",
          4595 => x"80",
          4596 => x"80",
          4597 => x"74",
          4598 => x"75",
          4599 => x"70",
          4600 => x"81",
          4601 => x"55",
          4602 => x"78",
          4603 => x"57",
          4604 => x"27",
          4605 => x"3f",
          4606 => x"1b",
          4607 => x"38",
          4608 => x"e7",
          4609 => x"bb",
          4610 => x"82",
          4611 => x"ab",
          4612 => x"80",
          4613 => x"2a",
          4614 => x"2e",
          4615 => x"fe",
          4616 => x"1b",
          4617 => x"3f",
          4618 => x"84",
          4619 => x"08",
          4620 => x"56",
          4621 => x"85",
          4622 => x"77",
          4623 => x"81",
          4624 => x"18",
          4625 => x"84",
          4626 => x"81",
          4627 => x"76",
          4628 => x"56",
          4629 => x"38",
          4630 => x"56",
          4631 => x"81",
          4632 => x"38",
          4633 => x"84",
          4634 => x"08",
          4635 => x"75",
          4636 => x"75",
          4637 => x"81",
          4638 => x"1c",
          4639 => x"33",
          4640 => x"81",
          4641 => x"1c",
          4642 => x"84",
          4643 => x"81",
          4644 => x"75",
          4645 => x"08",
          4646 => x"58",
          4647 => x"8b",
          4648 => x"55",
          4649 => x"70",
          4650 => x"74",
          4651 => x"33",
          4652 => x"34",
          4653 => x"75",
          4654 => x"04",
          4655 => x"07",
          4656 => x"74",
          4657 => x"3f",
          4658 => x"84",
          4659 => x"bd",
          4660 => x"7c",
          4661 => x"3f",
          4662 => x"81",
          4663 => x"08",
          4664 => x"19",
          4665 => x"27",
          4666 => x"82",
          4667 => x"08",
          4668 => x"90",
          4669 => x"51",
          4670 => x"58",
          4671 => x"79",
          4672 => x"57",
          4673 => x"05",
          4674 => x"76",
          4675 => x"59",
          4676 => x"ff",
          4677 => x"08",
          4678 => x"2e",
          4679 => x"76",
          4680 => x"81",
          4681 => x"1c",
          4682 => x"84",
          4683 => x"81",
          4684 => x"75",
          4685 => x"1f",
          4686 => x"5f",
          4687 => x"1c",
          4688 => x"1c",
          4689 => x"29",
          4690 => x"76",
          4691 => x"10",
          4692 => x"56",
          4693 => x"55",
          4694 => x"76",
          4695 => x"85",
          4696 => x"58",
          4697 => x"ff",
          4698 => x"1f",
          4699 => x"81",
          4700 => x"83",
          4701 => x"e1",
          4702 => x"bb",
          4703 => x"05",
          4704 => x"39",
          4705 => x"1c",
          4706 => x"d0",
          4707 => x"08",
          4708 => x"83",
          4709 => x"08",
          4710 => x"60",
          4711 => x"82",
          4712 => x"81",
          4713 => x"1c",
          4714 => x"52",
          4715 => x"77",
          4716 => x"08",
          4717 => x"e5",
          4718 => x"fb",
          4719 => x"80",
          4720 => x"7c",
          4721 => x"81",
          4722 => x"81",
          4723 => x"bb",
          4724 => x"bc",
          4725 => x"34",
          4726 => x"55",
          4727 => x"82",
          4728 => x"38",
          4729 => x"39",
          4730 => x"2e",
          4731 => x"1a",
          4732 => x"56",
          4733 => x"fd",
          4734 => x"1d",
          4735 => x"33",
          4736 => x"81",
          4737 => x"05",
          4738 => x"ce",
          4739 => x"0d",
          4740 => x"80",
          4741 => x"80",
          4742 => x"ff",
          4743 => x"60",
          4744 => x"5b",
          4745 => x"77",
          4746 => x"5b",
          4747 => x"d0",
          4748 => x"58",
          4749 => x"38",
          4750 => x"5d",
          4751 => x"30",
          4752 => x"5a",
          4753 => x"80",
          4754 => x"1f",
          4755 => x"70",
          4756 => x"a0",
          4757 => x"bc",
          4758 => x"72",
          4759 => x"8b",
          4760 => x"38",
          4761 => x"81",
          4762 => x"59",
          4763 => x"ff",
          4764 => x"80",
          4765 => x"53",
          4766 => x"bf",
          4767 => x"17",
          4768 => x"34",
          4769 => x"53",
          4770 => x"9c",
          4771 => x"1e",
          4772 => x"11",
          4773 => x"71",
          4774 => x"72",
          4775 => x"64",
          4776 => x"33",
          4777 => x"40",
          4778 => x"23",
          4779 => x"88",
          4780 => x"23",
          4781 => x"fe",
          4782 => x"ff",
          4783 => x"52",
          4784 => x"90",
          4785 => x"ff",
          4786 => x"ad",
          4787 => x"74",
          4788 => x"97",
          4789 => x"0b",
          4790 => x"75",
          4791 => x"fd",
          4792 => x"76",
          4793 => x"80",
          4794 => x"f9",
          4795 => x"58",
          4796 => x"cd",
          4797 => x"57",
          4798 => x"7c",
          4799 => x"14",
          4800 => x"99",
          4801 => x"11",
          4802 => x"38",
          4803 => x"5e",
          4804 => x"70",
          4805 => x"78",
          4806 => x"81",
          4807 => x"5e",
          4808 => x"38",
          4809 => x"cc",
          4810 => x"70",
          4811 => x"fc",
          4812 => x"08",
          4813 => x"33",
          4814 => x"38",
          4815 => x"df",
          4816 => x"98",
          4817 => x"96",
          4818 => x"75",
          4819 => x"16",
          4820 => x"81",
          4821 => x"df",
          4822 => x"81",
          4823 => x"8b",
          4824 => x"23",
          4825 => x"06",
          4826 => x"27",
          4827 => x"55",
          4828 => x"2e",
          4829 => x"b2",
          4830 => x"a0",
          4831 => x"56",
          4832 => x"75",
          4833 => x"70",
          4834 => x"ee",
          4835 => x"81",
          4836 => x"fd",
          4837 => x"23",
          4838 => x"52",
          4839 => x"fe",
          4840 => x"80",
          4841 => x"73",
          4842 => x"2e",
          4843 => x"80",
          4844 => x"dd",
          4845 => x"70",
          4846 => x"72",
          4847 => x"33",
          4848 => x"74",
          4849 => x"83",
          4850 => x"3f",
          4851 => x"06",
          4852 => x"73",
          4853 => x"04",
          4854 => x"06",
          4855 => x"38",
          4856 => x"34",
          4857 => x"84",
          4858 => x"93",
          4859 => x"32",
          4860 => x"41",
          4861 => x"38",
          4862 => x"55",
          4863 => x"72",
          4864 => x"25",
          4865 => x"38",
          4866 => x"2b",
          4867 => x"76",
          4868 => x"59",
          4869 => x"78",
          4870 => x"32",
          4871 => x"56",
          4872 => x"38",
          4873 => x"dd",
          4874 => x"76",
          4875 => x"80",
          4876 => x"72",
          4877 => x"82",
          4878 => x"53",
          4879 => x"80",
          4880 => x"70",
          4881 => x"38",
          4882 => x"17",
          4883 => x"14",
          4884 => x"09",
          4885 => x"1d",
          4886 => x"56",
          4887 => x"72",
          4888 => x"22",
          4889 => x"80",
          4890 => x"83",
          4891 => x"70",
          4892 => x"2e",
          4893 => x"72",
          4894 => x"59",
          4895 => x"07",
          4896 => x"54",
          4897 => x"7c",
          4898 => x"2e",
          4899 => x"77",
          4900 => x"8b",
          4901 => x"18",
          4902 => x"81",
          4903 => x"38",
          4904 => x"2e",
          4905 => x"e3",
          4906 => x"2e",
          4907 => x"74",
          4908 => x"2a",
          4909 => x"81",
          4910 => x"79",
          4911 => x"06",
          4912 => x"88",
          4913 => x"51",
          4914 => x"ab",
          4915 => x"08",
          4916 => x"84",
          4917 => x"f7",
          4918 => x"79",
          4919 => x"2a",
          4920 => x"7b",
          4921 => x"16",
          4922 => x"81",
          4923 => x"40",
          4924 => x"38",
          4925 => x"83",
          4926 => x"22",
          4927 => x"fc",
          4928 => x"2e",
          4929 => x"10",
          4930 => x"a0",
          4931 => x"26",
          4932 => x"81",
          4933 => x"73",
          4934 => x"77",
          4935 => x"3f",
          4936 => x"56",
          4937 => x"38",
          4938 => x"fa",
          4939 => x"2a",
          4940 => x"83",
          4941 => x"06",
          4942 => x"d2",
          4943 => x"33",
          4944 => x"82",
          4945 => x"08",
          4946 => x"22",
          4947 => x"76",
          4948 => x"ab",
          4949 => x"5a",
          4950 => x"fc",
          4951 => x"8c",
          4952 => x"79",
          4953 => x"0b",
          4954 => x"81",
          4955 => x"80",
          4956 => x"bb",
          4957 => x"80",
          4958 => x"27",
          4959 => x"7b",
          4960 => x"7d",
          4961 => x"39",
          4962 => x"74",
          4963 => x"84",
          4964 => x"2a",
          4965 => x"c4",
          4966 => x"94",
          4967 => x"26",
          4968 => x"85",
          4969 => x"ac",
          4970 => x"59",
          4971 => x"75",
          4972 => x"70",
          4973 => x"ee",
          4974 => x"80",
          4975 => x"99",
          4976 => x"81",
          4977 => x"59",
          4978 => x"07",
          4979 => x"83",
          4980 => x"7b",
          4981 => x"81",
          4982 => x"39",
          4983 => x"ac",
          4984 => x"78",
          4985 => x"7a",
          4986 => x"5b",
          4987 => x"d2",
          4988 => x"15",
          4989 => x"07",
          4990 => x"fd",
          4991 => x"88",
          4992 => x"1b",
          4993 => x"79",
          4994 => x"79",
          4995 => x"76",
          4996 => x"a3",
          4997 => x"81",
          4998 => x"0b",
          4999 => x"04",
          5000 => x"05",
          5001 => x"80",
          5002 => x"5b",
          5003 => x"79",
          5004 => x"26",
          5005 => x"38",
          5006 => x"c7",
          5007 => x"76",
          5008 => x"84",
          5009 => x"8c",
          5010 => x"76",
          5011 => x"33",
          5012 => x"81",
          5013 => x"84",
          5014 => x"81",
          5015 => x"96",
          5016 => x"84",
          5017 => x"81",
          5018 => x"a4",
          5019 => x"06",
          5020 => x"7f",
          5021 => x"38",
          5022 => x"58",
          5023 => x"83",
          5024 => x"7a",
          5025 => x"b8",
          5026 => x"58",
          5027 => x"08",
          5028 => x"59",
          5029 => x"99",
          5030 => x"18",
          5031 => x"83",
          5032 => x"a5",
          5033 => x"ba",
          5034 => x"38",
          5035 => x"38",
          5036 => x"38",
          5037 => x"33",
          5038 => x"84",
          5039 => x"38",
          5040 => x"33",
          5041 => x"a4",
          5042 => x"82",
          5043 => x"2b",
          5044 => x"88",
          5045 => x"45",
          5046 => x"0c",
          5047 => x"80",
          5048 => x"ff",
          5049 => x"81",
          5050 => x"06",
          5051 => x"5a",
          5052 => x"59",
          5053 => x"18",
          5054 => x"80",
          5055 => x"71",
          5056 => x"18",
          5057 => x"8d",
          5058 => x"17",
          5059 => x"2b",
          5060 => x"d8",
          5061 => x"71",
          5062 => x"14",
          5063 => x"33",
          5064 => x"42",
          5065 => x"18",
          5066 => x"8d",
          5067 => x"7d",
          5068 => x"75",
          5069 => x"7a",
          5070 => x"bb",
          5071 => x"80",
          5072 => x"08",
          5073 => x"38",
          5074 => x"83",
          5075 => x"85",
          5076 => x"9c",
          5077 => x"1d",
          5078 => x"1a",
          5079 => x"87",
          5080 => x"7b",
          5081 => x"ac",
          5082 => x"2e",
          5083 => x"2a",
          5084 => x"ff",
          5085 => x"a0",
          5086 => x"94",
          5087 => x"ff",
          5088 => x"2e",
          5089 => x"e2",
          5090 => x"e2",
          5091 => x"e2",
          5092 => x"98",
          5093 => x"84",
          5094 => x"84",
          5095 => x"76",
          5096 => x"57",
          5097 => x"82",
          5098 => x"5d",
          5099 => x"80",
          5100 => x"5c",
          5101 => x"81",
          5102 => x"5b",
          5103 => x"77",
          5104 => x"81",
          5105 => x"58",
          5106 => x"70",
          5107 => x"70",
          5108 => x"09",
          5109 => x"38",
          5110 => x"07",
          5111 => x"7a",
          5112 => x"84",
          5113 => x"98",
          5114 => x"80",
          5115 => x"81",
          5116 => x"38",
          5117 => x"33",
          5118 => x"81",
          5119 => x"eb",
          5120 => x"07",
          5121 => x"75",
          5122 => x"3d",
          5123 => x"16",
          5124 => x"a5",
          5125 => x"17",
          5126 => x"07",
          5127 => x"88",
          5128 => x"52",
          5129 => x"70",
          5130 => x"17",
          5131 => x"38",
          5132 => x"70",
          5133 => x"71",
          5134 => x"1c",
          5135 => x"08",
          5136 => x"fb",
          5137 => x"0b",
          5138 => x"7a",
          5139 => x"53",
          5140 => x"ff",
          5141 => x"76",
          5142 => x"74",
          5143 => x"38",
          5144 => x"2b",
          5145 => x"d4",
          5146 => x"80",
          5147 => x"81",
          5148 => x"eb",
          5149 => x"07",
          5150 => x"81",
          5151 => x"81",
          5152 => x"f9",
          5153 => x"09",
          5154 => x"76",
          5155 => x"f8",
          5156 => x"5a",
          5157 => x"a8",
          5158 => x"e6",
          5159 => x"05",
          5160 => x"33",
          5161 => x"56",
          5162 => x"75",
          5163 => x"8a",
          5164 => x"7b",
          5165 => x"81",
          5166 => x"1b",
          5167 => x"85",
          5168 => x"82",
          5169 => x"fa",
          5170 => x"97",
          5171 => x"2e",
          5172 => x"18",
          5173 => x"b7",
          5174 => x"97",
          5175 => x"18",
          5176 => x"70",
          5177 => x"05",
          5178 => x"5b",
          5179 => x"d1",
          5180 => x"0b",
          5181 => x"5a",
          5182 => x"7a",
          5183 => x"31",
          5184 => x"80",
          5185 => x"e1",
          5186 => x"59",
          5187 => x"39",
          5188 => x"33",
          5189 => x"81",
          5190 => x"81",
          5191 => x"78",
          5192 => x"7a",
          5193 => x"38",
          5194 => x"81",
          5195 => x"84",
          5196 => x"ff",
          5197 => x"79",
          5198 => x"84",
          5199 => x"71",
          5200 => x"d4",
          5201 => x"38",
          5202 => x"33",
          5203 => x"81",
          5204 => x"75",
          5205 => x"42",
          5206 => x"d2",
          5207 => x"84",
          5208 => x"33",
          5209 => x"81",
          5210 => x"75",
          5211 => x"5c",
          5212 => x"f2",
          5213 => x"84",
          5214 => x"33",
          5215 => x"81",
          5216 => x"75",
          5217 => x"84",
          5218 => x"33",
          5219 => x"81",
          5220 => x"75",
          5221 => x"59",
          5222 => x"5b",
          5223 => x"dc",
          5224 => x"dc",
          5225 => x"e4",
          5226 => x"18",
          5227 => x"f8",
          5228 => x"f2",
          5229 => x"53",
          5230 => x"52",
          5231 => x"84",
          5232 => x"a4",
          5233 => x"34",
          5234 => x"40",
          5235 => x"82",
          5236 => x"8d",
          5237 => x"a0",
          5238 => x"91",
          5239 => x"e6",
          5240 => x"80",
          5241 => x"71",
          5242 => x"7d",
          5243 => x"61",
          5244 => x"11",
          5245 => x"71",
          5246 => x"72",
          5247 => x"ac",
          5248 => x"43",
          5249 => x"75",
          5250 => x"82",
          5251 => x"f2",
          5252 => x"83",
          5253 => x"f5",
          5254 => x"b4",
          5255 => x"78",
          5256 => x"e7",
          5257 => x"02",
          5258 => x"93",
          5259 => x"40",
          5260 => x"70",
          5261 => x"55",
          5262 => x"73",
          5263 => x"38",
          5264 => x"24",
          5265 => x"e2",
          5266 => x"80",
          5267 => x"54",
          5268 => x"34",
          5269 => x"7c",
          5270 => x"3d",
          5271 => x"3f",
          5272 => x"bb",
          5273 => x"0b",
          5274 => x"04",
          5275 => x"06",
          5276 => x"38",
          5277 => x"05",
          5278 => x"38",
          5279 => x"5f",
          5280 => x"70",
          5281 => x"05",
          5282 => x"55",
          5283 => x"70",
          5284 => x"16",
          5285 => x"16",
          5286 => x"30",
          5287 => x"2e",
          5288 => x"be",
          5289 => x"72",
          5290 => x"54",
          5291 => x"84",
          5292 => x"99",
          5293 => x"83",
          5294 => x"54",
          5295 => x"02",
          5296 => x"5a",
          5297 => x"74",
          5298 => x"05",
          5299 => x"ed",
          5300 => x"84",
          5301 => x"80",
          5302 => x"84",
          5303 => x"6d",
          5304 => x"9a",
          5305 => x"bb",
          5306 => x"78",
          5307 => x"ca",
          5308 => x"76",
          5309 => x"07",
          5310 => x"2a",
          5311 => x"d1",
          5312 => x"33",
          5313 => x"42",
          5314 => x"86",
          5315 => x"80",
          5316 => x"17",
          5317 => x"66",
          5318 => x"67",
          5319 => x"80",
          5320 => x"7c",
          5321 => x"80",
          5322 => x"19",
          5323 => x"0b",
          5324 => x"83",
          5325 => x"38",
          5326 => x"59",
          5327 => x"38",
          5328 => x"38",
          5329 => x"39",
          5330 => x"2b",
          5331 => x"38",
          5332 => x"fe",
          5333 => x"80",
          5334 => x"06",
          5335 => x"81",
          5336 => x"89",
          5337 => x"95",
          5338 => x"75",
          5339 => x"07",
          5340 => x"0c",
          5341 => x"33",
          5342 => x"73",
          5343 => x"83",
          5344 => x"0c",
          5345 => x"33",
          5346 => x"81",
          5347 => x"75",
          5348 => x"43",
          5349 => x"56",
          5350 => x"90",
          5351 => x"80",
          5352 => x"1b",
          5353 => x"57",
          5354 => x"34",
          5355 => x"85",
          5356 => x"fc",
          5357 => x"80",
          5358 => x"0c",
          5359 => x"1c",
          5360 => x"30",
          5361 => x"78",
          5362 => x"76",
          5363 => x"db",
          5364 => x"bb",
          5365 => x"bb",
          5366 => x"57",
          5367 => x"38",
          5368 => x"80",
          5369 => x"95",
          5370 => x"74",
          5371 => x"80",
          5372 => x"80",
          5373 => x"80",
          5374 => x"7a",
          5375 => x"16",
          5376 => x"71",
          5377 => x"0c",
          5378 => x"33",
          5379 => x"81",
          5380 => x"75",
          5381 => x"45",
          5382 => x"58",
          5383 => x"23",
          5384 => x"1b",
          5385 => x"0b",
          5386 => x"80",
          5387 => x"51",
          5388 => x"79",
          5389 => x"38",
          5390 => x"ff",
          5391 => x"5d",
          5392 => x"cb",
          5393 => x"fb",
          5394 => x"2e",
          5395 => x"75",
          5396 => x"84",
          5397 => x"fe",
          5398 => x"76",
          5399 => x"17",
          5400 => x"74",
          5401 => x"26",
          5402 => x"5f",
          5403 => x"2e",
          5404 => x"7d",
          5405 => x"81",
          5406 => x"16",
          5407 => x"bb",
          5408 => x"57",
          5409 => x"56",
          5410 => x"7b",
          5411 => x"0c",
          5412 => x"34",
          5413 => x"39",
          5414 => x"98",
          5415 => x"5d",
          5416 => x"80",
          5417 => x"17",
          5418 => x"66",
          5419 => x"67",
          5420 => x"80",
          5421 => x"7c",
          5422 => x"38",
          5423 => x"76",
          5424 => x"59",
          5425 => x"fe",
          5426 => x"59",
          5427 => x"8a",
          5428 => x"08",
          5429 => x"d8",
          5430 => x"1c",
          5431 => x"52",
          5432 => x"3f",
          5433 => x"e2",
          5434 => x"da",
          5435 => x"b8",
          5436 => x"58",
          5437 => x"08",
          5438 => x"38",
          5439 => x"b4",
          5440 => x"bb",
          5441 => x"08",
          5442 => x"55",
          5443 => x"cf",
          5444 => x"17",
          5445 => x"33",
          5446 => x"fd",
          5447 => x"80",
          5448 => x"fd",
          5449 => x"65",
          5450 => x"0c",
          5451 => x"78",
          5452 => x"75",
          5453 => x"86",
          5454 => x"7a",
          5455 => x"74",
          5456 => x"91",
          5457 => x"90",
          5458 => x"76",
          5459 => x"08",
          5460 => x"79",
          5461 => x"2e",
          5462 => x"5c",
          5463 => x"22",
          5464 => x"58",
          5465 => x"88",
          5466 => x"c3",
          5467 => x"74",
          5468 => x"08",
          5469 => x"5c",
          5470 => x"8a",
          5471 => x"08",
          5472 => x"93",
          5473 => x"57",
          5474 => x"1c",
          5475 => x"7c",
          5476 => x"52",
          5477 => x"3f",
          5478 => x"90",
          5479 => x"80",
          5480 => x"2b",
          5481 => x"7f",
          5482 => x"70",
          5483 => x"fe",
          5484 => x"84",
          5485 => x"bb",
          5486 => x"5a",
          5487 => x"75",
          5488 => x"33",
          5489 => x"5b",
          5490 => x"75",
          5491 => x"ff",
          5492 => x"81",
          5493 => x"06",
          5494 => x"81",
          5495 => x"33",
          5496 => x"84",
          5497 => x"0c",
          5498 => x"06",
          5499 => x"77",
          5500 => x"7a",
          5501 => x"80",
          5502 => x"05",
          5503 => x"34",
          5504 => x"c1",
          5505 => x"78",
          5506 => x"56",
          5507 => x"19",
          5508 => x"3f",
          5509 => x"39",
          5510 => x"3f",
          5511 => x"74",
          5512 => x"57",
          5513 => x"31",
          5514 => x"84",
          5515 => x"58",
          5516 => x"33",
          5517 => x"15",
          5518 => x"75",
          5519 => x"81",
          5520 => x"da",
          5521 => x"1a",
          5522 => x"90",
          5523 => x"34",
          5524 => x"3d",
          5525 => x"66",
          5526 => x"0c",
          5527 => x"78",
          5528 => x"75",
          5529 => x"86",
          5530 => x"79",
          5531 => x"74",
          5532 => x"91",
          5533 => x"90",
          5534 => x"58",
          5535 => x"a9",
          5536 => x"57",
          5537 => x"5b",
          5538 => x"83",
          5539 => x"7f",
          5540 => x"2a",
          5541 => x"82",
          5542 => x"80",
          5543 => x"83",
          5544 => x"38",
          5545 => x"85",
          5546 => x"90",
          5547 => x"80",
          5548 => x"08",
          5549 => x"5d",
          5550 => x"8a",
          5551 => x"08",
          5552 => x"a6",
          5553 => x"5c",
          5554 => x"1d",
          5555 => x"7d",
          5556 => x"52",
          5557 => x"3f",
          5558 => x"9c",
          5559 => x"27",
          5560 => x"77",
          5561 => x"75",
          5562 => x"81",
          5563 => x"ef",
          5564 => x"5d",
          5565 => x"58",
          5566 => x"0c",
          5567 => x"71",
          5568 => x"5a",
          5569 => x"38",
          5570 => x"fd",
          5571 => x"80",
          5572 => x"80",
          5573 => x"3d",
          5574 => x"91",
          5575 => x"2e",
          5576 => x"8c",
          5577 => x"7b",
          5578 => x"51",
          5579 => x"08",
          5580 => x"7b",
          5581 => x"84",
          5582 => x"27",
          5583 => x"a8",
          5584 => x"2e",
          5585 => x"33",
          5586 => x"16",
          5587 => x"ff",
          5588 => x"fe",
          5589 => x"51",
          5590 => x"08",
          5591 => x"38",
          5592 => x"76",
          5593 => x"84",
          5594 => x"08",
          5595 => x"9c",
          5596 => x"18",
          5597 => x"bb",
          5598 => x"80",
          5599 => x"7f",
          5600 => x"51",
          5601 => x"08",
          5602 => x"74",
          5603 => x"81",
          5604 => x"bb",
          5605 => x"0b",
          5606 => x"84",
          5607 => x"0d",
          5608 => x"9f",
          5609 => x"97",
          5610 => x"8f",
          5611 => x"5a",
          5612 => x"80",
          5613 => x"ee",
          5614 => x"81",
          5615 => x"de",
          5616 => x"24",
          5617 => x"58",
          5618 => x"38",
          5619 => x"5c",
          5620 => x"81",
          5621 => x"16",
          5622 => x"f8",
          5623 => x"85",
          5624 => x"17",
          5625 => x"a4",
          5626 => x"56",
          5627 => x"88",
          5628 => x"5d",
          5629 => x"88",
          5630 => x"17",
          5631 => x"74",
          5632 => x"08",
          5633 => x"5b",
          5634 => x"56",
          5635 => x"59",
          5636 => x"80",
          5637 => x"18",
          5638 => x"80",
          5639 => x"18",
          5640 => x"34",
          5641 => x"bb",
          5642 => x"06",
          5643 => x"55",
          5644 => x"0d",
          5645 => x"b8",
          5646 => x"5b",
          5647 => x"bb",
          5648 => x"fe",
          5649 => x"17",
          5650 => x"31",
          5651 => x"a0",
          5652 => x"16",
          5653 => x"06",
          5654 => x"08",
          5655 => x"81",
          5656 => x"79",
          5657 => x"55",
          5658 => x"56",
          5659 => x"55",
          5660 => x"7a",
          5661 => x"75",
          5662 => x"78",
          5663 => x"0b",
          5664 => x"34",
          5665 => x"0b",
          5666 => x"34",
          5667 => x"7b",
          5668 => x"84",
          5669 => x"5b",
          5670 => x"39",
          5671 => x"3f",
          5672 => x"74",
          5673 => x"57",
          5674 => x"08",
          5675 => x"33",
          5676 => x"55",
          5677 => x"90",
          5678 => x"90",
          5679 => x"56",
          5680 => x"06",
          5681 => x"3d",
          5682 => x"3f",
          5683 => x"84",
          5684 => x"2e",
          5685 => x"2e",
          5686 => x"2e",
          5687 => x"22",
          5688 => x"80",
          5689 => x"38",
          5690 => x"0c",
          5691 => x"51",
          5692 => x"08",
          5693 => x"75",
          5694 => x"0d",
          5695 => x"80",
          5696 => x"57",
          5697 => x"ba",
          5698 => x"ba",
          5699 => x"51",
          5700 => x"e2",
          5701 => x"0c",
          5702 => x"bb",
          5703 => x"33",
          5704 => x"53",
          5705 => x"19",
          5706 => x"54",
          5707 => x"0b",
          5708 => x"79",
          5709 => x"33",
          5710 => x"9f",
          5711 => x"89",
          5712 => x"53",
          5713 => x"26",
          5714 => x"06",
          5715 => x"55",
          5716 => x"85",
          5717 => x"32",
          5718 => x"76",
          5719 => x"92",
          5720 => x"83",
          5721 => x"fe",
          5722 => x"77",
          5723 => x"3d",
          5724 => x"52",
          5725 => x"bb",
          5726 => x"80",
          5727 => x"0c",
          5728 => x"52",
          5729 => x"3f",
          5730 => x"84",
          5731 => x"05",
          5732 => x"77",
          5733 => x"33",
          5734 => x"75",
          5735 => x"11",
          5736 => x"07",
          5737 => x"79",
          5738 => x"0c",
          5739 => x"0d",
          5740 => x"09",
          5741 => x"84",
          5742 => x"95",
          5743 => x"2b",
          5744 => x"1b",
          5745 => x"98",
          5746 => x"0c",
          5747 => x"0d",
          5748 => x"08",
          5749 => x"80",
          5750 => x"e5",
          5751 => x"84",
          5752 => x"c8",
          5753 => x"61",
          5754 => x"58",
          5755 => x"80",
          5756 => x"98",
          5757 => x"ff",
          5758 => x"59",
          5759 => x"60",
          5760 => x"16",
          5761 => x"84",
          5762 => x"83",
          5763 => x"16",
          5764 => x"88",
          5765 => x"85",
          5766 => x"17",
          5767 => x"3d",
          5768 => x"71",
          5769 => x"40",
          5770 => x"da",
          5771 => x"52",
          5772 => x"bb",
          5773 => x"82",
          5774 => x"aa",
          5775 => x"84",
          5776 => x"3d",
          5777 => x"71",
          5778 => x"58",
          5779 => x"fd",
          5780 => x"bb",
          5781 => x"a1",
          5782 => x"bb",
          5783 => x"78",
          5784 => x"c8",
          5785 => x"52",
          5786 => x"7f",
          5787 => x"2e",
          5788 => x"81",
          5789 => x"f5",
          5790 => x"81",
          5791 => x"7e",
          5792 => x"e6",
          5793 => x"59",
          5794 => x"76",
          5795 => x"08",
          5796 => x"da",
          5797 => x"77",
          5798 => x"84",
          5799 => x"e6",
          5800 => x"59",
          5801 => x"38",
          5802 => x"5f",
          5803 => x"7a",
          5804 => x"7a",
          5805 => x"33",
          5806 => x"17",
          5807 => x"7c",
          5808 => x"2e",
          5809 => x"59",
          5810 => x"0c",
          5811 => x"33",
          5812 => x"90",
          5813 => x"fd",
          5814 => x"33",
          5815 => x"79",
          5816 => x"80",
          5817 => x"84",
          5818 => x"08",
          5819 => x"39",
          5820 => x"16",
          5821 => x"ff",
          5822 => x"84",
          5823 => x"08",
          5824 => x"17",
          5825 => x"55",
          5826 => x"38",
          5827 => x"09",
          5828 => x"b4",
          5829 => x"7d",
          5830 => x"f7",
          5831 => x"18",
          5832 => x"af",
          5833 => x"33",
          5834 => x"70",
          5835 => x"5a",
          5836 => x"e8",
          5837 => x"08",
          5838 => x"7c",
          5839 => x"27",
          5840 => x"18",
          5841 => x"70",
          5842 => x"d4",
          5843 => x"7c",
          5844 => x"e4",
          5845 => x"7f",
          5846 => x"9f",
          5847 => x"97",
          5848 => x"8f",
          5849 => x"5b",
          5850 => x"80",
          5851 => x"fb",
          5852 => x"f3",
          5853 => x"26",
          5854 => x"80",
          5855 => x"7b",
          5856 => x"5c",
          5857 => x"77",
          5858 => x"3f",
          5859 => x"54",
          5860 => x"3f",
          5861 => x"da",
          5862 => x"19",
          5863 => x"58",
          5864 => x"38",
          5865 => x"78",
          5866 => x"0c",
          5867 => x"06",
          5868 => x"cc",
          5869 => x"b2",
          5870 => x"bb",
          5871 => x"ff",
          5872 => x"83",
          5873 => x"08",
          5874 => x"0c",
          5875 => x"59",
          5876 => x"78",
          5877 => x"a9",
          5878 => x"fe",
          5879 => x"82",
          5880 => x"29",
          5881 => x"11",
          5882 => x"b3",
          5883 => x"08",
          5884 => x"8c",
          5885 => x"07",
          5886 => x"ff",
          5887 => x"38",
          5888 => x"81",
          5889 => x"2b",
          5890 => x"25",
          5891 => x"52",
          5892 => x"86",
          5893 => x"38",
          5894 => x"74",
          5895 => x"77",
          5896 => x"ff",
          5897 => x"80",
          5898 => x"18",
          5899 => x"0c",
          5900 => x"70",
          5901 => x"fd",
          5902 => x"59",
          5903 => x"06",
          5904 => x"fe",
          5905 => x"88",
          5906 => x"c7",
          5907 => x"2e",
          5908 => x"9c",
          5909 => x"0c",
          5910 => x"51",
          5911 => x"08",
          5912 => x"51",
          5913 => x"08",
          5914 => x"74",
          5915 => x"75",
          5916 => x"84",
          5917 => x"08",
          5918 => x"08",
          5919 => x"84",
          5920 => x"0c",
          5921 => x"34",
          5922 => x"3d",
          5923 => x"89",
          5924 => x"53",
          5925 => x"84",
          5926 => x"84",
          5927 => x"2e",
          5928 => x"73",
          5929 => x"04",
          5930 => x"ff",
          5931 => x"55",
          5932 => x"ab",
          5933 => x"80",
          5934 => x"70",
          5935 => x"80",
          5936 => x"9b",
          5937 => x"2b",
          5938 => x"55",
          5939 => x"88",
          5940 => x"84",
          5941 => x"9a",
          5942 => x"74",
          5943 => x"ff",
          5944 => x"39",
          5945 => x"39",
          5946 => x"98",
          5947 => x"88",
          5948 => x"fa",
          5949 => x"80",
          5950 => x"80",
          5951 => x"80",
          5952 => x"16",
          5953 => x"38",
          5954 => x"73",
          5955 => x"88",
          5956 => x"ff",
          5957 => x"81",
          5958 => x"08",
          5959 => x"7a",
          5960 => x"2e",
          5961 => x"2e",
          5962 => x"2e",
          5963 => x"22",
          5964 => x"38",
          5965 => x"80",
          5966 => x"38",
          5967 => x"3f",
          5968 => x"84",
          5969 => x"84",
          5970 => x"ff",
          5971 => x"ff",
          5972 => x"84",
          5973 => x"2c",
          5974 => x"54",
          5975 => x"0d",
          5976 => x"ff",
          5977 => x"ff",
          5978 => x"84",
          5979 => x"2c",
          5980 => x"54",
          5981 => x"97",
          5982 => x"bb",
          5983 => x"14",
          5984 => x"bb",
          5985 => x"d8",
          5986 => x"d2",
          5987 => x"53",
          5988 => x"56",
          5989 => x"55",
          5990 => x"38",
          5991 => x"0d",
          5992 => x"9a",
          5993 => x"bb",
          5994 => x"05",
          5995 => x"74",
          5996 => x"38",
          5997 => x"3f",
          5998 => x"0d",
          5999 => x"95",
          6000 => x"68",
          6001 => x"05",
          6002 => x"84",
          6003 => x"08",
          6004 => x"9c",
          6005 => x"59",
          6006 => x"38",
          6007 => x"0c",
          6008 => x"08",
          6009 => x"82",
          6010 => x"bb",
          6011 => x"c1",
          6012 => x"56",
          6013 => x"38",
          6014 => x"81",
          6015 => x"17",
          6016 => x"a8",
          6017 => x"85",
          6018 => x"18",
          6019 => x"cc",
          6020 => x"82",
          6021 => x"11",
          6022 => x"71",
          6023 => x"72",
          6024 => x"ff",
          6025 => x"70",
          6026 => x"83",
          6027 => x"43",
          6028 => x"56",
          6029 => x"7a",
          6030 => x"07",
          6031 => x"bb",
          6032 => x"54",
          6033 => x"53",
          6034 => x"97",
          6035 => x"fe",
          6036 => x"18",
          6037 => x"31",
          6038 => x"a0",
          6039 => x"17",
          6040 => x"06",
          6041 => x"08",
          6042 => x"81",
          6043 => x"77",
          6044 => x"92",
          6045 => x"ff",
          6046 => x"ff",
          6047 => x"08",
          6048 => x"84",
          6049 => x"07",
          6050 => x"5a",
          6051 => x"26",
          6052 => x"18",
          6053 => x"77",
          6054 => x"17",
          6055 => x"71",
          6056 => x"25",
          6057 => x"1f",
          6058 => x"78",
          6059 => x"5a",
          6060 => x"7a",
          6061 => x"17",
          6062 => x"34",
          6063 => x"e7",
          6064 => x"57",
          6065 => x"56",
          6066 => x"55",
          6067 => x"22",
          6068 => x"2e",
          6069 => x"76",
          6070 => x"76",
          6071 => x"81",
          6072 => x"74",
          6073 => x"08",
          6074 => x"dd",
          6075 => x"08",
          6076 => x"89",
          6077 => x"d8",
          6078 => x"0c",
          6079 => x"80",
          6080 => x"76",
          6081 => x"80",
          6082 => x"08",
          6083 => x"33",
          6084 => x"bb",
          6085 => x"81",
          6086 => x"75",
          6087 => x"04",
          6088 => x"38",
          6089 => x"3f",
          6090 => x"84",
          6091 => x"bb",
          6092 => x"84",
          6093 => x"38",
          6094 => x"85",
          6095 => x"d8",
          6096 => x"19",
          6097 => x"ff",
          6098 => x"84",
          6099 => x"18",
          6100 => x"a0",
          6101 => x"fe",
          6102 => x"81",
          6103 => x"78",
          6104 => x"0b",
          6105 => x"80",
          6106 => x"98",
          6107 => x"83",
          6108 => x"81",
          6109 => x"2e",
          6110 => x"7a",
          6111 => x"08",
          6112 => x"08",
          6113 => x"55",
          6114 => x"81",
          6115 => x"18",
          6116 => x"2e",
          6117 => x"51",
          6118 => x"08",
          6119 => x"38",
          6120 => x"3f",
          6121 => x"84",
          6122 => x"bb",
          6123 => x"84",
          6124 => x"38",
          6125 => x"83",
          6126 => x"f6",
          6127 => x"19",
          6128 => x"90",
          6129 => x"17",
          6130 => x"34",
          6131 => x"38",
          6132 => x"59",
          6133 => x"39",
          6134 => x"fc",
          6135 => x"18",
          6136 => x"19",
          6137 => x"0b",
          6138 => x"39",
          6139 => x"5a",
          6140 => x"19",
          6141 => x"bb",
          6142 => x"57",
          6143 => x"53",
          6144 => x"3d",
          6145 => x"84",
          6146 => x"2e",
          6147 => x"a7",
          6148 => x"08",
          6149 => x"ac",
          6150 => x"84",
          6151 => x"93",
          6152 => x"59",
          6153 => x"98",
          6154 => x"02",
          6155 => x"5d",
          6156 => x"7d",
          6157 => x"12",
          6158 => x"41",
          6159 => x"80",
          6160 => x"57",
          6161 => x"56",
          6162 => x"38",
          6163 => x"08",
          6164 => x"8c",
          6165 => x"84",
          6166 => x"bb",
          6167 => x"ed",
          6168 => x"bb",
          6169 => x"bb",
          6170 => x"16",
          6171 => x"71",
          6172 => x"5d",
          6173 => x"84",
          6174 => x"fe",
          6175 => x"08",
          6176 => x"d3",
          6177 => x"cb",
          6178 => x"bb",
          6179 => x"30",
          6180 => x"7a",
          6181 => x"95",
          6182 => x"7b",
          6183 => x"26",
          6184 => x"d2",
          6185 => x"84",
          6186 => x"a7",
          6187 => x"19",
          6188 => x"76",
          6189 => x"7a",
          6190 => x"06",
          6191 => x"b8",
          6192 => x"f2",
          6193 => x"2e",
          6194 => x"b4",
          6195 => x"9c",
          6196 => x"0b",
          6197 => x"27",
          6198 => x"ff",
          6199 => x"56",
          6200 => x"96",
          6201 => x"fe",
          6202 => x"81",
          6203 => x"81",
          6204 => x"81",
          6205 => x"09",
          6206 => x"84",
          6207 => x"a8",
          6208 => x"59",
          6209 => x"eb",
          6210 => x"2e",
          6211 => x"54",
          6212 => x"53",
          6213 => x"f1",
          6214 => x"79",
          6215 => x"74",
          6216 => x"84",
          6217 => x"08",
          6218 => x"84",
          6219 => x"bb",
          6220 => x"80",
          6221 => x"d4",
          6222 => x"9c",
          6223 => x"58",
          6224 => x"38",
          6225 => x"33",
          6226 => x"79",
          6227 => x"80",
          6228 => x"f7",
          6229 => x"95",
          6230 => x"3d",
          6231 => x"05",
          6232 => x"3f",
          6233 => x"84",
          6234 => x"bb",
          6235 => x"43",
          6236 => x"ff",
          6237 => x"56",
          6238 => x"0b",
          6239 => x"04",
          6240 => x"81",
          6241 => x"33",
          6242 => x"86",
          6243 => x"74",
          6244 => x"83",
          6245 => x"57",
          6246 => x"87",
          6247 => x"80",
          6248 => x"2e",
          6249 => x"7d",
          6250 => x"5d",
          6251 => x"19",
          6252 => x"80",
          6253 => x"17",
          6254 => x"05",
          6255 => x"17",
          6256 => x"76",
          6257 => x"55",
          6258 => x"22",
          6259 => x"81",
          6260 => x"17",
          6261 => x"bb",
          6262 => x"58",
          6263 => x"81",
          6264 => x"70",
          6265 => x"ee",
          6266 => x"08",
          6267 => x"18",
          6268 => x"31",
          6269 => x"ee",
          6270 => x"2e",
          6271 => x"54",
          6272 => x"53",
          6273 => x"ee",
          6274 => x"7b",
          6275 => x"fd",
          6276 => x"fd",
          6277 => x"f3",
          6278 => x"84",
          6279 => x"38",
          6280 => x"8d",
          6281 => x"fd",
          6282 => x"51",
          6283 => x"08",
          6284 => x"11",
          6285 => x"7b",
          6286 => x"0c",
          6287 => x"84",
          6288 => x"ff",
          6289 => x"9f",
          6290 => x"74",
          6291 => x"76",
          6292 => x"38",
          6293 => x"75",
          6294 => x"56",
          6295 => x"b8",
          6296 => x"c3",
          6297 => x"1a",
          6298 => x"0b",
          6299 => x"80",
          6300 => x"ff",
          6301 => x"34",
          6302 => x"17",
          6303 => x"81",
          6304 => x"d8",
          6305 => x"70",
          6306 => x"05",
          6307 => x"38",
          6308 => x"34",
          6309 => x"5b",
          6310 => x"78",
          6311 => x"34",
          6312 => x"f0",
          6313 => x"34",
          6314 => x"bb",
          6315 => x"fd",
          6316 => x"08",
          6317 => x"97",
          6318 => x"80",
          6319 => x"58",
          6320 => x"2a",
          6321 => x"5a",
          6322 => x"55",
          6323 => x"81",
          6324 => x"ed",
          6325 => x"75",
          6326 => x"04",
          6327 => x"17",
          6328 => x"ed",
          6329 => x"2a",
          6330 => x"88",
          6331 => x"7d",
          6332 => x"1b",
          6333 => x"90",
          6334 => x"88",
          6335 => x"55",
          6336 => x"81",
          6337 => x"ec",
          6338 => x"ff",
          6339 => x"b4",
          6340 => x"80",
          6341 => x"5b",
          6342 => x"ba",
          6343 => x"75",
          6344 => x"b1",
          6345 => x"51",
          6346 => x"08",
          6347 => x"8a",
          6348 => x"3d",
          6349 => x"3d",
          6350 => x"ff",
          6351 => x"56",
          6352 => x"81",
          6353 => x"86",
          6354 => x"3d",
          6355 => x"70",
          6356 => x"05",
          6357 => x"38",
          6358 => x"58",
          6359 => x"77",
          6360 => x"55",
          6361 => x"77",
          6362 => x"84",
          6363 => x"d8",
          6364 => x"cb",
          6365 => x"b1",
          6366 => x"70",
          6367 => x"89",
          6368 => x"ff",
          6369 => x"2e",
          6370 => x"e6",
          6371 => x"5f",
          6372 => x"79",
          6373 => x"12",
          6374 => x"38",
          6375 => x"55",
          6376 => x"89",
          6377 => x"58",
          6378 => x"55",
          6379 => x"38",
          6380 => x"70",
          6381 => x"07",
          6382 => x"38",
          6383 => x"83",
          6384 => x"5a",
          6385 => x"fd",
          6386 => x"b1",
          6387 => x"51",
          6388 => x"08",
          6389 => x"38",
          6390 => x"2e",
          6391 => x"51",
          6392 => x"08",
          6393 => x"38",
          6394 => x"88",
          6395 => x"75",
          6396 => x"81",
          6397 => x"ef",
          6398 => x"19",
          6399 => x"81",
          6400 => x"a0",
          6401 => x"5d",
          6402 => x"33",
          6403 => x"75",
          6404 => x"08",
          6405 => x"19",
          6406 => x"07",
          6407 => x"83",
          6408 => x"18",
          6409 => x"27",
          6410 => x"71",
          6411 => x"75",
          6412 => x"5d",
          6413 => x"38",
          6414 => x"38",
          6415 => x"81",
          6416 => x"84",
          6417 => x"ff",
          6418 => x"7f",
          6419 => x"7b",
          6420 => x"79",
          6421 => x"6a",
          6422 => x"7b",
          6423 => x"58",
          6424 => x"5b",
          6425 => x"38",
          6426 => x"18",
          6427 => x"ed",
          6428 => x"18",
          6429 => x"3d",
          6430 => x"95",
          6431 => x"db",
          6432 => x"bb",
          6433 => x"5c",
          6434 => x"16",
          6435 => x"33",
          6436 => x"81",
          6437 => x"53",
          6438 => x"fe",
          6439 => x"80",
          6440 => x"76",
          6441 => x"38",
          6442 => x"81",
          6443 => x"7b",
          6444 => x"fe",
          6445 => x"55",
          6446 => x"98",
          6447 => x"e1",
          6448 => x"7f",
          6449 => x"84",
          6450 => x"0d",
          6451 => x"b1",
          6452 => x"19",
          6453 => x"07",
          6454 => x"39",
          6455 => x"fe",
          6456 => x"fe",
          6457 => x"b1",
          6458 => x"08",
          6459 => x"fe",
          6460 => x"84",
          6461 => x"db",
          6462 => x"34",
          6463 => x"84",
          6464 => x"17",
          6465 => x"33",
          6466 => x"fe",
          6467 => x"a0",
          6468 => x"16",
          6469 => x"58",
          6470 => x"08",
          6471 => x"33",
          6472 => x"5c",
          6473 => x"84",
          6474 => x"17",
          6475 => x"84",
          6476 => x"27",
          6477 => x"7c",
          6478 => x"38",
          6479 => x"08",
          6480 => x"51",
          6481 => x"e8",
          6482 => x"05",
          6483 => x"33",
          6484 => x"05",
          6485 => x"3f",
          6486 => x"84",
          6487 => x"bb",
          6488 => x"5a",
          6489 => x"ff",
          6490 => x"56",
          6491 => x"80",
          6492 => x"86",
          6493 => x"61",
          6494 => x"7a",
          6495 => x"73",
          6496 => x"83",
          6497 => x"3f",
          6498 => x"0c",
          6499 => x"67",
          6500 => x"52",
          6501 => x"84",
          6502 => x"08",
          6503 => x"84",
          6504 => x"66",
          6505 => x"96",
          6506 => x"84",
          6507 => x"cf",
          6508 => x"55",
          6509 => x"86",
          6510 => x"59",
          6511 => x"2a",
          6512 => x"2a",
          6513 => x"2a",
          6514 => x"81",
          6515 => x"e1",
          6516 => x"bb",
          6517 => x"3d",
          6518 => x"9a",
          6519 => x"ff",
          6520 => x"84",
          6521 => x"84",
          6522 => x"7a",
          6523 => x"06",
          6524 => x"30",
          6525 => x"7b",
          6526 => x"76",
          6527 => x"80",
          6528 => x"80",
          6529 => x"f6",
          6530 => x"74",
          6531 => x"38",
          6532 => x"81",
          6533 => x"84",
          6534 => x"ff",
          6535 => x"78",
          6536 => x"56",
          6537 => x"8b",
          6538 => x"83",
          6539 => x"83",
          6540 => x"2b",
          6541 => x"70",
          6542 => x"07",
          6543 => x"56",
          6544 => x"0d",
          6545 => x"8e",
          6546 => x"3f",
          6547 => x"84",
          6548 => x"84",
          6549 => x"80",
          6550 => x"77",
          6551 => x"70",
          6552 => x"dc",
          6553 => x"08",
          6554 => x"38",
          6555 => x"b4",
          6556 => x"bb",
          6557 => x"08",
          6558 => x"55",
          6559 => x"a0",
          6560 => x"17",
          6561 => x"33",
          6562 => x"81",
          6563 => x"16",
          6564 => x"bb",
          6565 => x"fe",
          6566 => x"f8",
          6567 => x"84",
          6568 => x"bb",
          6569 => x"5c",
          6570 => x"1b",
          6571 => x"81",
          6572 => x"8b",
          6573 => x"77",
          6574 => x"7b",
          6575 => x"a0",
          6576 => x"57",
          6577 => x"53",
          6578 => x"3d",
          6579 => x"84",
          6580 => x"a6",
          6581 => x"55",
          6582 => x"ff",
          6583 => x"3d",
          6584 => x"5b",
          6585 => x"b7",
          6586 => x"75",
          6587 => x"74",
          6588 => x"83",
          6589 => x"51",
          6590 => x"bb",
          6591 => x"bb",
          6592 => x"76",
          6593 => x"94",
          6594 => x"ff",
          6595 => x"81",
          6596 => x"99",
          6597 => x"ff",
          6598 => x"89",
          6599 => x"e9",
          6600 => x"81",
          6601 => x"f8",
          6602 => x"81",
          6603 => x"2a",
          6604 => x"34",
          6605 => x"05",
          6606 => x"70",
          6607 => x"58",
          6608 => x"8f",
          6609 => x"e5",
          6610 => x"38",
          6611 => x"33",
          6612 => x"06",
          6613 => x"38",
          6614 => x"3d",
          6615 => x"84",
          6616 => x"08",
          6617 => x"84",
          6618 => x"83",
          6619 => x"84",
          6620 => x"55",
          6621 => x"84",
          6622 => x"83",
          6623 => x"81",
          6624 => x"84",
          6625 => x"08",
          6626 => x"c4",
          6627 => x"76",
          6628 => x"81",
          6629 => x"ef",
          6630 => x"34",
          6631 => x"bb",
          6632 => x"39",
          6633 => x"56",
          6634 => x"84",
          6635 => x"80",
          6636 => x"75",
          6637 => x"ee",
          6638 => x"84",
          6639 => x"06",
          6640 => x"b8",
          6641 => x"80",
          6642 => x"38",
          6643 => x"09",
          6644 => x"76",
          6645 => x"51",
          6646 => x"08",
          6647 => x"59",
          6648 => x"be",
          6649 => x"57",
          6650 => x"9e",
          6651 => x"07",
          6652 => x"38",
          6653 => x"38",
          6654 => x"3f",
          6655 => x"84",
          6656 => x"55",
          6657 => x"55",
          6658 => x"55",
          6659 => x"ff",
          6660 => x"88",
          6661 => x"59",
          6662 => x"33",
          6663 => x"15",
          6664 => x"76",
          6665 => x"81",
          6666 => x"da",
          6667 => x"7a",
          6668 => x"34",
          6669 => x"bb",
          6670 => x"57",
          6671 => x"08",
          6672 => x"fe",
          6673 => x"79",
          6674 => x"84",
          6675 => x"18",
          6676 => x"a0",
          6677 => x"33",
          6678 => x"bb",
          6679 => x"5a",
          6680 => x"3f",
          6681 => x"84",
          6682 => x"ae",
          6683 => x"2e",
          6684 => x"54",
          6685 => x"53",
          6686 => x"d4",
          6687 => x"0d",
          6688 => x"05",
          6689 => x"80",
          6690 => x"80",
          6691 => x"80",
          6692 => x"18",
          6693 => x"c2",
          6694 => x"a5",
          6695 => x"9d",
          6696 => x"8c",
          6697 => x"33",
          6698 => x"74",
          6699 => x"11",
          6700 => x"54",
          6701 => x"ff",
          6702 => x"07",
          6703 => x"90",
          6704 => x"58",
          6705 => x"08",
          6706 => x"78",
          6707 => x"51",
          6708 => x"55",
          6709 => x"38",
          6710 => x"2e",
          6711 => x"ff",
          6712 => x"08",
          6713 => x"7d",
          6714 => x"81",
          6715 => x"73",
          6716 => x"04",
          6717 => x"3d",
          6718 => x"d0",
          6719 => x"06",
          6720 => x"08",
          6721 => x"2e",
          6722 => x"7c",
          6723 => x"74",
          6724 => x"77",
          6725 => x"84",
          6726 => x"08",
          6727 => x"17",
          6728 => x"7e",
          6729 => x"ff",
          6730 => x"8c",
          6731 => x"07",
          6732 => x"08",
          6733 => x"76",
          6734 => x"31",
          6735 => x"07",
          6736 => x"fe",
          6737 => x"74",
          6738 => x"54",
          6739 => x"39",
          6740 => x"bb",
          6741 => x"08",
          6742 => x"87",
          6743 => x"a2",
          6744 => x"80",
          6745 => x"05",
          6746 => x"75",
          6747 => x"38",
          6748 => x"e2",
          6749 => x"e5",
          6750 => x"05",
          6751 => x"84",
          6752 => x"ba",
          6753 => x"33",
          6754 => x"fe",
          6755 => x"81",
          6756 => x"83",
          6757 => x"2a",
          6758 => x"9f",
          6759 => x"52",
          6760 => x"bb",
          6761 => x"74",
          6762 => x"80",
          6763 => x"75",
          6764 => x"80",
          6765 => x"83",
          6766 => x"83",
          6767 => x"74",
          6768 => x"3d",
          6769 => x"59",
          6770 => x"ab",
          6771 => x"07",
          6772 => x"38",
          6773 => x"54",
          6774 => x"cd",
          6775 => x"08",
          6776 => x"33",
          6777 => x"2b",
          6778 => x"d4",
          6779 => x"38",
          6780 => x"11",
          6781 => x"e7",
          6782 => x"82",
          6783 => x"2b",
          6784 => x"88",
          6785 => x"1f",
          6786 => x"90",
          6787 => x"33",
          6788 => x"71",
          6789 => x"3d",
          6790 => x"45",
          6791 => x"8e",
          6792 => x"38",
          6793 => x"87",
          6794 => x"45",
          6795 => x"61",
          6796 => x"38",
          6797 => x"38",
          6798 => x"7a",
          6799 => x"7a",
          6800 => x"0b",
          6801 => x"80",
          6802 => x"38",
          6803 => x"17",
          6804 => x"2e",
          6805 => x"77",
          6806 => x"84",
          6807 => x"84",
          6808 => x"38",
          6809 => x"84",
          6810 => x"2a",
          6811 => x"15",
          6812 => x"7b",
          6813 => x"ff",
          6814 => x"4e",
          6815 => x"38",
          6816 => x"70",
          6817 => x"82",
          6818 => x"78",
          6819 => x"ff",
          6820 => x"62",
          6821 => x"2e",
          6822 => x"ff",
          6823 => x"82",
          6824 => x"18",
          6825 => x"38",
          6826 => x"76",
          6827 => x"84",
          6828 => x"fe",
          6829 => x"9f",
          6830 => x"7c",
          6831 => x"57",
          6832 => x"82",
          6833 => x"5d",
          6834 => x"80",
          6835 => x"08",
          6836 => x"5c",
          6837 => x"ff",
          6838 => x"26",
          6839 => x"06",
          6840 => x"99",
          6841 => x"ff",
          6842 => x"2a",
          6843 => x"06",
          6844 => x"7a",
          6845 => x"2a",
          6846 => x"2e",
          6847 => x"5f",
          6848 => x"7f",
          6849 => x"05",
          6850 => x"96",
          6851 => x"fe",
          6852 => x"84",
          6853 => x"38",
          6854 => x"75",
          6855 => x"59",
          6856 => x"39",
          6857 => x"7a",
          6858 => x"61",
          6859 => x"2e",
          6860 => x"4a",
          6861 => x"84",
          6862 => x"8b",
          6863 => x"27",
          6864 => x"bb",
          6865 => x"90",
          6866 => x"86",
          6867 => x"38",
          6868 => x"fd",
          6869 => x"80",
          6870 => x"15",
          6871 => x"e6",
          6872 => x"05",
          6873 => x"34",
          6874 => x"8b",
          6875 => x"8c",
          6876 => x"7b",
          6877 => x"8e",
          6878 => x"61",
          6879 => x"34",
          6880 => x"80",
          6881 => x"82",
          6882 => x"6c",
          6883 => x"ad",
          6884 => x"74",
          6885 => x"4c",
          6886 => x"95",
          6887 => x"80",
          6888 => x"05",
          6889 => x"61",
          6890 => x"67",
          6891 => x"4c",
          6892 => x"2a",
          6893 => x"08",
          6894 => x"85",
          6895 => x"80",
          6896 => x"05",
          6897 => x"7c",
          6898 => x"96",
          6899 => x"61",
          6900 => x"05",
          6901 => x"61",
          6902 => x"55",
          6903 => x"70",
          6904 => x"74",
          6905 => x"80",
          6906 => x"4b",
          6907 => x"53",
          6908 => x"3f",
          6909 => x"e7",
          6910 => x"87",
          6911 => x"76",
          6912 => x"55",
          6913 => x"62",
          6914 => x"ff",
          6915 => x"f8",
          6916 => x"7c",
          6917 => x"46",
          6918 => x"70",
          6919 => x"56",
          6920 => x"76",
          6921 => x"54",
          6922 => x"c5",
          6923 => x"e6",
          6924 => x"76",
          6925 => x"55",
          6926 => x"31",
          6927 => x"05",
          6928 => x"77",
          6929 => x"56",
          6930 => x"75",
          6931 => x"79",
          6932 => x"84",
          6933 => x"76",
          6934 => x"58",
          6935 => x"6c",
          6936 => x"58",
          6937 => x"7d",
          6938 => x"06",
          6939 => x"61",
          6940 => x"57",
          6941 => x"80",
          6942 => x"60",
          6943 => x"81",
          6944 => x"05",
          6945 => x"67",
          6946 => x"c1",
          6947 => x"3f",
          6948 => x"84",
          6949 => x"67",
          6950 => x"67",
          6951 => x"05",
          6952 => x"6b",
          6953 => x"90",
          6954 => x"61",
          6955 => x"45",
          6956 => x"90",
          6957 => x"34",
          6958 => x"cd",
          6959 => x"52",
          6960 => x"57",
          6961 => x"80",
          6962 => x"96",
          6963 => x"f7",
          6964 => x"bb",
          6965 => x"90",
          6966 => x"74",
          6967 => x"39",
          6968 => x"81",
          6969 => x"74",
          6970 => x"98",
          6971 => x"82",
          6972 => x"80",
          6973 => x"38",
          6974 => x"3f",
          6975 => x"87",
          6976 => x"5c",
          6977 => x"80",
          6978 => x"0a",
          6979 => x"f8",
          6980 => x"ff",
          6981 => x"d3",
          6982 => x"bf",
          6983 => x"81",
          6984 => x"38",
          6985 => x"a0",
          6986 => x"61",
          6987 => x"7a",
          6988 => x"57",
          6989 => x"39",
          6990 => x"61",
          6991 => x"c5",
          6992 => x"05",
          6993 => x"88",
          6994 => x"7c",
          6995 => x"34",
          6996 => x"05",
          6997 => x"61",
          6998 => x"34",
          6999 => x"b0",
          7000 => x"86",
          7001 => x"05",
          7002 => x"34",
          7003 => x"61",
          7004 => x"57",
          7005 => x"76",
          7006 => x"55",
          7007 => x"70",
          7008 => x"05",
          7009 => x"38",
          7010 => x"60",
          7011 => x"81",
          7012 => x"38",
          7013 => x"62",
          7014 => x"bb",
          7015 => x"fe",
          7016 => x"0b",
          7017 => x"84",
          7018 => x"7b",
          7019 => x"34",
          7020 => x"ff",
          7021 => x"ff",
          7022 => x"05",
          7023 => x"61",
          7024 => x"34",
          7025 => x"34",
          7026 => x"86",
          7027 => x"bf",
          7028 => x"80",
          7029 => x"17",
          7030 => x"d2",
          7031 => x"55",
          7032 => x"34",
          7033 => x"34",
          7034 => x"83",
          7035 => x"e5",
          7036 => x"05",
          7037 => x"34",
          7038 => x"e8",
          7039 => x"61",
          7040 => x"56",
          7041 => x"98",
          7042 => x"34",
          7043 => x"61",
          7044 => x"ee",
          7045 => x"34",
          7046 => x"34",
          7047 => x"79",
          7048 => x"81",
          7049 => x"bd",
          7050 => x"a6",
          7051 => x"5b",
          7052 => x"57",
          7053 => x"59",
          7054 => x"78",
          7055 => x"7b",
          7056 => x"8d",
          7057 => x"38",
          7058 => x"81",
          7059 => x"77",
          7060 => x"7a",
          7061 => x"84",
          7062 => x"f7",
          7063 => x"05",
          7064 => x"d5",
          7065 => x"24",
          7066 => x"8c",
          7067 => x"16",
          7068 => x"84",
          7069 => x"8b",
          7070 => x"54",
          7071 => x"51",
          7072 => x"70",
          7073 => x"30",
          7074 => x"0c",
          7075 => x"76",
          7076 => x"e3",
          7077 => x"8d",
          7078 => x"55",
          7079 => x"ff",
          7080 => x"08",
          7081 => x"38",
          7082 => x"38",
          7083 => x"77",
          7084 => x"24",
          7085 => x"19",
          7086 => x"24",
          7087 => x"55",
          7088 => x"51",
          7089 => x"08",
          7090 => x"ff",
          7091 => x"0d",
          7092 => x"75",
          7093 => x"ff",
          7094 => x"30",
          7095 => x"52",
          7096 => x"52",
          7097 => x"39",
          7098 => x"0d",
          7099 => x"05",
          7100 => x"72",
          7101 => x"ff",
          7102 => x"0c",
          7103 => x"73",
          7104 => x"81",
          7105 => x"38",
          7106 => x"2e",
          7107 => x"ff",
          7108 => x"8d",
          7109 => x"70",
          7110 => x"12",
          7111 => x"0c",
          7112 => x"0d",
          7113 => x"96",
          7114 => x"80",
          7115 => x"84",
          7116 => x"71",
          7117 => x"38",
          7118 => x"10",
          7119 => x"bb",
          7120 => x"fb",
          7121 => x"ff",
          7122 => x"ff",
          7123 => x"9f",
          7124 => x"82",
          7125 => x"80",
          7126 => x"53",
          7127 => x"05",
          7128 => x"56",
          7129 => x"70",
          7130 => x"73",
          7131 => x"22",
          7132 => x"79",
          7133 => x"2e",
          7134 => x"84",
          7135 => x"bc",
          7136 => x"ea",
          7137 => x"05",
          7138 => x"70",
          7139 => x"51",
          7140 => x"ff",
          7141 => x"16",
          7142 => x"e6",
          7143 => x"06",
          7144 => x"83",
          7145 => x"e0",
          7146 => x"51",
          7147 => x"ff",
          7148 => x"73",
          7149 => x"83",
          7150 => x"a6",
          7151 => x"70",
          7152 => x"00",
          7153 => x"ff",
          7154 => x"ff",
          7155 => x"19",
          7156 => x"19",
          7157 => x"19",
          7158 => x"19",
          7159 => x"19",
          7160 => x"19",
          7161 => x"18",
          7162 => x"18",
          7163 => x"18",
          7164 => x"18",
          7165 => x"1f",
          7166 => x"1f",
          7167 => x"1f",
          7168 => x"1f",
          7169 => x"1f",
          7170 => x"1f",
          7171 => x"1f",
          7172 => x"1f",
          7173 => x"1f",
          7174 => x"1f",
          7175 => x"1f",
          7176 => x"1f",
          7177 => x"1f",
          7178 => x"1f",
          7179 => x"1f",
          7180 => x"1f",
          7181 => x"1f",
          7182 => x"1f",
          7183 => x"1f",
          7184 => x"1f",
          7185 => x"1f",
          7186 => x"24",
          7187 => x"1f",
          7188 => x"1f",
          7189 => x"1f",
          7190 => x"1f",
          7191 => x"1f",
          7192 => x"1f",
          7193 => x"1f",
          7194 => x"1f",
          7195 => x"23",
          7196 => x"22",
          7197 => x"23",
          7198 => x"21",
          7199 => x"1f",
          7200 => x"1f",
          7201 => x"1f",
          7202 => x"1f",
          7203 => x"1f",
          7204 => x"1f",
          7205 => x"1f",
          7206 => x"1f",
          7207 => x"1f",
          7208 => x"1f",
          7209 => x"1f",
          7210 => x"1f",
          7211 => x"1f",
          7212 => x"1f",
          7213 => x"1f",
          7214 => x"1f",
          7215 => x"1f",
          7216 => x"1f",
          7217 => x"1f",
          7218 => x"1f",
          7219 => x"1f",
          7220 => x"1f",
          7221 => x"1f",
          7222 => x"1f",
          7223 => x"1f",
          7224 => x"1f",
          7225 => x"21",
          7226 => x"1f",
          7227 => x"1f",
          7228 => x"1f",
          7229 => x"1f",
          7230 => x"21",
          7231 => x"21",
          7232 => x"21",
          7233 => x"21",
          7234 => x"32",
          7235 => x"32",
          7236 => x"32",
          7237 => x"3a",
          7238 => x"36",
          7239 => x"34",
          7240 => x"36",
          7241 => x"36",
          7242 => x"39",
          7243 => x"39",
          7244 => x"37",
          7245 => x"34",
          7246 => x"36",
          7247 => x"36",
          7248 => x"47",
          7249 => x"47",
          7250 => x"47",
          7251 => x"48",
          7252 => x"48",
          7253 => x"48",
          7254 => x"48",
          7255 => x"48",
          7256 => x"48",
          7257 => x"48",
          7258 => x"48",
          7259 => x"48",
          7260 => x"48",
          7261 => x"48",
          7262 => x"48",
          7263 => x"48",
          7264 => x"48",
          7265 => x"48",
          7266 => x"49",
          7267 => x"49",
          7268 => x"48",
          7269 => x"48",
          7270 => x"48",
          7271 => x"48",
          7272 => x"48",
          7273 => x"48",
          7274 => x"48",
          7275 => x"48",
          7276 => x"54",
          7277 => x"56",
          7278 => x"55",
          7279 => x"54",
          7280 => x"53",
          7281 => x"58",
          7282 => x"53",
          7283 => x"53",
          7284 => x"53",
          7285 => x"58",
          7286 => x"53",
          7287 => x"53",
          7288 => x"53",
          7289 => x"53",
          7290 => x"53",
          7291 => x"53",
          7292 => x"53",
          7293 => x"53",
          7294 => x"53",
          7295 => x"53",
          7296 => x"53",
          7297 => x"53",
          7298 => x"54",
          7299 => x"53",
          7300 => x"53",
          7301 => x"54",
          7302 => x"54",
          7303 => x"59",
          7304 => x"59",
          7305 => x"59",
          7306 => x"59",
          7307 => x"59",
          7308 => x"59",
          7309 => x"59",
          7310 => x"59",
          7311 => x"59",
          7312 => x"59",
          7313 => x"59",
          7314 => x"59",
          7315 => x"59",
          7316 => x"59",
          7317 => x"59",
          7318 => x"5a",
          7319 => x"5a",
          7320 => x"5b",
          7321 => x"5b",
          7322 => x"5b",
          7323 => x"5b",
          7324 => x"5a",
          7325 => x"5a",
          7326 => x"5a",
          7327 => x"5a",
          7328 => x"62",
          7329 => x"62",
          7330 => x"62",
          7331 => x"62",
          7332 => x"62",
          7333 => x"62",
          7334 => x"62",
          7335 => x"62",
          7336 => x"62",
          7337 => x"62",
          7338 => x"64",
          7339 => x"62",
          7340 => x"62",
          7341 => x"5f",
          7342 => x"df",
          7343 => x"df",
          7344 => x"df",
          7345 => x"df",
          7346 => x"df",
          7347 => x"0b",
          7348 => x"0f",
          7349 => x"0b",
          7350 => x"0b",
          7351 => x"0b",
          7352 => x"0d",
          7353 => x"0f",
          7354 => x"0b",
          7355 => x"0b",
          7356 => x"0b",
          7357 => x"0b",
          7358 => x"0b",
          7359 => x"0b",
          7360 => x"0b",
          7361 => x"0b",
          7362 => x"0b",
          7363 => x"0b",
          7364 => x"0b",
          7365 => x"0b",
          7366 => x"0b",
          7367 => x"0b",
          7368 => x"0b",
          7369 => x"0b",
          7370 => x"0b",
          7371 => x"0b",
          7372 => x"0f",
          7373 => x"0b",
          7374 => x"0b",
          7375 => x"0b",
          7376 => x"0b",
          7377 => x"0b",
          7378 => x"0b",
          7379 => x"0b",
          7380 => x"0e",
          7381 => x"0e",
          7382 => x"0e",
          7383 => x"0e",
          7384 => x"0b",
          7385 => x"0b",
          7386 => x"0c",
          7387 => x"0b",
          7388 => x"0f",
          7389 => x"0c",
          7390 => x"0b",
          7391 => x"6e",
          7392 => x"6f",
          7393 => x"6e",
          7394 => x"6f",
          7395 => x"78",
          7396 => x"6c",
          7397 => x"6f",
          7398 => x"69",
          7399 => x"75",
          7400 => x"62",
          7401 => x"77",
          7402 => x"65",
          7403 => x"65",
          7404 => x"00",
          7405 => x"73",
          7406 => x"73",
          7407 => x"66",
          7408 => x"73",
          7409 => x"73",
          7410 => x"61",
          7411 => x"61",
          7412 => x"6c",
          7413 => x"00",
          7414 => x"6e",
          7415 => x"00",
          7416 => x"74",
          7417 => x"6f",
          7418 => x"00",
          7419 => x"6e",
          7420 => x"66",
          7421 => x"00",
          7422 => x"69",
          7423 => x"65",
          7424 => x"00",
          7425 => x"73",
          7426 => x"2e",
          7427 => x"74",
          7428 => x"74",
          7429 => x"63",
          7430 => x"00",
          7431 => x"20",
          7432 => x"2e",
          7433 => x"70",
          7434 => x"66",
          7435 => x"65",
          7436 => x"20",
          7437 => x"2e",
          7438 => x"6f",
          7439 => x"65",
          7440 => x"69",
          7441 => x"65",
          7442 => x"76",
          7443 => x"00",
          7444 => x"77",
          7445 => x"6f",
          7446 => x"00",
          7447 => x"61",
          7448 => x"76",
          7449 => x"00",
          7450 => x"6c",
          7451 => x"78",
          7452 => x"00",
          7453 => x"20",
          7454 => x"00",
          7455 => x"64",
          7456 => x"6d",
          7457 => x"20",
          7458 => x"75",
          7459 => x"20",
          7460 => x"75",
          7461 => x"73",
          7462 => x"65",
          7463 => x"74",
          7464 => x"72",
          7465 => x"73",
          7466 => x"00",
          7467 => x"73",
          7468 => x"6c",
          7469 => x"20",
          7470 => x"6c",
          7471 => x"2f",
          7472 => x"00",
          7473 => x"00",
          7474 => x"00",
          7475 => x"32",
          7476 => x"00",
          7477 => x"00",
          7478 => x"00",
          7479 => x"20",
          7480 => x"53",
          7481 => x"28",
          7482 => x"32",
          7483 => x"2e",
          7484 => x"50",
          7485 => x"25",
          7486 => x"20",
          7487 => x"00",
          7488 => x"20",
          7489 => x"64",
          7490 => x"20",
          7491 => x"20",
          7492 => x"6c",
          7493 => x"20",
          7494 => x"64",
          7495 => x"20",
          7496 => x"20",
          7497 => x"6c",
          7498 => x"55",
          7499 => x"75",
          7500 => x"6c",
          7501 => x"52",
          7502 => x"6e",
          7503 => x"00",
          7504 => x"52",
          7505 => x"72",
          7506 => x"52",
          7507 => x"6e",
          7508 => x"00",
          7509 => x"52",
          7510 => x"72",
          7511 => x"43",
          7512 => x"6e",
          7513 => x"00",
          7514 => x"52",
          7515 => x"72",
          7516 => x"32",
          7517 => x"75",
          7518 => x"6d",
          7519 => x"72",
          7520 => x"74",
          7521 => x"20",
          7522 => x"2e",
          7523 => x"6e",
          7524 => x"2e",
          7525 => x"74",
          7526 => x"61",
          7527 => x"53",
          7528 => x"74",
          7529 => x"20",
          7530 => x"69",
          7531 => x"64",
          7532 => x"2c",
          7533 => x"20",
          7534 => x"6e",
          7535 => x"00",
          7536 => x"3a",
          7537 => x"00",
          7538 => x"6d",
          7539 => x"00",
          7540 => x"6e",
          7541 => x"5c",
          7542 => x"00",
          7543 => x"65",
          7544 => x"2e",
          7545 => x"73",
          7546 => x"20",
          7547 => x"74",
          7548 => x"00",
          7549 => x"67",
          7550 => x"20",
          7551 => x"2e",
          7552 => x"6c",
          7553 => x"6e",
          7554 => x"20",
          7555 => x"00",
          7556 => x"69",
          7557 => x"20",
          7558 => x"20",
          7559 => x"38",
          7560 => x"58",
          7561 => x"38",
          7562 => x"2d",
          7563 => x"69",
          7564 => x"00",
          7565 => x"25",
          7566 => x"30",
          7567 => x"78",
          7568 => x"70",
          7569 => x"00",
          7570 => x"25",
          7571 => x"65",
          7572 => x"2e",
          7573 => x"6d",
          7574 => x"79",
          7575 => x"65",
          7576 => x"3a",
          7577 => x"00",
          7578 => x"20",
          7579 => x"65",
          7580 => x"6f",
          7581 => x"73",
          7582 => x"6e",
          7583 => x"3f",
          7584 => x"25",
          7585 => x"3a",
          7586 => x"0a",
          7587 => x"6e",
          7588 => x"69",
          7589 => x"44",
          7590 => x"69",
          7591 => x"74",
          7592 => x"64",
          7593 => x"00",
          7594 => x"55",
          7595 => x"56",
          7596 => x"64",
          7597 => x"20",
          7598 => x"00",
          7599 => x"55",
          7600 => x"20",
          7601 => x"64",
          7602 => x"20",
          7603 => x"00",
          7604 => x"61",
          7605 => x"74",
          7606 => x"73",
          7607 => x"20",
          7608 => x"00",
          7609 => x"00",
          7610 => x"55",
          7611 => x"20",
          7612 => x"20",
          7613 => x"20",
          7614 => x"00",
          7615 => x"73",
          7616 => x"63",
          7617 => x"20",
          7618 => x"20",
          7619 => x"4d",
          7620 => x"20",
          7621 => x"6e",
          7622 => x"20",
          7623 => x"72",
          7624 => x"25",
          7625 => x"00",
          7626 => x"52",
          7627 => x"6b",
          7628 => x"20",
          7629 => x"20",
          7630 => x"4d",
          7631 => x"20",
          7632 => x"20",
          7633 => x"20",
          7634 => x"00",
          7635 => x"20",
          7636 => x"20",
          7637 => x"4e",
          7638 => x"00",
          7639 => x"54",
          7640 => x"28",
          7641 => x"73",
          7642 => x"0a",
          7643 => x"4d",
          7644 => x"28",
          7645 => x"20",
          7646 => x"0a",
          7647 => x"20",
          7648 => x"28",
          7649 => x"20",
          7650 => x"0a",
          7651 => x"4d",
          7652 => x"28",
          7653 => x"38",
          7654 => x"20",
          7655 => x"20",
          7656 => x"58",
          7657 => x"0a",
          7658 => x"53",
          7659 => x"28",
          7660 => x"38",
          7661 => x"20",
          7662 => x"20",
          7663 => x"58",
          7664 => x"0a",
          7665 => x"20",
          7666 => x"28",
          7667 => x"38",
          7668 => x"66",
          7669 => x"20",
          7670 => x"00",
          7671 => x"6e",
          7672 => x"00",
          7673 => x"00",
          7674 => x"00",
          7675 => x"00",
          7676 => x"f1",
          7677 => x"00",
          7678 => x"00",
          7679 => x"f1",
          7680 => x"00",
          7681 => x"00",
          7682 => x"f1",
          7683 => x"00",
          7684 => x"00",
          7685 => x"f1",
          7686 => x"00",
          7687 => x"00",
          7688 => x"f1",
          7689 => x"00",
          7690 => x"00",
          7691 => x"f1",
          7692 => x"00",
          7693 => x"00",
          7694 => x"f1",
          7695 => x"00",
          7696 => x"00",
          7697 => x"f1",
          7698 => x"00",
          7699 => x"00",
          7700 => x"f0",
          7701 => x"00",
          7702 => x"00",
          7703 => x"f0",
          7704 => x"00",
          7705 => x"00",
          7706 => x"f0",
          7707 => x"00",
          7708 => x"00",
          7709 => x"44",
          7710 => x"42",
          7711 => x"36",
          7712 => x"34",
          7713 => x"33",
          7714 => x"31",
          7715 => x"00",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"73",
          7721 => x"61",
          7722 => x"0a",
          7723 => x"20",
          7724 => x"65",
          7725 => x"74",
          7726 => x"65",
          7727 => x"6c",
          7728 => x"73",
          7729 => x"73",
          7730 => x"00",
          7731 => x"79",
          7732 => x"40",
          7733 => x"00",
          7734 => x"20",
          7735 => x"69",
          7736 => x"72",
          7737 => x"65",
          7738 => x"79",
          7739 => x"6f",
          7740 => x"00",
          7741 => x"00",
          7742 => x"00",
          7743 => x"42",
          7744 => x"44",
          7745 => x"00",
          7746 => x"00",
          7747 => x"00",
          7748 => x"00",
          7749 => x"00",
          7750 => x"00",
          7751 => x"00",
          7752 => x"00",
          7753 => x"00",
          7754 => x"00",
          7755 => x"00",
          7756 => x"00",
          7757 => x"35",
          7758 => x"36",
          7759 => x"25",
          7760 => x"2c",
          7761 => x"64",
          7762 => x"00",
          7763 => x"64",
          7764 => x"25",
          7765 => x"3a",
          7766 => x"25",
          7767 => x"32",
          7768 => x"5b",
          7769 => x"00",
          7770 => x"20",
          7771 => x"00",
          7772 => x"78",
          7773 => x"00",
          7774 => x"78",
          7775 => x"00",
          7776 => x"78",
          7777 => x"20",
          7778 => x"66",
          7779 => x"00",
          7780 => x"3a",
          7781 => x"00",
          7782 => x"00",
          7783 => x"54",
          7784 => x"90",
          7785 => x"30",
          7786 => x"45",
          7787 => x"20",
          7788 => x"20",
          7789 => x"20",
          7790 => x"20",
          7791 => x"00",
          7792 => x"00",
          7793 => x"10",
          7794 => x"00",
          7795 => x"8f",
          7796 => x"8e",
          7797 => x"55",
          7798 => x"9e",
          7799 => x"a6",
          7800 => x"ae",
          7801 => x"b6",
          7802 => x"be",
          7803 => x"c6",
          7804 => x"ce",
          7805 => x"d6",
          7806 => x"de",
          7807 => x"e6",
          7808 => x"ee",
          7809 => x"f6",
          7810 => x"fe",
          7811 => x"5d",
          7812 => x"3f",
          7813 => x"00",
          7814 => x"02",
          7815 => x"00",
          7816 => x"00",
          7817 => x"00",
          7818 => x"00",
          7819 => x"00",
          7820 => x"00",
          7821 => x"00",
          7822 => x"00",
          7823 => x"00",
          7824 => x"00",
          7825 => x"00",
          7826 => x"00",
          7827 => x"23",
          7828 => x"00",
          7829 => x"25",
          7830 => x"25",
          7831 => x"25",
          7832 => x"25",
          7833 => x"25",
          7834 => x"25",
          7835 => x"25",
          7836 => x"25",
          7837 => x"25",
          7838 => x"25",
          7839 => x"25",
          7840 => x"25",
          7841 => x"00",
          7842 => x"03",
          7843 => x"03",
          7844 => x"03",
          7845 => x"00",
          7846 => x"23",
          7847 => x"22",
          7848 => x"00",
          7849 => x"03",
          7850 => x"03",
          7851 => x"01",
          7852 => x"01",
          7853 => x"01",
          7854 => x"02",
          7855 => x"01",
          7856 => x"01",
          7857 => x"01",
          7858 => x"01",
          7859 => x"01",
          7860 => x"01",
          7861 => x"01",
          7862 => x"01",
          7863 => x"01",
          7864 => x"01",
          7865 => x"01",
          7866 => x"01",
          7867 => x"01",
          7868 => x"01",
          7869 => x"01",
          7870 => x"01",
          7871 => x"01",
          7872 => x"01",
          7873 => x"01",
          7874 => x"00",
          7875 => x"01",
          7876 => x"01",
          7877 => x"01",
          7878 => x"02",
          7879 => x"02",
          7880 => x"02",
          7881 => x"01",
          7882 => x"01",
          7883 => x"01",
          7884 => x"02",
          7885 => x"01",
          7886 => x"02",
          7887 => x"2c",
          7888 => x"01",
          7889 => x"02",
          7890 => x"02",
          7891 => x"02",
          7892 => x"02",
          7893 => x"01",
          7894 => x"02",
          7895 => x"01",
          7896 => x"02",
          7897 => x"03",
          7898 => x"03",
          7899 => x"03",
          7900 => x"03",
          7901 => x"03",
          7902 => x"00",
          7903 => x"03",
          7904 => x"03",
          7905 => x"03",
          7906 => x"03",
          7907 => x"04",
          7908 => x"04",
          7909 => x"04",
          7910 => x"01",
          7911 => x"00",
          7912 => x"1e",
          7913 => x"1f",
          7914 => x"1f",
          7915 => x"1f",
          7916 => x"1f",
          7917 => x"1f",
          7918 => x"06",
          7919 => x"1f",
          7920 => x"1f",
          7921 => x"1f",
          7922 => x"1f",
          7923 => x"06",
          7924 => x"00",
          7925 => x"1f",
          7926 => x"1f",
          7927 => x"1f",
          7928 => x"00",
          7929 => x"21",
          7930 => x"00",
          7931 => x"2c",
          7932 => x"2c",
          7933 => x"2c",
          7934 => x"ff",
          7935 => x"00",
          7936 => x"01",
          7937 => x"00",
          7938 => x"01",
          7939 => x"00",
          7940 => x"03",
          7941 => x"00",
          7942 => x"03",
          7943 => x"00",
          7944 => x"03",
          7945 => x"00",
          7946 => x"04",
          7947 => x"00",
          7948 => x"04",
          7949 => x"00",
          7950 => x"04",
          7951 => x"00",
          7952 => x"04",
          7953 => x"00",
          7954 => x"04",
          7955 => x"00",
          7956 => x"04",
          7957 => x"00",
          7958 => x"04",
          7959 => x"00",
          7960 => x"05",
          7961 => x"00",
          7962 => x"05",
          7963 => x"00",
          7964 => x"05",
          7965 => x"00",
          7966 => x"05",
          7967 => x"00",
          7968 => x"07",
          7969 => x"00",
          7970 => x"07",
          7971 => x"00",
          7972 => x"08",
          7973 => x"00",
          7974 => x"08",
          7975 => x"00",
          7976 => x"08",
          7977 => x"00",
          7978 => x"08",
          7979 => x"00",
          7980 => x"08",
          7981 => x"00",
          7982 => x"08",
          7983 => x"00",
          7984 => x"09",
          7985 => x"00",
          7986 => x"09",
          7987 => x"00",
          7988 => x"09",
          7989 => x"00",
          7990 => x"09",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"00",
          7996 => x"00",
          7997 => x"00",
          7998 => x"78",
          7999 => x"e1",
          8000 => x"e1",
          8001 => x"01",
          8002 => x"10",
          8003 => x"00",
          8004 => x"00",
          8005 => x"00",
          8006 => x"00",
          8007 => x"00",
          8008 => x"00",
          8009 => x"00",
          8010 => x"00",
          8011 => x"00",
          8012 => x"00",
          8013 => x"00",
          8014 => x"00",
          8015 => x"f1",
          8016 => x"f1",
          8017 => x"f1",
          8018 => x"fd",
          8019 => x"3a",
          8020 => x"f0",
          8021 => x"77",
          8022 => x"6f",
          8023 => x"67",
          8024 => x"37",
          8025 => x"2c",
          8026 => x"3f",
          8027 => x"f0",
          8028 => x"f0",
          8029 => x"3b",
          8030 => x"f0",
          8031 => x"57",
          8032 => x"4f",
          8033 => x"47",
          8034 => x"37",
          8035 => x"2c",
          8036 => x"3f",
          8037 => x"f0",
          8038 => x"f0",
          8039 => x"2a",
          8040 => x"f0",
          8041 => x"57",
          8042 => x"4f",
          8043 => x"47",
          8044 => x"27",
          8045 => x"3c",
          8046 => x"3f",
          8047 => x"f0",
          8048 => x"f0",
          8049 => x"f0",
          8050 => x"f0",
          8051 => x"17",
          8052 => x"0f",
          8053 => x"07",
          8054 => x"f0",
          8055 => x"f0",
          8056 => x"f0",
          8057 => x"f0",
          8058 => x"f0",
          8059 => x"4d",
          8060 => x"f0",
          8061 => x"78",
          8062 => x"d5",
          8063 => x"4c",
          8064 => x"5f",
          8065 => x"d0",
          8066 => x"bb",
          8067 => x"f0",
          8068 => x"f0",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"01",
          9104 => x"f2",
          9105 => x"fa",
          9106 => x"c2",
          9107 => x"e5",
          9108 => x"62",
          9109 => x"6b",
          9110 => x"22",
          9111 => x"4f",
          9112 => x"02",
          9113 => x"0a",
          9114 => x"12",
          9115 => x"1a",
          9116 => x"82",
          9117 => x"8a",
          9118 => x"92",
          9119 => x"9a",
          9120 => x"00",
          9121 => x"00",
          9122 => x"00",
          9123 => x"00",
          9124 => x"00",
          9125 => x"00",
          9126 => x"00",
          9127 => x"00",
          9128 => x"00",
          9129 => x"00",
          9130 => x"00",
          9131 => x"00",
          9132 => x"00",
          9133 => x"00",
          9134 => x"00",
          9135 => x"00",
          9136 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"93",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"2d",
             6 => x"00",
             7 => x"00",
             8 => x"fd",
             9 => x"05",
            10 => x"ff",
            11 => x"00",
            12 => x"fd",
            13 => x"06",
            14 => x"2b",
            15 => x"0b",
            16 => x"09",
            17 => x"06",
            18 => x"0a",
            19 => x"00",
            20 => x"72",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"73",
            25 => x"81",
            26 => x"10",
            27 => x"51",
            28 => x"72",
            29 => x"04",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"0a",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"72",
            45 => x"0b",
            46 => x"00",
            47 => x"00",
            48 => x"72",
            49 => x"74",
            50 => x"07",
            51 => x"00",
            52 => x"71",
            53 => x"09",
            54 => x"2b",
            55 => x"04",
            56 => x"09",
            57 => x"05",
            58 => x"04",
            59 => x"00",
            60 => x"09",
            61 => x"05",
            62 => x"51",
            63 => x"00",
            64 => x"09",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"72",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"09",
            73 => x"53",
            74 => x"00",
            75 => x"00",
            76 => x"fc",
            77 => x"05",
            78 => x"ff",
            79 => x"00",
            80 => x"fc",
            81 => x"73",
            82 => x"0b",
            83 => x"00",
            84 => x"08",
            85 => x"0b",
            86 => x"08",
            87 => x"51",
            88 => x"08",
            89 => x"0b",
            90 => x"08",
            91 => x"51",
            92 => x"09",
            93 => x"06",
            94 => x"09",
            95 => x"51",
            96 => x"09",
            97 => x"81",
            98 => x"73",
            99 => x"07",
           100 => x"ff",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"81",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"84",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"0d",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"8c",
           134 => x"04",
           135 => x"0b",
           136 => x"8c",
           137 => x"04",
           138 => x"0b",
           139 => x"8d",
           140 => x"04",
           141 => x"0b",
           142 => x"8d",
           143 => x"04",
           144 => x"0b",
           145 => x"8e",
           146 => x"04",
           147 => x"0b",
           148 => x"8e",
           149 => x"04",
           150 => x"0b",
           151 => x"8f",
           152 => x"04",
           153 => x"0b",
           154 => x"8f",
           155 => x"04",
           156 => x"0b",
           157 => x"90",
           158 => x"04",
           159 => x"0b",
           160 => x"90",
           161 => x"04",
           162 => x"0b",
           163 => x"91",
           164 => x"04",
           165 => x"0b",
           166 => x"91",
           167 => x"04",
           168 => x"0b",
           169 => x"92",
           170 => x"04",
           171 => x"0b",
           172 => x"92",
           173 => x"04",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"00",
           193 => x"80",
           194 => x"80",
           195 => x"0c",
           196 => x"80",
           197 => x"0c",
           198 => x"80",
           199 => x"0c",
           200 => x"80",
           201 => x"0c",
           202 => x"80",
           203 => x"0c",
           204 => x"80",
           205 => x"0c",
           206 => x"80",
           207 => x"0c",
           208 => x"80",
           209 => x"0c",
           210 => x"80",
           211 => x"0c",
           212 => x"80",
           213 => x"0c",
           214 => x"80",
           215 => x"0c",
           216 => x"80",
           217 => x"0c",
           218 => x"08",
           219 => x"90",
           220 => x"90",
           221 => x"bb",
           222 => x"bb",
           223 => x"84",
           224 => x"84",
           225 => x"04",
           226 => x"2d",
           227 => x"90",
           228 => x"89",
           229 => x"80",
           230 => x"d4",
           231 => x"c0",
           232 => x"82",
           233 => x"80",
           234 => x"0c",
           235 => x"08",
           236 => x"90",
           237 => x"90",
           238 => x"bb",
           239 => x"bb",
           240 => x"84",
           241 => x"84",
           242 => x"04",
           243 => x"2d",
           244 => x"90",
           245 => x"b7",
           246 => x"80",
           247 => x"85",
           248 => x"c0",
           249 => x"82",
           250 => x"80",
           251 => x"0c",
           252 => x"08",
           253 => x"90",
           254 => x"90",
           255 => x"bb",
           256 => x"bb",
           257 => x"84",
           258 => x"84",
           259 => x"04",
           260 => x"2d",
           261 => x"90",
           262 => x"f0",
           263 => x"80",
           264 => x"e7",
           265 => x"c0",
           266 => x"82",
           267 => x"80",
           268 => x"0c",
           269 => x"08",
           270 => x"90",
           271 => x"90",
           272 => x"bb",
           273 => x"bb",
           274 => x"84",
           275 => x"84",
           276 => x"04",
           277 => x"2d",
           278 => x"90",
           279 => x"a2",
           280 => x"80",
           281 => x"b8",
           282 => x"c0",
           283 => x"81",
           284 => x"80",
           285 => x"0c",
           286 => x"08",
           287 => x"90",
           288 => x"90",
           289 => x"bb",
           290 => x"bb",
           291 => x"84",
           292 => x"84",
           293 => x"04",
           294 => x"2d",
           295 => x"90",
           296 => x"2d",
           297 => x"90",
           298 => x"c9",
           299 => x"80",
           300 => x"de",
           301 => x"c0",
           302 => x"81",
           303 => x"80",
           304 => x"0c",
           305 => x"08",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"51",
           311 => x"73",
           312 => x"10",
           313 => x"0c",
           314 => x"81",
           315 => x"71",
           316 => x"72",
           317 => x"84",
           318 => x"8e",
           319 => x"0c",
           320 => x"81",
           321 => x"3d",
           322 => x"52",
           323 => x"e8",
           324 => x"0d",
           325 => x"85",
           326 => x"73",
           327 => x"52",
           328 => x"d3",
           329 => x"70",
           330 => x"55",
           331 => x"38",
           332 => x"8e",
           333 => x"84",
           334 => x"84",
           335 => x"57",
           336 => x"30",
           337 => x"54",
           338 => x"75",
           339 => x"0c",
           340 => x"bb",
           341 => x"3d",
           342 => x"99",
           343 => x"8e",
           344 => x"3d",
           345 => x"54",
           346 => x"fd",
           347 => x"76",
           348 => x"0d",
           349 => x"42",
           350 => x"85",
           351 => x"81",
           352 => x"7b",
           353 => x"7b",
           354 => x"38",
           355 => x"72",
           356 => x"5f",
           357 => x"b0",
           358 => x"54",
           359 => x"a9",
           360 => x"81",
           361 => x"38",
           362 => x"57",
           363 => x"54",
           364 => x"0d",
           365 => x"10",
           366 => x"70",
           367 => x"29",
           368 => x"5a",
           369 => x"86",
           370 => x"bd",
           371 => x"fe",
           372 => x"2e",
           373 => x"74",
           374 => x"5a",
           375 => x"7c",
           376 => x"33",
           377 => x"39",
           378 => x"55",
           379 => x"40",
           380 => x"72",
           381 => x"10",
           382 => x"04",
           383 => x"73",
           384 => x"8a",
           385 => x"76",
           386 => x"ff",
           387 => x"60",
           388 => x"cf",
           389 => x"94",
           390 => x"3f",
           391 => x"84",
           392 => x"53",
           393 => x"84",
           394 => x"81",
           395 => x"90",
           396 => x"84",
           397 => x"bb",
           398 => x"40",
           399 => x"84",
           400 => x"70",
           401 => x"70",
           402 => x"9e",
           403 => x"80",
           404 => x"38",
           405 => x"80",
           406 => x"83",
           407 => x"80",
           408 => x"81",
           409 => x"86",
           410 => x"70",
           411 => x"5b",
           412 => x"85",
           413 => x"70",
           414 => x"59",
           415 => x"7a",
           416 => x"eb",
           417 => x"73",
           418 => x"06",
           419 => x"06",
           420 => x"2a",
           421 => x"38",
           422 => x"80",
           423 => x"54",
           424 => x"b0",
           425 => x"80",
           426 => x"90",
           427 => x"e5",
           428 => x"2e",
           429 => x"29",
           430 => x"5b",
           431 => x"7c",
           432 => x"79",
           433 => x"05",
           434 => x"80",
           435 => x"81",
           436 => x"b9",
           437 => x"38",
           438 => x"76",
           439 => x"84",
           440 => x"ff",
           441 => x"3f",
           442 => x"06",
           443 => x"80",
           444 => x"80",
           445 => x"90",
           446 => x"fc",
           447 => x"f4",
           448 => x"7a",
           449 => x"fa",
           450 => x"c0",
           451 => x"61",
           452 => x"cf",
           453 => x"fd",
           454 => x"80",
           455 => x"2b",
           456 => x"fc",
           457 => x"52",
           458 => x"2a",
           459 => x"c9",
           460 => x"fc",
           461 => x"54",
           462 => x"7c",
           463 => x"39",
           464 => x"5b",
           465 => x"ca",
           466 => x"57",
           467 => x"ff",
           468 => x"54",
           469 => x"38",
           470 => x"33",
           471 => x"fc",
           472 => x"84",
           473 => x"70",
           474 => x"7b",
           475 => x"57",
           476 => x"7f",
           477 => x"40",
           478 => x"38",
           479 => x"bb",
           480 => x"07",
           481 => x"38",
           482 => x"80",
           483 => x"38",
           484 => x"71",
           485 => x"5f",
           486 => x"f6",
           487 => x"ff",
           488 => x"5a",
           489 => x"7a",
           490 => x"76",
           491 => x"60",
           492 => x"5d",
           493 => x"75",
           494 => x"08",
           495 => x"90",
           496 => x"80",
           497 => x"88",
           498 => x"80",
           499 => x"90",
           500 => x"fa",
           501 => x"c4",
           502 => x"83",
           503 => x"06",
           504 => x"83",
           505 => x"5f",
           506 => x"d8",
           507 => x"90",
           508 => x"06",
           509 => x"38",
           510 => x"82",
           511 => x"80",
           512 => x"7c",
           513 => x"3f",
           514 => x"f7",
           515 => x"31",
           516 => x"f9",
           517 => x"c4",
           518 => x"82",
           519 => x"75",
           520 => x"08",
           521 => x"90",
           522 => x"82",
           523 => x"06",
           524 => x"3d",
           525 => x"52",
           526 => x"0d",
           527 => x"0b",
           528 => x"70",
           529 => x"51",
           530 => x"77",
           531 => x"74",
           532 => x"77",
           533 => x"52",
           534 => x"2d",
           535 => x"38",
           536 => x"33",
           537 => x"e6",
           538 => x"e8",
           539 => x"8a",
           540 => x"84",
           541 => x"ff",
           542 => x"0c",
           543 => x"78",
           544 => x"33",
           545 => x"06",
           546 => x"77",
           547 => x"70",
           548 => x"2e",
           549 => x"75",
           550 => x"04",
           551 => x"72",
           552 => x"51",
           553 => x"bb",
           554 => x"74",
           555 => x"72",
           556 => x"84",
           557 => x"3f",
           558 => x"78",
           559 => x"81",
           560 => x"ff",
           561 => x"81",
           562 => x"8c",
           563 => x"25",
           564 => x"34",
           565 => x"15",
           566 => x"76",
           567 => x"3d",
           568 => x"06",
           569 => x"ff",
           570 => x"8c",
           571 => x"76",
           572 => x"85",
           573 => x"81",
           574 => x"ff",
           575 => x"81",
           576 => x"2a",
           577 => x"c3",
           578 => x"71",
           579 => x"76",
           580 => x"17",
           581 => x"84",
           582 => x"74",
           583 => x"34",
           584 => x"0c",
           585 => x"87",
           586 => x"08",
           587 => x"52",
           588 => x"b9",
           589 => x"54",
           590 => x"85",
           591 => x"17",
           592 => x"0c",
           593 => x"53",
           594 => x"39",
           595 => x"54",
           596 => x"51",
           597 => x"70",
           598 => x"70",
           599 => x"73",
           600 => x"04",
           601 => x"55",
           602 => x"38",
           603 => x"2e",
           604 => x"33",
           605 => x"11",
           606 => x"84",
           607 => x"55",
           608 => x"75",
           609 => x"53",
           610 => x"70",
           611 => x"13",
           612 => x"11",
           613 => x"3d",
           614 => x"81",
           615 => x"ff",
           616 => x"0c",
           617 => x"0d",
           618 => x"70",
           619 => x"70",
           620 => x"73",
           621 => x"04",
           622 => x"55",
           623 => x"38",
           624 => x"70",
           625 => x"70",
           626 => x"85",
           627 => x"78",
           628 => x"a1",
           629 => x"57",
           630 => x"81",
           631 => x"80",
           632 => x"e1",
           633 => x"0c",
           634 => x"f1",
           635 => x"80",
           636 => x"81",
           637 => x"72",
           638 => x"0d",
           639 => x"3d",
           640 => x"53",
           641 => x"bb",
           642 => x"05",
           643 => x"bb",
           644 => x"80",
           645 => x"15",
           646 => x"52",
           647 => x"3f",
           648 => x"bb",
           649 => x"3d",
           650 => x"53",
           651 => x"70",
           652 => x"2e",
           653 => x"2e",
           654 => x"70",
           655 => x"84",
           656 => x"0d",
           657 => x"54",
           658 => x"70",
           659 => x"70",
           660 => x"85",
           661 => x"7a",
           662 => x"8b",
           663 => x"bb",
           664 => x"80",
           665 => x"3f",
           666 => x"80",
           667 => x"73",
           668 => x"81",
           669 => x"76",
           670 => x"56",
           671 => x"74",
           672 => x"78",
           673 => x"81",
           674 => x"ff",
           675 => x"55",
           676 => x"07",
           677 => x"3d",
           678 => x"fc",
           679 => x"07",
           680 => x"31",
           681 => x"06",
           682 => x"88",
           683 => x"f0",
           684 => x"2b",
           685 => x"53",
           686 => x"30",
           687 => x"77",
           688 => x"70",
           689 => x"06",
           690 => x"51",
           691 => x"53",
           692 => x"56",
           693 => x"0d",
           694 => x"54",
           695 => x"84",
           696 => x"31",
           697 => x"0d",
           698 => x"54",
           699 => x"76",
           700 => x"08",
           701 => x"8d",
           702 => x"84",
           703 => x"71",
           704 => x"71",
           705 => x"71",
           706 => x"57",
           707 => x"2e",
           708 => x"07",
           709 => x"ff",
           710 => x"72",
           711 => x"56",
           712 => x"da",
           713 => x"3d",
           714 => x"2c",
           715 => x"32",
           716 => x"32",
           717 => x"56",
           718 => x"3f",
           719 => x"31",
           720 => x"04",
           721 => x"80",
           722 => x"56",
           723 => x"06",
           724 => x"70",
           725 => x"38",
           726 => x"b0",
           727 => x"80",
           728 => x"8a",
           729 => x"c4",
           730 => x"e0",
           731 => x"d0",
           732 => x"90",
           733 => x"81",
           734 => x"81",
           735 => x"38",
           736 => x"79",
           737 => x"a0",
           738 => x"84",
           739 => x"81",
           740 => x"3d",
           741 => x"0c",
           742 => x"2e",
           743 => x"15",
           744 => x"73",
           745 => x"73",
           746 => x"a0",
           747 => x"80",
           748 => x"e1",
           749 => x"3d",
           750 => x"78",
           751 => x"fe",
           752 => x"0c",
           753 => x"7b",
           754 => x"77",
           755 => x"a0",
           756 => x"15",
           757 => x"73",
           758 => x"80",
           759 => x"38",
           760 => x"26",
           761 => x"a0",
           762 => x"74",
           763 => x"ff",
           764 => x"ff",
           765 => x"38",
           766 => x"54",
           767 => x"78",
           768 => x"13",
           769 => x"56",
           770 => x"38",
           771 => x"56",
           772 => x"bb",
           773 => x"70",
           774 => x"56",
           775 => x"fe",
           776 => x"70",
           777 => x"a6",
           778 => x"a0",
           779 => x"38",
           780 => x"89",
           781 => x"bb",
           782 => x"58",
           783 => x"55",
           784 => x"0b",
           785 => x"04",
           786 => x"08",
           787 => x"04",
           788 => x"26",
           789 => x"94",
           790 => x"ac",
           791 => x"04",
           792 => x"83",
           793 => x"ef",
           794 => x"cf",
           795 => x"0d",
           796 => x"3f",
           797 => x"51",
           798 => x"83",
           799 => x"3d",
           800 => x"f1",
           801 => x"ec",
           802 => x"04",
           803 => x"83",
           804 => x"ee",
           805 => x"d1",
           806 => x"0d",
           807 => x"3f",
           808 => x"51",
           809 => x"83",
           810 => x"3d",
           811 => x"99",
           812 => x"98",
           813 => x"04",
           814 => x"83",
           815 => x"ed",
           816 => x"d2",
           817 => x"0d",
           818 => x"3f",
           819 => x"0d",
           820 => x"84",
           821 => x"81",
           822 => x"07",
           823 => x"57",
           824 => x"57",
           825 => x"51",
           826 => x"81",
           827 => x"58",
           828 => x"08",
           829 => x"80",
           830 => x"3f",
           831 => x"7b",
           832 => x"57",
           833 => x"87",
           834 => x"e7",
           835 => x"87",
           836 => x"bb",
           837 => x"78",
           838 => x"3f",
           839 => x"3d",
           840 => x"c0",
           841 => x"59",
           842 => x"84",
           843 => x"9f",
           844 => x"84",
           845 => x"55",
           846 => x"19",
           847 => x"e8",
           848 => x"bb",
           849 => x"3f",
           850 => x"84",
           851 => x"de",
           852 => x"0d",
           853 => x"58",
           854 => x"7a",
           855 => x"08",
           856 => x"76",
           857 => x"84",
           858 => x"84",
           859 => x"84",
           860 => x"78",
           861 => x"84",
           862 => x"0d",
           863 => x"cf",
           864 => x"5f",
           865 => x"2e",
           866 => x"8c",
           867 => x"51",
           868 => x"27",
           869 => x"38",
           870 => x"18",
           871 => x"72",
           872 => x"c6",
           873 => x"53",
           874 => x"74",
           875 => x"dd",
           876 => x"80",
           877 => x"53",
           878 => x"81",
           879 => x"38",
           880 => x"ff",
           881 => x"38",
           882 => x"84",
           883 => x"d4",
           884 => x"c2",
           885 => x"3f",
           886 => x"51",
           887 => x"98",
           888 => x"a0",
           889 => x"82",
           890 => x"26",
           891 => x"84",
           892 => x"a8",
           893 => x"e6",
           894 => x"fc",
           895 => x"fe",
           896 => x"86",
           897 => x"53",
           898 => x"79",
           899 => x"72",
           900 => x"83",
           901 => x"14",
           902 => x"51",
           903 => x"38",
           904 => x"db",
           905 => x"08",
           906 => x"73",
           907 => x"53",
           908 => x"52",
           909 => x"84",
           910 => x"a0",
           911 => x"dd",
           912 => x"08",
           913 => x"16",
           914 => x"3f",
           915 => x"53",
           916 => x"38",
           917 => x"81",
           918 => x"db",
           919 => x"bb",
           920 => x"70",
           921 => x"70",
           922 => x"06",
           923 => x"72",
           924 => x"9b",
           925 => x"2b",
           926 => x"30",
           927 => x"07",
           928 => x"59",
           929 => x"a9",
           930 => x"bb",
           931 => x"3d",
           932 => x"aa",
           933 => x"83",
           934 => x"51",
           935 => x"81",
           936 => x"72",
           937 => x"71",
           938 => x"81",
           939 => x"72",
           940 => x"71",
           941 => x"81",
           942 => x"72",
           943 => x"71",
           944 => x"81",
           945 => x"88",
           946 => x"a9",
           947 => x"51",
           948 => x"9c",
           949 => x"a9",
           950 => x"51",
           951 => x"9c",
           952 => x"72",
           953 => x"2e",
           954 => x"e3",
           955 => x"3f",
           956 => x"2a",
           957 => x"2e",
           958 => x"9b",
           959 => x"d3",
           960 => x"86",
           961 => x"80",
           962 => x"81",
           963 => x"51",
           964 => x"3f",
           965 => x"52",
           966 => x"bd",
           967 => x"d5",
           968 => x"9a",
           969 => x"06",
           970 => x"38",
           971 => x"3f",
           972 => x"80",
           973 => x"70",
           974 => x"fd",
           975 => x"9a",
           976 => x"cb",
           977 => x"82",
           978 => x"80",
           979 => x"ca",
           980 => x"61",
           981 => x"60",
           982 => x"84",
           983 => x"59",
           984 => x"d6",
           985 => x"43",
           986 => x"7e",
           987 => x"51",
           988 => x"f8",
           989 => x"79",
           990 => x"2e",
           991 => x"5e",
           992 => x"70",
           993 => x"38",
           994 => x"81",
           995 => x"5d",
           996 => x"5c",
           997 => x"29",
           998 => x"5b",
           999 => x"84",
          1000 => x"08",
          1001 => x"84",
          1002 => x"7d",
          1003 => x"70",
          1004 => x"27",
          1005 => x"80",
          1006 => x"7e",
          1007 => x"08",
          1008 => x"8d",
          1009 => x"b8",
          1010 => x"3f",
          1011 => x"5c",
          1012 => x"84",
          1013 => x"84",
          1014 => x"38",
          1015 => x"82",
          1016 => x"8c",
          1017 => x"38",
          1018 => x"52",
          1019 => x"c0",
          1020 => x"67",
          1021 => x"90",
          1022 => x"3f",
          1023 => x"08",
          1024 => x"25",
          1025 => x"83",
          1026 => x"06",
          1027 => x"1b",
          1028 => x"ff",
          1029 => x"32",
          1030 => x"ff",
          1031 => x"96",
          1032 => x"c6",
          1033 => x"52",
          1034 => x"83",
          1035 => x"5b",
          1036 => x"83",
          1037 => x"82",
          1038 => x"80",
          1039 => x"ef",
          1040 => x"f8",
          1041 => x"84",
          1042 => x"84",
          1043 => x"0b",
          1044 => x"ff",
          1045 => x"81",
          1046 => x"de",
          1047 => x"0b",
          1048 => x"55",
          1049 => x"f8",
          1050 => x"70",
          1051 => x"39",
          1052 => x"59",
          1053 => x"78",
          1054 => x"79",
          1055 => x"52",
          1056 => x"7e",
          1057 => x"bd",
          1058 => x"09",
          1059 => x"9a",
          1060 => x"83",
          1061 => x"51",
          1062 => x"83",
          1063 => x"a0",
          1064 => x"7c",
          1065 => x"81",
          1066 => x"f9",
          1067 => x"51",
          1068 => x"81",
          1069 => x"d7",
          1070 => x"78",
          1071 => x"3f",
          1072 => x"3d",
          1073 => x"51",
          1074 => x"80",
          1075 => x"d7",
          1076 => x"79",
          1077 => x"fa",
          1078 => x"83",
          1079 => x"90",
          1080 => x"ff",
          1081 => x"bb",
          1082 => x"68",
          1083 => x"3f",
          1084 => x"f4",
          1085 => x"98",
          1086 => x"f9",
          1087 => x"53",
          1088 => x"84",
          1089 => x"59",
          1090 => x"b8",
          1091 => x"08",
          1092 => x"81",
          1093 => x"ae",
          1094 => x"87",
          1095 => x"59",
          1096 => x"53",
          1097 => x"84",
          1098 => x"38",
          1099 => x"80",
          1100 => x"84",
          1101 => x"22",
          1102 => x"cf",
          1103 => x"80",
          1104 => x"7e",
          1105 => x"f8",
          1106 => x"38",
          1107 => x"39",
          1108 => x"80",
          1109 => x"84",
          1110 => x"3d",
          1111 => x"51",
          1112 => x"80",
          1113 => x"f8",
          1114 => x"b4",
          1115 => x"f7",
          1116 => x"a6",
          1117 => x"27",
          1118 => x"33",
          1119 => x"38",
          1120 => x"78",
          1121 => x"3f",
          1122 => x"1b",
          1123 => x"84",
          1124 => x"e4",
          1125 => x"f7",
          1126 => x"53",
          1127 => x"84",
          1128 => x"38",
          1129 => x"80",
          1130 => x"84",
          1131 => x"d9",
          1132 => x"79",
          1133 => x"79",
          1134 => x"65",
          1135 => x"ff",
          1136 => x"e8",
          1137 => x"2e",
          1138 => x"11",
          1139 => x"3f",
          1140 => x"70",
          1141 => x"cc",
          1142 => x"80",
          1143 => x"7e",
          1144 => x"f6",
          1145 => x"38",
          1146 => x"59",
          1147 => x"68",
          1148 => x"11",
          1149 => x"3f",
          1150 => x"d8",
          1151 => x"33",
          1152 => x"3d",
          1153 => x"51",
          1154 => x"ff",
          1155 => x"ff",
          1156 => x"e6",
          1157 => x"2e",
          1158 => x"11",
          1159 => x"3f",
          1160 => x"88",
          1161 => x"ff",
          1162 => x"bb",
          1163 => x"08",
          1164 => x"3f",
          1165 => x"8f",
          1166 => x"05",
          1167 => x"8a",
          1168 => x"b8",
          1169 => x"3f",
          1170 => x"80",
          1171 => x"53",
          1172 => x"e9",
          1173 => x"2e",
          1174 => x"51",
          1175 => x"3d",
          1176 => x"51",
          1177 => x"91",
          1178 => x"80",
          1179 => x"08",
          1180 => x"ff",
          1181 => x"bb",
          1182 => x"33",
          1183 => x"83",
          1184 => x"f8",
          1185 => x"fc",
          1186 => x"a5",
          1187 => x"2e",
          1188 => x"70",
          1189 => x"06",
          1190 => x"38",
          1191 => x"83",
          1192 => x"55",
          1193 => x"51",
          1194 => x"d6",
          1195 => x"71",
          1196 => x"3d",
          1197 => x"51",
          1198 => x"80",
          1199 => x"0c",
          1200 => x"fe",
          1201 => x"e1",
          1202 => x"38",
          1203 => x"ce",
          1204 => x"23",
          1205 => x"53",
          1206 => x"84",
          1207 => x"38",
          1208 => x"7e",
          1209 => x"b8",
          1210 => x"05",
          1211 => x"08",
          1212 => x"3d",
          1213 => x"51",
          1214 => x"80",
          1215 => x"80",
          1216 => x"05",
          1217 => x"f0",
          1218 => x"f0",
          1219 => x"81",
          1220 => x"64",
          1221 => x"39",
          1222 => x"98",
          1223 => x"80",
          1224 => x"c8",
          1225 => x"7c",
          1226 => x"83",
          1227 => x"f0",
          1228 => x"ff",
          1229 => x"bb",
          1230 => x"59",
          1231 => x"82",
          1232 => x"39",
          1233 => x"2e",
          1234 => x"47",
          1235 => x"5c",
          1236 => x"c8",
          1237 => x"f8",
          1238 => x"b6",
          1239 => x"3f",
          1240 => x"8a",
          1241 => x"83",
          1242 => x"83",
          1243 => x"c6",
          1244 => x"80",
          1245 => x"47",
          1246 => x"5e",
          1247 => x"d8",
          1248 => x"8b",
          1249 => x"83",
          1250 => x"83",
          1251 => x"9b",
          1252 => x"b9",
          1253 => x"80",
          1254 => x"47",
          1255 => x"fc",
          1256 => x"f3",
          1257 => x"39",
          1258 => x"b4",
          1259 => x"56",
          1260 => x"da",
          1261 => x"2b",
          1262 => x"52",
          1263 => x"bb",
          1264 => x"94",
          1265 => x"80",
          1266 => x"bb",
          1267 => x"55",
          1268 => x"83",
          1269 => x"77",
          1270 => x"94",
          1271 => x"c0",
          1272 => x"81",
          1273 => x"a1",
          1274 => x"0b",
          1275 => x"72",
          1276 => x"bd",
          1277 => x"ba",
          1278 => x"c0",
          1279 => x"3f",
          1280 => x"94",
          1281 => x"d3",
          1282 => x"d3",
          1283 => x"3f",
          1284 => x"80",
          1285 => x"3f",
          1286 => x"51",
          1287 => x"04",
          1288 => x"56",
          1289 => x"81",
          1290 => x"06",
          1291 => x"06",
          1292 => x"81",
          1293 => x"2e",
          1294 => x"73",
          1295 => x"72",
          1296 => x"33",
          1297 => x"70",
          1298 => x"80",
          1299 => x"38",
          1300 => x"81",
          1301 => x"09",
          1302 => x"a2",
          1303 => x"07",
          1304 => x"38",
          1305 => x"71",
          1306 => x"84",
          1307 => x"2e",
          1308 => x"38",
          1309 => x"81",
          1310 => x"2e",
          1311 => x"15",
          1312 => x"2e",
          1313 => x"39",
          1314 => x"8b",
          1315 => x"86",
          1316 => x"52",
          1317 => x"84",
          1318 => x"bb",
          1319 => x"3d",
          1320 => x"52",
          1321 => x"98",
          1322 => x"82",
          1323 => x"84",
          1324 => x"26",
          1325 => x"84",
          1326 => x"86",
          1327 => x"26",
          1328 => x"86",
          1329 => x"38",
          1330 => x"87",
          1331 => x"87",
          1332 => x"c0",
          1333 => x"c0",
          1334 => x"c0",
          1335 => x"c0",
          1336 => x"c0",
          1337 => x"c0",
          1338 => x"a4",
          1339 => x"80",
          1340 => x"52",
          1341 => x"0d",
          1342 => x"c0",
          1343 => x"c0",
          1344 => x"87",
          1345 => x"1c",
          1346 => x"79",
          1347 => x"08",
          1348 => x"98",
          1349 => x"87",
          1350 => x"1c",
          1351 => x"7b",
          1352 => x"08",
          1353 => x"0c",
          1354 => x"83",
          1355 => x"57",
          1356 => x"55",
          1357 => x"53",
          1358 => x"d9",
          1359 => x"3d",
          1360 => x"05",
          1361 => x"72",
          1362 => x"84",
          1363 => x"52",
          1364 => x"38",
          1365 => x"bb",
          1366 => x"51",
          1367 => x"08",
          1368 => x"71",
          1369 => x"72",
          1370 => x"84",
          1371 => x"52",
          1372 => x"fd",
          1373 => x"88",
          1374 => x"3f",
          1375 => x"98",
          1376 => x"38",
          1377 => x"83",
          1378 => x"84",
          1379 => x"0d",
          1380 => x"33",
          1381 => x"70",
          1382 => x"94",
          1383 => x"06",
          1384 => x"38",
          1385 => x"51",
          1386 => x"06",
          1387 => x"93",
          1388 => x"73",
          1389 => x"80",
          1390 => x"c0",
          1391 => x"84",
          1392 => x"71",
          1393 => x"70",
          1394 => x"53",
          1395 => x"2a",
          1396 => x"38",
          1397 => x"2a",
          1398 => x"cf",
          1399 => x"8f",
          1400 => x"51",
          1401 => x"83",
          1402 => x"55",
          1403 => x"70",
          1404 => x"83",
          1405 => x"54",
          1406 => x"38",
          1407 => x"2a",
          1408 => x"80",
          1409 => x"81",
          1410 => x"81",
          1411 => x"8a",
          1412 => x"71",
          1413 => x"87",
          1414 => x"86",
          1415 => x"72",
          1416 => x"73",
          1417 => x"0c",
          1418 => x"70",
          1419 => x"72",
          1420 => x"2e",
          1421 => x"52",
          1422 => x"c0",
          1423 => x"81",
          1424 => x"d7",
          1425 => x"80",
          1426 => x"52",
          1427 => x"c0",
          1428 => x"87",
          1429 => x"0c",
          1430 => x"c8",
          1431 => x"f3",
          1432 => x"83",
          1433 => x"08",
          1434 => x"ac",
          1435 => x"9e",
          1436 => x"c0",
          1437 => x"87",
          1438 => x"0c",
          1439 => x"e8",
          1440 => x"f3",
          1441 => x"83",
          1442 => x"08",
          1443 => x"c0",
          1444 => x"87",
          1445 => x"0c",
          1446 => x"80",
          1447 => x"80",
          1448 => x"84",
          1449 => x"82",
          1450 => x"80",
          1451 => x"88",
          1452 => x"80",
          1453 => x"f4",
          1454 => x"90",
          1455 => x"52",
          1456 => x"52",
          1457 => x"87",
          1458 => x"80",
          1459 => x"83",
          1460 => x"34",
          1461 => x"70",
          1462 => x"70",
          1463 => x"83",
          1464 => x"9e",
          1465 => x"51",
          1466 => x"81",
          1467 => x"0b",
          1468 => x"80",
          1469 => x"2e",
          1470 => x"8b",
          1471 => x"08",
          1472 => x"52",
          1473 => x"71",
          1474 => x"c0",
          1475 => x"06",
          1476 => x"38",
          1477 => x"80",
          1478 => x"80",
          1479 => x"80",
          1480 => x"f4",
          1481 => x"90",
          1482 => x"52",
          1483 => x"71",
          1484 => x"90",
          1485 => x"53",
          1486 => x"0b",
          1487 => x"80",
          1488 => x"83",
          1489 => x"34",
          1490 => x"06",
          1491 => x"f4",
          1492 => x"90",
          1493 => x"70",
          1494 => x"83",
          1495 => x"08",
          1496 => x"34",
          1497 => x"82",
          1498 => x"51",
          1499 => x"33",
          1500 => x"a8",
          1501 => x"33",
          1502 => x"8b",
          1503 => x"f4",
          1504 => x"83",
          1505 => x"38",
          1506 => x"cc",
          1507 => x"84",
          1508 => x"73",
          1509 => x"55",
          1510 => x"33",
          1511 => x"87",
          1512 => x"f4",
          1513 => x"83",
          1514 => x"38",
          1515 => x"e1",
          1516 => x"3f",
          1517 => x"cc",
          1518 => x"ec",
          1519 => x"b5",
          1520 => x"83",
          1521 => x"83",
          1522 => x"f3",
          1523 => x"ff",
          1524 => x"56",
          1525 => x"fb",
          1526 => x"c0",
          1527 => x"bb",
          1528 => x"ff",
          1529 => x"55",
          1530 => x"55",
          1531 => x"83",
          1532 => x"52",
          1533 => x"84",
          1534 => x"31",
          1535 => x"83",
          1536 => x"87",
          1537 => x"56",
          1538 => x"93",
          1539 => x"c0",
          1540 => x"bb",
          1541 => x"ff",
          1542 => x"55",
          1543 => x"9f",
          1544 => x"3f",
          1545 => x"83",
          1546 => x"51",
          1547 => x"08",
          1548 => x"a6",
          1549 => x"db",
          1550 => x"db",
          1551 => x"f3",
          1552 => x"ff",
          1553 => x"56",
          1554 => x"93",
          1555 => x"c0",
          1556 => x"bb",
          1557 => x"ff",
          1558 => x"55",
          1559 => x"cb",
          1560 => x"b1",
          1561 => x"80",
          1562 => x"83",
          1563 => x"83",
          1564 => x"fc",
          1565 => x"51",
          1566 => x"33",
          1567 => x"d7",
          1568 => x"f1",
          1569 => x"80",
          1570 => x"f4",
          1571 => x"ff",
          1572 => x"56",
          1573 => x"39",
          1574 => x"d4",
          1575 => x"91",
          1576 => x"38",
          1577 => x"83",
          1578 => x"83",
          1579 => x"fb",
          1580 => x"08",
          1581 => x"83",
          1582 => x"83",
          1583 => x"fb",
          1584 => x"08",
          1585 => x"83",
          1586 => x"83",
          1587 => x"fa",
          1588 => x"08",
          1589 => x"83",
          1590 => x"83",
          1591 => x"fa",
          1592 => x"08",
          1593 => x"83",
          1594 => x"83",
          1595 => x"fa",
          1596 => x"08",
          1597 => x"83",
          1598 => x"83",
          1599 => x"f9",
          1600 => x"51",
          1601 => x"51",
          1602 => x"33",
          1603 => x"c4",
          1604 => x"33",
          1605 => x"10",
          1606 => x"08",
          1607 => x"ce",
          1608 => x"bc",
          1609 => x"0d",
          1610 => x"b6",
          1611 => x"cc",
          1612 => x"0d",
          1613 => x"9e",
          1614 => x"dc",
          1615 => x"0d",
          1616 => x"0b",
          1617 => x"f4",
          1618 => x"04",
          1619 => x"3d",
          1620 => x"80",
          1621 => x"87",
          1622 => x"ed",
          1623 => x"f4",
          1624 => x"76",
          1625 => x"84",
          1626 => x"c0",
          1627 => x"17",
          1628 => x"08",
          1629 => x"ff",
          1630 => x"34",
          1631 => x"9f",
          1632 => x"85",
          1633 => x"ec",
          1634 => x"87",
          1635 => x"38",
          1636 => x"bb",
          1637 => x"e3",
          1638 => x"76",
          1639 => x"52",
          1640 => x"ff",
          1641 => x"84",
          1642 => x"83",
          1643 => x"80",
          1644 => x"0d",
          1645 => x"ad",
          1646 => x"57",
          1647 => x"92",
          1648 => x"75",
          1649 => x"70",
          1650 => x"84",
          1651 => x"08",
          1652 => x"84",
          1653 => x"73",
          1654 => x"2e",
          1655 => x"06",
          1656 => x"80",
          1657 => x"3d",
          1658 => x"ff",
          1659 => x"c7",
          1660 => x"2e",
          1661 => x"76",
          1662 => x"08",
          1663 => x"c9",
          1664 => x"57",
          1665 => x"ff",
          1666 => x"76",
          1667 => x"70",
          1668 => x"2e",
          1669 => x"75",
          1670 => x"59",
          1671 => x"84",
          1672 => x"56",
          1673 => x"08",
          1674 => x"53",
          1675 => x"fa",
          1676 => x"ba",
          1677 => x"84",
          1678 => x"bb",
          1679 => x"84",
          1680 => x"80",
          1681 => x"16",
          1682 => x"f6",
          1683 => x"ff",
          1684 => x"0c",
          1685 => x"b6",
          1686 => x"08",
          1687 => x"5b",
          1688 => x"34",
          1689 => x"f4",
          1690 => x"74",
          1691 => x"56",
          1692 => x"77",
          1693 => x"78",
          1694 => x"77",
          1695 => x"b5",
          1696 => x"3f",
          1697 => x"98",
          1698 => x"d7",
          1699 => x"c0",
          1700 => x"84",
          1701 => x"97",
          1702 => x"10",
          1703 => x"70",
          1704 => x"5b",
          1705 => x"2e",
          1706 => x"a8",
          1707 => x"ff",
          1708 => x"80",
          1709 => x"16",
          1710 => x"83",
          1711 => x"62",
          1712 => x"08",
          1713 => x"2e",
          1714 => x"38",
          1715 => x"76",
          1716 => x"70",
          1717 => x"bc",
          1718 => x"71",
          1719 => x"df",
          1720 => x"58",
          1721 => x"b1",
          1722 => x"51",
          1723 => x"98",
          1724 => x"ff",
          1725 => x"7d",
          1726 => x"fe",
          1727 => x"38",
          1728 => x"0a",
          1729 => x"06",
          1730 => x"c0",
          1731 => x"51",
          1732 => x"33",
          1733 => x"83",
          1734 => x"43",
          1735 => x"76",
          1736 => x"39",
          1737 => x"38",
          1738 => x"39",
          1739 => x"84",
          1740 => x"34",
          1741 => x"55",
          1742 => x"10",
          1743 => x"08",
          1744 => x"0c",
          1745 => x"0b",
          1746 => x"e2",
          1747 => x"e3",
          1748 => x"51",
          1749 => x"33",
          1750 => x"34",
          1751 => x"70",
          1752 => x"5a",
          1753 => x"38",
          1754 => x"42",
          1755 => x"70",
          1756 => x"fc",
          1757 => x"38",
          1758 => x"10",
          1759 => x"58",
          1760 => x"e2",
          1761 => x"c4",
          1762 => x"74",
          1763 => x"08",
          1764 => x"84",
          1765 => x"b4",
          1766 => x"88",
          1767 => x"c8",
          1768 => x"c8",
          1769 => x"cc",
          1770 => x"75",
          1771 => x"7c",
          1772 => x"75",
          1773 => x"ff",
          1774 => x"38",
          1775 => x"70",
          1776 => x"7c",
          1777 => x"10",
          1778 => x"59",
          1779 => x"51",
          1780 => x"08",
          1781 => x"08",
          1782 => x"52",
          1783 => x"e2",
          1784 => x"56",
          1785 => x"e6",
          1786 => x"9c",
          1787 => x"51",
          1788 => x"08",
          1789 => x"84",
          1790 => x"84",
          1791 => x"55",
          1792 => x"81",
          1793 => x"57",
          1794 => x"84",
          1795 => x"76",
          1796 => x"33",
          1797 => x"e2",
          1798 => x"e2",
          1799 => x"27",
          1800 => x"52",
          1801 => x"34",
          1802 => x"b2",
          1803 => x"81",
          1804 => x"57",
          1805 => x"f9",
          1806 => x"e2",
          1807 => x"f9",
          1808 => x"e2",
          1809 => x"2c",
          1810 => x"61",
          1811 => x"e8",
          1812 => x"3f",
          1813 => x"70",
          1814 => x"57",
          1815 => x"38",
          1816 => x"ff",
          1817 => x"29",
          1818 => x"84",
          1819 => x"7b",
          1820 => x"08",
          1821 => x"74",
          1822 => x"05",
          1823 => x"5d",
          1824 => x"38",
          1825 => x"18",
          1826 => x"52",
          1827 => x"75",
          1828 => x"05",
          1829 => x"5c",
          1830 => x"38",
          1831 => x"34",
          1832 => x"51",
          1833 => x"0a",
          1834 => x"2c",
          1835 => x"79",
          1836 => x"39",
          1837 => x"2e",
          1838 => x"52",
          1839 => x"e2",
          1840 => x"e2",
          1841 => x"dd",
          1842 => x"41",
          1843 => x"52",
          1844 => x"e2",
          1845 => x"84",
          1846 => x"77",
          1847 => x"57",
          1848 => x"f4",
          1849 => x"9c",
          1850 => x"8b",
          1851 => x"06",
          1852 => x"53",
          1853 => x"bb",
          1854 => x"33",
          1855 => x"70",
          1856 => x"5b",
          1857 => x"33",
          1858 => x"70",
          1859 => x"38",
          1860 => x"2e",
          1861 => x"77",
          1862 => x"84",
          1863 => x"c4",
          1864 => x"3d",
          1865 => x"74",
          1866 => x"08",
          1867 => x"84",
          1868 => x"ae",
          1869 => x"88",
          1870 => x"c8",
          1871 => x"c8",
          1872 => x"cc",
          1873 => x"fe",
          1874 => x"80",
          1875 => x"39",
          1876 => x"06",
          1877 => x"38",
          1878 => x"79",
          1879 => x"77",
          1880 => x"08",
          1881 => x"84",
          1882 => x"98",
          1883 => x"5a",
          1884 => x"84",
          1885 => x"ad",
          1886 => x"98",
          1887 => x"33",
          1888 => x"f3",
          1889 => x"88",
          1890 => x"80",
          1891 => x"98",
          1892 => x"55",
          1893 => x"e6",
          1894 => x"bc",
          1895 => x"80",
          1896 => x"c4",
          1897 => x"ff",
          1898 => x"57",
          1899 => x"e8",
          1900 => x"8c",
          1901 => x"80",
          1902 => x"c4",
          1903 => x"fe",
          1904 => x"33",
          1905 => x"76",
          1906 => x"81",
          1907 => x"70",
          1908 => x"57",
          1909 => x"fe",
          1910 => x"81",
          1911 => x"74",
          1912 => x"08",
          1913 => x"84",
          1914 => x"ab",
          1915 => x"88",
          1916 => x"c8",
          1917 => x"c8",
          1918 => x"cc",
          1919 => x"8e",
          1920 => x"80",
          1921 => x"bb",
          1922 => x"e2",
          1923 => x"58",
          1924 => x"e2",
          1925 => x"38",
          1926 => x"42",
          1927 => x"5b",
          1928 => x"80",
          1929 => x"98",
          1930 => x"58",
          1931 => x"55",
          1932 => x"ff",
          1933 => x"79",
          1934 => x"61",
          1935 => x"84",
          1936 => x"c8",
          1937 => x"ff",
          1938 => x"ff",
          1939 => x"24",
          1940 => x"98",
          1941 => x"5a",
          1942 => x"e6",
          1943 => x"b4",
          1944 => x"80",
          1945 => x"c4",
          1946 => x"f0",
          1947 => x"88",
          1948 => x"80",
          1949 => x"98",
          1950 => x"42",
          1951 => x"83",
          1952 => x"3f",
          1953 => x"0c",
          1954 => x"c0",
          1955 => x"ec",
          1956 => x"83",
          1957 => x"80",
          1958 => x"7b",
          1959 => x"b4",
          1960 => x"80",
          1961 => x"c4",
          1962 => x"da",
          1963 => x"2b",
          1964 => x"5c",
          1965 => x"93",
          1966 => x"08",
          1967 => x"9c",
          1968 => x"bb",
          1969 => x"75",
          1970 => x"f4",
          1971 => x"74",
          1972 => x"81",
          1973 => x"51",
          1974 => x"f4",
          1975 => x"40",
          1976 => x"97",
          1977 => x"18",
          1978 => x"38",
          1979 => x"ce",
          1980 => x"c4",
          1981 => x"06",
          1982 => x"ff",
          1983 => x"c4",
          1984 => x"5d",
          1985 => x"e6",
          1986 => x"dc",
          1987 => x"51",
          1988 => x"08",
          1989 => x"84",
          1990 => x"84",
          1991 => x"55",
          1992 => x"3f",
          1993 => x"34",
          1994 => x"81",
          1995 => x"aa",
          1996 => x"84",
          1997 => x"80",
          1998 => x"08",
          1999 => x"84",
          2000 => x"a5",
          2001 => x"88",
          2002 => x"c8",
          2003 => x"c8",
          2004 => x"39",
          2005 => x"bb",
          2006 => x"bb",
          2007 => x"53",
          2008 => x"3f",
          2009 => x"e2",
          2010 => x"52",
          2011 => x"38",
          2012 => x"ff",
          2013 => x"52",
          2014 => x"e6",
          2015 => x"f4",
          2016 => x"5b",
          2017 => x"ff",
          2018 => x"80",
          2019 => x"84",
          2020 => x"0c",
          2021 => x"08",
          2022 => x"75",
          2023 => x"84",
          2024 => x"84",
          2025 => x"75",
          2026 => x"84",
          2027 => x"56",
          2028 => x"84",
          2029 => x"a4",
          2030 => x"a0",
          2031 => x"e8",
          2032 => x"3f",
          2033 => x"78",
          2034 => x"06",
          2035 => x"bf",
          2036 => x"2b",
          2037 => x"81",
          2038 => x"dd",
          2039 => x"0c",
          2040 => x"83",
          2041 => x"83",
          2042 => x"3f",
          2043 => x"83",
          2044 => x"5e",
          2045 => x"53",
          2046 => x"3f",
          2047 => x"81",
          2048 => x"83",
          2049 => x"f4",
          2050 => x"54",
          2051 => x"d9",
          2052 => x"8a",
          2053 => x"ec",
          2054 => x"0b",
          2055 => x"e2",
          2056 => x"b5",
          2057 => x"74",
          2058 => x"84",
          2059 => x"08",
          2060 => x"08",
          2061 => x"b7",
          2062 => x"84",
          2063 => x"06",
          2064 => x"51",
          2065 => x"08",
          2066 => x"25",
          2067 => x"ff",
          2068 => x"34",
          2069 => x"33",
          2070 => x"70",
          2071 => x"8a",
          2072 => x"83",
          2073 => x"57",
          2074 => x"84",
          2075 => x"70",
          2076 => x"08",
          2077 => x"ff",
          2078 => x"70",
          2079 => x"08",
          2080 => x"1d",
          2081 => x"7d",
          2082 => x"2e",
          2083 => x"e7",
          2084 => x"79",
          2085 => x"83",
          2086 => x"ff",
          2087 => x"e0",
          2088 => x"ff",
          2089 => x"3f",
          2090 => x"87",
          2091 => x"1b",
          2092 => x"e7",
          2093 => x"83",
          2094 => x"f4",
          2095 => x"e3",
          2096 => x"83",
          2097 => x"f4",
          2098 => x"74",
          2099 => x"39",
          2100 => x"39",
          2101 => x"39",
          2102 => x"3f",
          2103 => x"f2",
          2104 => x"02",
          2105 => x"53",
          2106 => x"81",
          2107 => x"83",
          2108 => x"38",
          2109 => x"b0",
          2110 => x"a0",
          2111 => x"83",
          2112 => x"34",
          2113 => x"b0",
          2114 => x"07",
          2115 => x"7f",
          2116 => x"94",
          2117 => x"0c",
          2118 => x"76",
          2119 => x"a2",
          2120 => x"d6",
          2121 => x"a0",
          2122 => x"70",
          2123 => x"72",
          2124 => x"c7",
          2125 => x"70",
          2126 => x"71",
          2127 => x"58",
          2128 => x"84",
          2129 => x"84",
          2130 => x"83",
          2131 => x"06",
          2132 => x"5e",
          2133 => x"38",
          2134 => x"81",
          2135 => x"81",
          2136 => x"62",
          2137 => x"5d",
          2138 => x"26",
          2139 => x"76",
          2140 => x"5f",
          2141 => x"fe",
          2142 => x"77",
          2143 => x"81",
          2144 => x"74",
          2145 => x"86",
          2146 => x"80",
          2147 => x"ff",
          2148 => x"ff",
          2149 => x"29",
          2150 => x"57",
          2151 => x"81",
          2152 => x"71",
          2153 => x"2e",
          2154 => x"b4",
          2155 => x"83",
          2156 => x"90",
          2157 => x"07",
          2158 => x"79",
          2159 => x"72",
          2160 => x"70",
          2161 => x"83",
          2162 => x"86",
          2163 => x"56",
          2164 => x"14",
          2165 => x"06",
          2166 => x"06",
          2167 => x"ff",
          2168 => x"5a",
          2169 => x"79",
          2170 => x"15",
          2171 => x"81",
          2172 => x"71",
          2173 => x"81",
          2174 => x"5b",
          2175 => x"38",
          2176 => x"16",
          2177 => x"e2",
          2178 => x"da",
          2179 => x"7b",
          2180 => x"0d",
          2181 => x"73",
          2182 => x"81",
          2183 => x"80",
          2184 => x"87",
          2185 => x"80",
          2186 => x"8a",
          2187 => x"75",
          2188 => x"3f",
          2189 => x"54",
          2190 => x"73",
          2191 => x"75",
          2192 => x"80",
          2193 => x"86",
          2194 => x"81",
          2195 => x"f3",
          2196 => x"07",
          2197 => x"84",
          2198 => x"84",
          2199 => x"f8",
          2200 => x"3d",
          2201 => x"05",
          2202 => x"5b",
          2203 => x"82",
          2204 => x"fa",
          2205 => x"71",
          2206 => x"83",
          2207 => x"71",
          2208 => x"06",
          2209 => x"53",
          2210 => x"fa",
          2211 => x"fa",
          2212 => x"05",
          2213 => x"06",
          2214 => x"8c",
          2215 => x"b4",
          2216 => x"ff",
          2217 => x"55",
          2218 => x"84",
          2219 => x"58",
          2220 => x"38",
          2221 => x"e0",
          2222 => x"72",
          2223 => x"81",
          2224 => x"b8",
          2225 => x"9f",
          2226 => x"84",
          2227 => x"e0",
          2228 => x"05",
          2229 => x"74",
          2230 => x"ff",
          2231 => x"75",
          2232 => x"ff",
          2233 => x"81",
          2234 => x"84",
          2235 => x"55",
          2236 => x"58",
          2237 => x"06",
          2238 => x"19",
          2239 => x"b9",
          2240 => x"e0",
          2241 => x"33",
          2242 => x"70",
          2243 => x"05",
          2244 => x"33",
          2245 => x"19",
          2246 => x"ce",
          2247 => x"0c",
          2248 => x"b4",
          2249 => x"ff",
          2250 => x"55",
          2251 => x"77",
          2252 => x"ff",
          2253 => x"56",
          2254 => x"fe",
          2255 => x"84",
          2256 => x"72",
          2257 => x"73",
          2258 => x"33",
          2259 => x"55",
          2260 => x"34",
          2261 => x"ff",
          2262 => x"38",
          2263 => x"75",
          2264 => x"53",
          2265 => x"0b",
          2266 => x"89",
          2267 => x"84",
          2268 => x"b8",
          2269 => x"3d",
          2270 => x"33",
          2271 => x"70",
          2272 => x"70",
          2273 => x"71",
          2274 => x"b5",
          2275 => x"86",
          2276 => x"b5",
          2277 => x"ff",
          2278 => x"38",
          2279 => x"34",
          2280 => x"3d",
          2281 => x"73",
          2282 => x"06",
          2283 => x"b4",
          2284 => x"72",
          2285 => x"55",
          2286 => x"70",
          2287 => x"0b",
          2288 => x"04",
          2289 => x"70",
          2290 => x"56",
          2291 => x"80",
          2292 => x"0d",
          2293 => x"84",
          2294 => x"51",
          2295 => x"72",
          2296 => x"bb",
          2297 => x"0b",
          2298 => x"33",
          2299 => x"52",
          2300 => x"12",
          2301 => x"d0",
          2302 => x"33",
          2303 => x"10",
          2304 => x"08",
          2305 => x"f0",
          2306 => x"70",
          2307 => x"51",
          2308 => x"9c",
          2309 => x"34",
          2310 => x"3d",
          2311 => x"9f",
          2312 => x"b0",
          2313 => x"83",
          2314 => x"80",
          2315 => x"34",
          2316 => x"fe",
          2317 => x"b0",
          2318 => x"fa",
          2319 => x"0c",
          2320 => x"33",
          2321 => x"83",
          2322 => x"fa",
          2323 => x"fa",
          2324 => x"b0",
          2325 => x"70",
          2326 => x"83",
          2327 => x"07",
          2328 => x"81",
          2329 => x"06",
          2330 => x"34",
          2331 => x"81",
          2332 => x"34",
          2333 => x"81",
          2334 => x"83",
          2335 => x"fa",
          2336 => x"51",
          2337 => x"39",
          2338 => x"80",
          2339 => x"34",
          2340 => x"81",
          2341 => x"83",
          2342 => x"fa",
          2343 => x"51",
          2344 => x"39",
          2345 => x"51",
          2346 => x"39",
          2347 => x"82",
          2348 => x"fd",
          2349 => x"05",
          2350 => x"33",
          2351 => x"33",
          2352 => x"33",
          2353 => x"82",
          2354 => x"a5",
          2355 => x"7d",
          2356 => x"b8",
          2357 => x"7b",
          2358 => x"b5",
          2359 => x"2e",
          2360 => x"84",
          2361 => x"fc",
          2362 => x"a8",
          2363 => x"83",
          2364 => x"f8",
          2365 => x"84",
          2366 => x"53",
          2367 => x"80",
          2368 => x"80",
          2369 => x"fa",
          2370 => x"7c",
          2371 => x"04",
          2372 => x"0b",
          2373 => x"fa",
          2374 => x"34",
          2375 => x"ba",
          2376 => x"57",
          2377 => x"7b",
          2378 => x"94",
          2379 => x"84",
          2380 => x"27",
          2381 => x"05",
          2382 => x"51",
          2383 => x"81",
          2384 => x"5b",
          2385 => x"d3",
          2386 => x"84",
          2387 => x"fc",
          2388 => x"83",
          2389 => x"34",
          2390 => x"b8",
          2391 => x"34",
          2392 => x"0b",
          2393 => x"fa",
          2394 => x"90",
          2395 => x"83",
          2396 => x"80",
          2397 => x"be",
          2398 => x"fd",
          2399 => x"52",
          2400 => x"3f",
          2401 => x"5a",
          2402 => x"84",
          2403 => x"33",
          2404 => x"33",
          2405 => x"80",
          2406 => x"59",
          2407 => x"ff",
          2408 => x"59",
          2409 => x"81",
          2410 => x"38",
          2411 => x"81",
          2412 => x"82",
          2413 => x"fa",
          2414 => x"72",
          2415 => x"80",
          2416 => x"34",
          2417 => x"33",
          2418 => x"12",
          2419 => x"b6",
          2420 => x"71",
          2421 => x"33",
          2422 => x"b8",
          2423 => x"fa",
          2424 => x"72",
          2425 => x"83",
          2426 => x"34",
          2427 => x"55",
          2428 => x"b8",
          2429 => x"ff",
          2430 => x"84",
          2431 => x"8c",
          2432 => x"80",
          2433 => x"bb",
          2434 => x"8d",
          2435 => x"f7",
          2436 => x"fe",
          2437 => x"96",
          2438 => x"ff",
          2439 => x"53",
          2440 => x"75",
          2441 => x"38",
          2442 => x"ba",
          2443 => x"54",
          2444 => x"76",
          2445 => x"13",
          2446 => x"73",
          2447 => x"83",
          2448 => x"52",
          2449 => x"84",
          2450 => x"75",
          2451 => x"ca",
          2452 => x"ff",
          2453 => x"38",
          2454 => x"76",
          2455 => x"fa",
          2456 => x"ff",
          2457 => x"53",
          2458 => x"39",
          2459 => x"52",
          2460 => x"39",
          2461 => x"fe",
          2462 => x"f3",
          2463 => x"59",
          2464 => x"82",
          2465 => x"84",
          2466 => x"38",
          2467 => x"89",
          2468 => x"33",
          2469 => x"33",
          2470 => x"84",
          2471 => x"80",
          2472 => x"fa",
          2473 => x"71",
          2474 => x"83",
          2475 => x"33",
          2476 => x"83",
          2477 => x"80",
          2478 => x"81",
          2479 => x"fa",
          2480 => x"40",
          2481 => x"84",
          2482 => x"81",
          2483 => x"81",
          2484 => x"79",
          2485 => x"83",
          2486 => x"84",
          2487 => x"2e",
          2488 => x"fd",
          2489 => x"78",
          2490 => x"0b",
          2491 => x"33",
          2492 => x"33",
          2493 => x"84",
          2494 => x"80",
          2495 => x"fa",
          2496 => x"71",
          2497 => x"83",
          2498 => x"33",
          2499 => x"fa",
          2500 => x"34",
          2501 => x"06",
          2502 => x"33",
          2503 => x"58",
          2504 => x"99",
          2505 => x"81",
          2506 => x"ca",
          2507 => x"0b",
          2508 => x"04",
          2509 => x"9b",
          2510 => x"09",
          2511 => x"83",
          2512 => x"84",
          2513 => x"2e",
          2514 => x"89",
          2515 => x"33",
          2516 => x"84",
          2517 => x"77",
          2518 => x"ba",
          2519 => x"84",
          2520 => x"2e",
          2521 => x"80",
          2522 => x"b4",
          2523 => x"29",
          2524 => x"19",
          2525 => x"84",
          2526 => x"83",
          2527 => x"41",
          2528 => x"1f",
          2529 => x"29",
          2530 => x"86",
          2531 => x"f8",
          2532 => x"b2",
          2533 => x"29",
          2534 => x"fa",
          2535 => x"34",
          2536 => x"52",
          2537 => x"83",
          2538 => x"b8",
          2539 => x"81",
          2540 => x"71",
          2541 => x"83",
          2542 => x"7e",
          2543 => x"83",
          2544 => x"5c",
          2545 => x"81",
          2546 => x"fc",
          2547 => x"b5",
          2548 => x"ba",
          2549 => x"34",
          2550 => x"0b",
          2551 => x"ba",
          2552 => x"0c",
          2553 => x"33",
          2554 => x"33",
          2555 => x"33",
          2556 => x"ba",
          2557 => x"0c",
          2558 => x"2e",
          2559 => x"fa",
          2560 => x"81",
          2561 => x"81",
          2562 => x"c7",
          2563 => x"5c",
          2564 => x"ff",
          2565 => x"5c",
          2566 => x"2e",
          2567 => x"ff",
          2568 => x"57",
          2569 => x"ff",
          2570 => x"ff",
          2571 => x"5b",
          2572 => x"80",
          2573 => x"fa",
          2574 => x"71",
          2575 => x"0b",
          2576 => x"b4",
          2577 => x"56",
          2578 => x"80",
          2579 => x"81",
          2580 => x"fa",
          2581 => x"5d",
          2582 => x"7f",
          2583 => x"70",
          2584 => x"26",
          2585 => x"5a",
          2586 => x"77",
          2587 => x"33",
          2588 => x"56",
          2589 => x"d8",
          2590 => x"78",
          2591 => x"84",
          2592 => x"bf",
          2593 => x"38",
          2594 => x"58",
          2595 => x"b5",
          2596 => x"3f",
          2597 => x"3d",
          2598 => x"b8",
          2599 => x"fa",
          2600 => x"75",
          2601 => x"83",
          2602 => x"29",
          2603 => x"f9",
          2604 => x"5b",
          2605 => x"80",
          2606 => x"ff",
          2607 => x"29",
          2608 => x"33",
          2609 => x"b8",
          2610 => x"fa",
          2611 => x"41",
          2612 => x"1c",
          2613 => x"29",
          2614 => x"86",
          2615 => x"f8",
          2616 => x"b2",
          2617 => x"29",
          2618 => x"fa",
          2619 => x"60",
          2620 => x"58",
          2621 => x"b8",
          2622 => x"ff",
          2623 => x"81",
          2624 => x"7b",
          2625 => x"b4",
          2626 => x"b5",
          2627 => x"ff",
          2628 => x"29",
          2629 => x"84",
          2630 => x"1b",
          2631 => x"b5",
          2632 => x"29",
          2633 => x"83",
          2634 => x"33",
          2635 => x"fa",
          2636 => x"34",
          2637 => x"06",
          2638 => x"33",
          2639 => x"40",
          2640 => x"d6",
          2641 => x"ff",
          2642 => x"d6",
          2643 => x"df",
          2644 => x"80",
          2645 => x"0d",
          2646 => x"84",
          2647 => x"fa",
          2648 => x"ff",
          2649 => x"84",
          2650 => x"84",
          2651 => x"b6",
          2652 => x"33",
          2653 => x"b8",
          2654 => x"5b",
          2655 => x"ba",
          2656 => x"d8",
          2657 => x"bb",
          2658 => x"84",
          2659 => x"75",
          2660 => x"fe",
          2661 => x"61",
          2662 => x"39",
          2663 => x"b9",
          2664 => x"b4",
          2665 => x"b5",
          2666 => x"84",
          2667 => x"83",
          2668 => x"41",
          2669 => x"7f",
          2670 => x"b8",
          2671 => x"fa",
          2672 => x"43",
          2673 => x"34",
          2674 => x"1b",
          2675 => x"86",
          2676 => x"f8",
          2677 => x"b2",
          2678 => x"29",
          2679 => x"fa",
          2680 => x"81",
          2681 => x"60",
          2682 => x"f9",
          2683 => x"1a",
          2684 => x"0b",
          2685 => x"33",
          2686 => x"84",
          2687 => x"38",
          2688 => x"80",
          2689 => x"0d",
          2690 => x"b4",
          2691 => x"b5",
          2692 => x"83",
          2693 => x"fa",
          2694 => x"fa",
          2695 => x"fa",
          2696 => x"9e",
          2697 => x"80",
          2698 => x"22",
          2699 => x"ff",
          2700 => x"05",
          2701 => x"54",
          2702 => x"3d",
          2703 => x"76",
          2704 => x"84",
          2705 => x"33",
          2706 => x"fe",
          2707 => x"51",
          2708 => x"80",
          2709 => x"79",
          2710 => x"fe",
          2711 => x"05",
          2712 => x"26",
          2713 => x"c8",
          2714 => x"ba",
          2715 => x"a4",
          2716 => x"d9",
          2717 => x"9f",
          2718 => x"5c",
          2719 => x"39",
          2720 => x"2e",
          2721 => x"ff",
          2722 => x"f8",
          2723 => x"fd",
          2724 => x"fd",
          2725 => x"34",
          2726 => x"06",
          2727 => x"38",
          2728 => x"34",
          2729 => x"b5",
          2730 => x"f7",
          2731 => x"25",
          2732 => x"83",
          2733 => x"ba",
          2734 => x"e0",
          2735 => x"d9",
          2736 => x"9f",
          2737 => x"5a",
          2738 => x"39",
          2739 => x"2e",
          2740 => x"41",
          2741 => x"b6",
          2742 => x"b5",
          2743 => x"29",
          2744 => x"fa",
          2745 => x"60",
          2746 => x"83",
          2747 => x"06",
          2748 => x"80",
          2749 => x"f9",
          2750 => x"85",
          2751 => x"38",
          2752 => x"2e",
          2753 => x"0b",
          2754 => x"84",
          2755 => x"90",
          2756 => x"fa",
          2757 => x"f8",
          2758 => x"7d",
          2759 => x"fa",
          2760 => x"85",
          2761 => x"38",
          2762 => x"33",
          2763 => x"ff",
          2764 => x"83",
          2765 => x"34",
          2766 => x"fe",
          2767 => x"85",
          2768 => x"c7",
          2769 => x"70",
          2770 => x"fe",
          2771 => x"ff",
          2772 => x"58",
          2773 => x"33",
          2774 => x"84",
          2775 => x"83",
          2776 => x"ff",
          2777 => x"39",
          2778 => x"27",
          2779 => x"ff",
          2780 => x"d9",
          2781 => x"84",
          2782 => x"ff",
          2783 => x"5c",
          2784 => x"79",
          2785 => x"06",
          2786 => x"83",
          2787 => x"34",
          2788 => x"40",
          2789 => x"56",
          2790 => x"39",
          2791 => x"2e",
          2792 => x"84",
          2793 => x"26",
          2794 => x"84",
          2795 => x"83",
          2796 => x"86",
          2797 => x"22",
          2798 => x"83",
          2799 => x"46",
          2800 => x"2e",
          2801 => x"06",
          2802 => x"24",
          2803 => x"56",
          2804 => x"16",
          2805 => x"81",
          2806 => x"80",
          2807 => x"f7",
          2808 => x"38",
          2809 => x"34",
          2810 => x"22",
          2811 => x"90",
          2812 => x"81",
          2813 => x"5b",
          2814 => x"86",
          2815 => x"7f",
          2816 => x"42",
          2817 => x"d6",
          2818 => x"e0",
          2819 => x"33",
          2820 => x"70",
          2821 => x"05",
          2822 => x"33",
          2823 => x"1d",
          2824 => x"f7",
          2825 => x"84",
          2826 => x"05",
          2827 => x"33",
          2828 => x"18",
          2829 => x"33",
          2830 => x"58",
          2831 => x"e6",
          2832 => x"80",
          2833 => x"ba",
          2834 => x"ce",
          2835 => x"ff",
          2836 => x"40",
          2837 => x"ba",
          2838 => x"81",
          2839 => x"33",
          2840 => x"b4",
          2841 => x"2e",
          2842 => x"40",
          2843 => x"81",
          2844 => x"fe",
          2845 => x"07",
          2846 => x"10",
          2847 => x"c7",
          2848 => x"86",
          2849 => x"58",
          2850 => x"83",
          2851 => x"fa",
          2852 => x"2b",
          2853 => x"79",
          2854 => x"27",
          2855 => x"59",
          2856 => x"0c",
          2857 => x"f8",
          2858 => x"7e",
          2859 => x"83",
          2860 => x"05",
          2861 => x"8c",
          2862 => x"29",
          2863 => x"57",
          2864 => x"83",
          2865 => x"59",
          2866 => x"79",
          2867 => x"17",
          2868 => x"a0",
          2869 => x"70",
          2870 => x"75",
          2871 => x"ff",
          2872 => x"fe",
          2873 => x"80",
          2874 => x"06",
          2875 => x"7b",
          2876 => x"38",
          2877 => x"81",
          2878 => x"f5",
          2879 => x"5e",
          2880 => x"83",
          2881 => x"83",
          2882 => x"42",
          2883 => x"fa",
          2884 => x"fa",
          2885 => x"06",
          2886 => x"b0",
          2887 => x"75",
          2888 => x"fa",
          2889 => x"56",
          2890 => x"83",
          2891 => x"07",
          2892 => x"39",
          2893 => x"90",
          2894 => x"ff",
          2895 => x"b0",
          2896 => x"59",
          2897 => x"33",
          2898 => x"b0",
          2899 => x"33",
          2900 => x"83",
          2901 => x"fa",
          2902 => x"07",
          2903 => x"ea",
          2904 => x"06",
          2905 => x"b0",
          2906 => x"33",
          2907 => x"83",
          2908 => x"fa",
          2909 => x"56",
          2910 => x"39",
          2911 => x"84",
          2912 => x"fe",
          2913 => x"fa",
          2914 => x"b0",
          2915 => x"33",
          2916 => x"b0",
          2917 => x"33",
          2918 => x"b0",
          2919 => x"33",
          2920 => x"b0",
          2921 => x"33",
          2922 => x"75",
          2923 => x"83",
          2924 => x"07",
          2925 => x"ba",
          2926 => x"80",
          2927 => x"ff",
          2928 => x"b4",
          2929 => x"b5",
          2930 => x"83",
          2931 => x"80",
          2932 => x"ba",
          2933 => x"0c",
          2934 => x"b5",
          2935 => x"ff",
          2936 => x"39",
          2937 => x"11",
          2938 => x"3f",
          2939 => x"bb",
          2940 => x"0b",
          2941 => x"bb",
          2942 => x"83",
          2943 => x"ba",
          2944 => x"84",
          2945 => x"06",
          2946 => x"ba",
          2947 => x"84",
          2948 => x"b5",
          2949 => x"3f",
          2950 => x"06",
          2951 => x"80",
          2952 => x"81",
          2953 => x"8a",
          2954 => x"39",
          2955 => x"09",
          2956 => x"57",
          2957 => x"d9",
          2958 => x"60",
          2959 => x"b5",
          2960 => x"33",
          2961 => x"72",
          2962 => x"83",
          2963 => x"f7",
          2964 => x"78",
          2965 => x"bb",
          2966 => x"ff",
          2967 => x"a6",
          2968 => x"f8",
          2969 => x"b5",
          2970 => x"a0",
          2971 => x"5f",
          2972 => x"ff",
          2973 => x"44",
          2974 => x"f5",
          2975 => x"11",
          2976 => x"38",
          2977 => x"27",
          2978 => x"83",
          2979 => x"ff",
          2980 => x"df",
          2981 => x"76",
          2982 => x"75",
          2983 => x"06",
          2984 => x"5a",
          2985 => x"31",
          2986 => x"71",
          2987 => x"c7",
          2988 => x"7c",
          2989 => x"71",
          2990 => x"79",
          2991 => x"d6",
          2992 => x"84",
          2993 => x"05",
          2994 => x"33",
          2995 => x"18",
          2996 => x"33",
          2997 => x"58",
          2998 => x"e0",
          2999 => x"33",
          3000 => x"70",
          3001 => x"05",
          3002 => x"33",
          3003 => x"1d",
          3004 => x"ff",
          3005 => x"b6",
          3006 => x"33",
          3007 => x"b8",
          3008 => x"b8",
          3009 => x"e9",
          3010 => x"f7",
          3011 => x"5c",
          3012 => x"76",
          3013 => x"81",
          3014 => x"7a",
          3015 => x"fa",
          3016 => x"81",
          3017 => x"80",
          3018 => x"75",
          3019 => x"83",
          3020 => x"f8",
          3021 => x"7f",
          3022 => x"c5",
          3023 => x"f4",
          3024 => x"81",
          3025 => x"44",
          3026 => x"81",
          3027 => x"ff",
          3028 => x"fd",
          3029 => x"fa",
          3030 => x"31",
          3031 => x"90",
          3032 => x"26",
          3033 => x"05",
          3034 => x"70",
          3035 => x"f4",
          3036 => x"58",
          3037 => x"81",
          3038 => x"38",
          3039 => x"75",
          3040 => x"80",
          3041 => x"39",
          3042 => x"39",
          3043 => x"8e",
          3044 => x"f1",
          3045 => x"5a",
          3046 => x"80",
          3047 => x"39",
          3048 => x"84",
          3049 => x"2e",
          3050 => x"80",
          3051 => x"0d",
          3052 => x"3f",
          3053 => x"3d",
          3054 => x"05",
          3055 => x"33",
          3056 => x"11",
          3057 => x"2e",
          3058 => x"83",
          3059 => x"bb",
          3060 => x"f8",
          3061 => x"2e",
          3062 => x"71",
          3063 => x"5d",
          3064 => x"ff",
          3065 => x"81",
          3066 => x"32",
          3067 => x"5c",
          3068 => x"38",
          3069 => x"33",
          3070 => x"12",
          3071 => x"b2",
          3072 => x"05",
          3073 => x"89",
          3074 => x"2e",
          3075 => x"87",
          3076 => x"c0",
          3077 => x"08",
          3078 => x"8e",
          3079 => x"b4",
          3080 => x"06",
          3081 => x"38",
          3082 => x"70",
          3083 => x"33",
          3084 => x"c1",
          3085 => x"38",
          3086 => x"81",
          3087 => x"85",
          3088 => x"34",
          3089 => x"ae",
          3090 => x"06",
          3091 => x"38",
          3092 => x"70",
          3093 => x"f8",
          3094 => x"86",
          3095 => x"54",
          3096 => x"81",
          3097 => x"81",
          3098 => x"38",
          3099 => x"0b",
          3100 => x"08",
          3101 => x"e0",
          3102 => x"42",
          3103 => x"16",
          3104 => x"38",
          3105 => x"80",
          3106 => x"16",
          3107 => x"38",
          3108 => x"81",
          3109 => x"73",
          3110 => x"cc",
          3111 => x"da",
          3112 => x"81",
          3113 => x"cc",
          3114 => x"80",
          3115 => x"05",
          3116 => x"73",
          3117 => x"87",
          3118 => x"0c",
          3119 => x"57",
          3120 => x"76",
          3121 => x"e0",
          3122 => x"26",
          3123 => x"c9",
          3124 => x"f9",
          3125 => x"38",
          3126 => x"08",
          3127 => x"38",
          3128 => x"54",
          3129 => x"73",
          3130 => x"9c",
          3131 => x"ff",
          3132 => x"83",
          3133 => x"80",
          3134 => x"fc",
          3135 => x"72",
          3136 => x"2e",
          3137 => x"81",
          3138 => x"fe",
          3139 => x"59",
          3140 => x"2e",
          3141 => x"81",
          3142 => x"80",
          3143 => x"87",
          3144 => x"72",
          3145 => x"9c",
          3146 => x"76",
          3147 => x"71",
          3148 => x"80",
          3149 => x"10",
          3150 => x"78",
          3151 => x"5b",
          3152 => x"08",
          3153 => x"39",
          3154 => x"38",
          3155 => x"39",
          3156 => x"2e",
          3157 => x"fa",
          3158 => x"e8",
          3159 => x"80",
          3160 => x"8a",
          3161 => x"f9",
          3162 => x"38",
          3163 => x"f9",
          3164 => x"7c",
          3165 => x"81",
          3166 => x"e2",
          3167 => x"80",
          3168 => x"33",
          3169 => x"ff",
          3170 => x"78",
          3171 => x"04",
          3172 => x"f6",
          3173 => x"83",
          3174 => x"7a",
          3175 => x"39",
          3176 => x"ff",
          3177 => x"0b",
          3178 => x"39",
          3179 => x"ff",
          3180 => x"16",
          3181 => x"38",
          3182 => x"2e",
          3183 => x"f8",
          3184 => x"98",
          3185 => x"fb",
          3186 => x"83",
          3187 => x"59",
          3188 => x"b8",
          3189 => x"f8",
          3190 => x"72",
          3191 => x"34",
          3192 => x"f8",
          3193 => x"83",
          3194 => x"5d",
          3195 => x"9c",
          3196 => x"fc",
          3197 => x"fc",
          3198 => x"06",
          3199 => x"76",
          3200 => x"80",
          3201 => x"75",
          3202 => x"fb",
          3203 => x"0b",
          3204 => x"83",
          3205 => x"34",
          3206 => x"83",
          3207 => x"38",
          3208 => x"ff",
          3209 => x"ff",
          3210 => x"79",
          3211 => x"fa",
          3212 => x"15",
          3213 => x"80",
          3214 => x"b8",
          3215 => x"ff",
          3216 => x"80",
          3217 => x"59",
          3218 => x"ff",
          3219 => x"39",
          3220 => x"08",
          3221 => x"9d",
          3222 => x"83",
          3223 => x"80",
          3224 => x"82",
          3225 => x"0b",
          3226 => x"a3",
          3227 => x"90",
          3228 => x"0b",
          3229 => x"0b",
          3230 => x"80",
          3231 => x"83",
          3232 => x"05",
          3233 => x"87",
          3234 => x"2e",
          3235 => x"98",
          3236 => x"87",
          3237 => x"87",
          3238 => x"70",
          3239 => x"71",
          3240 => x"98",
          3241 => x"87",
          3242 => x"98",
          3243 => x"38",
          3244 => x"08",
          3245 => x"71",
          3246 => x"98",
          3247 => x"38",
          3248 => x"81",
          3249 => x"98",
          3250 => x"fe",
          3251 => x"76",
          3252 => x"04",
          3253 => x"3d",
          3254 => x"84",
          3255 => x"0b",
          3256 => x"87",
          3257 => x"2a",
          3258 => x"15",
          3259 => x"15",
          3260 => x"15",
          3261 => x"90",
          3262 => x"f5",
          3263 => x"85",
          3264 => x"fe",
          3265 => x"90",
          3266 => x"08",
          3267 => x"90",
          3268 => x"52",
          3269 => x"72",
          3270 => x"c0",
          3271 => x"27",
          3272 => x"38",
          3273 => x"55",
          3274 => x"55",
          3275 => x"c0",
          3276 => x"53",
          3277 => x"c0",
          3278 => x"f6",
          3279 => x"9c",
          3280 => x"38",
          3281 => x"c0",
          3282 => x"83",
          3283 => x"70",
          3284 => x"2e",
          3285 => x"52",
          3286 => x"81",
          3287 => x"c6",
          3288 => x"52",
          3289 => x"81",
          3290 => x"53",
          3291 => x"84",
          3292 => x"81",
          3293 => x"0d",
          3294 => x"0d",
          3295 => x"56",
          3296 => x"77",
          3297 => x"70",
          3298 => x"57",
          3299 => x"51",
          3300 => x"52",
          3301 => x"34",
          3302 => x"11",
          3303 => x"70",
          3304 => x"05",
          3305 => x"34",
          3306 => x"90",
          3307 => x"f5",
          3308 => x"85",
          3309 => x"fe",
          3310 => x"90",
          3311 => x"08",
          3312 => x"90",
          3313 => x"52",
          3314 => x"72",
          3315 => x"c0",
          3316 => x"27",
          3317 => x"38",
          3318 => x"55",
          3319 => x"55",
          3320 => x"c0",
          3321 => x"53",
          3322 => x"c0",
          3323 => x"f6",
          3324 => x"9c",
          3325 => x"38",
          3326 => x"c0",
          3327 => x"83",
          3328 => x"70",
          3329 => x"2e",
          3330 => x"71",
          3331 => x"ff",
          3332 => x"81",
          3333 => x"3d",
          3334 => x"3d",
          3335 => x"d0",
          3336 => x"08",
          3337 => x"80",
          3338 => x"c0",
          3339 => x"56",
          3340 => x"98",
          3341 => x"08",
          3342 => x"15",
          3343 => x"52",
          3344 => x"fe",
          3345 => x"08",
          3346 => x"c8",
          3347 => x"c0",
          3348 => x"ce",
          3349 => x"08",
          3350 => x"70",
          3351 => x"87",
          3352 => x"73",
          3353 => x"db",
          3354 => x"72",
          3355 => x"53",
          3356 => x"52",
          3357 => x"ff",
          3358 => x"39",
          3359 => x"fe",
          3360 => x"f9",
          3361 => x"71",
          3362 => x"06",
          3363 => x"81",
          3364 => x"2b",
          3365 => x"33",
          3366 => x"5c",
          3367 => x"52",
          3368 => x"af",
          3369 => x"12",
          3370 => x"07",
          3371 => x"71",
          3372 => x"53",
          3373 => x"24",
          3374 => x"14",
          3375 => x"07",
          3376 => x"56",
          3377 => x"ff",
          3378 => x"ba",
          3379 => x"85",
          3380 => x"88",
          3381 => x"84",
          3382 => x"ba",
          3383 => x"13",
          3384 => x"ba",
          3385 => x"73",
          3386 => x"16",
          3387 => x"2b",
          3388 => x"2a",
          3389 => x"75",
          3390 => x"86",
          3391 => x"2b",
          3392 => x"16",
          3393 => x"07",
          3394 => x"53",
          3395 => x"85",
          3396 => x"16",
          3397 => x"8b",
          3398 => x"5a",
          3399 => x"13",
          3400 => x"2a",
          3401 => x"34",
          3402 => x"08",
          3403 => x"88",
          3404 => x"88",
          3405 => x"34",
          3406 => x"08",
          3407 => x"71",
          3408 => x"05",
          3409 => x"2b",
          3410 => x"06",
          3411 => x"53",
          3412 => x"82",
          3413 => x"ba",
          3414 => x"12",
          3415 => x"07",
          3416 => x"71",
          3417 => x"70",
          3418 => x"57",
          3419 => x"14",
          3420 => x"82",
          3421 => x"2b",
          3422 => x"33",
          3423 => x"90",
          3424 => x"57",
          3425 => x"38",
          3426 => x"2b",
          3427 => x"2a",
          3428 => x"81",
          3429 => x"17",
          3430 => x"2b",
          3431 => x"14",
          3432 => x"07",
          3433 => x"58",
          3434 => x"75",
          3435 => x"f9",
          3436 => x"58",
          3437 => x"80",
          3438 => x"3f",
          3439 => x"0b",
          3440 => x"84",
          3441 => x"76",
          3442 => x"ed",
          3443 => x"75",
          3444 => x"ba",
          3445 => x"81",
          3446 => x"08",
          3447 => x"87",
          3448 => x"ba",
          3449 => x"07",
          3450 => x"2a",
          3451 => x"34",
          3452 => x"22",
          3453 => x"08",
          3454 => x"15",
          3455 => x"ee",
          3456 => x"53",
          3457 => x"fb",
          3458 => x"ff",
          3459 => x"ff",
          3460 => x"33",
          3461 => x"70",
          3462 => x"ff",
          3463 => x"75",
          3464 => x"12",
          3465 => x"ff",
          3466 => x"ff",
          3467 => x"5c",
          3468 => x"70",
          3469 => x"58",
          3470 => x"88",
          3471 => x"73",
          3472 => x"74",
          3473 => x"11",
          3474 => x"2b",
          3475 => x"56",
          3476 => x"83",
          3477 => x"26",
          3478 => x"2e",
          3479 => x"88",
          3480 => x"11",
          3481 => x"2a",
          3482 => x"34",
          3483 => x"08",
          3484 => x"82",
          3485 => x"ba",
          3486 => x"12",
          3487 => x"2b",
          3488 => x"83",
          3489 => x"58",
          3490 => x"12",
          3491 => x"83",
          3492 => x"54",
          3493 => x"84",
          3494 => x"33",
          3495 => x"83",
          3496 => x"53",
          3497 => x"15",
          3498 => x"55",
          3499 => x"33",
          3500 => x"54",
          3501 => x"71",
          3502 => x"70",
          3503 => x"71",
          3504 => x"05",
          3505 => x"15",
          3506 => x"f4",
          3507 => x"11",
          3508 => x"07",
          3509 => x"70",
          3510 => x"84",
          3511 => x"70",
          3512 => x"04",
          3513 => x"8b",
          3514 => x"84",
          3515 => x"2b",
          3516 => x"53",
          3517 => x"85",
          3518 => x"19",
          3519 => x"8b",
          3520 => x"86",
          3521 => x"2b",
          3522 => x"52",
          3523 => x"34",
          3524 => x"08",
          3525 => x"88",
          3526 => x"88",
          3527 => x"34",
          3528 => x"08",
          3529 => x"f9",
          3530 => x"58",
          3531 => x"54",
          3532 => x"0c",
          3533 => x"91",
          3534 => x"84",
          3535 => x"f4",
          3536 => x"0b",
          3537 => x"53",
          3538 => x"cb",
          3539 => x"76",
          3540 => x"84",
          3541 => x"34",
          3542 => x"f4",
          3543 => x"0b",
          3544 => x"84",
          3545 => x"80",
          3546 => x"88",
          3547 => x"17",
          3548 => x"f0",
          3549 => x"f4",
          3550 => x"82",
          3551 => x"77",
          3552 => x"fe",
          3553 => x"41",
          3554 => x"59",
          3555 => x"38",
          3556 => x"80",
          3557 => x"60",
          3558 => x"2a",
          3559 => x"55",
          3560 => x"78",
          3561 => x"06",
          3562 => x"81",
          3563 => x"75",
          3564 => x"10",
          3565 => x"61",
          3566 => x"88",
          3567 => x"2c",
          3568 => x"43",
          3569 => x"42",
          3570 => x"15",
          3571 => x"07",
          3572 => x"81",
          3573 => x"2b",
          3574 => x"80",
          3575 => x"27",
          3576 => x"62",
          3577 => x"85",
          3578 => x"25",
          3579 => x"79",
          3580 => x"33",
          3581 => x"83",
          3582 => x"12",
          3583 => x"07",
          3584 => x"58",
          3585 => x"1e",
          3586 => x"8b",
          3587 => x"86",
          3588 => x"2b",
          3589 => x"14",
          3590 => x"07",
          3591 => x"5b",
          3592 => x"84",
          3593 => x"ba",
          3594 => x"85",
          3595 => x"2b",
          3596 => x"15",
          3597 => x"2a",
          3598 => x"57",
          3599 => x"34",
          3600 => x"81",
          3601 => x"ff",
          3602 => x"5e",
          3603 => x"34",
          3604 => x"11",
          3605 => x"71",
          3606 => x"81",
          3607 => x"88",
          3608 => x"55",
          3609 => x"34",
          3610 => x"33",
          3611 => x"83",
          3612 => x"83",
          3613 => x"88",
          3614 => x"55",
          3615 => x"1a",
          3616 => x"82",
          3617 => x"2b",
          3618 => x"2b",
          3619 => x"05",
          3620 => x"f4",
          3621 => x"1c",
          3622 => x"5f",
          3623 => x"54",
          3624 => x"0d",
          3625 => x"f4",
          3626 => x"23",
          3627 => x"ff",
          3628 => x"ba",
          3629 => x"0b",
          3630 => x"5d",
          3631 => x"1e",
          3632 => x"86",
          3633 => x"84",
          3634 => x"ff",
          3635 => x"ff",
          3636 => x"5b",
          3637 => x"18",
          3638 => x"10",
          3639 => x"05",
          3640 => x"0b",
          3641 => x"57",
          3642 => x"82",
          3643 => x"fe",
          3644 => x"84",
          3645 => x"95",
          3646 => x"f4",
          3647 => x"44",
          3648 => x"71",
          3649 => x"70",
          3650 => x"63",
          3651 => x"84",
          3652 => x"57",
          3653 => x"19",
          3654 => x"70",
          3655 => x"07",
          3656 => x"74",
          3657 => x"88",
          3658 => x"5d",
          3659 => x"ff",
          3660 => x"84",
          3661 => x"34",
          3662 => x"f4",
          3663 => x"3f",
          3664 => x"31",
          3665 => x"fa",
          3666 => x"76",
          3667 => x"17",
          3668 => x"07",
          3669 => x"81",
          3670 => x"2b",
          3671 => x"45",
          3672 => x"ff",
          3673 => x"38",
          3674 => x"83",
          3675 => x"fc",
          3676 => x"f4",
          3677 => x"0b",
          3678 => x"53",
          3679 => x"c3",
          3680 => x"7e",
          3681 => x"84",
          3682 => x"34",
          3683 => x"f4",
          3684 => x"0b",
          3685 => x"84",
          3686 => x"80",
          3687 => x"88",
          3688 => x"88",
          3689 => x"84",
          3690 => x"84",
          3691 => x"43",
          3692 => x"83",
          3693 => x"24",
          3694 => x"06",
          3695 => x"fc",
          3696 => x"38",
          3697 => x"73",
          3698 => x"04",
          3699 => x"33",
          3700 => x"7a",
          3701 => x"71",
          3702 => x"05",
          3703 => x"88",
          3704 => x"45",
          3705 => x"56",
          3706 => x"85",
          3707 => x"17",
          3708 => x"8b",
          3709 => x"86",
          3710 => x"2b",
          3711 => x"48",
          3712 => x"05",
          3713 => x"ba",
          3714 => x"33",
          3715 => x"06",
          3716 => x"7b",
          3717 => x"ba",
          3718 => x"83",
          3719 => x"2b",
          3720 => x"33",
          3721 => x"5e",
          3722 => x"76",
          3723 => x"ba",
          3724 => x"12",
          3725 => x"07",
          3726 => x"33",
          3727 => x"40",
          3728 => x"78",
          3729 => x"84",
          3730 => x"33",
          3731 => x"66",
          3732 => x"52",
          3733 => x"fe",
          3734 => x"1e",
          3735 => x"5c",
          3736 => x"0b",
          3737 => x"84",
          3738 => x"7f",
          3739 => x"a5",
          3740 => x"76",
          3741 => x"ba",
          3742 => x"81",
          3743 => x"08",
          3744 => x"87",
          3745 => x"ba",
          3746 => x"07",
          3747 => x"2a",
          3748 => x"34",
          3749 => x"22",
          3750 => x"08",
          3751 => x"1c",
          3752 => x"51",
          3753 => x"39",
          3754 => x"8b",
          3755 => x"84",
          3756 => x"2b",
          3757 => x"43",
          3758 => x"63",
          3759 => x"08",
          3760 => x"33",
          3761 => x"74",
          3762 => x"71",
          3763 => x"5f",
          3764 => x"64",
          3765 => x"34",
          3766 => x"81",
          3767 => x"ff",
          3768 => x"58",
          3769 => x"34",
          3770 => x"33",
          3771 => x"83",
          3772 => x"12",
          3773 => x"2b",
          3774 => x"88",
          3775 => x"5d",
          3776 => x"83",
          3777 => x"1f",
          3778 => x"2b",
          3779 => x"33",
          3780 => x"81",
          3781 => x"5d",
          3782 => x"60",
          3783 => x"83",
          3784 => x"86",
          3785 => x"2b",
          3786 => x"18",
          3787 => x"07",
          3788 => x"41",
          3789 => x"1e",
          3790 => x"84",
          3791 => x"2b",
          3792 => x"14",
          3793 => x"07",
          3794 => x"5a",
          3795 => x"34",
          3796 => x"f4",
          3797 => x"71",
          3798 => x"70",
          3799 => x"75",
          3800 => x"f4",
          3801 => x"33",
          3802 => x"74",
          3803 => x"88",
          3804 => x"f8",
          3805 => x"54",
          3806 => x"7f",
          3807 => x"84",
          3808 => x"81",
          3809 => x"2b",
          3810 => x"33",
          3811 => x"06",
          3812 => x"5b",
          3813 => x"81",
          3814 => x"1f",
          3815 => x"8b",
          3816 => x"86",
          3817 => x"2b",
          3818 => x"14",
          3819 => x"07",
          3820 => x"5c",
          3821 => x"77",
          3822 => x"84",
          3823 => x"33",
          3824 => x"83",
          3825 => x"87",
          3826 => x"88",
          3827 => x"41",
          3828 => x"16",
          3829 => x"33",
          3830 => x"81",
          3831 => x"5c",
          3832 => x"1a",
          3833 => x"82",
          3834 => x"2b",
          3835 => x"33",
          3836 => x"70",
          3837 => x"5a",
          3838 => x"1a",
          3839 => x"70",
          3840 => x"71",
          3841 => x"33",
          3842 => x"70",
          3843 => x"5a",
          3844 => x"83",
          3845 => x"1f",
          3846 => x"88",
          3847 => x"83",
          3848 => x"84",
          3849 => x"ba",
          3850 => x"05",
          3851 => x"44",
          3852 => x"87",
          3853 => x"2b",
          3854 => x"1d",
          3855 => x"2a",
          3856 => x"61",
          3857 => x"34",
          3858 => x"11",
          3859 => x"71",
          3860 => x"33",
          3861 => x"70",
          3862 => x"59",
          3863 => x"7a",
          3864 => x"08",
          3865 => x"88",
          3866 => x"88",
          3867 => x"34",
          3868 => x"08",
          3869 => x"71",
          3870 => x"05",
          3871 => x"2b",
          3872 => x"06",
          3873 => x"5c",
          3874 => x"82",
          3875 => x"ba",
          3876 => x"12",
          3877 => x"07",
          3878 => x"71",
          3879 => x"70",
          3880 => x"59",
          3881 => x"1e",
          3882 => x"f3",
          3883 => x"a1",
          3884 => x"bb",
          3885 => x"53",
          3886 => x"fe",
          3887 => x"3f",
          3888 => x"38",
          3889 => x"7a",
          3890 => x"76",
          3891 => x"8a",
          3892 => x"3d",
          3893 => x"84",
          3894 => x"08",
          3895 => x"52",
          3896 => x"bd",
          3897 => x"3d",
          3898 => x"ba",
          3899 => x"f0",
          3900 => x"84",
          3901 => x"84",
          3902 => x"81",
          3903 => x"08",
          3904 => x"85",
          3905 => x"76",
          3906 => x"34",
          3907 => x"22",
          3908 => x"83",
          3909 => x"51",
          3910 => x"89",
          3911 => x"10",
          3912 => x"f8",
          3913 => x"81",
          3914 => x"80",
          3915 => x"ff",
          3916 => x"81",
          3917 => x"bb",
          3918 => x"84",
          3919 => x"0d",
          3920 => x"71",
          3921 => x"bb",
          3922 => x"06",
          3923 => x"80",
          3924 => x"53",
          3925 => x"0d",
          3926 => x"02",
          3927 => x"57",
          3928 => x"38",
          3929 => x"81",
          3930 => x"73",
          3931 => x"0c",
          3932 => x"ca",
          3933 => x"06",
          3934 => x"c0",
          3935 => x"79",
          3936 => x"80",
          3937 => x"81",
          3938 => x"0c",
          3939 => x"81",
          3940 => x"56",
          3941 => x"39",
          3942 => x"8c",
          3943 => x"59",
          3944 => x"84",
          3945 => x"06",
          3946 => x"58",
          3947 => x"78",
          3948 => x"3f",
          3949 => x"55",
          3950 => x"98",
          3951 => x"78",
          3952 => x"06",
          3953 => x"54",
          3954 => x"8b",
          3955 => x"19",
          3956 => x"79",
          3957 => x"fc",
          3958 => x"05",
          3959 => x"53",
          3960 => x"87",
          3961 => x"72",
          3962 => x"38",
          3963 => x"81",
          3964 => x"71",
          3965 => x"38",
          3966 => x"86",
          3967 => x"0c",
          3968 => x"0d",
          3969 => x"84",
          3970 => x"71",
          3971 => x"53",
          3972 => x"81",
          3973 => x"2e",
          3974 => x"55",
          3975 => x"08",
          3976 => x"87",
          3977 => x"82",
          3978 => x"38",
          3979 => x"38",
          3980 => x"58",
          3981 => x"56",
          3982 => x"a8",
          3983 => x"81",
          3984 => x"18",
          3985 => x"84",
          3986 => x"78",
          3987 => x"04",
          3988 => x"18",
          3989 => x"fc",
          3990 => x"08",
          3991 => x"84",
          3992 => x"18",
          3993 => x"1a",
          3994 => x"56",
          3995 => x"82",
          3996 => x"81",
          3997 => x"1b",
          3998 => x"fc",
          3999 => x"75",
          4000 => x"38",
          4001 => x"09",
          4002 => x"5a",
          4003 => x"70",
          4004 => x"76",
          4005 => x"19",
          4006 => x"34",
          4007 => x"b9",
          4008 => x"34",
          4009 => x"f2",
          4010 => x"0b",
          4011 => x"84",
          4012 => x"9f",
          4013 => x"84",
          4014 => x"7a",
          4015 => x"56",
          4016 => x"2a",
          4017 => x"18",
          4018 => x"7a",
          4019 => x"34",
          4020 => x"19",
          4021 => x"a7",
          4022 => x"70",
          4023 => x"53",
          4024 => x"e8",
          4025 => x"80",
          4026 => x"3f",
          4027 => x"b7",
          4028 => x"60",
          4029 => x"76",
          4030 => x"26",
          4031 => x"84",
          4032 => x"33",
          4033 => x"38",
          4034 => x"81",
          4035 => x"81",
          4036 => x"08",
          4037 => x"08",
          4038 => x"5c",
          4039 => x"de",
          4040 => x"52",
          4041 => x"84",
          4042 => x"ff",
          4043 => x"7a",
          4044 => x"17",
          4045 => x"2a",
          4046 => x"59",
          4047 => x"80",
          4048 => x"5d",
          4049 => x"b5",
          4050 => x"52",
          4051 => x"84",
          4052 => x"ff",
          4053 => x"79",
          4054 => x"17",
          4055 => x"07",
          4056 => x"5d",
          4057 => x"76",
          4058 => x"8f",
          4059 => x"18",
          4060 => x"2e",
          4061 => x"71",
          4062 => x"81",
          4063 => x"53",
          4064 => x"f7",
          4065 => x"2e",
          4066 => x"b4",
          4067 => x"10",
          4068 => x"81",
          4069 => x"07",
          4070 => x"3d",
          4071 => x"06",
          4072 => x"18",
          4073 => x"2e",
          4074 => x"71",
          4075 => x"81",
          4076 => x"53",
          4077 => x"f6",
          4078 => x"2e",
          4079 => x"b4",
          4080 => x"82",
          4081 => x"05",
          4082 => x"90",
          4083 => x"33",
          4084 => x"71",
          4085 => x"84",
          4086 => x"5a",
          4087 => x"b4",
          4088 => x"81",
          4089 => x"81",
          4090 => x"09",
          4091 => x"84",
          4092 => x"a8",
          4093 => x"5b",
          4094 => x"84",
          4095 => x"2e",
          4096 => x"54",
          4097 => x"53",
          4098 => x"98",
          4099 => x"54",
          4100 => x"53",
          4101 => x"3f",
          4102 => x"81",
          4103 => x"08",
          4104 => x"18",
          4105 => x"27",
          4106 => x"82",
          4107 => x"08",
          4108 => x"17",
          4109 => x"18",
          4110 => x"5a",
          4111 => x"81",
          4112 => x"08",
          4113 => x"18",
          4114 => x"5e",
          4115 => x"38",
          4116 => x"09",
          4117 => x"b4",
          4118 => x"7b",
          4119 => x"3f",
          4120 => x"b4",
          4121 => x"81",
          4122 => x"81",
          4123 => x"09",
          4124 => x"84",
          4125 => x"a8",
          4126 => x"5b",
          4127 => x"91",
          4128 => x"2e",
          4129 => x"54",
          4130 => x"53",
          4131 => x"90",
          4132 => x"54",
          4133 => x"53",
          4134 => x"f8",
          4135 => x"f9",
          4136 => x"0d",
          4137 => x"58",
          4138 => x"1a",
          4139 => x"74",
          4140 => x"81",
          4141 => x"38",
          4142 => x"0d",
          4143 => x"05",
          4144 => x"5c",
          4145 => x"19",
          4146 => x"09",
          4147 => x"77",
          4148 => x"51",
          4149 => x"80",
          4150 => x"77",
          4151 => x"b0",
          4152 => x"05",
          4153 => x"76",
          4154 => x"79",
          4155 => x"34",
          4156 => x"0d",
          4157 => x"fe",
          4158 => x"08",
          4159 => x"58",
          4160 => x"83",
          4161 => x"2e",
          4162 => x"54",
          4163 => x"33",
          4164 => x"08",
          4165 => x"5a",
          4166 => x"fe",
          4167 => x"06",
          4168 => x"70",
          4169 => x"0a",
          4170 => x"7d",
          4171 => x"1d",
          4172 => x"1d",
          4173 => x"1d",
          4174 => x"e8",
          4175 => x"2a",
          4176 => x"59",
          4177 => x"80",
          4178 => x"5d",
          4179 => x"d4",
          4180 => x"52",
          4181 => x"84",
          4182 => x"ff",
          4183 => x"7b",
          4184 => x"ff",
          4185 => x"81",
          4186 => x"80",
          4187 => x"f0",
          4188 => x"56",
          4189 => x"1a",
          4190 => x"05",
          4191 => x"5f",
          4192 => x"54",
          4193 => x"1a",
          4194 => x"58",
          4195 => x"81",
          4196 => x"08",
          4197 => x"a8",
          4198 => x"bb",
          4199 => x"7a",
          4200 => x"74",
          4201 => x"75",
          4202 => x"ee",
          4203 => x"2e",
          4204 => x"b4",
          4205 => x"83",
          4206 => x"2a",
          4207 => x"2a",
          4208 => x"06",
          4209 => x"0b",
          4210 => x"54",
          4211 => x"1a",
          4212 => x"5a",
          4213 => x"81",
          4214 => x"08",
          4215 => x"a8",
          4216 => x"bb",
          4217 => x"77",
          4218 => x"55",
          4219 => x"bd",
          4220 => x"52",
          4221 => x"7b",
          4222 => x"53",
          4223 => x"52",
          4224 => x"bb",
          4225 => x"fd",
          4226 => x"1a",
          4227 => x"08",
          4228 => x"08",
          4229 => x"fc",
          4230 => x"82",
          4231 => x"81",
          4232 => x"19",
          4233 => x"fc",
          4234 => x"19",
          4235 => x"ed",
          4236 => x"08",
          4237 => x"38",
          4238 => x"b4",
          4239 => x"a0",
          4240 => x"5f",
          4241 => x"38",
          4242 => x"09",
          4243 => x"7c",
          4244 => x"51",
          4245 => x"39",
          4246 => x"81",
          4247 => x"58",
          4248 => x"fe",
          4249 => x"06",
          4250 => x"76",
          4251 => x"f9",
          4252 => x"7b",
          4253 => x"05",
          4254 => x"2b",
          4255 => x"07",
          4256 => x"34",
          4257 => x"34",
          4258 => x"34",
          4259 => x"34",
          4260 => x"7e",
          4261 => x"8a",
          4262 => x"2e",
          4263 => x"27",
          4264 => x"56",
          4265 => x"76",
          4266 => x"81",
          4267 => x"89",
          4268 => x"b2",
          4269 => x"3f",
          4270 => x"d0",
          4271 => x"81",
          4272 => x"09",
          4273 => x"70",
          4274 => x"82",
          4275 => x"06",
          4276 => x"bb",
          4277 => x"57",
          4278 => x"58",
          4279 => x"a4",
          4280 => x"08",
          4281 => x"55",
          4282 => x"38",
          4283 => x"26",
          4284 => x"81",
          4285 => x"83",
          4286 => x"ef",
          4287 => x"08",
          4288 => x"84",
          4289 => x"80",
          4290 => x"08",
          4291 => x"85",
          4292 => x"9a",
          4293 => x"27",
          4294 => x"27",
          4295 => x"fe",
          4296 => x"38",
          4297 => x"f5",
          4298 => x"84",
          4299 => x"07",
          4300 => x"c4",
          4301 => x"1a",
          4302 => x"1a",
          4303 => x"38",
          4304 => x"33",
          4305 => x"75",
          4306 => x"3d",
          4307 => x"0c",
          4308 => x"08",
          4309 => x"ff",
          4310 => x"51",
          4311 => x"55",
          4312 => x"84",
          4313 => x"ff",
          4314 => x"81",
          4315 => x"7a",
          4316 => x"f0",
          4317 => x"9f",
          4318 => x"90",
          4319 => x"80",
          4320 => x"26",
          4321 => x"82",
          4322 => x"79",
          4323 => x"19",
          4324 => x"08",
          4325 => x"38",
          4326 => x"73",
          4327 => x"19",
          4328 => x"0c",
          4329 => x"bb",
          4330 => x"17",
          4331 => x"38",
          4332 => x"59",
          4333 => x"08",
          4334 => x"80",
          4335 => x"17",
          4336 => x"05",
          4337 => x"91",
          4338 => x"3f",
          4339 => x"84",
          4340 => x"84",
          4341 => x"9c",
          4342 => x"73",
          4343 => x"54",
          4344 => x"39",
          4345 => x"3d",
          4346 => x"08",
          4347 => x"57",
          4348 => x"80",
          4349 => x"55",
          4350 => x"79",
          4351 => x"81",
          4352 => x"a9",
          4353 => x"57",
          4354 => x"77",
          4355 => x"78",
          4356 => x"56",
          4357 => x"0d",
          4358 => x"22",
          4359 => x"7b",
          4360 => x"9c",
          4361 => x"56",
          4362 => x"d0",
          4363 => x"ff",
          4364 => x"bb",
          4365 => x"80",
          4366 => x"52",
          4367 => x"84",
          4368 => x"08",
          4369 => x"84",
          4370 => x"38",
          4371 => x"2e",
          4372 => x"83",
          4373 => x"38",
          4374 => x"59",
          4375 => x"38",
          4376 => x"1b",
          4377 => x"0c",
          4378 => x"55",
          4379 => x"ff",
          4380 => x"8a",
          4381 => x"80",
          4382 => x"52",
          4383 => x"84",
          4384 => x"16",
          4385 => x"84",
          4386 => x"0d",
          4387 => x"b8",
          4388 => x"56",
          4389 => x"80",
          4390 => x"1a",
          4391 => x"31",
          4392 => x"e8",
          4393 => x"2e",
          4394 => x"54",
          4395 => x"53",
          4396 => x"c8",
          4397 => x"55",
          4398 => x"76",
          4399 => x"94",
          4400 => x"fe",
          4401 => x"27",
          4402 => x"71",
          4403 => x"0c",
          4404 => x"bb",
          4405 => x"3d",
          4406 => x"08",
          4407 => x"08",
          4408 => x"d2",
          4409 => x"58",
          4410 => x"38",
          4411 => x"78",
          4412 => x"81",
          4413 => x"19",
          4414 => x"84",
          4415 => x"81",
          4416 => x"76",
          4417 => x"33",
          4418 => x"38",
          4419 => x"ff",
          4420 => x"76",
          4421 => x"32",
          4422 => x"25",
          4423 => x"93",
          4424 => x"61",
          4425 => x"2e",
          4426 => x"52",
          4427 => x"84",
          4428 => x"b2",
          4429 => x"dc",
          4430 => x"3d",
          4431 => x"53",
          4432 => x"a8",
          4433 => x"78",
          4434 => x"84",
          4435 => x"19",
          4436 => x"84",
          4437 => x"27",
          4438 => x"60",
          4439 => x"38",
          4440 => x"08",
          4441 => x"51",
          4442 => x"39",
          4443 => x"e7",
          4444 => x"7a",
          4445 => x"77",
          4446 => x"7f",
          4447 => x"7d",
          4448 => x"5d",
          4449 => x"2e",
          4450 => x"39",
          4451 => x"7a",
          4452 => x"04",
          4453 => x"33",
          4454 => x"cb",
          4455 => x"9a",
          4456 => x"56",
          4457 => x"70",
          4458 => x"51",
          4459 => x"84",
          4460 => x"71",
          4461 => x"56",
          4462 => x"81",
          4463 => x"61",
          4464 => x"81",
          4465 => x"27",
          4466 => x"81",
          4467 => x"38",
          4468 => x"79",
          4469 => x"ff",
          4470 => x"fd",
          4471 => x"ca",
          4472 => x"7c",
          4473 => x"81",
          4474 => x"70",
          4475 => x"70",
          4476 => x"59",
          4477 => x"81",
          4478 => x"84",
          4479 => x"ef",
          4480 => x"80",
          4481 => x"bb",
          4482 => x"82",
          4483 => x"ff",
          4484 => x"98",
          4485 => x"08",
          4486 => x"33",
          4487 => x"81",
          4488 => x"53",
          4489 => x"dc",
          4490 => x"2e",
          4491 => x"b4",
          4492 => x"38",
          4493 => x"76",
          4494 => x"33",
          4495 => x"58",
          4496 => x"2e",
          4497 => x"06",
          4498 => x"74",
          4499 => x"e5",
          4500 => x"58",
          4501 => x"80",
          4502 => x"33",
          4503 => x"ff",
          4504 => x"74",
          4505 => x"33",
          4506 => x"0b",
          4507 => x"05",
          4508 => x"33",
          4509 => x"42",
          4510 => x"75",
          4511 => x"ff",
          4512 => x"51",
          4513 => x"5a",
          4514 => x"8f",
          4515 => x"3d",
          4516 => x"53",
          4517 => x"80",
          4518 => x"78",
          4519 => x"84",
          4520 => x"1b",
          4521 => x"84",
          4522 => x"27",
          4523 => x"79",
          4524 => x"38",
          4525 => x"08",
          4526 => x"51",
          4527 => x"39",
          4528 => x"33",
          4529 => x"60",
          4530 => x"06",
          4531 => x"19",
          4532 => x"1f",
          4533 => x"5f",
          4534 => x"55",
          4535 => x"92",
          4536 => x"bb",
          4537 => x"fe",
          4538 => x"38",
          4539 => x"0c",
          4540 => x"7e",
          4541 => x"8c",
          4542 => x"33",
          4543 => x"76",
          4544 => x"06",
          4545 => x"77",
          4546 => x"79",
          4547 => x"88",
          4548 => x"2e",
          4549 => x"ff",
          4550 => x"3f",
          4551 => x"05",
          4552 => x"56",
          4553 => x"84",
          4554 => x"38",
          4555 => x"27",
          4556 => x"2a",
          4557 => x"92",
          4558 => x"10",
          4559 => x"fe",
          4560 => x"06",
          4561 => x"84",
          4562 => x"76",
          4563 => x"81",
          4564 => x"0d",
          4565 => x"81",
          4566 => x"56",
          4567 => x"08",
          4568 => x"2e",
          4569 => x"70",
          4570 => x"95",
          4571 => x"7b",
          4572 => x"57",
          4573 => x"ff",
          4574 => x"db",
          4575 => x"76",
          4576 => x"0b",
          4577 => x"40",
          4578 => x"8b",
          4579 => x"81",
          4580 => x"58",
          4581 => x"85",
          4582 => x"22",
          4583 => x"74",
          4584 => x"81",
          4585 => x"70",
          4586 => x"81",
          4587 => x"2e",
          4588 => x"57",
          4589 => x"38",
          4590 => x"02",
          4591 => x"76",
          4592 => x"27",
          4593 => x"34",
          4594 => x"59",
          4595 => x"59",
          4596 => x"56",
          4597 => x"55",
          4598 => x"56",
          4599 => x"1a",
          4600 => x"09",
          4601 => x"a0",
          4602 => x"3d",
          4603 => x"33",
          4604 => x"76",
          4605 => x"8f",
          4606 => x"81",
          4607 => x"91",
          4608 => x"82",
          4609 => x"84",
          4610 => x"06",
          4611 => x"33",
          4612 => x"05",
          4613 => x"81",
          4614 => x"80",
          4615 => x"51",
          4616 => x"08",
          4617 => x"8c",
          4618 => x"bb",
          4619 => x"84",
          4620 => x"08",
          4621 => x"2e",
          4622 => x"7f",
          4623 => x"38",
          4624 => x"81",
          4625 => x"bb",
          4626 => x"56",
          4627 => x"56",
          4628 => x"33",
          4629 => x"c9",
          4630 => x"07",
          4631 => x"38",
          4632 => x"89",
          4633 => x"3f",
          4634 => x"84",
          4635 => x"58",
          4636 => x"58",
          4637 => x"7f",
          4638 => x"b4",
          4639 => x"1c",
          4640 => x"38",
          4641 => x"81",
          4642 => x"bb",
          4643 => x"57",
          4644 => x"58",
          4645 => x"1f",
          4646 => x"05",
          4647 => x"38",
          4648 => x"58",
          4649 => x"77",
          4650 => x"55",
          4651 => x"1f",
          4652 => x"1b",
          4653 => x"56",
          4654 => x"0d",
          4655 => x"72",
          4656 => x"38",
          4657 => x"c2",
          4658 => x"bb",
          4659 => x"fe",
          4660 => x"53",
          4661 => x"80",
          4662 => x"09",
          4663 => x"84",
          4664 => x"a8",
          4665 => x"08",
          4666 => x"60",
          4667 => x"84",
          4668 => x"2b",
          4669 => x"7d",
          4670 => x"08",
          4671 => x"38",
          4672 => x"8b",
          4673 => x"29",
          4674 => x"57",
          4675 => x"19",
          4676 => x"81",
          4677 => x"1e",
          4678 => x"77",
          4679 => x"7a",
          4680 => x"38",
          4681 => x"81",
          4682 => x"bb",
          4683 => x"57",
          4684 => x"58",
          4685 => x"9c",
          4686 => x"5c",
          4687 => x"8b",
          4688 => x"9a",
          4689 => x"8d",
          4690 => x"59",
          4691 => x"78",
          4692 => x"58",
          4693 => x"05",
          4694 => x"34",
          4695 => x"76",
          4696 => x"18",
          4697 => x"83",
          4698 => x"10",
          4699 => x"2e",
          4700 => x"0b",
          4701 => x"e9",
          4702 => x"84",
          4703 => x"ff",
          4704 => x"eb",
          4705 => x"b8",
          4706 => x"59",
          4707 => x"84",
          4708 => x"08",
          4709 => x"1d",
          4710 => x"41",
          4711 => x"38",
          4712 => x"09",
          4713 => x"b4",
          4714 => x"78",
          4715 => x"3f",
          4716 => x"1f",
          4717 => x"81",
          4718 => x"38",
          4719 => x"76",
          4720 => x"39",
          4721 => x"39",
          4722 => x"52",
          4723 => x"84",
          4724 => x"06",
          4725 => x"1d",
          4726 => x"31",
          4727 => x"38",
          4728 => x"aa",
          4729 => x"f8",
          4730 => x"80",
          4731 => x"75",
          4732 => x"59",
          4733 => x"fa",
          4734 => x"a0",
          4735 => x"1c",
          4736 => x"39",
          4737 => x"08",
          4738 => x"51",
          4739 => x"3d",
          4740 => x"5c",
          4741 => x"08",
          4742 => x"08",
          4743 => x"71",
          4744 => x"58",
          4745 => x"38",
          4746 => x"1b",
          4747 => x"80",
          4748 => x"06",
          4749 => x"83",
          4750 => x"22",
          4751 => x"7a",
          4752 => x"06",
          4753 => x"57",
          4754 => x"89",
          4755 => x"16",
          4756 => x"74",
          4757 => x"81",
          4758 => x"70",
          4759 => x"77",
          4760 => x"8b",
          4761 => x"34",
          4762 => x"05",
          4763 => x"27",
          4764 => x"55",
          4765 => x"33",
          4766 => x"38",
          4767 => x"7c",
          4768 => x"17",
          4769 => x"55",
          4770 => x"34",
          4771 => x"88",
          4772 => x"83",
          4773 => x"2b",
          4774 => x"70",
          4775 => x"07",
          4776 => x"17",
          4777 => x"5b",
          4778 => x"1e",
          4779 => x"71",
          4780 => x"1e",
          4781 => x"55",
          4782 => x"81",
          4783 => x"b5",
          4784 => x"81",
          4785 => x"83",
          4786 => x"27",
          4787 => x"38",
          4788 => x"74",
          4789 => x"80",
          4790 => x"19",
          4791 => x"79",
          4792 => x"30",
          4793 => x"72",
          4794 => x"80",
          4795 => x"05",
          4796 => x"5b",
          4797 => x"5a",
          4798 => x"38",
          4799 => x"89",
          4800 => x"78",
          4801 => x"8c",
          4802 => x"b4",
          4803 => x"06",
          4804 => x"14",
          4805 => x"73",
          4806 => x"16",
          4807 => x"33",
          4808 => x"b7",
          4809 => x"53",
          4810 => x"25",
          4811 => x"58",
          4812 => x"70",
          4813 => x"70",
          4814 => x"83",
          4815 => x"81",
          4816 => x"38",
          4817 => x"33",
          4818 => x"9f",
          4819 => x"8c",
          4820 => x"70",
          4821 => x"81",
          4822 => x"2e",
          4823 => x"27",
          4824 => x"76",
          4825 => x"ff",
          4826 => x"73",
          4827 => x"5b",
          4828 => x"dc",
          4829 => x"26",
          4830 => x"e6",
          4831 => x"54",
          4832 => x"73",
          4833 => x"33",
          4834 => x"73",
          4835 => x"7a",
          4836 => x"80",
          4837 => x"7d",
          4838 => x"05",
          4839 => x"2e",
          4840 => x"73",
          4841 => x"25",
          4842 => x"80",
          4843 => x"54",
          4844 => x"2e",
          4845 => x"30",
          4846 => x"57",
          4847 => x"73",
          4848 => x"55",
          4849 => x"39",
          4850 => x"ae",
          4851 => x"ff",
          4852 => x"54",
          4853 => x"0d",
          4854 => x"ff",
          4855 => x"e3",
          4856 => x"1d",
          4857 => x"3f",
          4858 => x"0c",
          4859 => x"dc",
          4860 => x"07",
          4861 => x"a1",
          4862 => x"33",
          4863 => x"38",
          4864 => x"80",
          4865 => x"e1",
          4866 => x"82",
          4867 => x"38",
          4868 => x"17",
          4869 => x"17",
          4870 => x"a0",
          4871 => x"42",
          4872 => x"84",
          4873 => x"76",
          4874 => x"80",
          4875 => x"38",
          4876 => x"06",
          4877 => x"2e",
          4878 => x"06",
          4879 => x"76",
          4880 => x"05",
          4881 => x"9d",
          4882 => x"ff",
          4883 => x"fe",
          4884 => x"2e",
          4885 => x"a0",
          4886 => x"05",
          4887 => x"38",
          4888 => x"70",
          4889 => x"74",
          4890 => x"2e",
          4891 => x"30",
          4892 => x"77",
          4893 => x"38",
          4894 => x"81",
          4895 => x"72",
          4896 => x"51",
          4897 => x"38",
          4898 => x"77",
          4899 => x"75",
          4900 => x"5b",
          4901 => x"77",
          4902 => x"22",
          4903 => x"95",
          4904 => x"e5",
          4905 => x"82",
          4906 => x"8c",
          4907 => x"55",
          4908 => x"81",
          4909 => x"7d",
          4910 => x"38",
          4911 => x"81",
          4912 => x"79",
          4913 => x"7b",
          4914 => x"08",
          4915 => x"84",
          4916 => x"bb",
          4917 => x"fb",
          4918 => x"5a",
          4919 => x"82",
          4920 => x"38",
          4921 => x"8c",
          4922 => x"39",
          4923 => x"22",
          4924 => x"f0",
          4925 => x"79",
          4926 => x"18",
          4927 => x"06",
          4928 => x"ae",
          4929 => x"76",
          4930 => x"0b",
          4931 => x"73",
          4932 => x"70",
          4933 => x"8a",
          4934 => x"58",
          4935 => x"bf",
          4936 => x"33",
          4937 => x"d6",
          4938 => x"77",
          4939 => x"84",
          4940 => x"2e",
          4941 => x"ff",
          4942 => x"80",
          4943 => x"62",
          4944 => x"2e",
          4945 => x"7b",
          4946 => x"77",
          4947 => x"38",
          4948 => x"fb",
          4949 => x"56",
          4950 => x"81",
          4951 => x"77",
          4952 => x"38",
          4953 => x"85",
          4954 => x"09",
          4955 => x"ff",
          4956 => x"84",
          4957 => x"74",
          4958 => x"75",
          4959 => x"78",
          4960 => x"07",
          4961 => x"a4",
          4962 => x"52",
          4963 => x"bb",
          4964 => x"87",
          4965 => x"2e",
          4966 => x"e7",
          4967 => x"ff",
          4968 => x"81",
          4969 => x"e6",
          4970 => x"54",
          4971 => x"73",
          4972 => x"33",
          4973 => x"73",
          4974 => x"78",
          4975 => x"73",
          4976 => x"70",
          4977 => x"15",
          4978 => x"81",
          4979 => x"70",
          4980 => x"53",
          4981 => x"34",
          4982 => x"fc",
          4983 => x"e6",
          4984 => x"53",
          4985 => x"df",
          4986 => x"5b",
          4987 => x"5b",
          4988 => x"cc",
          4989 => x"2b",
          4990 => x"57",
          4991 => x"75",
          4992 => x"81",
          4993 => x"74",
          4994 => x"39",
          4995 => x"5a",
          4996 => x"fa",
          4997 => x"2a",
          4998 => x"85",
          4999 => x"0d",
          5000 => x"88",
          5001 => x"5e",
          5002 => x"59",
          5003 => x"38",
          5004 => x"9f",
          5005 => x"d0",
          5006 => x"85",
          5007 => x"80",
          5008 => x"10",
          5009 => x"5a",
          5010 => x"38",
          5011 => x"77",
          5012 => x"38",
          5013 => x"3f",
          5014 => x"70",
          5015 => x"86",
          5016 => x"5d",
          5017 => x"34",
          5018 => x"bb",
          5019 => x"ff",
          5020 => x"58",
          5021 => x"8d",
          5022 => x"8a",
          5023 => x"7a",
          5024 => x"0c",
          5025 => x"53",
          5026 => x"52",
          5027 => x"84",
          5028 => x"81",
          5029 => x"78",
          5030 => x"b6",
          5031 => x"56",
          5032 => x"85",
          5033 => x"84",
          5034 => x"bf",
          5035 => x"cd",
          5036 => x"c5",
          5037 => x"18",
          5038 => x"7c",
          5039 => x"ad",
          5040 => x"18",
          5041 => x"75",
          5042 => x"33",
          5043 => x"88",
          5044 => x"07",
          5045 => x"5a",
          5046 => x"18",
          5047 => x"34",
          5048 => x"81",
          5049 => x"7c",
          5050 => x"ff",
          5051 => x"33",
          5052 => x"77",
          5053 => x"ff",
          5054 => x"38",
          5055 => x"33",
          5056 => x"88",
          5057 => x"5a",
          5058 => x"cc",
          5059 => x"88",
          5060 => x"80",
          5061 => x"33",
          5062 => x"81",
          5063 => x"75",
          5064 => x"42",
          5065 => x"c6",
          5066 => x"58",
          5067 => x"38",
          5068 => x"79",
          5069 => x"74",
          5070 => x"84",
          5071 => x"08",
          5072 => x"84",
          5073 => x"83",
          5074 => x"26",
          5075 => x"26",
          5076 => x"70",
          5077 => x"7b",
          5078 => x"b0",
          5079 => x"8a",
          5080 => x"58",
          5081 => x"16",
          5082 => x"82",
          5083 => x"81",
          5084 => x"83",
          5085 => x"78",
          5086 => x"0b",
          5087 => x"0c",
          5088 => x"83",
          5089 => x"84",
          5090 => x"84",
          5091 => x"84",
          5092 => x"0b",
          5093 => x"bb",
          5094 => x"0b",
          5095 => x"04",
          5096 => x"06",
          5097 => x"38",
          5098 => x"05",
          5099 => x"38",
          5100 => x"40",
          5101 => x"70",
          5102 => x"05",
          5103 => x"56",
          5104 => x"70",
          5105 => x"17",
          5106 => x"17",
          5107 => x"30",
          5108 => x"2e",
          5109 => x"be",
          5110 => x"72",
          5111 => x"55",
          5112 => x"1c",
          5113 => x"ff",
          5114 => x"78",
          5115 => x"2a",
          5116 => x"c5",
          5117 => x"78",
          5118 => x"09",
          5119 => x"81",
          5120 => x"7b",
          5121 => x"38",
          5122 => x"93",
          5123 => x"fa",
          5124 => x"2e",
          5125 => x"80",
          5126 => x"2b",
          5127 => x"07",
          5128 => x"07",
          5129 => x"7a",
          5130 => x"90",
          5131 => x"be",
          5132 => x"30",
          5133 => x"3d",
          5134 => x"b6",
          5135 => x"78",
          5136 => x"80",
          5137 => x"ff",
          5138 => x"56",
          5139 => x"7a",
          5140 => x"51",
          5141 => x"08",
          5142 => x"56",
          5143 => x"bf",
          5144 => x"88",
          5145 => x"82",
          5146 => x"38",
          5147 => x"75",
          5148 => x"81",
          5149 => x"7a",
          5150 => x"75",
          5151 => x"77",
          5152 => x"ba",
          5153 => x"2e",
          5154 => x"81",
          5155 => x"2e",
          5156 => x"5a",
          5157 => x"f8",
          5158 => x"83",
          5159 => x"81",
          5160 => x"40",
          5161 => x"52",
          5162 => x"38",
          5163 => x"81",
          5164 => x"58",
          5165 => x"70",
          5166 => x"ff",
          5167 => x"2e",
          5168 => x"38",
          5169 => x"7c",
          5170 => x"0c",
          5171 => x"80",
          5172 => x"8a",
          5173 => x"ff",
          5174 => x"0c",
          5175 => x"ee",
          5176 => x"78",
          5177 => x"81",
          5178 => x"1b",
          5179 => x"83",
          5180 => x"85",
          5181 => x"5c",
          5182 => x"33",
          5183 => x"71",
          5184 => x"77",
          5185 => x"2e",
          5186 => x"83",
          5187 => x"c6",
          5188 => x"18",
          5189 => x"75",
          5190 => x"38",
          5191 => x"08",
          5192 => x"5b",
          5193 => x"9b",
          5194 => x"52",
          5195 => x"3f",
          5196 => x"38",
          5197 => x"0c",
          5198 => x"34",
          5199 => x"33",
          5200 => x"82",
          5201 => x"fc",
          5202 => x"12",
          5203 => x"07",
          5204 => x"2b",
          5205 => x"45",
          5206 => x"a4",
          5207 => x"38",
          5208 => x"12",
          5209 => x"07",
          5210 => x"2b",
          5211 => x"5b",
          5212 => x"e4",
          5213 => x"38",
          5214 => x"12",
          5215 => x"07",
          5216 => x"2b",
          5217 => x"5d",
          5218 => x"12",
          5219 => x"07",
          5220 => x"2b",
          5221 => x"0c",
          5222 => x"45",
          5223 => x"e2",
          5224 => x"e2",
          5225 => x"e2",
          5226 => x"98",
          5227 => x"24",
          5228 => x"56",
          5229 => x"08",
          5230 => x"33",
          5231 => x"bb",
          5232 => x"81",
          5233 => x"18",
          5234 => x"31",
          5235 => x"38",
          5236 => x"81",
          5237 => x"fd",
          5238 => x"f3",
          5239 => x"83",
          5240 => x"39",
          5241 => x"33",
          5242 => x"58",
          5243 => x"42",
          5244 => x"83",
          5245 => x"2b",
          5246 => x"70",
          5247 => x"07",
          5248 => x"5a",
          5249 => x"39",
          5250 => x"38",
          5251 => x"2e",
          5252 => x"5a",
          5253 => x"79",
          5254 => x"54",
          5255 => x"53",
          5256 => x"ad",
          5257 => x"0d",
          5258 => x"43",
          5259 => x"5a",
          5260 => x"78",
          5261 => x"26",
          5262 => x"38",
          5263 => x"d9",
          5264 => x"74",
          5265 => x"84",
          5266 => x"73",
          5267 => x"62",
          5268 => x"74",
          5269 => x"54",
          5270 => x"93",
          5271 => x"81",
          5272 => x"84",
          5273 => x"8b",
          5274 => x"0d",
          5275 => x"ff",
          5276 => x"91",
          5277 => x"d0",
          5278 => x"f7",
          5279 => x"5e",
          5280 => x"79",
          5281 => x"81",
          5282 => x"57",
          5283 => x"15",
          5284 => x"9f",
          5285 => x"e0",
          5286 => x"74",
          5287 => x"76",
          5288 => x"ff",
          5289 => x"70",
          5290 => x"57",
          5291 => x"1b",
          5292 => x"ff",
          5293 => x"7a",
          5294 => x"0c",
          5295 => x"6c",
          5296 => x"56",
          5297 => x"38",
          5298 => x"cc",
          5299 => x"59",
          5300 => x"57",
          5301 => x"38",
          5302 => x"bb",
          5303 => x"40",
          5304 => x"e1",
          5305 => x"84",
          5306 => x"38",
          5307 => x"81",
          5308 => x"38",
          5309 => x"88",
          5310 => x"83",
          5311 => x"81",
          5312 => x"12",
          5313 => x"33",
          5314 => x"2e",
          5315 => x"34",
          5316 => x"90",
          5317 => x"34",
          5318 => x"7e",
          5319 => x"34",
          5320 => x"5d",
          5321 => x"58",
          5322 => x"9d",
          5323 => x"80",
          5324 => x"0b",
          5325 => x"e2",
          5326 => x"08",
          5327 => x"89",
          5328 => x"ec",
          5329 => x"a3",
          5330 => x"98",
          5331 => x"b8",
          5332 => x"7c",
          5333 => x"02",
          5334 => x"81",
          5335 => x"78",
          5336 => x"2e",
          5337 => x"82",
          5338 => x"56",
          5339 => x"c0",
          5340 => x"1c",
          5341 => x"11",
          5342 => x"07",
          5343 => x"7b",
          5344 => x"1b",
          5345 => x"12",
          5346 => x"07",
          5347 => x"2b",
          5348 => x"0c",
          5349 => x"59",
          5350 => x"78",
          5351 => x"34",
          5352 => x"94",
          5353 => x"7c",
          5354 => x"58",
          5355 => x"78",
          5356 => x"2e",
          5357 => x"74",
          5358 => x"1b",
          5359 => x"88",
          5360 => x"76",
          5361 => x"55",
          5362 => x"70",
          5363 => x"83",
          5364 => x"ac",
          5365 => x"84",
          5366 => x"82",
          5367 => x"b6",
          5368 => x"02",
          5369 => x"7d",
          5370 => x"55",
          5371 => x"57",
          5372 => x"57",
          5373 => x"57",
          5374 => x"76",
          5375 => x"95",
          5376 => x"2b",
          5377 => x"1d",
          5378 => x"12",
          5379 => x"07",
          5380 => x"2b",
          5381 => x"0c",
          5382 => x"5b",
          5383 => x"1b",
          5384 => x"91",
          5385 => x"80",
          5386 => x"84",
          5387 => x"7b",
          5388 => x"08",
          5389 => x"c0",
          5390 => x"51",
          5391 => x"08",
          5392 => x"80",
          5393 => x"2e",
          5394 => x"ff",
          5395 => x"52",
          5396 => x"bb",
          5397 => x"08",
          5398 => x"58",
          5399 => x"94",
          5400 => x"55",
          5401 => x"7d",
          5402 => x"72",
          5403 => x"7e",
          5404 => x"77",
          5405 => x"38",
          5406 => x"81",
          5407 => x"84",
          5408 => x"ff",
          5409 => x"7e",
          5410 => x"57",
          5411 => x"7a",
          5412 => x"17",
          5413 => x"9e",
          5414 => x"71",
          5415 => x"07",
          5416 => x"34",
          5417 => x"90",
          5418 => x"34",
          5419 => x"7e",
          5420 => x"34",
          5421 => x"5d",
          5422 => x"d6",
          5423 => x"0c",
          5424 => x"06",
          5425 => x"7e",
          5426 => x"40",
          5427 => x"38",
          5428 => x"1b",
          5429 => x"f9",
          5430 => x"9c",
          5431 => x"7b",
          5432 => x"e9",
          5433 => x"f7",
          5434 => x"f7",
          5435 => x"53",
          5436 => x"52",
          5437 => x"84",
          5438 => x"ce",
          5439 => x"34",
          5440 => x"84",
          5441 => x"17",
          5442 => x"33",
          5443 => x"fd",
          5444 => x"a0",
          5445 => x"16",
          5446 => x"5c",
          5447 => x"57",
          5448 => x"5c",
          5449 => x"63",
          5450 => x"7e",
          5451 => x"38",
          5452 => x"38",
          5453 => x"38",
          5454 => x"5b",
          5455 => x"55",
          5456 => x"38",
          5457 => x"38",
          5458 => x"56",
          5459 => x"19",
          5460 => x"56",
          5461 => x"80",
          5462 => x"06",
          5463 => x"11",
          5464 => x"5d",
          5465 => x"38",
          5466 => x"83",
          5467 => x"38",
          5468 => x"19",
          5469 => x"05",
          5470 => x"38",
          5471 => x"1a",
          5472 => x"83",
          5473 => x"5c",
          5474 => x"7a",
          5475 => x"75",
          5476 => x"7c",
          5477 => x"81",
          5478 => x"38",
          5479 => x"56",
          5480 => x"89",
          5481 => x"18",
          5482 => x"19",
          5483 => x"79",
          5484 => x"bb",
          5485 => x"84",
          5486 => x"74",
          5487 => x"56",
          5488 => x"19",
          5489 => x"5d",
          5490 => x"54",
          5491 => x"51",
          5492 => x"08",
          5493 => x"ff",
          5494 => x"58",
          5495 => x"18",
          5496 => x"bb",
          5497 => x"1a",
          5498 => x"ff",
          5499 => x"79",
          5500 => x"7d",
          5501 => x"76",
          5502 => x"81",
          5503 => x"5a",
          5504 => x"fe",
          5505 => x"33",
          5506 => x"16",
          5507 => x"98",
          5508 => x"bc",
          5509 => x"a4",
          5510 => x"a7",
          5511 => x"55",
          5512 => x"56",
          5513 => x"77",
          5514 => x"38",
          5515 => x"1b",
          5516 => x"57",
          5517 => x"ff",
          5518 => x"38",
          5519 => x"70",
          5520 => x"74",
          5521 => x"91",
          5522 => x"0c",
          5523 => x"1a",
          5524 => x"90",
          5525 => x"64",
          5526 => x"7f",
          5527 => x"38",
          5528 => x"38",
          5529 => x"38",
          5530 => x"5a",
          5531 => x"55",
          5532 => x"38",
          5533 => x"38",
          5534 => x"06",
          5535 => x"82",
          5536 => x"5d",
          5537 => x"09",
          5538 => x"76",
          5539 => x"38",
          5540 => x"89",
          5541 => x"76",
          5542 => x"74",
          5543 => x"2e",
          5544 => x"d8",
          5545 => x"08",
          5546 => x"58",
          5547 => x"57",
          5548 => x"19",
          5549 => x"05",
          5550 => x"38",
          5551 => x"1a",
          5552 => x"83",
          5553 => x"5b",
          5554 => x"79",
          5555 => x"75",
          5556 => x"7d",
          5557 => x"80",
          5558 => x"38",
          5559 => x"7a",
          5560 => x"1a",
          5561 => x"55",
          5562 => x"70",
          5563 => x"74",
          5564 => x"06",
          5565 => x"2b",
          5566 => x"60",
          5567 => x"70",
          5568 => x"59",
          5569 => x"83",
          5570 => x"7a",
          5571 => x"77",
          5572 => x"34",
          5573 => x"91",
          5574 => x"0c",
          5575 => x"7c",
          5576 => x"76",
          5577 => x"54",
          5578 => x"33",
          5579 => x"84",
          5580 => x"57",
          5581 => x"06",
          5582 => x"78",
          5583 => x"16",
          5584 => x"80",
          5585 => x"58",
          5586 => x"ff",
          5587 => x"33",
          5588 => x"34",
          5589 => x"78",
          5590 => x"84",
          5591 => x"fd",
          5592 => x"39",
          5593 => x"3f",
          5594 => x"84",
          5595 => x"54",
          5596 => x"81",
          5597 => x"84",
          5598 => x"33",
          5599 => x"34",
          5600 => x"33",
          5601 => x"84",
          5602 => x"38",
          5603 => x"39",
          5604 => x"84",
          5605 => x"82",
          5606 => x"bb",
          5607 => x"3d",
          5608 => x"2e",
          5609 => x"2e",
          5610 => x"2e",
          5611 => x"22",
          5612 => x"38",
          5613 => x"81",
          5614 => x"2a",
          5615 => x"81",
          5616 => x"76",
          5617 => x"08",
          5618 => x"b8",
          5619 => x"5b",
          5620 => x"06",
          5621 => x"b8",
          5622 => x"95",
          5623 => x"2e",
          5624 => x"b4",
          5625 => x"38",
          5626 => x"07",
          5627 => x"08",
          5628 => x"06",
          5629 => x"7a",
          5630 => x"9c",
          5631 => x"5b",
          5632 => x"18",
          5633 => x"2a",
          5634 => x"2a",
          5635 => x"2a",
          5636 => x"34",
          5637 => x"98",
          5638 => x"34",
          5639 => x"93",
          5640 => x"1c",
          5641 => x"84",
          5642 => x"bf",
          5643 => x"75",
          5644 => x"3d",
          5645 => x"53",
          5646 => x"52",
          5647 => x"84",
          5648 => x"06",
          5649 => x"83",
          5650 => x"08",
          5651 => x"74",
          5652 => x"82",
          5653 => x"81",
          5654 => x"16",
          5655 => x"52",
          5656 => x"3f",
          5657 => x"2a",
          5658 => x"2a",
          5659 => x"08",
          5660 => x"5b",
          5661 => x"56",
          5662 => x"59",
          5663 => x"80",
          5664 => x"18",
          5665 => x"80",
          5666 => x"18",
          5667 => x"34",
          5668 => x"bb",
          5669 => x"06",
          5670 => x"a7",
          5671 => x"9f",
          5672 => x"55",
          5673 => x"56",
          5674 => x"18",
          5675 => x"11",
          5676 => x"81",
          5677 => x"38",
          5678 => x"78",
          5679 => x"58",
          5680 => x"81",
          5681 => x"f9",
          5682 => x"a6",
          5683 => x"bb",
          5684 => x"80",
          5685 => x"80",
          5686 => x"80",
          5687 => x"16",
          5688 => x"38",
          5689 => x"84",
          5690 => x"84",
          5691 => x"33",
          5692 => x"84",
          5693 => x"73",
          5694 => x"3d",
          5695 => x"75",
          5696 => x"05",
          5697 => x"71",
          5698 => x"71",
          5699 => x"33",
          5700 => x"84",
          5701 => x"84",
          5702 => x"84",
          5703 => x"78",
          5704 => x"53",
          5705 => x"82",
          5706 => x"59",
          5707 => x"80",
          5708 => x"08",
          5709 => x"58",
          5710 => x"ff",
          5711 => x"26",
          5712 => x"06",
          5713 => x"99",
          5714 => x"ff",
          5715 => x"2a",
          5716 => x"06",
          5717 => x"76",
          5718 => x"2a",
          5719 => x"2e",
          5720 => x"58",
          5721 => x"51",
          5722 => x"38",
          5723 => x"ea",
          5724 => x"05",
          5725 => x"84",
          5726 => x"08",
          5727 => x"84",
          5728 => x"68",
          5729 => x"d3",
          5730 => x"bb",
          5731 => x"d7",
          5732 => x"80",
          5733 => x"05",
          5734 => x"59",
          5735 => x"9b",
          5736 => x"2b",
          5737 => x"58",
          5738 => x"19",
          5739 => x"3d",
          5740 => x"2e",
          5741 => x"0b",
          5742 => x"04",
          5743 => x"98",
          5744 => x"98",
          5745 => x"7e",
          5746 => x"84",
          5747 => x"3d",
          5748 => x"3d",
          5749 => x"53",
          5750 => x"80",
          5751 => x"bb",
          5752 => x"83",
          5753 => x"7f",
          5754 => x"0c",
          5755 => x"79",
          5756 => x"3d",
          5757 => x"51",
          5758 => x"08",
          5759 => x"38",
          5760 => x"b4",
          5761 => x"bb",
          5762 => x"7d",
          5763 => x"b8",
          5764 => x"8d",
          5765 => x"2e",
          5766 => x"b4",
          5767 => x"df",
          5768 => x"33",
          5769 => x"5d",
          5770 => x"82",
          5771 => x"80",
          5772 => x"84",
          5773 => x"08",
          5774 => x"ff",
          5775 => x"59",
          5776 => x"df",
          5777 => x"33",
          5778 => x"42",
          5779 => x"81",
          5780 => x"84",
          5781 => x"a6",
          5782 => x"84",
          5783 => x"38",
          5784 => x"81",
          5785 => x"05",
          5786 => x"78",
          5787 => x"80",
          5788 => x"17",
          5789 => x"7c",
          5790 => x"26",
          5791 => x"38",
          5792 => x"80",
          5793 => x"19",
          5794 => x"34",
          5795 => x"3d",
          5796 => x"80",
          5797 => x"38",
          5798 => x"0b",
          5799 => x"83",
          5800 => x"43",
          5801 => x"8d",
          5802 => x"57",
          5803 => x"5b",
          5804 => x"76",
          5805 => x"7e",
          5806 => x"81",
          5807 => x"ba",
          5808 => x"ff",
          5809 => x"91",
          5810 => x"84",
          5811 => x"16",
          5812 => x"71",
          5813 => x"5e",
          5814 => x"17",
          5815 => x"07",
          5816 => x"5d",
          5817 => x"3f",
          5818 => x"84",
          5819 => x"b1",
          5820 => x"b8",
          5821 => x"5e",
          5822 => x"bb",
          5823 => x"84",
          5824 => x"a8",
          5825 => x"5a",
          5826 => x"83",
          5827 => x"2e",
          5828 => x"54",
          5829 => x"53",
          5830 => x"89",
          5831 => x"ff",
          5832 => x"58",
          5833 => x"e0",
          5834 => x"05",
          5835 => x"5e",
          5836 => x"fd",
          5837 => x"3d",
          5838 => x"33",
          5839 => x"60",
          5840 => x"08",
          5841 => x"7c",
          5842 => x"26",
          5843 => x"80",
          5844 => x"80",
          5845 => x"7d",
          5846 => x"2e",
          5847 => x"2e",
          5848 => x"2e",
          5849 => x"22",
          5850 => x"38",
          5851 => x"82",
          5852 => x"82",
          5853 => x"78",
          5854 => x"56",
          5855 => x"38",
          5856 => x"52",
          5857 => x"38",
          5858 => x"93",
          5859 => x"79",
          5860 => x"83",
          5861 => x"82",
          5862 => x"94",
          5863 => x"08",
          5864 => x"92",
          5865 => x"78",
          5866 => x"19",
          5867 => x"81",
          5868 => x"82",
          5869 => x"9b",
          5870 => x"84",
          5871 => x"75",
          5872 => x"27",
          5873 => x"16",
          5874 => x"18",
          5875 => x"08",
          5876 => x"0c",
          5877 => x"2e",
          5878 => x"08",
          5879 => x"27",
          5880 => x"71",
          5881 => x"2a",
          5882 => x"82",
          5883 => x"17",
          5884 => x"75",
          5885 => x"c0",
          5886 => x"83",
          5887 => x"ab",
          5888 => x"2e",
          5889 => x"98",
          5890 => x"80",
          5891 => x"77",
          5892 => x"ff",
          5893 => x"a5",
          5894 => x"55",
          5895 => x"53",
          5896 => x"58",
          5897 => x"08",
          5898 => x"91",
          5899 => x"84",
          5900 => x"33",
          5901 => x"75",
          5902 => x"57",
          5903 => x"81",
          5904 => x"0c",
          5905 => x"0c",
          5906 => x"80",
          5907 => x"80",
          5908 => x"79",
          5909 => x"84",
          5910 => x"76",
          5911 => x"84",
          5912 => x"33",
          5913 => x"84",
          5914 => x"38",
          5915 => x"39",
          5916 => x"3f",
          5917 => x"84",
          5918 => x"84",
          5919 => x"bb",
          5920 => x"18",
          5921 => x"18",
          5922 => x"8d",
          5923 => x"56",
          5924 => x"80",
          5925 => x"3d",
          5926 => x"bb",
          5927 => x"80",
          5928 => x"54",
          5929 => x"0d",
          5930 => x"51",
          5931 => x"08",
          5932 => x"38",
          5933 => x"59",
          5934 => x"33",
          5935 => x"79",
          5936 => x"08",
          5937 => x"88",
          5938 => x"5a",
          5939 => x"77",
          5940 => x"22",
          5941 => x"ff",
          5942 => x"55",
          5943 => x"2e",
          5944 => x"fe",
          5945 => x"f6",
          5946 => x"71",
          5947 => x"07",
          5948 => x"39",
          5949 => x"74",
          5950 => x"72",
          5951 => x"71",
          5952 => x"84",
          5953 => x"94",
          5954 => x"38",
          5955 => x"0c",
          5956 => x"51",
          5957 => x"08",
          5958 => x"75",
          5959 => x"0d",
          5960 => x"80",
          5961 => x"80",
          5962 => x"80",
          5963 => x"16",
          5964 => x"97",
          5965 => x"75",
          5966 => x"f3",
          5967 => x"ae",
          5968 => x"bb",
          5969 => x"bb",
          5970 => x"51",
          5971 => x"51",
          5972 => x"08",
          5973 => x"9f",
          5974 => x"57",
          5975 => x"3d",
          5976 => x"53",
          5977 => x"51",
          5978 => x"08",
          5979 => x"9f",
          5980 => x"57",
          5981 => x"ff",
          5982 => x"84",
          5983 => x"81",
          5984 => x"84",
          5985 => x"fe",
          5986 => x"fe",
          5987 => x"80",
          5988 => x"52",
          5989 => x"08",
          5990 => x"8a",
          5991 => x"3d",
          5992 => x"b6",
          5993 => x"84",
          5994 => x"cb",
          5995 => x"80",
          5996 => x"d1",
          5997 => x"ae",
          5998 => x"3d",
          5999 => x"0c",
          6000 => x"66",
          6001 => x"ec",
          6002 => x"3f",
          6003 => x"84",
          6004 => x"08",
          6005 => x"08",
          6006 => x"8d",
          6007 => x"84",
          6008 => x"84",
          6009 => x"2e",
          6010 => x"84",
          6011 => x"80",
          6012 => x"5d",
          6013 => x"ef",
          6014 => x"7c",
          6015 => x"b8",
          6016 => x"fd",
          6017 => x"2e",
          6018 => x"b4",
          6019 => x"80",
          6020 => x"2e",
          6021 => x"83",
          6022 => x"2b",
          6023 => x"70",
          6024 => x"80",
          6025 => x"30",
          6026 => x"05",
          6027 => x"41",
          6028 => x"5e",
          6029 => x"0c",
          6030 => x"81",
          6031 => x"84",
          6032 => x"81",
          6033 => x"70",
          6034 => x"fd",
          6035 => x"08",
          6036 => x"83",
          6037 => x"08",
          6038 => x"74",
          6039 => x"82",
          6040 => x"81",
          6041 => x"17",
          6042 => x"52",
          6043 => x"3f",
          6044 => x"42",
          6045 => x"51",
          6046 => x"08",
          6047 => x"84",
          6048 => x"bb",
          6049 => x"08",
          6050 => x"62",
          6051 => x"76",
          6052 => x"94",
          6053 => x"58",
          6054 => x"77",
          6055 => x"33",
          6056 => x"80",
          6057 => x"ff",
          6058 => x"55",
          6059 => x"77",
          6060 => x"5a",
          6061 => x"84",
          6062 => x"18",
          6063 => x"5a",
          6064 => x"89",
          6065 => x"08",
          6066 => x"33",
          6067 => x"16",
          6068 => x"79",
          6069 => x"5b",
          6070 => x"57",
          6071 => x"70",
          6072 => x"56",
          6073 => x"18",
          6074 => x"80",
          6075 => x"18",
          6076 => x"27",
          6077 => x"80",
          6078 => x"19",
          6079 => x"78",
          6080 => x"34",
          6081 => x"79",
          6082 => x"18",
          6083 => x"11",
          6084 => x"84",
          6085 => x"38",
          6086 => x"56",
          6087 => x"0d",
          6088 => x"ff",
          6089 => x"94",
          6090 => x"bb",
          6091 => x"84",
          6092 => x"38",
          6093 => x"f5",
          6094 => x"ff",
          6095 => x"82",
          6096 => x"94",
          6097 => x"27",
          6098 => x"0c",
          6099 => x"84",
          6100 => x"ff",
          6101 => x"51",
          6102 => x"08",
          6103 => x"74",
          6104 => x"80",
          6105 => x"57",
          6106 => x"39",
          6107 => x"fe",
          6108 => x"2e",
          6109 => x"81",
          6110 => x"38",
          6111 => x"1a",
          6112 => x"84",
          6113 => x"57",
          6114 => x"27",
          6115 => x"9c",
          6116 => x"80",
          6117 => x"76",
          6118 => x"84",
          6119 => x"e3",
          6120 => x"9c",
          6121 => x"bb",
          6122 => x"84",
          6123 => x"38",
          6124 => x"8f",
          6125 => x"ff",
          6126 => x"80",
          6127 => x"94",
          6128 => x"27",
          6129 => x"84",
          6130 => x"18",
          6131 => x"a1",
          6132 => x"33",
          6133 => x"bb",
          6134 => x"57",
          6135 => x"90",
          6136 => x"90",
          6137 => x"82",
          6138 => x"f6",
          6139 => x"33",
          6140 => x"90",
          6141 => x"84",
          6142 => x"81",
          6143 => x"82",
          6144 => x"a8",
          6145 => x"bb",
          6146 => x"80",
          6147 => x"0c",
          6148 => x"3d",
          6149 => x"ff",
          6150 => x"56",
          6151 => x"81",
          6152 => x"06",
          6153 => x"76",
          6154 => x"38",
          6155 => x"06",
          6156 => x"38",
          6157 => x"9a",
          6158 => x"33",
          6159 => x"2e",
          6160 => x"06",
          6161 => x"87",
          6162 => x"83",
          6163 => x"84",
          6164 => x"ff",
          6165 => x"56",
          6166 => x"84",
          6167 => x"91",
          6168 => x"84",
          6169 => x"84",
          6170 => x"95",
          6171 => x"2b",
          6172 => x"5d",
          6173 => x"08",
          6174 => x"08",
          6175 => x"3d",
          6176 => x"80",
          6177 => x"8b",
          6178 => x"84",
          6179 => x"75",
          6180 => x"5a",
          6181 => x"2e",
          6182 => x"81",
          6183 => x"7b",
          6184 => x"fd",
          6185 => x"3f",
          6186 => x"0c",
          6187 => x"98",
          6188 => x"08",
          6189 => x"33",
          6190 => x"81",
          6191 => x"53",
          6192 => x"fe",
          6193 => x"80",
          6194 => x"75",
          6195 => x"38",
          6196 => x"81",
          6197 => x"7c",
          6198 => x"51",
          6199 => x"08",
          6200 => x"ff",
          6201 => x"06",
          6202 => x"39",
          6203 => x"52",
          6204 => x"3f",
          6205 => x"2e",
          6206 => x"bb",
          6207 => x"08",
          6208 => x"08",
          6209 => x"fe",
          6210 => x"82",
          6211 => x"81",
          6212 => x"05",
          6213 => x"fe",
          6214 => x"39",
          6215 => x"38",
          6216 => x"3f",
          6217 => x"84",
          6218 => x"bb",
          6219 => x"84",
          6220 => x"38",
          6221 => x"fd",
          6222 => x"38",
          6223 => x"08",
          6224 => x"b0",
          6225 => x"17",
          6226 => x"34",
          6227 => x"38",
          6228 => x"fd",
          6229 => x"fd",
          6230 => x"e3",
          6231 => x"bc",
          6232 => x"f9",
          6233 => x"bb",
          6234 => x"84",
          6235 => x"7d",
          6236 => x"5a",
          6237 => x"08",
          6238 => x"88",
          6239 => x"0d",
          6240 => x"09",
          6241 => x"05",
          6242 => x"58",
          6243 => x"5f",
          6244 => x"ff",
          6245 => x"75",
          6246 => x"38",
          6247 => x"2e",
          6248 => x"ff",
          6249 => x"38",
          6250 => x"33",
          6251 => x"fe",
          6252 => x"56",
          6253 => x"8a",
          6254 => x"08",
          6255 => x"b8",
          6256 => x"80",
          6257 => x"15",
          6258 => x"17",
          6259 => x"38",
          6260 => x"81",
          6261 => x"84",
          6262 => x"18",
          6263 => x"39",
          6264 => x"17",
          6265 => x"fe",
          6266 => x"84",
          6267 => x"83",
          6268 => x"08",
          6269 => x"fe",
          6270 => x"82",
          6271 => x"75",
          6272 => x"05",
          6273 => x"fe",
          6274 => x"56",
          6275 => x"27",
          6276 => x"27",
          6277 => x"fe",
          6278 => x"5a",
          6279 => x"96",
          6280 => x"fd",
          6281 => x"2e",
          6282 => x"76",
          6283 => x"84",
          6284 => x"fe",
          6285 => x"77",
          6286 => x"18",
          6287 => x"7b",
          6288 => x"26",
          6289 => x"0c",
          6290 => x"55",
          6291 => x"56",
          6292 => x"f0",
          6293 => x"a0",
          6294 => x"16",
          6295 => x"0b",
          6296 => x"80",
          6297 => x"ce",
          6298 => x"a1",
          6299 => x"0b",
          6300 => x"ff",
          6301 => x"17",
          6302 => x"d3",
          6303 => x"2e",
          6304 => x"80",
          6305 => x"74",
          6306 => x"81",
          6307 => x"ef",
          6308 => x"17",
          6309 => x"06",
          6310 => x"34",
          6311 => x"17",
          6312 => x"80",
          6313 => x"1c",
          6314 => x"84",
          6315 => x"08",
          6316 => x"84",
          6317 => x"08",
          6318 => x"34",
          6319 => x"6a",
          6320 => x"88",
          6321 => x"33",
          6322 => x"69",
          6323 => x"57",
          6324 => x"fe",
          6325 => x"56",
          6326 => x"0d",
          6327 => x"ec",
          6328 => x"80",
          6329 => x"90",
          6330 => x"7a",
          6331 => x"34",
          6332 => x"b8",
          6333 => x"7b",
          6334 => x"77",
          6335 => x"69",
          6336 => x"57",
          6337 => x"fe",
          6338 => x"56",
          6339 => x"3d",
          6340 => x"79",
          6341 => x"05",
          6342 => x"75",
          6343 => x"38",
          6344 => x"53",
          6345 => x"3d",
          6346 => x"84",
          6347 => x"2e",
          6348 => x"b1",
          6349 => x"b2",
          6350 => x"59",
          6351 => x"08",
          6352 => x"02",
          6353 => x"5d",
          6354 => x"92",
          6355 => x"75",
          6356 => x"81",
          6357 => x"ef",
          6358 => x"58",
          6359 => x"33",
          6360 => x"15",
          6361 => x"52",
          6362 => x"bb",
          6363 => x"85",
          6364 => x"81",
          6365 => x"0c",
          6366 => x"11",
          6367 => x"74",
          6368 => x"81",
          6369 => x"7a",
          6370 => x"83",
          6371 => x"5f",
          6372 => x"33",
          6373 => x"9f",
          6374 => x"89",
          6375 => x"57",
          6376 => x"26",
          6377 => x"06",
          6378 => x"59",
          6379 => x"85",
          6380 => x"32",
          6381 => x"7a",
          6382 => x"95",
          6383 => x"7b",
          6384 => x"7e",
          6385 => x"24",
          6386 => x"53",
          6387 => x"3d",
          6388 => x"84",
          6389 => x"b2",
          6390 => x"08",
          6391 => x"77",
          6392 => x"84",
          6393 => x"92",
          6394 => x"02",
          6395 => x"5a",
          6396 => x"70",
          6397 => x"79",
          6398 => x"8b",
          6399 => x"2a",
          6400 => x"75",
          6401 => x"7f",
          6402 => x"18",
          6403 => x"5c",
          6404 => x"3d",
          6405 => x"9b",
          6406 => x"2b",
          6407 => x"7d",
          6408 => x"9c",
          6409 => x"7d",
          6410 => x"76",
          6411 => x"5e",
          6412 => x"7a",
          6413 => x"aa",
          6414 => x"bc",
          6415 => x"52",
          6416 => x"3f",
          6417 => x"38",
          6418 => x"0c",
          6419 => x"56",
          6420 => x"5a",
          6421 => x"38",
          6422 => x"56",
          6423 => x"2a",
          6424 => x"33",
          6425 => x"93",
          6426 => x"ec",
          6427 => x"80",
          6428 => x"83",
          6429 => x"b2",
          6430 => x"2e",
          6431 => x"fb",
          6432 => x"84",
          6433 => x"16",
          6434 => x"b4",
          6435 => x"16",
          6436 => x"09",
          6437 => x"76",
          6438 => x"51",
          6439 => x"08",
          6440 => x"58",
          6441 => x"aa",
          6442 => x"34",
          6443 => x"08",
          6444 => x"51",
          6445 => x"08",
          6446 => x"ff",
          6447 => x"f9",
          6448 => x"38",
          6449 => x"bb",
          6450 => x"3d",
          6451 => x"0c",
          6452 => x"94",
          6453 => x"2b",
          6454 => x"8d",
          6455 => x"fb",
          6456 => x"2e",
          6457 => x"0c",
          6458 => x"16",
          6459 => x"51",
          6460 => x"bb",
          6461 => x"fe",
          6462 => x"17",
          6463 => x"31",
          6464 => x"a0",
          6465 => x"16",
          6466 => x"06",
          6467 => x"08",
          6468 => x"81",
          6469 => x"79",
          6470 => x"17",
          6471 => x"18",
          6472 => x"81",
          6473 => x"38",
          6474 => x"b4",
          6475 => x"bb",
          6476 => x"08",
          6477 => x"5d",
          6478 => x"81",
          6479 => x"18",
          6480 => x"33",
          6481 => x"fb",
          6482 => x"df",
          6483 => x"05",
          6484 => x"cc",
          6485 => x"91",
          6486 => x"bb",
          6487 => x"84",
          6488 => x"78",
          6489 => x"51",
          6490 => x"08",
          6491 => x"02",
          6492 => x"54",
          6493 => x"06",
          6494 => x"06",
          6495 => x"55",
          6496 => x"0b",
          6497 => x"d3",
          6498 => x"84",
          6499 => x"0d",
          6500 => x"05",
          6501 => x"3f",
          6502 => x"84",
          6503 => x"bb",
          6504 => x"5a",
          6505 => x"ff",
          6506 => x"55",
          6507 => x"80",
          6508 => x"86",
          6509 => x"22",
          6510 => x"59",
          6511 => x"88",
          6512 => x"90",
          6513 => x"98",
          6514 => x"57",
          6515 => x"fe",
          6516 => x"84",
          6517 => x"e8",
          6518 => x"53",
          6519 => x"51",
          6520 => x"08",
          6521 => x"bb",
          6522 => x"57",
          6523 => x"76",
          6524 => x"76",
          6525 => x"5b",
          6526 => x"70",
          6527 => x"81",
          6528 => x"56",
          6529 => x"82",
          6530 => x"55",
          6531 => x"98",
          6532 => x"52",
          6533 => x"3f",
          6534 => x"38",
          6535 => x"0c",
          6536 => x"33",
          6537 => x"2e",
          6538 => x"2e",
          6539 => x"05",
          6540 => x"90",
          6541 => x"33",
          6542 => x"71",
          6543 => x"59",
          6544 => x"3d",
          6545 => x"52",
          6546 => x"c4",
          6547 => x"bb",
          6548 => x"76",
          6549 => x"38",
          6550 => x"39",
          6551 => x"16",
          6552 => x"fe",
          6553 => x"84",
          6554 => x"e8",
          6555 => x"34",
          6556 => x"84",
          6557 => x"17",
          6558 => x"33",
          6559 => x"fe",
          6560 => x"a0",
          6561 => x"16",
          6562 => x"59",
          6563 => x"81",
          6564 => x"84",
          6565 => x"38",
          6566 => x"fe",
          6567 => x"57",
          6568 => x"84",
          6569 => x"66",
          6570 => x"7c",
          6571 => x"34",
          6572 => x"38",
          6573 => x"34",
          6574 => x"18",
          6575 => x"79",
          6576 => x"79",
          6577 => x"82",
          6578 => x"a2",
          6579 => x"bb",
          6580 => x"82",
          6581 => x"57",
          6582 => x"34",
          6583 => x"a3",
          6584 => x"06",
          6585 => x"81",
          6586 => x"5c",
          6587 => x"55",
          6588 => x"74",
          6589 => x"74",
          6590 => x"84",
          6591 => x"84",
          6592 => x"57",
          6593 => x"e8",
          6594 => x"81",
          6595 => x"2e",
          6596 => x"2e",
          6597 => x"81",
          6598 => x"2e",
          6599 => x"06",
          6600 => x"78",
          6601 => x"81",
          6602 => x"38",
          6603 => x"88",
          6604 => x"5d",
          6605 => x"81",
          6606 => x"08",
          6607 => x"58",
          6608 => x"38",
          6609 => x"81",
          6610 => x"99",
          6611 => x"70",
          6612 => x"81",
          6613 => x"ed",
          6614 => x"95",
          6615 => x"3f",
          6616 => x"84",
          6617 => x"75",
          6618 => x"04",
          6619 => x"3f",
          6620 => x"06",
          6621 => x"75",
          6622 => x"04",
          6623 => x"39",
          6624 => x"3f",
          6625 => x"84",
          6626 => x"82",
          6627 => x"55",
          6628 => x"70",
          6629 => x"74",
          6630 => x"1e",
          6631 => x"84",
          6632 => x"87",
          6633 => x"86",
          6634 => x"08",
          6635 => x"38",
          6636 => x"38",
          6637 => x"fe",
          6638 => x"57",
          6639 => x"81",
          6640 => x"08",
          6641 => x"57",
          6642 => x"b2",
          6643 => x"2e",
          6644 => x"54",
          6645 => x"33",
          6646 => x"84",
          6647 => x"81",
          6648 => x"78",
          6649 => x"33",
          6650 => x"81",
          6651 => x"78",
          6652 => x"d7",
          6653 => x"a5",
          6654 => x"da",
          6655 => x"bb",
          6656 => x"87",
          6657 => x"76",
          6658 => x"57",
          6659 => x"34",
          6660 => x"56",
          6661 => x"7e",
          6662 => x"58",
          6663 => x"ff",
          6664 => x"38",
          6665 => x"70",
          6666 => x"74",
          6667 => x"e5",
          6668 => x"1e",
          6669 => x"84",
          6670 => x"81",
          6671 => x"18",
          6672 => x"51",
          6673 => x"08",
          6674 => x"38",
          6675 => x"b4",
          6676 => x"7b",
          6677 => x"18",
          6678 => x"84",
          6679 => x"74",
          6680 => x"8a",
          6681 => x"bb",
          6682 => x"fe",
          6683 => x"80",
          6684 => x"81",
          6685 => x"05",
          6686 => x"fe",
          6687 => x"3d",
          6688 => x"cb",
          6689 => x"76",
          6690 => x"74",
          6691 => x"73",
          6692 => x"84",
          6693 => x"81",
          6694 => x"81",
          6695 => x"81",
          6696 => x"38",
          6697 => x"17",
          6698 => x"5d",
          6699 => x"8a",
          6700 => x"7c",
          6701 => x"3f",
          6702 => x"72",
          6703 => x"05",
          6704 => x"55",
          6705 => x"19",
          6706 => x"77",
          6707 => x"76",
          6708 => x"7f",
          6709 => x"83",
          6710 => x"81",
          6711 => x"08",
          6712 => x"84",
          6713 => x"78",
          6714 => x"09",
          6715 => x"54",
          6716 => x"0d",
          6717 => x"90",
          6718 => x"fe",
          6719 => x"81",
          6720 => x"77",
          6721 => x"80",
          6722 => x"58",
          6723 => x"54",
          6724 => x"53",
          6725 => x"3f",
          6726 => x"84",
          6727 => x"ff",
          6728 => x"7e",
          6729 => x"2e",
          6730 => x"79",
          6731 => x"c0",
          6732 => x"15",
          6733 => x"5a",
          6734 => x"7d",
          6735 => x"81",
          6736 => x"54",
          6737 => x"39",
          6738 => x"82",
          6739 => x"c0",
          6740 => x"84",
          6741 => x"3d",
          6742 => x"81",
          6743 => x"0b",
          6744 => x"79",
          6745 => x"81",
          6746 => x"56",
          6747 => x"ed",
          6748 => x"84",
          6749 => x"84",
          6750 => x"cc",
          6751 => x"2e",
          6752 => x"84",
          6753 => x"12",
          6754 => x"51",
          6755 => x"08",
          6756 => x"56",
          6757 => x"82",
          6758 => x"84",
          6759 => x"83",
          6760 => x"84",
          6761 => x"55",
          6762 => x"82",
          6763 => x"15",
          6764 => x"7e",
          6765 => x"26",
          6766 => x"26",
          6767 => x"55",
          6768 => x"a6",
          6769 => x"77",
          6770 => x"85",
          6771 => x"77",
          6772 => x"b0",
          6773 => x"81",
          6774 => x"fe",
          6775 => x"84",
          6776 => x"05",
          6777 => x"88",
          6778 => x"82",
          6779 => x"f8",
          6780 => x"b2",
          6781 => x"82",
          6782 => x"33",
          6783 => x"88",
          6784 => x"07",
          6785 => x"ba",
          6786 => x"71",
          6787 => x"14",
          6788 => x"33",
          6789 => x"a3",
          6790 => x"54",
          6791 => x"4d",
          6792 => x"90",
          6793 => x"82",
          6794 => x"06",
          6795 => x"38",
          6796 => x"89",
          6797 => x"f4",
          6798 => x"43",
          6799 => x"38",
          6800 => x"81",
          6801 => x"74",
          6802 => x"98",
          6803 => x"82",
          6804 => x"80",
          6805 => x"38",
          6806 => x"3f",
          6807 => x"55",
          6808 => x"96",
          6809 => x"10",
          6810 => x"72",
          6811 => x"ff",
          6812 => x"47",
          6813 => x"11",
          6814 => x"58",
          6815 => x"b8",
          6816 => x"16",
          6817 => x"26",
          6818 => x"31",
          6819 => x"fc",
          6820 => x"40",
          6821 => x"82",
          6822 => x"83",
          6823 => x"27",
          6824 => x"77",
          6825 => x"ef",
          6826 => x"57",
          6827 => x"0d",
          6828 => x"fb",
          6829 => x"0c",
          6830 => x"04",
          6831 => x"06",
          6832 => x"38",
          6833 => x"05",
          6834 => x"38",
          6835 => x"7d",
          6836 => x"05",
          6837 => x"33",
          6838 => x"99",
          6839 => x"ff",
          6840 => x"64",
          6841 => x"81",
          6842 => x"9f",
          6843 => x"81",
          6844 => x"75",
          6845 => x"9f",
          6846 => x"80",
          6847 => x"1f",
          6848 => x"38",
          6849 => x"f8",
          6850 => x"cb",
          6851 => x"08",
          6852 => x"06",
          6853 => x"83",
          6854 => x"7e",
          6855 => x"31",
          6856 => x"d2",
          6857 => x"7b",
          6858 => x"39",
          6859 => x"80",
          6860 => x"30",
          6861 => x"bb",
          6862 => x"7a",
          6863 => x"7b",
          6864 => x"84",
          6865 => x"bb",
          6866 => x"2e",
          6867 => x"8b",
          6868 => x"7a",
          6869 => x"55",
          6870 => x"ff",
          6871 => x"83",
          6872 => x"81",
          6873 => x"58",
          6874 => x"60",
          6875 => x"61",
          6876 => x"34",
          6877 => x"61",
          6878 => x"7b",
          6879 => x"05",
          6880 => x"48",
          6881 => x"2a",
          6882 => x"34",
          6883 => x"86",
          6884 => x"55",
          6885 => x"2a",
          6886 => x"61",
          6887 => x"34",
          6888 => x"9a",
          6889 => x"7e",
          6890 => x"48",
          6891 => x"2a",
          6892 => x"98",
          6893 => x"90",
          6894 => x"2e",
          6895 => x"34",
          6896 => x"a9",
          6897 => x"34",
          6898 => x"61",
          6899 => x"6a",
          6900 => x"a4",
          6901 => x"93",
          6902 => x"57",
          6903 => x"76",
          6904 => x"55",
          6905 => x"49",
          6906 => x"05",
          6907 => x"7e",
          6908 => x"c8",
          6909 => x"fa",
          6910 => x"2e",
          6911 => x"80",
          6912 => x"15",
          6913 => x"5b",
          6914 => x"ff",
          6915 => x"38",
          6916 => x"2a",
          6917 => x"05",
          6918 => x"64",
          6919 => x"2a",
          6920 => x"59",
          6921 => x"78",
          6922 => x"fe",
          6923 => x"85",
          6924 => x"80",
          6925 => x"15",
          6926 => x"7a",
          6927 => x"81",
          6928 => x"38",
          6929 => x"66",
          6930 => x"38",
          6931 => x"52",
          6932 => x"bb",
          6933 => x"76",
          6934 => x"8c",
          6935 => x"58",
          6936 => x"84",
          6937 => x"58",
          6938 => x"81",
          6939 => x"80",
          6940 => x"05",
          6941 => x"38",
          6942 => x"34",
          6943 => x"34",
          6944 => x"82",
          6945 => x"77",
          6946 => x"fd",
          6947 => x"8b",
          6948 => x"bb",
          6949 => x"76",
          6950 => x"08",
          6951 => x"c6",
          6952 => x"34",
          6953 => x"bb",
          6954 => x"62",
          6955 => x"2a",
          6956 => x"62",
          6957 => x"05",
          6958 => x"83",
          6959 => x"60",
          6960 => x"81",
          6961 => x"38",
          6962 => x"c4",
          6963 => x"08",
          6964 => x"84",
          6965 => x"bb",
          6966 => x"39",
          6967 => x"c4",
          6968 => x"57",
          6969 => x"58",
          6970 => x"26",
          6971 => x"10",
          6972 => x"74",
          6973 => x"ee",
          6974 => x"b3",
          6975 => x"84",
          6976 => x"a0",
          6977 => x"fc",
          6978 => x"f0",
          6979 => x"57",
          6980 => x"83",
          6981 => x"f8",
          6982 => x"f4",
          6983 => x"68",
          6984 => x"af",
          6985 => x"61",
          6986 => x"68",
          6987 => x"5b",
          6988 => x"2a",
          6989 => x"c6",
          6990 => x"80",
          6991 => x"80",
          6992 => x"c6",
          6993 => x"7c",
          6994 => x"34",
          6995 => x"05",
          6996 => x"a7",
          6997 => x"80",
          6998 => x"05",
          6999 => x"61",
          7000 => x"34",
          7001 => x"b3",
          7002 => x"05",
          7003 => x"93",
          7004 => x"59",
          7005 => x"33",
          7006 => x"15",
          7007 => x"76",
          7008 => x"81",
          7009 => x"da",
          7010 => x"53",
          7011 => x"3f",
          7012 => x"b0",
          7013 => x"77",
          7014 => x"84",
          7015 => x"51",
          7016 => x"81",
          7017 => x"0d",
          7018 => x"34",
          7019 => x"4c",
          7020 => x"34",
          7021 => x"34",
          7022 => x"86",
          7023 => x"ff",
          7024 => x"05",
          7025 => x"65",
          7026 => x"54",
          7027 => x"fe",
          7028 => x"57",
          7029 => x"ff",
          7030 => x"80",
          7031 => x"7b",
          7032 => x"57",
          7033 => x"57",
          7034 => x"61",
          7035 => x"83",
          7036 => x"e6",
          7037 => x"05",
          7038 => x"83",
          7039 => x"78",
          7040 => x"2a",
          7041 => x"7a",
          7042 => x"05",
          7043 => x"76",
          7044 => x"83",
          7045 => x"05",
          7046 => x"6b",
          7047 => x"52",
          7048 => x"54",
          7049 => x"fe",
          7050 => x"f7",
          7051 => x"5b",
          7052 => x"57",
          7053 => x"3d",
          7054 => x"53",
          7055 => x"3f",
          7056 => x"38",
          7057 => x"90",
          7058 => x"34",
          7059 => x"38",
          7060 => x"34",
          7061 => x"74",
          7062 => x"04",
          7063 => x"b3",
          7064 => x"80",
          7065 => x"76",
          7066 => x"17",
          7067 => x"81",
          7068 => x"74",
          7069 => x"0c",
          7070 => x"05",
          7071 => x"08",
          7072 => x"32",
          7073 => x"70",
          7074 => x"1b",
          7075 => x"52",
          7076 => x"39",
          7077 => x"33",
          7078 => x"57",
          7079 => x"34",
          7080 => x"3d",
          7081 => x"f7",
          7082 => x"c0",
          7083 => x"59",
          7084 => x"bb",
          7085 => x"81",
          7086 => x"75",
          7087 => x"11",
          7088 => x"08",
          7089 => x"84",
          7090 => x"38",
          7091 => x"3d",
          7092 => x"55",
          7093 => x"51",
          7094 => x"70",
          7095 => x"30",
          7096 => x"8d",
          7097 => x"81",
          7098 => x"3d",
          7099 => x"84",
          7100 => x"52",
          7101 => x"83",
          7102 => x"84",
          7103 => x"ff",
          7104 => x"09",
          7105 => x"e4",
          7106 => x"71",
          7107 => x"ff",
          7108 => x"26",
          7109 => x"05",
          7110 => x"80",
          7111 => x"84",
          7112 => x"3d",
          7113 => x"05",
          7114 => x"70",
          7115 => x"72",
          7116 => x"04",
          7117 => x"ef",
          7118 => x"70",
          7119 => x"84",
          7120 => x"04",
          7121 => x"ff",
          7122 => x"ff",
          7123 => x"75",
          7124 => x"70",
          7125 => x"70",
          7126 => x"56",
          7127 => x"82",
          7128 => x"54",
          7129 => x"54",
          7130 => x"38",
          7131 => x"52",
          7132 => x"75",
          7133 => x"80",
          7134 => x"bb",
          7135 => x"ee",
          7136 => x"26",
          7137 => x"f0",
          7138 => x"16",
          7139 => x"75",
          7140 => x"83",
          7141 => x"88",
          7142 => x"51",
          7143 => x"ff",
          7144 => x"70",
          7145 => x"39",
          7146 => x"57",
          7147 => x"ff",
          7148 => x"75",
          7149 => x"70",
          7150 => x"ff",
          7151 => x"05",
          7152 => x"00",
          7153 => x"00",
          7154 => x"ff",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"00",
          7372 => x"00",
          7373 => x"00",
          7374 => x"00",
          7375 => x"00",
          7376 => x"00",
          7377 => x"00",
          7378 => x"00",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"00",
          7383 => x"00",
          7384 => x"00",
          7385 => x"00",
          7386 => x"00",
          7387 => x"00",
          7388 => x"00",
          7389 => x"00",
          7390 => x"00",
          7391 => x"69",
          7392 => x"69",
          7393 => x"69",
          7394 => x"6c",
          7395 => x"65",
          7396 => x"63",
          7397 => x"63",
          7398 => x"64",
          7399 => x"64",
          7400 => x"65",
          7401 => x"65",
          7402 => x"69",
          7403 => x"66",
          7404 => x"00",
          7405 => x"65",
          7406 => x"65",
          7407 => x"6e",
          7408 => x"65",
          7409 => x"6c",
          7410 => x"62",
          7411 => x"62",
          7412 => x"69",
          7413 => x"64",
          7414 => x"77",
          7415 => x"2e",
          7416 => x"65",
          7417 => x"63",
          7418 => x"00",
          7419 => x"61",
          7420 => x"20",
          7421 => x"00",
          7422 => x"66",
          7423 => x"6d",
          7424 => x"00",
          7425 => x"69",
          7426 => x"64",
          7427 => x"75",
          7428 => x"61",
          7429 => x"6e",
          7430 => x"00",
          7431 => x"74",
          7432 => x"64",
          7433 => x"6d",
          7434 => x"20",
          7435 => x"74",
          7436 => x"64",
          7437 => x"6b",
          7438 => x"6e",
          7439 => x"6c",
          7440 => x"72",
          7441 => x"62",
          7442 => x"6e",
          7443 => x"00",
          7444 => x"20",
          7445 => x"72",
          7446 => x"2e",
          7447 => x"68",
          7448 => x"6e",
          7449 => x"00",
          7450 => x"61",
          7451 => x"65",
          7452 => x"00",
          7453 => x"73",
          7454 => x"2e",
          7455 => x"69",
          7456 => x"61",
          7457 => x"6f",
          7458 => x"6f",
          7459 => x"6f",
          7460 => x"6f",
          7461 => x"69",
          7462 => x"72",
          7463 => x"6e",
          7464 => x"65",
          7465 => x"69",
          7466 => x"72",
          7467 => x"73",
          7468 => x"25",
          7469 => x"73",
          7470 => x"25",
          7471 => x"73",
          7472 => x"00",
          7473 => x"00",
          7474 => x"00",
          7475 => x"30",
          7476 => x"7c",
          7477 => x"20",
          7478 => x"00",
          7479 => x"20",
          7480 => x"4f",
          7481 => x"20",
          7482 => x"2f",
          7483 => x"31",
          7484 => x"5a",
          7485 => x"20",
          7486 => x"73",
          7487 => x"0a",
          7488 => x"20",
          7489 => x"41",
          7490 => x"20",
          7491 => x"20",
          7492 => x"38",
          7493 => x"20",
          7494 => x"64",
          7495 => x"20",
          7496 => x"20",
          7497 => x"38",
          7498 => x"50",
          7499 => x"72",
          7500 => x"64",
          7501 => x"41",
          7502 => x"69",
          7503 => x"74",
          7504 => x"20",
          7505 => x"72",
          7506 => x"41",
          7507 => x"69",
          7508 => x"74",
          7509 => x"20",
          7510 => x"72",
          7511 => x"4f",
          7512 => x"69",
          7513 => x"74",
          7514 => x"20",
          7515 => x"72",
          7516 => x"53",
          7517 => x"72",
          7518 => x"69",
          7519 => x"65",
          7520 => x"65",
          7521 => x"70",
          7522 => x"2e",
          7523 => x"69",
          7524 => x"72",
          7525 => x"75",
          7526 => x"62",
          7527 => x"4f",
          7528 => x"73",
          7529 => x"64",
          7530 => x"74",
          7531 => x"73",
          7532 => x"30",
          7533 => x"65",
          7534 => x"61",
          7535 => x"00",
          7536 => x"64",
          7537 => x"3a",
          7538 => x"6f",
          7539 => x"00",
          7540 => x"69",
          7541 => x"73",
          7542 => x"00",
          7543 => x"72",
          7544 => x"67",
          7545 => x"65",
          7546 => x"67",
          7547 => x"61",
          7548 => x"00",
          7549 => x"6e",
          7550 => x"40",
          7551 => x"2e",
          7552 => x"61",
          7553 => x"72",
          7554 => x"65",
          7555 => x"00",
          7556 => x"74",
          7557 => x"65",
          7558 => x"78",
          7559 => x"30",
          7560 => x"6c",
          7561 => x"30",
          7562 => x"58",
          7563 => x"72",
          7564 => x"00",
          7565 => x"28",
          7566 => x"25",
          7567 => x"38",
          7568 => x"6f",
          7569 => x"2e",
          7570 => x"20",
          7571 => x"6c",
          7572 => x"2e",
          7573 => x"75",
          7574 => x"72",
          7575 => x"6c",
          7576 => x"64",
          7577 => x"00",
          7578 => x"79",
          7579 => x"74",
          7580 => x"6e",
          7581 => x"65",
          7582 => x"61",
          7583 => x"3f",
          7584 => x"2f",
          7585 => x"64",
          7586 => x"64",
          7587 => x"6f",
          7588 => x"74",
          7589 => x"0a",
          7590 => x"20",
          7591 => x"6e",
          7592 => x"64",
          7593 => x"3a",
          7594 => x"50",
          7595 => x"20",
          7596 => x"41",
          7597 => x"3d",
          7598 => x"00",
          7599 => x"50",
          7600 => x"79",
          7601 => x"41",
          7602 => x"3d",
          7603 => x"00",
          7604 => x"74",
          7605 => x"72",
          7606 => x"73",
          7607 => x"3d",
          7608 => x"00",
          7609 => x"00",
          7610 => x"50",
          7611 => x"20",
          7612 => x"20",
          7613 => x"3d",
          7614 => x"00",
          7615 => x"79",
          7616 => x"6f",
          7617 => x"20",
          7618 => x"3d",
          7619 => x"64",
          7620 => x"20",
          7621 => x"6f",
          7622 => x"4d",
          7623 => x"46",
          7624 => x"2e",
          7625 => x"0a",
          7626 => x"44",
          7627 => x"63",
          7628 => x"20",
          7629 => x"3d",
          7630 => x"64",
          7631 => x"20",
          7632 => x"20",
          7633 => x"20",
          7634 => x"00",
          7635 => x"42",
          7636 => x"20",
          7637 => x"4f",
          7638 => x"00",
          7639 => x"4e",
          7640 => x"20",
          7641 => x"6c",
          7642 => x"2e",
          7643 => x"49",
          7644 => x"20",
          7645 => x"20",
          7646 => x"2e",
          7647 => x"44",
          7648 => x"20",
          7649 => x"73",
          7650 => x"2e",
          7651 => x"41",
          7652 => x"20",
          7653 => x"30",
          7654 => x"20",
          7655 => x"20",
          7656 => x"38",
          7657 => x"2e",
          7658 => x"4e",
          7659 => x"20",
          7660 => x"30",
          7661 => x"20",
          7662 => x"20",
          7663 => x"38",
          7664 => x"2e",
          7665 => x"42",
          7666 => x"20",
          7667 => x"30",
          7668 => x"28",
          7669 => x"43",
          7670 => x"29",
          7671 => x"77",
          7672 => x"00",
          7673 => x"00",
          7674 => x"6d",
          7675 => x"00",
          7676 => x"00",
          7677 => x"00",
          7678 => x"00",
          7679 => x"00",
          7680 => x"00",
          7681 => x"00",
          7682 => x"00",
          7683 => x"00",
          7684 => x"00",
          7685 => x"00",
          7686 => x"00",
          7687 => x"00",
          7688 => x"00",
          7689 => x"00",
          7690 => x"00",
          7691 => x"00",
          7692 => x"00",
          7693 => x"00",
          7694 => x"00",
          7695 => x"00",
          7696 => x"00",
          7697 => x"00",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"00",
          7703 => x"00",
          7704 => x"00",
          7705 => x"00",
          7706 => x"00",
          7707 => x"00",
          7708 => x"00",
          7709 => x"5b",
          7710 => x"5b",
          7711 => x"5b",
          7712 => x"5b",
          7713 => x"5b",
          7714 => x"5b",
          7715 => x"00",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"69",
          7721 => x"65",
          7722 => x"78",
          7723 => x"74",
          7724 => x"72",
          7725 => x"73",
          7726 => x"6c",
          7727 => x"62",
          7728 => x"69",
          7729 => x"69",
          7730 => x"00",
          7731 => x"72",
          7732 => x"72",
          7733 => x"00",
          7734 => x"20",
          7735 => x"61",
          7736 => x"20",
          7737 => x"68",
          7738 => x"72",
          7739 => x"74",
          7740 => x"00",
          7741 => x"00",
          7742 => x"00",
          7743 => x"5b",
          7744 => x"5b",
          7745 => x"00",
          7746 => x"00",
          7747 => x"00",
          7748 => x"00",
          7749 => x"00",
          7750 => x"00",
          7751 => x"00",
          7752 => x"00",
          7753 => x"00",
          7754 => x"00",
          7755 => x"00",
          7756 => x"00",
          7757 => x"5b",
          7758 => x"5b",
          7759 => x"3a",
          7760 => x"64",
          7761 => x"25",
          7762 => x"00",
          7763 => x"25",
          7764 => x"3a",
          7765 => x"64",
          7766 => x"3a",
          7767 => x"30",
          7768 => x"63",
          7769 => x"00",
          7770 => x"74",
          7771 => x"3a",
          7772 => x"32",
          7773 => x"00",
          7774 => x"32",
          7775 => x"00",
          7776 => x"32",
          7777 => x"6f",
          7778 => x"65",
          7779 => x"00",
          7780 => x"2a",
          7781 => x"00",
          7782 => x"5d",
          7783 => x"41",
          7784 => x"fe",
          7785 => x"2e",
          7786 => x"4d",
          7787 => x"54",
          7788 => x"4f",
          7789 => x"20",
          7790 => x"20",
          7791 => x"00",
          7792 => x"00",
          7793 => x"0e",
          7794 => x"00",
          7795 => x"41",
          7796 => x"49",
          7797 => x"4f",
          7798 => x"9d",
          7799 => x"a5",
          7800 => x"ad",
          7801 => x"b5",
          7802 => x"bd",
          7803 => x"c5",
          7804 => x"cd",
          7805 => x"d5",
          7806 => x"dd",
          7807 => x"e5",
          7808 => x"ed",
          7809 => x"f5",
          7810 => x"fd",
          7811 => x"5b",
          7812 => x"3e",
          7813 => x"01",
          7814 => x"00",
          7815 => x"01",
          7816 => x"10",
          7817 => x"c7",
          7818 => x"e4",
          7819 => x"ea",
          7820 => x"ee",
          7821 => x"c9",
          7822 => x"f6",
          7823 => x"ff",
          7824 => x"a3",
          7825 => x"e1",
          7826 => x"f1",
          7827 => x"bf",
          7828 => x"bc",
          7829 => x"91",
          7830 => x"24",
          7831 => x"55",
          7832 => x"5d",
          7833 => x"14",
          7834 => x"00",
          7835 => x"5a",
          7836 => x"60",
          7837 => x"68",
          7838 => x"58",
          7839 => x"6a",
          7840 => x"84",
          7841 => x"b1",
          7842 => x"a3",
          7843 => x"a6",
          7844 => x"1e",
          7845 => x"61",
          7846 => x"20",
          7847 => x"b0",
          7848 => x"7f",
          7849 => x"61",
          7850 => x"f8",
          7851 => x"78",
          7852 => x"06",
          7853 => x"2e",
          7854 => x"4d",
          7855 => x"82",
          7856 => x"87",
          7857 => x"8b",
          7858 => x"8f",
          7859 => x"93",
          7860 => x"97",
          7861 => x"9b",
          7862 => x"9f",
          7863 => x"a2",
          7864 => x"a7",
          7865 => x"ab",
          7866 => x"af",
          7867 => x"b3",
          7868 => x"b7",
          7869 => x"bb",
          7870 => x"f7",
          7871 => x"c3",
          7872 => x"c7",
          7873 => x"cb",
          7874 => x"dd",
          7875 => x"12",
          7876 => x"f4",
          7877 => x"22",
          7878 => x"65",
          7879 => x"66",
          7880 => x"41",
          7881 => x"40",
          7882 => x"89",
          7883 => x"5a",
          7884 => x"5e",
          7885 => x"62",
          7886 => x"66",
          7887 => x"6a",
          7888 => x"6e",
          7889 => x"9d",
          7890 => x"76",
          7891 => x"7a",
          7892 => x"7e",
          7893 => x"82",
          7894 => x"86",
          7895 => x"b1",
          7896 => x"8e",
          7897 => x"b7",
          7898 => x"fe",
          7899 => x"86",
          7900 => x"b1",
          7901 => x"a3",
          7902 => x"cc",
          7903 => x"8f",
          7904 => x"0a",
          7905 => x"f5",
          7906 => x"f9",
          7907 => x"20",
          7908 => x"22",
          7909 => x"0e",
          7910 => x"d0",
          7911 => x"00",
          7912 => x"63",
          7913 => x"5a",
          7914 => x"06",
          7915 => x"08",
          7916 => x"07",
          7917 => x"54",
          7918 => x"60",
          7919 => x"ba",
          7920 => x"ca",
          7921 => x"f8",
          7922 => x"fa",
          7923 => x"90",
          7924 => x"b0",
          7925 => x"b2",
          7926 => x"c3",
          7927 => x"02",
          7928 => x"f3",
          7929 => x"01",
          7930 => x"84",
          7931 => x"1a",
          7932 => x"02",
          7933 => x"02",
          7934 => x"26",
          7935 => x"00",
          7936 => x"02",
          7937 => x"00",
          7938 => x"04",
          7939 => x"00",
          7940 => x"14",
          7941 => x"00",
          7942 => x"2b",
          7943 => x"00",
          7944 => x"30",
          7945 => x"00",
          7946 => x"3c",
          7947 => x"00",
          7948 => x"3d",
          7949 => x"00",
          7950 => x"3f",
          7951 => x"00",
          7952 => x"40",
          7953 => x"00",
          7954 => x"41",
          7955 => x"00",
          7956 => x"42",
          7957 => x"00",
          7958 => x"43",
          7959 => x"00",
          7960 => x"50",
          7961 => x"00",
          7962 => x"51",
          7963 => x"00",
          7964 => x"54",
          7965 => x"00",
          7966 => x"55",
          7967 => x"00",
          7968 => x"79",
          7969 => x"00",
          7970 => x"78",
          7971 => x"00",
          7972 => x"82",
          7973 => x"00",
          7974 => x"83",
          7975 => x"00",
          7976 => x"85",
          7977 => x"00",
          7978 => x"87",
          7979 => x"00",
          7980 => x"88",
          7981 => x"00",
          7982 => x"89",
          7983 => x"00",
          7984 => x"8c",
          7985 => x"00",
          7986 => x"8d",
          7987 => x"00",
          7988 => x"8e",
          7989 => x"00",
          7990 => x"8f",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"01",
          7995 => x"01",
          7996 => x"00",
          7997 => x"00",
          7998 => x"00",
          7999 => x"f5",
          8000 => x"f5",
          8001 => x"01",
          8002 => x"01",
          8003 => x"00",
          8004 => x"00",
          8005 => x"00",
          8006 => x"00",
          8007 => x"00",
          8008 => x"00",
          8009 => x"00",
          8010 => x"00",
          8011 => x"00",
          8012 => x"00",
          8013 => x"00",
          8014 => x"00",
          8015 => x"00",
          8016 => x"00",
          8017 => x"00",
          8018 => x"01",
          8019 => x"3b",
          8020 => x"f0",
          8021 => x"76",
          8022 => x"6e",
          8023 => x"66",
          8024 => x"36",
          8025 => x"39",
          8026 => x"f2",
          8027 => x"f0",
          8028 => x"f0",
          8029 => x"3a",
          8030 => x"f0",
          8031 => x"56",
          8032 => x"4e",
          8033 => x"46",
          8034 => x"36",
          8035 => x"39",
          8036 => x"f2",
          8037 => x"f0",
          8038 => x"f0",
          8039 => x"2b",
          8040 => x"f0",
          8041 => x"56",
          8042 => x"4e",
          8043 => x"46",
          8044 => x"26",
          8045 => x"29",
          8046 => x"f8",
          8047 => x"f0",
          8048 => x"f0",
          8049 => x"f0",
          8050 => x"f0",
          8051 => x"16",
          8052 => x"0e",
          8053 => x"06",
          8054 => x"f0",
          8055 => x"1f",
          8056 => x"f0",
          8057 => x"f0",
          8058 => x"f0",
          8059 => x"b5",
          8060 => x"f0",
          8061 => x"a6",
          8062 => x"33",
          8063 => x"43",
          8064 => x"1e",
          8065 => x"a3",
          8066 => x"c4",
          8067 => x"f0",
          8068 => x"f0",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"01",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"e0",
          9105 => x"f9",
          9106 => x"c1",
          9107 => x"e4",
          9108 => x"61",
          9109 => x"69",
          9110 => x"21",
          9111 => x"29",
          9112 => x"01",
          9113 => x"09",
          9114 => x"11",
          9115 => x"19",
          9116 => x"81",
          9117 => x"89",
          9118 => x"91",
          9119 => x"99",
          9120 => x"00",
          9121 => x"00",
          9122 => x"00",
          9123 => x"00",
          9124 => x"00",
          9125 => x"00",
          9126 => x"00",
          9127 => x"00",
          9128 => x"00",
          9129 => x"00",
          9130 => x"00",
          9131 => x"00",
          9132 => x"00",
          9133 => x"00",
          9134 => x"00",
          9135 => x"02",
          9136 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"00",
             3 => x"00",
             4 => x"88",
             5 => x"08",
             6 => x"04",
             7 => x"00",
             8 => x"71",
             9 => x"81",
            10 => x"ff",
            11 => x"00",
            12 => x"71",
            13 => x"83",
            14 => x"2b",
            15 => x"0b",
            16 => x"72",
            17 => x"09",
            18 => x"07",
            19 => x"00",
            20 => x"72",
            21 => x"51",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"09",
            26 => x"0a",
            27 => x"51",
            28 => x"72",
            29 => x"51",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"72",
            45 => x"0b",
            46 => x"00",
            47 => x"00",
            48 => x"72",
            49 => x"09",
            50 => x"06",
            51 => x"00",
            52 => x"71",
            53 => x"06",
            54 => x"0b",
            55 => x"51",
            56 => x"72",
            57 => x"81",
            58 => x"51",
            59 => x"00",
            60 => x"72",
            61 => x"81",
            62 => x"53",
            63 => x"00",
            64 => x"71",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"72",
            69 => x"04",
            70 => x"00",
            71 => x"00",
            72 => x"72",
            73 => x"07",
            74 => x"00",
            75 => x"00",
            76 => x"71",
            77 => x"81",
            78 => x"81",
            79 => x"00",
            80 => x"71",
            81 => x"84",
            82 => x"06",
            83 => x"00",
            84 => x"88",
            85 => x"0b",
            86 => x"88",
            87 => x"0c",
            88 => x"88",
            89 => x"0b",
            90 => x"88",
            91 => x"0c",
            92 => x"72",
            93 => x"81",
            94 => x"73",
            95 => x"07",
            96 => x"72",
            97 => x"09",
            98 => x"06",
            99 => x"06",
           100 => x"05",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"04",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"71",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"04",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"02",
           117 => x"04",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"02",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"0b",
           134 => x"96",
           135 => x"0b",
           136 => x"0b",
           137 => x"d6",
           138 => x"0b",
           139 => x"0b",
           140 => x"96",
           141 => x"0b",
           142 => x"0b",
           143 => x"d7",
           144 => x"0b",
           145 => x"0b",
           146 => x"9b",
           147 => x"0b",
           148 => x"0b",
           149 => x"df",
           150 => x"0b",
           151 => x"0b",
           152 => x"a3",
           153 => x"0b",
           154 => x"0b",
           155 => x"e7",
           156 => x"0b",
           157 => x"0b",
           158 => x"ab",
           159 => x"0b",
           160 => x"0b",
           161 => x"ef",
           162 => x"0b",
           163 => x"0b",
           164 => x"b3",
           165 => x"0b",
           166 => x"0b",
           167 => x"f7",
           168 => x"0b",
           169 => x"0b",
           170 => x"bb",
           171 => x"0b",
           172 => x"0b",
           173 => x"fe",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"04",
           193 => x"0c",
           194 => x"08",
           195 => x"90",
           196 => x"08",
           197 => x"90",
           198 => x"08",
           199 => x"90",
           200 => x"08",
           201 => x"90",
           202 => x"08",
           203 => x"90",
           204 => x"08",
           205 => x"90",
           206 => x"08",
           207 => x"90",
           208 => x"08",
           209 => x"90",
           210 => x"08",
           211 => x"90",
           212 => x"08",
           213 => x"90",
           214 => x"08",
           215 => x"90",
           216 => x"08",
           217 => x"90",
           218 => x"90",
           219 => x"bb",
           220 => x"bb",
           221 => x"84",
           222 => x"84",
           223 => x"04",
           224 => x"2d",
           225 => x"90",
           226 => x"f6",
           227 => x"80",
           228 => x"e3",
           229 => x"c0",
           230 => x"82",
           231 => x"80",
           232 => x"0c",
           233 => x"08",
           234 => x"90",
           235 => x"90",
           236 => x"bb",
           237 => x"bb",
           238 => x"84",
           239 => x"84",
           240 => x"04",
           241 => x"2d",
           242 => x"90",
           243 => x"e2",
           244 => x"80",
           245 => x"f4",
           246 => x"c0",
           247 => x"83",
           248 => x"80",
           249 => x"0c",
           250 => x"08",
           251 => x"90",
           252 => x"90",
           253 => x"bb",
           254 => x"bb",
           255 => x"84",
           256 => x"84",
           257 => x"04",
           258 => x"2d",
           259 => x"90",
           260 => x"d9",
           261 => x"80",
           262 => x"e3",
           263 => x"c0",
           264 => x"82",
           265 => x"80",
           266 => x"0c",
           267 => x"08",
           268 => x"90",
           269 => x"90",
           270 => x"bb",
           271 => x"bb",
           272 => x"84",
           273 => x"84",
           274 => x"04",
           275 => x"2d",
           276 => x"90",
           277 => x"a1",
           278 => x"80",
           279 => x"ba",
           280 => x"c0",
           281 => x"83",
           282 => x"80",
           283 => x"0c",
           284 => x"08",
           285 => x"90",
           286 => x"90",
           287 => x"bb",
           288 => x"bb",
           289 => x"84",
           290 => x"84",
           291 => x"04",
           292 => x"2d",
           293 => x"90",
           294 => x"b5",
           295 => x"80",
           296 => x"9a",
           297 => x"80",
           298 => x"dc",
           299 => x"c0",
           300 => x"81",
           301 => x"80",
           302 => x"0c",
           303 => x"08",
           304 => x"90",
           305 => x"90",
           306 => x"04",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"53",
           311 => x"06",
           312 => x"05",
           313 => x"06",
           314 => x"72",
           315 => x"05",
           316 => x"53",
           317 => x"04",
           318 => x"27",
           319 => x"53",
           320 => x"8c",
           321 => x"fc",
           322 => x"05",
           323 => x"e6",
           324 => x"3d",
           325 => x"7c",
           326 => x"80",
           327 => x"80",
           328 => x"80",
           329 => x"32",
           330 => x"51",
           331 => x"b7",
           332 => x"51",
           333 => x"53",
           334 => x"38",
           335 => x"05",
           336 => x"70",
           337 => x"54",
           338 => x"80",
           339 => x"84",
           340 => x"84",
           341 => x"f5",
           342 => x"05",
           343 => x"58",
           344 => x"8d",
           345 => x"19",
           346 => x"04",
           347 => x"53",
           348 => x"3d",
           349 => x"65",
           350 => x"0c",
           351 => x"32",
           352 => x"72",
           353 => x"38",
           354 => x"c5",
           355 => x"5c",
           356 => x"17",
           357 => x"76",
           358 => x"51",
           359 => x"2e",
           360 => x"32",
           361 => x"9e",
           362 => x"33",
           363 => x"08",
           364 => x"3d",
           365 => x"10",
           366 => x"2b",
           367 => x"0a",
           368 => x"52",
           369 => x"81",
           370 => x"ff",
           371 => x"76",
           372 => x"a5",
           373 => x"73",
           374 => x"58",
           375 => x"39",
           376 => x"7b",
           377 => x"8d",
           378 => x"54",
           379 => x"06",
           380 => x"53",
           381 => x"10",
           382 => x"08",
           383 => x"d8",
           384 => x"51",
           385 => x"5b",
           386 => x"80",
           387 => x"7f",
           388 => x"ff",
           389 => x"bb",
           390 => x"9a",
           391 => x"06",
           392 => x"56",
           393 => x"bb",
           394 => x"70",
           395 => x"51",
           396 => x"56",
           397 => x"84",
           398 => x"06",
           399 => x"77",
           400 => x"05",
           401 => x"2a",
           402 => x"2e",
           403 => x"f8",
           404 => x"8b",
           405 => x"80",
           406 => x"7a",
           407 => x"72",
           408 => x"70",
           409 => x"24",
           410 => x"06",
           411 => x"56",
           412 => x"2e",
           413 => x"2b",
           414 => x"56",
           415 => x"38",
           416 => x"85",
           417 => x"54",
           418 => x"81",
           419 => x"81",
           420 => x"88",
           421 => x"b2",
           422 => x"fc",
           423 => x"40",
           424 => x"52",
           425 => x"84",
           426 => x"70",
           427 => x"24",
           428 => x"80",
           429 => x"0a",
           430 => x"2c",
           431 => x"38",
           432 => x"78",
           433 => x"0a",
           434 => x"74",
           435 => x"70",
           436 => x"81",
           437 => x"d8",
           438 => x"38",
           439 => x"7d",
           440 => x"52",
           441 => x"a5",
           442 => x"81",
           443 => x"7a",
           444 => x"84",
           445 => x"70",
           446 => x"25",
           447 => x"86",
           448 => x"5b",
           449 => x"76",
           450 => x"80",
           451 => x"60",
           452 => x"ff",
           453 => x"fb",
           454 => x"fe",
           455 => x"98",
           456 => x"29",
           457 => x"5e",
           458 => x"87",
           459 => x"fe",
           460 => x"29",
           461 => x"5a",
           462 => x"38",
           463 => x"e2",
           464 => x"06",
           465 => x"fe",
           466 => x"05",
           467 => x"39",
           468 => x"5b",
           469 => x"ab",
           470 => x"57",
           471 => x"75",
           472 => x"78",
           473 => x"05",
           474 => x"e3",
           475 => x"56",
           476 => x"39",
           477 => x"53",
           478 => x"df",
           479 => x"84",
           480 => x"84",
           481 => x"89",
           482 => x"5b",
           483 => x"f9",
           484 => x"05",
           485 => x"41",
           486 => x"87",
           487 => x"ff",
           488 => x"54",
           489 => x"39",
           490 => x"5b",
           491 => x"7f",
           492 => x"06",
           493 => x"38",
           494 => x"84",
           495 => x"31",
           496 => x"81",
           497 => x"f7",
           498 => x"84",
           499 => x"70",
           500 => x"25",
           501 => x"83",
           502 => x"51",
           503 => x"81",
           504 => x"51",
           505 => x"06",
           506 => x"fa",
           507 => x"31",
           508 => x"80",
           509 => x"90",
           510 => x"51",
           511 => x"73",
           512 => x"39",
           513 => x"e5",
           514 => x"2e",
           515 => x"74",
           516 => x"53",
           517 => x"82",
           518 => x"51",
           519 => x"52",
           520 => x"84",
           521 => x"31",
           522 => x"7a",
           523 => x"bf",
           524 => x"fe",
           525 => x"75",
           526 => x"3d",
           527 => x"80",
           528 => x"33",
           529 => x"06",
           530 => x"72",
           531 => x"38",
           532 => x"72",
           533 => x"08",
           534 => x"72",
           535 => x"83",
           536 => x"56",
           537 => x"84",
           538 => x"e6",
           539 => x"52",
           540 => x"2d",
           541 => x"38",
           542 => x"84",
           543 => x"0d",
           544 => x"16",
           545 => x"81",
           546 => x"72",
           547 => x"73",
           548 => x"77",
           549 => x"56",
           550 => x"0d",
           551 => x"53",
           552 => x"72",
           553 => x"84",
           554 => x"ff",
           555 => x"57",
           556 => x"0d",
           557 => x"85",
           558 => x"0d",
           559 => x"2a",
           560 => x"57",
           561 => x"2a",
           562 => x"38",
           563 => x"08",
           564 => x"76",
           565 => x"8c",
           566 => x"0c",
           567 => x"88",
           568 => x"ff",
           569 => x"2d",
           570 => x"38",
           571 => x"0c",
           572 => x"77",
           573 => x"70",
           574 => x"56",
           575 => x"2a",
           576 => x"82",
           577 => x"80",
           578 => x"53",
           579 => x"13",
           580 => x"8c",
           581 => x"73",
           582 => x"04",
           583 => x"17",
           584 => x"17",
           585 => x"0c",
           586 => x"16",
           587 => x"08",
           588 => x"ff",
           589 => x"07",
           590 => x"2e",
           591 => x"85",
           592 => x"84",
           593 => x"07",
           594 => x"ec",
           595 => x"54",
           596 => x"33",
           597 => x"72",
           598 => x"72",
           599 => x"38",
           600 => x"0d",
           601 => x"7a",
           602 => x"9d",
           603 => x"80",
           604 => x"53",
           605 => x"ff",
           606 => x"bb",
           607 => x"12",
           608 => x"14",
           609 => x"53",
           610 => x"51",
           611 => x"ff",
           612 => x"ff",
           613 => x"fe",
           614 => x"70",
           615 => x"38",
           616 => x"84",
           617 => x"3d",
           618 => x"72",
           619 => x"72",
           620 => x"38",
           621 => x"0d",
           622 => x"79",
           623 => x"93",
           624 => x"73",
           625 => x"51",
           626 => x"0c",
           627 => x"76",
           628 => x"2e",
           629 => x"05",
           630 => x"09",
           631 => x"71",
           632 => x"72",
           633 => x"84",
           634 => x"2e",
           635 => x"72",
           636 => x"52",
           637 => x"72",
           638 => x"3d",
           639 => x"86",
           640 => x"79",
           641 => x"84",
           642 => x"81",
           643 => x"84",
           644 => x"08",
           645 => x"08",
           646 => x"75",
           647 => x"b1",
           648 => x"84",
           649 => x"fd",
           650 => x"55",
           651 => x"72",
           652 => x"80",
           653 => x"ff",
           654 => x"13",
           655 => x"bb",
           656 => x"3d",
           657 => x"54",
           658 => x"72",
           659 => x"51",
           660 => x"0c",
           661 => x"78",
           662 => x"2e",
           663 => x"84",
           664 => x"73",
           665 => x"e3",
           666 => x"53",
           667 => x"38",
           668 => x"38",
           669 => x"31",
           670 => x"80",
           671 => x"10",
           672 => x"07",
           673 => x"70",
           674 => x"31",
           675 => x"58",
           676 => x"76",
           677 => x"88",
           678 => x"70",
           679 => x"72",
           680 => x"71",
           681 => x"80",
           682 => x"2b",
           683 => x"81",
           684 => x"82",
           685 => x"55",
           686 => x"70",
           687 => x"31",
           688 => x"32",
           689 => x"31",
           690 => x"0c",
           691 => x"5a",
           692 => x"56",
           693 => x"3d",
           694 => x"70",
           695 => x"3f",
           696 => x"71",
           697 => x"3d",
           698 => x"58",
           699 => x"38",
           700 => x"84",
           701 => x"2e",
           702 => x"72",
           703 => x"53",
           704 => x"53",
           705 => x"74",
           706 => x"2b",
           707 => x"76",
           708 => x"2a",
           709 => x"31",
           710 => x"7b",
           711 => x"5c",
           712 => x"74",
           713 => x"88",
           714 => x"9f",
           715 => x"7b",
           716 => x"73",
           717 => x"31",
           718 => x"b4",
           719 => x"75",
           720 => x"0d",
           721 => x"57",
           722 => x"33",
           723 => x"81",
           724 => x"0c",
           725 => x"f3",
           726 => x"73",
           727 => x"58",
           728 => x"38",
           729 => x"80",
           730 => x"38",
           731 => x"53",
           732 => x"53",
           733 => x"70",
           734 => x"27",
           735 => x"83",
           736 => x"70",
           737 => x"73",
           738 => x"2e",
           739 => x"0c",
           740 => x"8b",
           741 => x"79",
           742 => x"b0",
           743 => x"81",
           744 => x"55",
           745 => x"58",
           746 => x"56",
           747 => x"53",
           748 => x"fe",
           749 => x"8b",
           750 => x"70",
           751 => x"56",
           752 => x"84",
           753 => x"0d",
           754 => x"0c",
           755 => x"73",
           756 => x"81",
           757 => x"55",
           758 => x"2e",
           759 => x"83",
           760 => x"89",
           761 => x"56",
           762 => x"e0",
           763 => x"81",
           764 => x"81",
           765 => x"8f",
           766 => x"54",
           767 => x"72",
           768 => x"29",
           769 => x"33",
           770 => x"be",
           771 => x"30",
           772 => x"84",
           773 => x"81",
           774 => x"56",
           775 => x"06",
           776 => x"0c",
           777 => x"2e",
           778 => x"2e",
           779 => x"c6",
           780 => x"58",
           781 => x"84",
           782 => x"82",
           783 => x"33",
           784 => x"80",
           785 => x"0d",
           786 => x"84",
           787 => x"0c",
           788 => x"93",
           789 => x"bf",
           790 => x"cf",
           791 => x"0d",
           792 => x"3f",
           793 => x"51",
           794 => x"83",
           795 => x"3d",
           796 => x"92",
           797 => x"94",
           798 => x"04",
           799 => x"83",
           800 => x"ee",
           801 => x"d0",
           802 => x"0d",
           803 => x"3f",
           804 => x"51",
           805 => x"83",
           806 => x"3d",
           807 => x"ba",
           808 => x"e4",
           809 => x"04",
           810 => x"83",
           811 => x"ee",
           812 => x"d2",
           813 => x"0d",
           814 => x"3f",
           815 => x"51",
           816 => x"83",
           817 => x"3d",
           818 => x"e2",
           819 => x"3d",
           820 => x"05",
           821 => x"0b",
           822 => x"7b",
           823 => x"78",
           824 => x"81",
           825 => x"06",
           826 => x"38",
           827 => x"52",
           828 => x"84",
           829 => x"2e",
           830 => x"98",
           831 => x"25",
           832 => x"53",
           833 => x"38",
           834 => x"87",
           835 => x"78",
           836 => x"84",
           837 => x"53",
           838 => x"d7",
           839 => x"96",
           840 => x"87",
           841 => x"08",
           842 => x"54",
           843 => x"82",
           844 => x"57",
           845 => x"7a",
           846 => x"74",
           847 => x"87",
           848 => x"84",
           849 => x"9c",
           850 => x"d3",
           851 => x"51",
           852 => x"3d",
           853 => x"33",
           854 => x"52",
           855 => x"84",
           856 => x"38",
           857 => x"bb",
           858 => x"04",
           859 => x"54",
           860 => x"51",
           861 => x"bb",
           862 => x"3d",
           863 => x"80",
           864 => x"41",
           865 => x"80",
           866 => x"d3",
           867 => x"94",
           868 => x"79",
           869 => x"ed",
           870 => x"73",
           871 => x"38",
           872 => x"dd",
           873 => x"08",
           874 => x"78",
           875 => x"51",
           876 => x"27",
           877 => x"55",
           878 => x"38",
           879 => x"83",
           880 => x"81",
           881 => x"88",
           882 => x"38",
           883 => x"eb",
           884 => x"26",
           885 => x"ca",
           886 => x"80",
           887 => x"08",
           888 => x"76",
           889 => x"2e",
           890 => x"78",
           891 => x"bb",
           892 => x"d3",
           893 => x"84",
           894 => x"ea",
           895 => x"38",
           896 => x"dc",
           897 => x"08",
           898 => x"73",
           899 => x"53",
           900 => x"52",
           901 => x"82",
           902 => x"a0",
           903 => x"dd",
           904 => x"51",
           905 => x"e8",
           906 => x"3f",
           907 => x"18",
           908 => x"08",
           909 => x"3f",
           910 => x"54",
           911 => x"26",
           912 => x"e8",
           913 => x"81",
           914 => x"a6",
           915 => x"06",
           916 => x"ec",
           917 => x"09",
           918 => x"fc",
           919 => x"84",
           920 => x"2c",
           921 => x"32",
           922 => x"07",
           923 => x"53",
           924 => x"51",
           925 => x"98",
           926 => x"70",
           927 => x"72",
           928 => x"58",
           929 => x"ff",
           930 => x"84",
           931 => x"fe",
           932 => x"53",
           933 => x"3f",
           934 => x"80",
           935 => x"70",
           936 => x"38",
           937 => x"52",
           938 => x"70",
           939 => x"38",
           940 => x"52",
           941 => x"70",
           942 => x"38",
           943 => x"52",
           944 => x"70",
           945 => x"72",
           946 => x"38",
           947 => x"81",
           948 => x"51",
           949 => x"3f",
           950 => x"81",
           951 => x"51",
           952 => x"3f",
           953 => x"80",
           954 => x"9b",
           955 => x"f4",
           956 => x"87",
           957 => x"80",
           958 => x"51",
           959 => x"9b",
           960 => x"72",
           961 => x"71",
           962 => x"39",
           963 => x"b8",
           964 => x"94",
           965 => x"51",
           966 => x"ff",
           967 => x"83",
           968 => x"51",
           969 => x"81",
           970 => x"94",
           971 => x"dc",
           972 => x"3f",
           973 => x"2a",
           974 => x"2e",
           975 => x"51",
           976 => x"9a",
           977 => x"72",
           978 => x"71",
           979 => x"39",
           980 => x"ff",
           981 => x"52",
           982 => x"bb",
           983 => x"40",
           984 => x"83",
           985 => x"3d",
           986 => x"3f",
           987 => x"7e",
           988 => x"ef",
           989 => x"59",
           990 => x"81",
           991 => x"06",
           992 => x"67",
           993 => x"e0",
           994 => x"09",
           995 => x"33",
           996 => x"80",
           997 => x"90",
           998 => x"52",
           999 => x"08",
          1000 => x"7b",
          1001 => x"bb",
          1002 => x"5e",
          1003 => x"1c",
          1004 => x"7c",
          1005 => x"7b",
          1006 => x"52",
          1007 => x"84",
          1008 => x"2e",
          1009 => x"48",
          1010 => x"a9",
          1011 => x"06",
          1012 => x"38",
          1013 => x"3f",
          1014 => x"f3",
          1015 => x"7a",
          1016 => x"24",
          1017 => x"e8",
          1018 => x"80",
          1019 => x"f3",
          1020 => x"56",
          1021 => x"53",
          1022 => x"ae",
          1023 => x"84",
          1024 => x"80",
          1025 => x"7a",
          1026 => x"7a",
          1027 => x"81",
          1028 => x"7a",
          1029 => x"81",
          1030 => x"61",
          1031 => x"81",
          1032 => x"d3",
          1033 => x"80",
          1034 => x"0b",
          1035 => x"06",
          1036 => x"53",
          1037 => x"51",
          1038 => x"08",
          1039 => x"83",
          1040 => x"80",
          1041 => x"3f",
          1042 => x"38",
          1043 => x"3f",
          1044 => x"81",
          1045 => x"09",
          1046 => x"84",
          1047 => x"82",
          1048 => x"80",
          1049 => x"80",
          1050 => x"67",
          1051 => x"90",
          1052 => x"33",
          1053 => x"38",
          1054 => x"5a",
          1055 => x"88",
          1056 => x"53",
          1057 => x"86",
          1058 => x"2e",
          1059 => x"70",
          1060 => x"39",
          1061 => x"7d",
          1062 => x"39",
          1063 => x"d7",
          1064 => x"52",
          1065 => x"39",
          1066 => x"9a",
          1067 => x"83",
          1068 => x"39",
          1069 => x"83",
          1070 => x"59",
          1071 => x"fa",
          1072 => x"b8",
          1073 => x"05",
          1074 => x"08",
          1075 => x"83",
          1076 => x"5a",
          1077 => x"2e",
          1078 => x"52",
          1079 => x"fa",
          1080 => x"53",
          1081 => x"84",
          1082 => x"38",
          1083 => x"af",
          1084 => x"fe",
          1085 => x"e9",
          1086 => x"2e",
          1087 => x"11",
          1088 => x"3f",
          1089 => x"64",
          1090 => x"d8",
          1091 => x"e4",
          1092 => x"d0",
          1093 => x"78",
          1094 => x"26",
          1095 => x"46",
          1096 => x"11",
          1097 => x"3f",
          1098 => x"f9",
          1099 => x"ff",
          1100 => x"bb",
          1101 => x"78",
          1102 => x"51",
          1103 => x"53",
          1104 => x"3f",
          1105 => x"2e",
          1106 => x"ca",
          1107 => x"cf",
          1108 => x"ff",
          1109 => x"bb",
          1110 => x"b8",
          1111 => x"05",
          1112 => x"08",
          1113 => x"fe",
          1114 => x"e9",
          1115 => x"2e",
          1116 => x"ce",
          1117 => x"7c",
          1118 => x"7a",
          1119 => x"95",
          1120 => x"53",
          1121 => x"ff",
          1122 => x"81",
          1123 => x"ff",
          1124 => x"e8",
          1125 => x"2e",
          1126 => x"11",
          1127 => x"3f",
          1128 => x"89",
          1129 => x"ff",
          1130 => x"bb",
          1131 => x"83",
          1132 => x"5a",
          1133 => x"5c",
          1134 => x"34",
          1135 => x"3d",
          1136 => x"51",
          1137 => x"80",
          1138 => x"fc",
          1139 => x"ed",
          1140 => x"68",
          1141 => x"51",
          1142 => x"53",
          1143 => x"3f",
          1144 => x"2e",
          1145 => x"97",
          1146 => x"68",
          1147 => x"34",
          1148 => x"fc",
          1149 => x"9d",
          1150 => x"f5",
          1151 => x"05",
          1152 => x"b8",
          1153 => x"05",
          1154 => x"08",
          1155 => x"3d",
          1156 => x"51",
          1157 => x"80",
          1158 => x"fc",
          1159 => x"cd",
          1160 => x"f5",
          1161 => x"53",
          1162 => x"84",
          1163 => x"84",
          1164 => x"a7",
          1165 => x"27",
          1166 => x"84",
          1167 => x"38",
          1168 => x"39",
          1169 => x"b1",
          1170 => x"ff",
          1171 => x"81",
          1172 => x"51",
          1173 => x"80",
          1174 => x"08",
          1175 => x"b8",
          1176 => x"05",
          1177 => x"08",
          1178 => x"79",
          1179 => x"c0",
          1180 => x"53",
          1181 => x"84",
          1182 => x"88",
          1183 => x"38",
          1184 => x"fe",
          1185 => x"e4",
          1186 => x"2e",
          1187 => x"88",
          1188 => x"32",
          1189 => x"7e",
          1190 => x"88",
          1191 => x"46",
          1192 => x"80",
          1193 => x"68",
          1194 => x"51",
          1195 => x"64",
          1196 => x"b8",
          1197 => x"05",
          1198 => x"08",
          1199 => x"71",
          1200 => x"3d",
          1201 => x"51",
          1202 => x"c6",
          1203 => x"80",
          1204 => x"40",
          1205 => x"11",
          1206 => x"3f",
          1207 => x"91",
          1208 => x"22",
          1209 => x"45",
          1210 => x"80",
          1211 => x"84",
          1212 => x"b8",
          1213 => x"05",
          1214 => x"08",
          1215 => x"02",
          1216 => x"81",
          1217 => x"fe",
          1218 => x"e0",
          1219 => x"2e",
          1220 => x"5d",
          1221 => x"e1",
          1222 => x"f3",
          1223 => x"54",
          1224 => x"51",
          1225 => x"52",
          1226 => x"39",
          1227 => x"f0",
          1228 => x"53",
          1229 => x"84",
          1230 => x"64",
          1231 => x"70",
          1232 => x"e7",
          1233 => x"80",
          1234 => x"08",
          1235 => x"33",
          1236 => x"f3",
          1237 => x"d9",
          1238 => x"f7",
          1239 => x"ba",
          1240 => x"f4",
          1241 => x"38",
          1242 => x"39",
          1243 => x"f9",
          1244 => x"78",
          1245 => x"08",
          1246 => x"33",
          1247 => x"f3",
          1248 => x"f4",
          1249 => x"38",
          1250 => x"39",
          1251 => x"2e",
          1252 => x"fb",
          1253 => x"7c",
          1254 => x"08",
          1255 => x"08",
          1256 => x"83",
          1257 => x"b5",
          1258 => x"bb",
          1259 => x"08",
          1260 => x"51",
          1261 => x"90",
          1262 => x"80",
          1263 => x"84",
          1264 => x"c0",
          1265 => x"84",
          1266 => x"84",
          1267 => x"57",
          1268 => x"da",
          1269 => x"07",
          1270 => x"c0",
          1271 => x"87",
          1272 => x"5c",
          1273 => x"05",
          1274 => x"e4",
          1275 => x"70",
          1276 => x"b8",
          1277 => x"3f",
          1278 => x"d3",
          1279 => x"8f",
          1280 => x"55",
          1281 => x"83",
          1282 => x"83",
          1283 => x"b2",
          1284 => x"3f",
          1285 => x"df",
          1286 => x"a8",
          1287 => x"80",
          1288 => x"56",
          1289 => x"2e",
          1290 => x"ff",
          1291 => x"81",
          1292 => x"70",
          1293 => x"a0",
          1294 => x"54",
          1295 => x"52",
          1296 => x"72",
          1297 => x"54",
          1298 => x"70",
          1299 => x"86",
          1300 => x"73",
          1301 => x"2e",
          1302 => x"70",
          1303 => x"76",
          1304 => x"88",
          1305 => x"34",
          1306 => x"bb",
          1307 => x"80",
          1308 => x"be",
          1309 => x"70",
          1310 => x"a2",
          1311 => x"81",
          1312 => x"81",
          1313 => x"dc",
          1314 => x"08",
          1315 => x"0c",
          1316 => x"05",
          1317 => x"bb",
          1318 => x"84",
          1319 => x"fc",
          1320 => x"05",
          1321 => x"81",
          1322 => x"54",
          1323 => x"38",
          1324 => x"97",
          1325 => x"54",
          1326 => x"38",
          1327 => x"bb",
          1328 => x"55",
          1329 => x"d9",
          1330 => x"73",
          1331 => x"0b",
          1332 => x"87",
          1333 => x"87",
          1334 => x"87",
          1335 => x"87",
          1336 => x"87",
          1337 => x"87",
          1338 => x"98",
          1339 => x"0c",
          1340 => x"80",
          1341 => x"3d",
          1342 => x"87",
          1343 => x"87",
          1344 => x"23",
          1345 => x"82",
          1346 => x"5a",
          1347 => x"b0",
          1348 => x"c0",
          1349 => x"34",
          1350 => x"86",
          1351 => x"5c",
          1352 => x"a0",
          1353 => x"7d",
          1354 => x"7b",
          1355 => x"33",
          1356 => x"33",
          1357 => x"33",
          1358 => x"83",
          1359 => x"8f",
          1360 => x"93",
          1361 => x"38",
          1362 => x"bb",
          1363 => x"51",
          1364 => x"86",
          1365 => x"84",
          1366 => x"72",
          1367 => x"84",
          1368 => x"52",
          1369 => x"38",
          1370 => x"bb",
          1371 => x"51",
          1372 => x"39",
          1373 => x"71",
          1374 => x"fb",
          1375 => x"70",
          1376 => x"eb",
          1377 => x"52",
          1378 => x"bb",
          1379 => x"3d",
          1380 => x"bc",
          1381 => x"55",
          1382 => x"c0",
          1383 => x"81",
          1384 => x"8c",
          1385 => x"51",
          1386 => x"81",
          1387 => x"71",
          1388 => x"38",
          1389 => x"94",
          1390 => x"87",
          1391 => x"74",
          1392 => x"04",
          1393 => x"51",
          1394 => x"06",
          1395 => x"93",
          1396 => x"c0",
          1397 => x"96",
          1398 => x"70",
          1399 => x"02",
          1400 => x"2a",
          1401 => x"34",
          1402 => x"78",
          1403 => x"57",
          1404 => x"15",
          1405 => x"06",
          1406 => x"ff",
          1407 => x"96",
          1408 => x"70",
          1409 => x"70",
          1410 => x"72",
          1411 => x"2e",
          1412 => x"52",
          1413 => x"51",
          1414 => x"2e",
          1415 => x"73",
          1416 => x"57",
          1417 => x"84",
          1418 => x"2a",
          1419 => x"38",
          1420 => x"80",
          1421 => x"06",
          1422 => x"87",
          1423 => x"70",
          1424 => x"38",
          1425 => x"9e",
          1426 => x"52",
          1427 => x"87",
          1428 => x"0c",
          1429 => x"c4",
          1430 => x"f3",
          1431 => x"83",
          1432 => x"08",
          1433 => x"a0",
          1434 => x"9e",
          1435 => x"c0",
          1436 => x"87",
          1437 => x"0c",
          1438 => x"e4",
          1439 => x"f3",
          1440 => x"83",
          1441 => x"08",
          1442 => x"80",
          1443 => x"87",
          1444 => x"0c",
          1445 => x"fc",
          1446 => x"f4",
          1447 => x"34",
          1448 => x"70",
          1449 => x"70",
          1450 => x"34",
          1451 => x"70",
          1452 => x"70",
          1453 => x"83",
          1454 => x"9e",
          1455 => x"51",
          1456 => x"81",
          1457 => x"0b",
          1458 => x"80",
          1459 => x"2e",
          1460 => x"88",
          1461 => x"08",
          1462 => x"52",
          1463 => x"71",
          1464 => x"c0",
          1465 => x"06",
          1466 => x"38",
          1467 => x"80",
          1468 => x"84",
          1469 => x"80",
          1470 => x"f4",
          1471 => x"90",
          1472 => x"52",
          1473 => x"52",
          1474 => x"87",
          1475 => x"80",
          1476 => x"83",
          1477 => x"34",
          1478 => x"70",
          1479 => x"70",
          1480 => x"83",
          1481 => x"9e",
          1482 => x"52",
          1483 => x"52",
          1484 => x"9e",
          1485 => x"2a",
          1486 => x"80",
          1487 => x"84",
          1488 => x"2e",
          1489 => x"91",
          1490 => x"f0",
          1491 => x"83",
          1492 => x"9e",
          1493 => x"52",
          1494 => x"71",
          1495 => x"90",
          1496 => x"94",
          1497 => x"fd",
          1498 => x"94",
          1499 => x"84",
          1500 => x"da",
          1501 => x"86",
          1502 => x"f4",
          1503 => x"83",
          1504 => x"38",
          1505 => x"f5",
          1506 => x"84",
          1507 => x"75",
          1508 => x"54",
          1509 => x"33",
          1510 => x"85",
          1511 => x"f4",
          1512 => x"83",
          1513 => x"38",
          1514 => x"ea",
          1515 => x"81",
          1516 => x"92",
          1517 => x"da",
          1518 => x"f3",
          1519 => x"ff",
          1520 => x"52",
          1521 => x"3f",
          1522 => x"83",
          1523 => x"51",
          1524 => x"08",
          1525 => x"c9",
          1526 => x"84",
          1527 => x"84",
          1528 => x"51",
          1529 => x"33",
          1530 => x"33",
          1531 => x"04",
          1532 => x"c0",
          1533 => x"bb",
          1534 => x"71",
          1535 => x"52",
          1536 => x"3f",
          1537 => x"08",
          1538 => x"c9",
          1539 => x"84",
          1540 => x"84",
          1541 => x"51",
          1542 => x"33",
          1543 => x"ff",
          1544 => x"b2",
          1545 => x"3f",
          1546 => x"cc",
          1547 => x"ec",
          1548 => x"b3",
          1549 => x"83",
          1550 => x"83",
          1551 => x"83",
          1552 => x"51",
          1553 => x"08",
          1554 => x"c8",
          1555 => x"84",
          1556 => x"84",
          1557 => x"51",
          1558 => x"33",
          1559 => x"fe",
          1560 => x"bf",
          1561 => x"73",
          1562 => x"39",
          1563 => x"3f",
          1564 => x"2e",
          1565 => x"94",
          1566 => x"8c",
          1567 => x"38",
          1568 => x"be",
          1569 => x"73",
          1570 => x"83",
          1571 => x"51",
          1572 => x"33",
          1573 => x"d2",
          1574 => x"dd",
          1575 => x"f4",
          1576 => x"ed",
          1577 => x"52",
          1578 => x"3f",
          1579 => x"2e",
          1580 => x"d0",
          1581 => x"52",
          1582 => x"3f",
          1583 => x"2e",
          1584 => x"c8",
          1585 => x"52",
          1586 => x"3f",
          1587 => x"2e",
          1588 => x"c0",
          1589 => x"52",
          1590 => x"3f",
          1591 => x"2e",
          1592 => x"d8",
          1593 => x"52",
          1594 => x"3f",
          1595 => x"2e",
          1596 => x"e0",
          1597 => x"52",
          1598 => x"3f",
          1599 => x"2e",
          1600 => x"a0",
          1601 => x"a8",
          1602 => x"86",
          1603 => x"38",
          1604 => x"05",
          1605 => x"71",
          1606 => x"71",
          1607 => x"af",
          1608 => x"df",
          1609 => x"3d",
          1610 => x"af",
          1611 => x"df",
          1612 => x"3d",
          1613 => x"af",
          1614 => x"df",
          1615 => x"3d",
          1616 => x"80",
          1617 => x"83",
          1618 => x"0c",
          1619 => x"ad",
          1620 => x"58",
          1621 => x"82",
          1622 => x"80",
          1623 => x"83",
          1624 => x"52",
          1625 => x"bb",
          1626 => x"51",
          1627 => x"81",
          1628 => x"84",
          1629 => x"08",
          1630 => x"74",
          1631 => x"07",
          1632 => x"2e",
          1633 => x"f4",
          1634 => x"82",
          1635 => x"8f",
          1636 => x"84",
          1637 => x"83",
          1638 => x"78",
          1639 => x"76",
          1640 => x"51",
          1641 => x"56",
          1642 => x"52",
          1643 => x"3f",
          1644 => x"3d",
          1645 => x"08",
          1646 => x"33",
          1647 => x"81",
          1648 => x"56",
          1649 => x"05",
          1650 => x"3f",
          1651 => x"73",
          1652 => x"bb",
          1653 => x"54",
          1654 => x"82",
          1655 => x"ff",
          1656 => x"38",
          1657 => x"aa",
          1658 => x"3d",
          1659 => x"51",
          1660 => x"80",
          1661 => x"52",
          1662 => x"84",
          1663 => x"2e",
          1664 => x"06",
          1665 => x"38",
          1666 => x"56",
          1667 => x"15",
          1668 => x"a0",
          1669 => x"75",
          1670 => x"3d",
          1671 => x"bb",
          1672 => x"52",
          1673 => x"84",
          1674 => x"08",
          1675 => x"cf",
          1676 => x"2e",
          1677 => x"3f",
          1678 => x"84",
          1679 => x"bb",
          1680 => x"55",
          1681 => x"81",
          1682 => x"aa",
          1683 => x"06",
          1684 => x"84",
          1685 => x"0d",
          1686 => x"3d",
          1687 => x"42",
          1688 => x"3d",
          1689 => x"83",
          1690 => x"55",
          1691 => x"06",
          1692 => x"38",
          1693 => x"70",
          1694 => x"38",
          1695 => x"3d",
          1696 => x"fb",
          1697 => x"70",
          1698 => x"81",
          1699 => x"e2",
          1700 => x"2c",
          1701 => x"70",
          1702 => x"10",
          1703 => x"15",
          1704 => x"52",
          1705 => x"79",
          1706 => x"81",
          1707 => x"81",
          1708 => x"42",
          1709 => x"10",
          1710 => x"0b",
          1711 => x"77",
          1712 => x"15",
          1713 => x"75",
          1714 => x"c2",
          1715 => x"57",
          1716 => x"1b",
          1717 => x"e2",
          1718 => x"2c",
          1719 => x"83",
          1720 => x"5e",
          1721 => x"81",
          1722 => x"80",
          1723 => x"08",
          1724 => x"79",
          1725 => x"38",
          1726 => x"2d",
          1727 => x"99",
          1728 => x"80",
          1729 => x"ff",
          1730 => x"80",
          1731 => x"2b",
          1732 => x"16",
          1733 => x"38",
          1734 => x"33",
          1735 => x"38",
          1736 => x"d1",
          1737 => x"8a",
          1738 => x"90",
          1739 => x"76",
          1740 => x"bc",
          1741 => x"63",
          1742 => x"74",
          1743 => x"76",
          1744 => x"60",
          1745 => x"80",
          1746 => x"84",
          1747 => x"fc",
          1748 => x"88",
          1749 => x"c8",
          1750 => x"c8",
          1751 => x"33",
          1752 => x"33",
          1753 => x"b4",
          1754 => x"15",
          1755 => x"16",
          1756 => x"3f",
          1757 => x"bd",
          1758 => x"10",
          1759 => x"57",
          1760 => x"84",
          1761 => x"e2",
          1762 => x"56",
          1763 => x"e8",
          1764 => x"3f",
          1765 => x"ff",
          1766 => x"52",
          1767 => x"e2",
          1768 => x"e2",
          1769 => x"74",
          1770 => x"3f",
          1771 => x"39",
          1772 => x"56",
          1773 => x"81",
          1774 => x"90",
          1775 => x"05",
          1776 => x"38",
          1777 => x"10",
          1778 => x"57",
          1779 => x"75",
          1780 => x"84",
          1781 => x"84",
          1782 => x"75",
          1783 => x"84",
          1784 => x"56",
          1785 => x"84",
          1786 => x"b3",
          1787 => x"a0",
          1788 => x"e8",
          1789 => x"3f",
          1790 => x"74",
          1791 => x"06",
          1792 => x"70",
          1793 => x"5c",
          1794 => x"38",
          1795 => x"57",
          1796 => x"70",
          1797 => x"84",
          1798 => x"84",
          1799 => x"78",
          1800 => x"08",
          1801 => x"c8",
          1802 => x"ff",
          1803 => x"70",
          1804 => x"5a",
          1805 => x"38",
          1806 => x"84",
          1807 => x"2e",
          1808 => x"84",
          1809 => x"98",
          1810 => x"59",
          1811 => x"e6",
          1812 => x"cd",
          1813 => x"2b",
          1814 => x"5a",
          1815 => x"c4",
          1816 => x"51",
          1817 => x"0a",
          1818 => x"2c",
          1819 => x"74",
          1820 => x"e8",
          1821 => x"3f",
          1822 => x"0a",
          1823 => x"33",
          1824 => x"b9",
          1825 => x"81",
          1826 => x"08",
          1827 => x"3f",
          1828 => x"0a",
          1829 => x"33",
          1830 => x"e6",
          1831 => x"78",
          1832 => x"33",
          1833 => x"80",
          1834 => x"98",
          1835 => x"55",
          1836 => x"b6",
          1837 => x"80",
          1838 => x"08",
          1839 => x"84",
          1840 => x"84",
          1841 => x"55",
          1842 => x"05",
          1843 => x"08",
          1844 => x"84",
          1845 => x"3f",
          1846 => x"58",
          1847 => x"33",
          1848 => x"83",
          1849 => x"f4",
          1850 => x"74",
          1851 => x"fc",
          1852 => x"70",
          1853 => x"84",
          1854 => x"f4",
          1855 => x"05",
          1856 => x"52",
          1857 => x"f4",
          1858 => x"05",
          1859 => x"cf",
          1860 => x"80",
          1861 => x"58",
          1862 => x"0b",
          1863 => x"e2",
          1864 => x"b5",
          1865 => x"55",
          1866 => x"e8",
          1867 => x"3f",
          1868 => x"ff",
          1869 => x"52",
          1870 => x"e2",
          1871 => x"e2",
          1872 => x"74",
          1873 => x"9e",
          1874 => x"34",
          1875 => x"e4",
          1876 => x"ff",
          1877 => x"d4",
          1878 => x"5a",
          1879 => x"58",
          1880 => x"e8",
          1881 => x"3f",
          1882 => x"70",
          1883 => x"52",
          1884 => x"38",
          1885 => x"ff",
          1886 => x"70",
          1887 => x"c4",
          1888 => x"24",
          1889 => x"52",
          1890 => x"81",
          1891 => x"70",
          1892 => x"51",
          1893 => x"84",
          1894 => x"ac",
          1895 => x"81",
          1896 => x"e2",
          1897 => x"25",
          1898 => x"16",
          1899 => x"e6",
          1900 => x"ac",
          1901 => x"81",
          1902 => x"e2",
          1903 => x"25",
          1904 => x"17",
          1905 => x"52",
          1906 => x"75",
          1907 => x"05",
          1908 => x"44",
          1909 => x"38",
          1910 => x"0b",
          1911 => x"55",
          1912 => x"e8",
          1913 => x"3f",
          1914 => x"ff",
          1915 => x"52",
          1916 => x"e2",
          1917 => x"e2",
          1918 => x"74",
          1919 => x"9c",
          1920 => x"34",
          1921 => x"84",
          1922 => x"84",
          1923 => x"58",
          1924 => x"84",
          1925 => x"ae",
          1926 => x"57",
          1927 => x"16",
          1928 => x"81",
          1929 => x"70",
          1930 => x"57",
          1931 => x"18",
          1932 => x"81",
          1933 => x"33",
          1934 => x"76",
          1935 => x"75",
          1936 => x"e2",
          1937 => x"81",
          1938 => x"81",
          1939 => x"76",
          1940 => x"70",
          1941 => x"57",
          1942 => x"84",
          1943 => x"a9",
          1944 => x"81",
          1945 => x"e2",
          1946 => x"25",
          1947 => x"52",
          1948 => x"81",
          1949 => x"70",
          1950 => x"57",
          1951 => x"f0",
          1952 => x"c8",
          1953 => x"ec",
          1954 => x"e2",
          1955 => x"f4",
          1956 => x"75",
          1957 => x"38",
          1958 => x"52",
          1959 => x"a8",
          1960 => x"81",
          1961 => x"e2",
          1962 => x"24",
          1963 => x"98",
          1964 => x"06",
          1965 => x"ef",
          1966 => x"ec",
          1967 => x"f4",
          1968 => x"74",
          1969 => x"56",
          1970 => x"83",
          1971 => x"55",
          1972 => x"51",
          1973 => x"08",
          1974 => x"83",
          1975 => x"40",
          1976 => x"db",
          1977 => x"84",
          1978 => x"ac",
          1979 => x"aa",
          1980 => x"e2",
          1981 => x"ff",
          1982 => x"51",
          1983 => x"e2",
          1984 => x"57",
          1985 => x"84",
          1986 => x"a6",
          1987 => x"a0",
          1988 => x"e8",
          1989 => x"3f",
          1990 => x"78",
          1991 => x"06",
          1992 => x"e7",
          1993 => x"c4",
          1994 => x"06",
          1995 => x"ff",
          1996 => x"33",
          1997 => x"74",
          1998 => x"e8",
          1999 => x"3f",
          2000 => x"ff",
          2001 => x"52",
          2002 => x"e2",
          2003 => x"e2",
          2004 => x"c7",
          2005 => x"84",
          2006 => x"84",
          2007 => x"05",
          2008 => x"a9",
          2009 => x"84",
          2010 => x"58",
          2011 => x"f2",
          2012 => x"51",
          2013 => x"08",
          2014 => x"84",
          2015 => x"a4",
          2016 => x"05",
          2017 => x"81",
          2018 => x"34",
          2019 => x"0b",
          2020 => x"84",
          2021 => x"9c",
          2022 => x"38",
          2023 => x"bb",
          2024 => x"bb",
          2025 => x"53",
          2026 => x"3f",
          2027 => x"33",
          2028 => x"38",
          2029 => x"ff",
          2030 => x"52",
          2031 => x"e6",
          2032 => x"ed",
          2033 => x"59",
          2034 => x"ff",
          2035 => x"d7",
          2036 => x"82",
          2037 => x"05",
          2038 => x"80",
          2039 => x"79",
          2040 => x"10",
          2041 => x"43",
          2042 => x"b7",
          2043 => x"10",
          2044 => x"5e",
          2045 => x"75",
          2046 => x"f9",
          2047 => x"70",
          2048 => x"27",
          2049 => x"34",
          2050 => x"05",
          2051 => x"81",
          2052 => x"52",
          2053 => x"f4",
          2054 => x"80",
          2055 => x"84",
          2056 => x"0c",
          2057 => x"52",
          2058 => x"bb",
          2059 => x"84",
          2060 => x"ec",
          2061 => x"82",
          2062 => x"5a",
          2063 => x"81",
          2064 => x"08",
          2065 => x"84",
          2066 => x"08",
          2067 => x"08",
          2068 => x"76",
          2069 => x"f4",
          2070 => x"05",
          2071 => x"81",
          2072 => x"06",
          2073 => x"53",
          2074 => x"bb",
          2075 => x"33",
          2076 => x"70",
          2077 => x"59",
          2078 => x"33",
          2079 => x"70",
          2080 => x"81",
          2081 => x"93",
          2082 => x"ff",
          2083 => x"77",
          2084 => x"53",
          2085 => x"3f",
          2086 => x"81",
          2087 => x"80",
          2088 => x"34",
          2089 => x"90",
          2090 => x"2b",
          2091 => x"81",
          2092 => x"d9",
          2093 => x"0c",
          2094 => x"83",
          2095 => x"83",
          2096 => x"3f",
          2097 => x"83",
          2098 => x"42",
          2099 => x"86",
          2100 => x"df",
          2101 => x"f1",
          2102 => x"c2",
          2103 => x"39",
          2104 => x"33",
          2105 => x"5b",
          2106 => x"72",
          2107 => x"25",
          2108 => x"a8",
          2109 => x"c7",
          2110 => x"9f",
          2111 => x"75",
          2112 => x"b5",
          2113 => x"fa",
          2114 => x"2b",
          2115 => x"7a",
          2116 => x"27",
          2117 => x"56",
          2118 => x"0c",
          2119 => x"27",
          2120 => x"99",
          2121 => x"55",
          2122 => x"74",
          2123 => x"53",
          2124 => x"86",
          2125 => x"33",
          2126 => x"33",
          2127 => x"41",
          2128 => x"0b",
          2129 => x"06",
          2130 => x"06",
          2131 => x"ff",
          2132 => x"58",
          2133 => x"87",
          2134 => x"79",
          2135 => x"7c",
          2136 => x"06",
          2137 => x"14",
          2138 => x"74",
          2139 => x"74",
          2140 => x"59",
          2141 => x"2e",
          2142 => x"72",
          2143 => x"70",
          2144 => x"33",
          2145 => x"39",
          2146 => x"b0",
          2147 => x"81",
          2148 => x"81",
          2149 => x"74",
          2150 => x"5e",
          2151 => x"73",
          2152 => x"71",
          2153 => x"80",
          2154 => x"fa",
          2155 => x"34",
          2156 => x"71",
          2157 => x"71",
          2158 => x"76",
          2159 => x"39",
          2160 => x"33",
          2161 => x"11",
          2162 => x"11",
          2163 => x"5b",
          2164 => x"70",
          2165 => x"ff",
          2166 => x"ff",
          2167 => x"ff",
          2168 => x"5e",
          2169 => x"57",
          2170 => x"31",
          2171 => x"7d",
          2172 => x"71",
          2173 => x"62",
          2174 => x"5f",
          2175 => x"85",
          2176 => x"31",
          2177 => x"fd",
          2178 => x"fd",
          2179 => x"31",
          2180 => x"3d",
          2181 => x"8a",
          2182 => x"34",
          2183 => x"55",
          2184 => x"34",
          2185 => x"34",
          2186 => x"54",
          2187 => x"80",
          2188 => x"d8",
          2189 => x"54",
          2190 => x"f8",
          2191 => x"72",
          2192 => x"06",
          2193 => x"34",
          2194 => x"06",
          2195 => x"81",
          2196 => x"88",
          2197 => x"0b",
          2198 => x"bb",
          2199 => x"b8",
          2200 => x"f7",
          2201 => x"84",
          2202 => x"33",
          2203 => x"26",
          2204 => x"83",
          2205 => x"72",
          2206 => x"11",
          2207 => x"59",
          2208 => x"ff",
          2209 => x"58",
          2210 => x"83",
          2211 => x"83",
          2212 => x"76",
          2213 => x"ff",
          2214 => x"82",
          2215 => x"fa",
          2216 => x"83",
          2217 => x"5c",
          2218 => x"38",
          2219 => x"54",
          2220 => x"ac",
          2221 => x"55",
          2222 => x"34",
          2223 => x"70",
          2224 => x"84",
          2225 => x"9f",
          2226 => x"33",
          2227 => x"0b",
          2228 => x"81",
          2229 => x"9f",
          2230 => x"33",
          2231 => x"23",
          2232 => x"83",
          2233 => x"26",
          2234 => x"05",
          2235 => x"58",
          2236 => x"80",
          2237 => x"ff",
          2238 => x"29",
          2239 => x"27",
          2240 => x"e0",
          2241 => x"13",
          2242 => x"73",
          2243 => x"81",
          2244 => x"f8",
          2245 => x"29",
          2246 => x"26",
          2247 => x"84",
          2248 => x"fa",
          2249 => x"83",
          2250 => x"5c",
          2251 => x"38",
          2252 => x"81",
          2253 => x"33",
          2254 => x"06",
          2255 => x"05",
          2256 => x"78",
          2257 => x"73",
          2258 => x"b0",
          2259 => x"31",
          2260 => x"16",
          2261 => x"34",
          2262 => x"8a",
          2263 => x"75",
          2264 => x"13",
          2265 => x"80",
          2266 => x"fe",
          2267 => x"59",
          2268 => x"84",
          2269 => x"fc",
          2270 => x"05",
          2271 => x"38",
          2272 => x"51",
          2273 => x"51",
          2274 => x"fa",
          2275 => x"0c",
          2276 => x"fa",
          2277 => x"81",
          2278 => x"e2",
          2279 => x"b4",
          2280 => x"86",
          2281 => x"70",
          2282 => x"72",
          2283 => x"fa",
          2284 => x"33",
          2285 => x"11",
          2286 => x"38",
          2287 => x"80",
          2288 => x"0d",
          2289 => x"31",
          2290 => x"54",
          2291 => x"34",
          2292 => x"3d",
          2293 => x"05",
          2294 => x"55",
          2295 => x"53",
          2296 => x"84",
          2297 => x"80",
          2298 => x"b4",
          2299 => x"56",
          2300 => x"81",
          2301 => x"fe",
          2302 => x"05",
          2303 => x"70",
          2304 => x"70",
          2305 => x"80",
          2306 => x"06",
          2307 => x"53",
          2308 => x"06",
          2309 => x"b0",
          2310 => x"83",
          2311 => x"81",
          2312 => x"fa",
          2313 => x"0c",
          2314 => x"33",
          2315 => x"b0",
          2316 => x"81",
          2317 => x"fa",
          2318 => x"83",
          2319 => x"84",
          2320 => x"b0",
          2321 => x"70",
          2322 => x"83",
          2323 => x"83",
          2324 => x"fa",
          2325 => x"51",
          2326 => x"39",
          2327 => x"83",
          2328 => x"ff",
          2329 => x"f9",
          2330 => x"b0",
          2331 => x"33",
          2332 => x"b0",
          2333 => x"33",
          2334 => x"70",
          2335 => x"83",
          2336 => x"07",
          2337 => x"ba",
          2338 => x"06",
          2339 => x"b0",
          2340 => x"33",
          2341 => x"70",
          2342 => x"83",
          2343 => x"07",
          2344 => x"82",
          2345 => x"06",
          2346 => x"f2",
          2347 => x"06",
          2348 => x"34",
          2349 => x"bf",
          2350 => x"05",
          2351 => x"b3",
          2352 => x"fa",
          2353 => x"78",
          2354 => x"24",
          2355 => x"38",
          2356 => x"84",
          2357 => x"34",
          2358 => x"fa",
          2359 => x"83",
          2360 => x"0b",
          2361 => x"b8",
          2362 => x"34",
          2363 => x"0b",
          2364 => x"b8",
          2365 => x"56",
          2366 => x"7c",
          2367 => x"ff",
          2368 => x"34",
          2369 => x"83",
          2370 => x"23",
          2371 => x"0d",
          2372 => x"81",
          2373 => x"83",
          2374 => x"b5",
          2375 => x"84",
          2376 => x"33",
          2377 => x"55",
          2378 => x"e5",
          2379 => x"0b",
          2380 => x"79",
          2381 => x"d8",
          2382 => x"ac",
          2383 => x"70",
          2384 => x"52",
          2385 => x"83",
          2386 => x"7d",
          2387 => x"b8",
          2388 => x"7b",
          2389 => x"b5",
          2390 => x"84",
          2391 => x"fc",
          2392 => x"a8",
          2393 => x"83",
          2394 => x"ff",
          2395 => x"52",
          2396 => x"3f",
          2397 => x"90",
          2398 => x"27",
          2399 => x"33",
          2400 => x"87",
          2401 => x"5a",
          2402 => x"02",
          2403 => x"f8",
          2404 => x"b4",
          2405 => x"a0",
          2406 => x"51",
          2407 => x"83",
          2408 => x"52",
          2409 => x"2e",
          2410 => x"f9",
          2411 => x"75",
          2412 => x"2e",
          2413 => x"83",
          2414 => x"72",
          2415 => x"b9",
          2416 => x"14",
          2417 => x"b5",
          2418 => x"29",
          2419 => x"fa",
          2420 => x"73",
          2421 => x"b0",
          2422 => x"84",
          2423 => x"83",
          2424 => x"72",
          2425 => x"57",
          2426 => x"14",
          2427 => x"59",
          2428 => x"84",
          2429 => x"38",
          2430 => x"34",
          2431 => x"2e",
          2432 => x"76",
          2433 => x"84",
          2434 => x"75",
          2435 => x"80",
          2436 => x"06",
          2437 => x"f1",
          2438 => x"34",
          2439 => x"33",
          2440 => x"34",
          2441 => x"89",
          2442 => x"fd",
          2443 => x"06",
          2444 => x"38",
          2445 => x"81",
          2446 => x"83",
          2447 => x"74",
          2448 => x"75",
          2449 => x"0b",
          2450 => x"04",
          2451 => x"fd",
          2452 => x"81",
          2453 => x"83",
          2454 => x"34",
          2455 => x"83",
          2456 => x"55",
          2457 => x"73",
          2458 => x"a0",
          2459 => x"81",
          2460 => x"90",
          2461 => x"3f",
          2462 => x"80",
          2463 => x"57",
          2464 => x"75",
          2465 => x"2e",
          2466 => x"d1",
          2467 => x"78",
          2468 => x"f8",
          2469 => x"b5",
          2470 => x"5c",
          2471 => x"a0",
          2472 => x"83",
          2473 => x"72",
          2474 => x"78",
          2475 => x"b4",
          2476 => x"5a",
          2477 => x"b0",
          2478 => x"70",
          2479 => x"83",
          2480 => x"42",
          2481 => x"33",
          2482 => x"70",
          2483 => x"26",
          2484 => x"5a",
          2485 => x"75",
          2486 => x"bb",
          2487 => x"b7",
          2488 => x"81",
          2489 => x"38",
          2490 => x"80",
          2491 => x"f8",
          2492 => x"b5",
          2493 => x"40",
          2494 => x"a0",
          2495 => x"83",
          2496 => x"72",
          2497 => x"78",
          2498 => x"b4",
          2499 => x"83",
          2500 => x"1b",
          2501 => x"ff",
          2502 => x"b5",
          2503 => x"43",
          2504 => x"84",
          2505 => x"77",
          2506 => x"fe",
          2507 => x"80",
          2508 => x"0d",
          2509 => x"78",
          2510 => x"2e",
          2511 => x"0b",
          2512 => x"bb",
          2513 => x"9b",
          2514 => x"75",
          2515 => x"84",
          2516 => x"ba",
          2517 => x"34",
          2518 => x"84",
          2519 => x"bb",
          2520 => x"9b",
          2521 => x"ba",
          2522 => x"fa",
          2523 => x"72",
          2524 => x"80",
          2525 => x"34",
          2526 => x"33",
          2527 => x"12",
          2528 => x"b6",
          2529 => x"71",
          2530 => x"33",
          2531 => x"b8",
          2532 => x"fa",
          2533 => x"72",
          2534 => x"83",
          2535 => x"05",
          2536 => x"81",
          2537 => x"0b",
          2538 => x"84",
          2539 => x"70",
          2540 => x"73",
          2541 => x"05",
          2542 => x"72",
          2543 => x"06",
          2544 => x"5a",
          2545 => x"78",
          2546 => x"76",
          2547 => x"fa",
          2548 => x"84",
          2549 => x"85",
          2550 => x"80",
          2551 => x"84",
          2552 => x"84",
          2553 => x"b4",
          2554 => x"b5",
          2555 => x"b3",
          2556 => x"84",
          2557 => x"84",
          2558 => x"ff",
          2559 => x"83",
          2560 => x"70",
          2561 => x"70",
          2562 => x"86",
          2563 => x"22",
          2564 => x"83",
          2565 => x"44",
          2566 => x"81",
          2567 => x"06",
          2568 => x"75",
          2569 => x"81",
          2570 => x"81",
          2571 => x"40",
          2572 => x"a0",
          2573 => x"83",
          2574 => x"72",
          2575 => x"a0",
          2576 => x"fa",
          2577 => x"5a",
          2578 => x"b0",
          2579 => x"70",
          2580 => x"83",
          2581 => x"43",
          2582 => x"33",
          2583 => x"1a",
          2584 => x"7b",
          2585 => x"33",
          2586 => x"58",
          2587 => x"b5",
          2588 => x"05",
          2589 => x"95",
          2590 => x"38",
          2591 => x"ba",
          2592 => x"ff",
          2593 => x"c8",
          2594 => x"05",
          2595 => x"fa",
          2596 => x"9f",
          2597 => x"9c",
          2598 => x"84",
          2599 => x"83",
          2600 => x"72",
          2601 => x"05",
          2602 => x"7b",
          2603 => x"83",
          2604 => x"59",
          2605 => x"38",
          2606 => x"81",
          2607 => x"72",
          2608 => x"a0",
          2609 => x"84",
          2610 => x"83",
          2611 => x"5e",
          2612 => x"b6",
          2613 => x"71",
          2614 => x"33",
          2615 => x"b8",
          2616 => x"fa",
          2617 => x"72",
          2618 => x"83",
          2619 => x"34",
          2620 => x"5b",
          2621 => x"84",
          2622 => x"38",
          2623 => x"34",
          2624 => x"59",
          2625 => x"fa",
          2626 => x"fa",
          2627 => x"81",
          2628 => x"72",
          2629 => x"5b",
          2630 => x"80",
          2631 => x"fa",
          2632 => x"71",
          2633 => x"0b",
          2634 => x"b4",
          2635 => x"83",
          2636 => x"1a",
          2637 => x"ff",
          2638 => x"b5",
          2639 => x"5a",
          2640 => x"99",
          2641 => x"81",
          2642 => x"fe",
          2643 => x"fe",
          2644 => x"0c",
          2645 => x"3d",
          2646 => x"59",
          2647 => x"83",
          2648 => x"58",
          2649 => x"0b",
          2650 => x"bb",
          2651 => x"fa",
          2652 => x"1b",
          2653 => x"84",
          2654 => x"5b",
          2655 => x"84",
          2656 => x"53",
          2657 => x"84",
          2658 => x"38",
          2659 => x"5a",
          2660 => x"83",
          2661 => x"22",
          2662 => x"cf",
          2663 => x"84",
          2664 => x"fa",
          2665 => x"fa",
          2666 => x"39",
          2667 => x"33",
          2668 => x"05",
          2669 => x"33",
          2670 => x"84",
          2671 => x"83",
          2672 => x"5a",
          2673 => x"18",
          2674 => x"29",
          2675 => x"60",
          2676 => x"b8",
          2677 => x"fa",
          2678 => x"72",
          2679 => x"83",
          2680 => x"34",
          2681 => x"58",
          2682 => x"b8",
          2683 => x"ff",
          2684 => x"80",
          2685 => x"fb",
          2686 => x"38",
          2687 => x"b4",
          2688 => x"3f",
          2689 => x"3d",
          2690 => x"fa",
          2691 => x"fa",
          2692 => x"76",
          2693 => x"83",
          2694 => x"83",
          2695 => x"83",
          2696 => x"ff",
          2697 => x"7a",
          2698 => x"d8",
          2699 => x"06",
          2700 => x"81",
          2701 => x"05",
          2702 => x"94",
          2703 => x"3f",
          2704 => x"bb",
          2705 => x"88",
          2706 => x"24",
          2707 => x"e8",
          2708 => x"39",
          2709 => x"58",
          2710 => x"27",
          2711 => x"d8",
          2712 => x"b1",
          2713 => x"83",
          2714 => x"84",
          2715 => x"8f",
          2716 => x"ba",
          2717 => x"70",
          2718 => x"5e",
          2719 => x"e7",
          2720 => x"80",
          2721 => x"33",
          2722 => x"b8",
          2723 => x"27",
          2724 => x"34",
          2725 => x"b5",
          2726 => x"ff",
          2727 => x"a7",
          2728 => x"b4",
          2729 => x"fa",
          2730 => x"b8",
          2731 => x"76",
          2732 => x"75",
          2733 => x"84",
          2734 => x"8d",
          2735 => x"ba",
          2736 => x"70",
          2737 => x"42",
          2738 => x"cf",
          2739 => x"80",
          2740 => x"22",
          2741 => x"fc",
          2742 => x"fa",
          2743 => x"71",
          2744 => x"83",
          2745 => x"71",
          2746 => x"06",
          2747 => x"80",
          2748 => x"82",
          2749 => x"83",
          2750 => x"ba",
          2751 => x"e7",
          2752 => x"99",
          2753 => x"81",
          2754 => x"39",
          2755 => x"2e",
          2756 => x"83",
          2757 => x"b8",
          2758 => x"75",
          2759 => x"83",
          2760 => x"ba",
          2761 => x"c8",
          2762 => x"b4",
          2763 => x"33",
          2764 => x"25",
          2765 => x"b4",
          2766 => x"51",
          2767 => x"ba",
          2768 => x"8b",
          2769 => x"05",
          2770 => x"51",
          2771 => x"81",
          2772 => x"58",
          2773 => x"85",
          2774 => x"38",
          2775 => x"26",
          2776 => x"81",
          2777 => x"97",
          2778 => x"77",
          2779 => x"33",
          2780 => x"ba",
          2781 => x"06",
          2782 => x"06",
          2783 => x"5c",
          2784 => x"5a",
          2785 => x"ff",
          2786 => x"27",
          2787 => x"b4",
          2788 => x"57",
          2789 => x"7a",
          2790 => x"af",
          2791 => x"80",
          2792 => x"33",
          2793 => x"7f",
          2794 => x"33",
          2795 => x"06",
          2796 => x"11",
          2797 => x"b2",
          2798 => x"70",
          2799 => x"33",
          2800 => x"81",
          2801 => x"ff",
          2802 => x"7c",
          2803 => x"33",
          2804 => x"ff",
          2805 => x"7c",
          2806 => x"57",
          2807 => x"b8",
          2808 => x"ee",
          2809 => x"b4",
          2810 => x"b2",
          2811 => x"26",
          2812 => x"7e",
          2813 => x"5e",
          2814 => x"5b",
          2815 => x"06",
          2816 => x"1d",
          2817 => x"f7",
          2818 => x"e0",
          2819 => x"1f",
          2820 => x"76",
          2821 => x"81",
          2822 => x"f8",
          2823 => x"29",
          2824 => x"27",
          2825 => x"5f",
          2826 => x"81",
          2827 => x"58",
          2828 => x"81",
          2829 => x"f7",
          2830 => x"5e",
          2831 => x"f6",
          2832 => x"75",
          2833 => x"84",
          2834 => x"f6",
          2835 => x"33",
          2836 => x"59",
          2837 => x"84",
          2838 => x"09",
          2839 => x"b5",
          2840 => x"fa",
          2841 => x"ff",
          2842 => x"33",
          2843 => x"7e",
          2844 => x"f5",
          2845 => x"27",
          2846 => x"10",
          2847 => x"86",
          2848 => x"5a",
          2849 => x"06",
          2850 => x"79",
          2851 => x"83",
          2852 => x"90",
          2853 => x"07",
          2854 => x"7a",
          2855 => x"05",
          2856 => x"58",
          2857 => x"b8",
          2858 => x"5f",
          2859 => x"06",
          2860 => x"64",
          2861 => x"26",
          2862 => x"7b",
          2863 => x"1d",
          2864 => x"38",
          2865 => x"18",
          2866 => x"34",
          2867 => x"81",
          2868 => x"38",
          2869 => x"78",
          2870 => x"57",
          2871 => x"39",
          2872 => x"58",
          2873 => x"70",
          2874 => x"f0",
          2875 => x"57",
          2876 => x"be",
          2877 => x"34",
          2878 => x"56",
          2879 => x"33",
          2880 => x"34",
          2881 => x"33",
          2882 => x"33",
          2883 => x"83",
          2884 => x"83",
          2885 => x"ff",
          2886 => x"fa",
          2887 => x"56",
          2888 => x"83",
          2889 => x"07",
          2890 => x"39",
          2891 => x"81",
          2892 => x"c3",
          2893 => x"06",
          2894 => x"34",
          2895 => x"fa",
          2896 => x"06",
          2897 => x"b0",
          2898 => x"fa",
          2899 => x"b0",
          2900 => x"75",
          2901 => x"83",
          2902 => x"e0",
          2903 => x"fe",
          2904 => x"cf",
          2905 => x"fa",
          2906 => x"b0",
          2907 => x"75",
          2908 => x"83",
          2909 => x"07",
          2910 => x"b3",
          2911 => x"06",
          2912 => x"34",
          2913 => x"81",
          2914 => x"fa",
          2915 => x"b0",
          2916 => x"fa",
          2917 => x"b0",
          2918 => x"fa",
          2919 => x"b0",
          2920 => x"fa",
          2921 => x"b0",
          2922 => x"56",
          2923 => x"39",
          2924 => x"b0",
          2925 => x"fd",
          2926 => x"34",
          2927 => x"ec",
          2928 => x"fa",
          2929 => x"fa",
          2930 => x"78",
          2931 => x"ba",
          2932 => x"84",
          2933 => x"84",
          2934 => x"fa",
          2935 => x"81",
          2936 => x"cf",
          2937 => x"dc",
          2938 => x"b5",
          2939 => x"84",
          2940 => x"80",
          2941 => x"84",
          2942 => x"77",
          2943 => x"84",
          2944 => x"7a",
          2945 => x"fe",
          2946 => x"84",
          2947 => x"ba",
          2948 => x"fa",
          2949 => x"97",
          2950 => x"ff",
          2951 => x"39",
          2952 => x"52",
          2953 => x"39",
          2954 => x"8f",
          2955 => x"70",
          2956 => x"5f",
          2957 => x"51",
          2958 => x"75",
          2959 => x"fa",
          2960 => x"b4",
          2961 => x"2c",
          2962 => x"39",
          2963 => x"b8",
          2964 => x"75",
          2965 => x"f3",
          2966 => x"81",
          2967 => x"ee",
          2968 => x"b8",
          2969 => x"fa",
          2970 => x"c7",
          2971 => x"5f",
          2972 => x"ff",
          2973 => x"5b",
          2974 => x"81",
          2975 => x"ff",
          2976 => x"89",
          2977 => x"76",
          2978 => x"75",
          2979 => x"06",
          2980 => x"83",
          2981 => x"76",
          2982 => x"56",
          2983 => x"ff",
          2984 => x"80",
          2985 => x"77",
          2986 => x"71",
          2987 => x"86",
          2988 => x"80",
          2989 => x"06",
          2990 => x"5d",
          2991 => x"99",
          2992 => x"5e",
          2993 => x"81",
          2994 => x"58",
          2995 => x"81",
          2996 => x"f7",
          2997 => x"5d",
          2998 => x"e0",
          2999 => x"1e",
          3000 => x"76",
          3001 => x"81",
          3002 => x"f8",
          3003 => x"29",
          3004 => x"26",
          3005 => x"fa",
          3006 => x"1c",
          3007 => x"84",
          3008 => x"84",
          3009 => x"fd",
          3010 => x"b8",
          3011 => x"11",
          3012 => x"38",
          3013 => x"77",
          3014 => x"80",
          3015 => x"83",
          3016 => x"70",
          3017 => x"56",
          3018 => x"56",
          3019 => x"39",
          3020 => x"b8",
          3021 => x"75",
          3022 => x"ef",
          3023 => x"06",
          3024 => x"70",
          3025 => x"7a",
          3026 => x"09",
          3027 => x"39",
          3028 => x"34",
          3029 => x"83",
          3030 => x"7b",
          3031 => x"f2",
          3032 => x"7a",
          3033 => x"81",
          3034 => x"77",
          3035 => x"26",
          3036 => x"05",
          3037 => x"70",
          3038 => x"d4",
          3039 => x"56",
          3040 => x"39",
          3041 => x"ad",
          3042 => x"84",
          3043 => x"f1",
          3044 => x"34",
          3045 => x"33",
          3046 => x"34",
          3047 => x"a7",
          3048 => x"33",
          3049 => x"80",
          3050 => x"3f",
          3051 => x"3d",
          3052 => x"ab",
          3053 => x"85",
          3054 => x"bf",
          3055 => x"88",
          3056 => x"e8",
          3057 => x"80",
          3058 => x"75",
          3059 => x"84",
          3060 => x"83",
          3061 => x"80",
          3062 => x"30",
          3063 => x"56",
          3064 => x"0c",
          3065 => x"09",
          3066 => x"83",
          3067 => x"07",
          3068 => x"c4",
          3069 => x"b5",
          3070 => x"29",
          3071 => x"fa",
          3072 => x"29",
          3073 => x"f9",
          3074 => x"81",
          3075 => x"73",
          3076 => x"87",
          3077 => x"88",
          3078 => x"87",
          3079 => x"f6",
          3080 => x"ff",
          3081 => x"cf",
          3082 => x"33",
          3083 => x"16",
          3084 => x"85",
          3085 => x"b4",
          3086 => x"75",
          3087 => x"2e",
          3088 => x"15",
          3089 => x"f8",
          3090 => x"ff",
          3091 => x"b3",
          3092 => x"2b",
          3093 => x"83",
          3094 => x"70",
          3095 => x"51",
          3096 => x"38",
          3097 => x"09",
          3098 => x"e4",
          3099 => x"80",
          3100 => x"e4",
          3101 => x"f8",
          3102 => x"5d",
          3103 => x"b8",
          3104 => x"8d",
          3105 => x"73",
          3106 => x"c2",
          3107 => x"8b",
          3108 => x"73",
          3109 => x"54",
          3110 => x"f8",
          3111 => x"81",
          3112 => x"72",
          3113 => x"f8",
          3114 => x"84",
          3115 => x"e8",
          3116 => x"54",
          3117 => x"0b",
          3118 => x"d8",
          3119 => x"06",
          3120 => x"38",
          3121 => x"f8",
          3122 => x"9c",
          3123 => x"83",
          3124 => x"83",
          3125 => x"91",
          3126 => x"9c",
          3127 => x"dc",
          3128 => x"54",
          3129 => x"54",
          3130 => x"98",
          3131 => x"81",
          3132 => x"38",
          3133 => x"b9",
          3134 => x"54",
          3135 => x"53",
          3136 => x"81",
          3137 => x"34",
          3138 => x"58",
          3139 => x"83",
          3140 => x"77",
          3141 => x"7d",
          3142 => x"2e",
          3143 => x"59",
          3144 => x"54",
          3145 => x"2e",
          3146 => x"06",
          3147 => x"27",
          3148 => x"54",
          3149 => x"10",
          3150 => x"2b",
          3151 => x"33",
          3152 => x"9c",
          3153 => x"ea",
          3154 => x"a8",
          3155 => x"a0",
          3156 => x"ff",
          3157 => x"b8",
          3158 => x"83",
          3159 => x"70",
          3160 => x"7d",
          3161 => x"06",
          3162 => x"c6",
          3163 => x"83",
          3164 => x"78",
          3165 => x"70",
          3166 => x"27",
          3167 => x"72",
          3168 => x"fc",
          3169 => x"81",
          3170 => x"3f",
          3171 => x"0d",
          3172 => x"f9",
          3173 => x"38",
          3174 => x"5b",
          3175 => x"c9",
          3176 => x"34",
          3177 => x"ff",
          3178 => x"b1",
          3179 => x"81",
          3180 => x"cc",
          3181 => x"8a",
          3182 => x"81",
          3183 => x"83",
          3184 => x"c0",
          3185 => x"27",
          3186 => x"08",
          3187 => x"06",
          3188 => x"f8",
          3189 => x"83",
          3190 => x"53",
          3191 => x"de",
          3192 => x"83",
          3193 => x"70",
          3194 => x"33",
          3195 => x"fa",
          3196 => x"06",
          3197 => x"2e",
          3198 => x"81",
          3199 => x"ef",
          3200 => x"39",
          3201 => x"54",
          3202 => x"b8",
          3203 => x"80",
          3204 => x"76",
          3205 => x"fa",
          3206 => x"53",
          3207 => x"83",
          3208 => x"f6",
          3209 => x"81",
          3210 => x"80",
          3211 => x"83",
          3212 => x"ff",
          3213 => x"38",
          3214 => x"84",
          3215 => x"56",
          3216 => x"38",
          3217 => x"ff",
          3218 => x"51",
          3219 => x"aa",
          3220 => x"14",
          3221 => x"dd",
          3222 => x"34",
          3223 => x"39",
          3224 => x"3f",
          3225 => x"80",
          3226 => x"02",
          3227 => x"f5",
          3228 => x"85",
          3229 => x"fe",
          3230 => x"90",
          3231 => x"08",
          3232 => x"90",
          3233 => x"52",
          3234 => x"72",
          3235 => x"c0",
          3236 => x"27",
          3237 => x"38",
          3238 => x"55",
          3239 => x"55",
          3240 => x"c0",
          3241 => x"53",
          3242 => x"c0",
          3243 => x"f6",
          3244 => x"9c",
          3245 => x"38",
          3246 => x"c0",
          3247 => x"83",
          3248 => x"70",
          3249 => x"2e",
          3250 => x"71",
          3251 => x"38",
          3252 => x"0d",
          3253 => x"88",
          3254 => x"02",
          3255 => x"80",
          3256 => x"2b",
          3257 => x"98",
          3258 => x"83",
          3259 => x"84",
          3260 => x"85",
          3261 => x"f5",
          3262 => x"83",
          3263 => x"34",
          3264 => x"56",
          3265 => x"87",
          3266 => x"9c",
          3267 => x"ce",
          3268 => x"08",
          3269 => x"70",
          3270 => x"87",
          3271 => x"73",
          3272 => x"db",
          3273 => x"ff",
          3274 => x"71",
          3275 => x"87",
          3276 => x"05",
          3277 => x"87",
          3278 => x"2e",
          3279 => x"98",
          3280 => x"87",
          3281 => x"87",
          3282 => x"26",
          3283 => x"16",
          3284 => x"80",
          3285 => x"06",
          3286 => x"70",
          3287 => x"80",
          3288 => x"52",
          3289 => x"70",
          3290 => x"05",
          3291 => x"76",
          3292 => x"04",
          3293 => x"3d",
          3294 => x"3d",
          3295 => x"33",
          3296 => x"08",
          3297 => x"06",
          3298 => x"55",
          3299 => x"2a",
          3300 => x"2a",
          3301 => x"15",
          3302 => x"c6",
          3303 => x"51",
          3304 => x"81",
          3305 => x"54",
          3306 => x"f5",
          3307 => x"83",
          3308 => x"34",
          3309 => x"56",
          3310 => x"87",
          3311 => x"9c",
          3312 => x"ce",
          3313 => x"08",
          3314 => x"70",
          3315 => x"87",
          3316 => x"73",
          3317 => x"db",
          3318 => x"ff",
          3319 => x"71",
          3320 => x"87",
          3321 => x"05",
          3322 => x"87",
          3323 => x"2e",
          3324 => x"98",
          3325 => x"87",
          3326 => x"87",
          3327 => x"26",
          3328 => x"16",
          3329 => x"80",
          3330 => x"52",
          3331 => x"81",
          3332 => x"38",
          3333 => x"88",
          3334 => x"fb",
          3335 => x"80",
          3336 => x"90",
          3337 => x"34",
          3338 => x"87",
          3339 => x"08",
          3340 => x"c0",
          3341 => x"9c",
          3342 => x"81",
          3343 => x"52",
          3344 => x"81",
          3345 => x"a4",
          3346 => x"80",
          3347 => x"80",
          3348 => x"80",
          3349 => x"9c",
          3350 => x"51",
          3351 => x"33",
          3352 => x"73",
          3353 => x"2e",
          3354 => x"51",
          3355 => x"71",
          3356 => x"57",
          3357 => x"81",
          3358 => x"ff",
          3359 => x"51",
          3360 => x"04",
          3361 => x"7a",
          3362 => x"ff",
          3363 => x"33",
          3364 => x"83",
          3365 => x"12",
          3366 => x"07",
          3367 => x"59",
          3368 => x"81",
          3369 => x"83",
          3370 => x"2b",
          3371 => x"33",
          3372 => x"57",
          3373 => x"71",
          3374 => x"85",
          3375 => x"2b",
          3376 => x"54",
          3377 => x"81",
          3378 => x"84",
          3379 => x"33",
          3380 => x"70",
          3381 => x"77",
          3382 => x"84",
          3383 => x"86",
          3384 => x"84",
          3385 => x"34",
          3386 => x"08",
          3387 => x"88",
          3388 => x"88",
          3389 => x"34",
          3390 => x"04",
          3391 => x"8b",
          3392 => x"84",
          3393 => x"2b",
          3394 => x"51",
          3395 => x"72",
          3396 => x"70",
          3397 => x"71",
          3398 => x"5a",
          3399 => x"87",
          3400 => x"88",
          3401 => x"13",
          3402 => x"f4",
          3403 => x"71",
          3404 => x"70",
          3405 => x"72",
          3406 => x"f4",
          3407 => x"33",
          3408 => x"74",
          3409 => x"88",
          3410 => x"f8",
          3411 => x"52",
          3412 => x"77",
          3413 => x"84",
          3414 => x"81",
          3415 => x"2b",
          3416 => x"33",
          3417 => x"06",
          3418 => x"5a",
          3419 => x"81",
          3420 => x"17",
          3421 => x"8b",
          3422 => x"70",
          3423 => x"71",
          3424 => x"5a",
          3425 => x"e4",
          3426 => x"88",
          3427 => x"88",
          3428 => x"77",
          3429 => x"70",
          3430 => x"8b",
          3431 => x"82",
          3432 => x"2b",
          3433 => x"52",
          3434 => x"34",
          3435 => x"04",
          3436 => x"08",
          3437 => x"77",
          3438 => x"90",
          3439 => x"f4",
          3440 => x"0b",
          3441 => x"53",
          3442 => x"d1",
          3443 => x"76",
          3444 => x"84",
          3445 => x"34",
          3446 => x"f4",
          3447 => x"0b",
          3448 => x"84",
          3449 => x"80",
          3450 => x"88",
          3451 => x"17",
          3452 => x"f0",
          3453 => x"f4",
          3454 => x"82",
          3455 => x"fe",
          3456 => x"80",
          3457 => x"38",
          3458 => x"83",
          3459 => x"ff",
          3460 => x"11",
          3461 => x"07",
          3462 => x"ff",
          3463 => x"38",
          3464 => x"81",
          3465 => x"81",
          3466 => x"ff",
          3467 => x"5c",
          3468 => x"38",
          3469 => x"55",
          3470 => x"71",
          3471 => x"38",
          3472 => x"77",
          3473 => x"78",
          3474 => x"88",
          3475 => x"56",
          3476 => x"2e",
          3477 => x"73",
          3478 => x"80",
          3479 => x"82",
          3480 => x"78",
          3481 => x"88",
          3482 => x"74",
          3483 => x"f4",
          3484 => x"71",
          3485 => x"84",
          3486 => x"81",
          3487 => x"83",
          3488 => x"7e",
          3489 => x"5c",
          3490 => x"82",
          3491 => x"72",
          3492 => x"18",
          3493 => x"34",
          3494 => x"11",
          3495 => x"71",
          3496 => x"5c",
          3497 => x"85",
          3498 => x"16",
          3499 => x"12",
          3500 => x"2a",
          3501 => x"34",
          3502 => x"08",
          3503 => x"33",
          3504 => x"74",
          3505 => x"86",
          3506 => x"ba",
          3507 => x"84",
          3508 => x"2b",
          3509 => x"59",
          3510 => x"34",
          3511 => x"51",
          3512 => x"0d",
          3513 => x"71",
          3514 => x"05",
          3515 => x"88",
          3516 => x"59",
          3517 => x"76",
          3518 => x"70",
          3519 => x"71",
          3520 => x"05",
          3521 => x"88",
          3522 => x"5f",
          3523 => x"1a",
          3524 => x"f4",
          3525 => x"71",
          3526 => x"70",
          3527 => x"77",
          3528 => x"f4",
          3529 => x"39",
          3530 => x"08",
          3531 => x"77",
          3532 => x"84",
          3533 => x"fb",
          3534 => x"bb",
          3535 => x"ff",
          3536 => x"80",
          3537 => x"80",
          3538 => x"fe",
          3539 => x"55",
          3540 => x"34",
          3541 => x"15",
          3542 => x"ba",
          3543 => x"81",
          3544 => x"08",
          3545 => x"80",
          3546 => x"70",
          3547 => x"88",
          3548 => x"ba",
          3549 => x"ba",
          3550 => x"76",
          3551 => x"34",
          3552 => x"38",
          3553 => x"67",
          3554 => x"08",
          3555 => x"aa",
          3556 => x"7f",
          3557 => x"84",
          3558 => x"83",
          3559 => x"06",
          3560 => x"7f",
          3561 => x"ff",
          3562 => x"33",
          3563 => x"70",
          3564 => x"70",
          3565 => x"2b",
          3566 => x"71",
          3567 => x"90",
          3568 => x"54",
          3569 => x"5f",
          3570 => x"82",
          3571 => x"2b",
          3572 => x"33",
          3573 => x"90",
          3574 => x"56",
          3575 => x"62",
          3576 => x"77",
          3577 => x"2e",
          3578 => x"62",
          3579 => x"61",
          3580 => x"70",
          3581 => x"71",
          3582 => x"81",
          3583 => x"2b",
          3584 => x"5b",
          3585 => x"76",
          3586 => x"71",
          3587 => x"11",
          3588 => x"8b",
          3589 => x"84",
          3590 => x"2b",
          3591 => x"52",
          3592 => x"77",
          3593 => x"84",
          3594 => x"33",
          3595 => x"83",
          3596 => x"87",
          3597 => x"88",
          3598 => x"41",
          3599 => x"16",
          3600 => x"33",
          3601 => x"81",
          3602 => x"5c",
          3603 => x"1a",
          3604 => x"82",
          3605 => x"2b",
          3606 => x"33",
          3607 => x"70",
          3608 => x"5a",
          3609 => x"1a",
          3610 => x"70",
          3611 => x"71",
          3612 => x"33",
          3613 => x"70",
          3614 => x"5a",
          3615 => x"83",
          3616 => x"1f",
          3617 => x"88",
          3618 => x"83",
          3619 => x"84",
          3620 => x"ba",
          3621 => x"05",
          3622 => x"44",
          3623 => x"7e",
          3624 => x"3d",
          3625 => x"ba",
          3626 => x"f0",
          3627 => x"84",
          3628 => x"84",
          3629 => x"81",
          3630 => x"08",
          3631 => x"85",
          3632 => x"60",
          3633 => x"34",
          3634 => x"22",
          3635 => x"83",
          3636 => x"5a",
          3637 => x"89",
          3638 => x"10",
          3639 => x"f8",
          3640 => x"81",
          3641 => x"08",
          3642 => x"2e",
          3643 => x"2e",
          3644 => x"3f",
          3645 => x"0c",
          3646 => x"ba",
          3647 => x"5e",
          3648 => x"33",
          3649 => x"06",
          3650 => x"40",
          3651 => x"61",
          3652 => x"2a",
          3653 => x"83",
          3654 => x"1f",
          3655 => x"2b",
          3656 => x"06",
          3657 => x"70",
          3658 => x"5b",
          3659 => x"81",
          3660 => x"34",
          3661 => x"7b",
          3662 => x"ba",
          3663 => x"88",
          3664 => x"75",
          3665 => x"54",
          3666 => x"06",
          3667 => x"82",
          3668 => x"2b",
          3669 => x"33",
          3670 => x"90",
          3671 => x"58",
          3672 => x"38",
          3673 => x"83",
          3674 => x"77",
          3675 => x"27",
          3676 => x"ff",
          3677 => x"80",
          3678 => x"80",
          3679 => x"fe",
          3680 => x"5a",
          3681 => x"34",
          3682 => x"1a",
          3683 => x"ba",
          3684 => x"81",
          3685 => x"08",
          3686 => x"80",
          3687 => x"70",
          3688 => x"64",
          3689 => x"34",
          3690 => x"10",
          3691 => x"42",
          3692 => x"61",
          3693 => x"7a",
          3694 => x"ff",
          3695 => x"38",
          3696 => x"bd",
          3697 => x"54",
          3698 => x"0d",
          3699 => x"12",
          3700 => x"07",
          3701 => x"33",
          3702 => x"7e",
          3703 => x"71",
          3704 => x"44",
          3705 => x"45",
          3706 => x"64",
          3707 => x"70",
          3708 => x"71",
          3709 => x"05",
          3710 => x"88",
          3711 => x"42",
          3712 => x"86",
          3713 => x"84",
          3714 => x"12",
          3715 => x"ff",
          3716 => x"5d",
          3717 => x"84",
          3718 => x"33",
          3719 => x"83",
          3720 => x"15",
          3721 => x"2a",
          3722 => x"54",
          3723 => x"84",
          3724 => x"81",
          3725 => x"2b",
          3726 => x"15",
          3727 => x"2a",
          3728 => x"55",
          3729 => x"34",
          3730 => x"11",
          3731 => x"07",
          3732 => x"42",
          3733 => x"51",
          3734 => x"08",
          3735 => x"06",
          3736 => x"f4",
          3737 => x"0b",
          3738 => x"53",
          3739 => x"bf",
          3740 => x"7f",
          3741 => x"84",
          3742 => x"34",
          3743 => x"f4",
          3744 => x"0b",
          3745 => x"84",
          3746 => x"80",
          3747 => x"88",
          3748 => x"1f",
          3749 => x"f0",
          3750 => x"f4",
          3751 => x"82",
          3752 => x"7e",
          3753 => x"c0",
          3754 => x"71",
          3755 => x"05",
          3756 => x"88",
          3757 => x"5e",
          3758 => x"34",
          3759 => x"f4",
          3760 => x"12",
          3761 => x"07",
          3762 => x"33",
          3763 => x"41",
          3764 => x"79",
          3765 => x"05",
          3766 => x"33",
          3767 => x"81",
          3768 => x"42",
          3769 => x"19",
          3770 => x"70",
          3771 => x"71",
          3772 => x"81",
          3773 => x"83",
          3774 => x"63",
          3775 => x"40",
          3776 => x"7b",
          3777 => x"70",
          3778 => x"8b",
          3779 => x"70",
          3780 => x"07",
          3781 => x"48",
          3782 => x"60",
          3783 => x"61",
          3784 => x"39",
          3785 => x"8b",
          3786 => x"84",
          3787 => x"2b",
          3788 => x"52",
          3789 => x"85",
          3790 => x"19",
          3791 => x"8b",
          3792 => x"86",
          3793 => x"2b",
          3794 => x"52",
          3795 => x"05",
          3796 => x"ba",
          3797 => x"33",
          3798 => x"06",
          3799 => x"77",
          3800 => x"ba",
          3801 => x"12",
          3802 => x"07",
          3803 => x"71",
          3804 => x"ff",
          3805 => x"56",
          3806 => x"55",
          3807 => x"34",
          3808 => x"33",
          3809 => x"83",
          3810 => x"12",
          3811 => x"ff",
          3812 => x"58",
          3813 => x"76",
          3814 => x"70",
          3815 => x"71",
          3816 => x"11",
          3817 => x"8b",
          3818 => x"84",
          3819 => x"2b",
          3820 => x"52",
          3821 => x"57",
          3822 => x"34",
          3823 => x"11",
          3824 => x"71",
          3825 => x"33",
          3826 => x"70",
          3827 => x"57",
          3828 => x"87",
          3829 => x"70",
          3830 => x"07",
          3831 => x"5a",
          3832 => x"81",
          3833 => x"1f",
          3834 => x"8b",
          3835 => x"73",
          3836 => x"07",
          3837 => x"5f",
          3838 => x"81",
          3839 => x"1f",
          3840 => x"2b",
          3841 => x"14",
          3842 => x"07",
          3843 => x"5f",
          3844 => x"75",
          3845 => x"70",
          3846 => x"71",
          3847 => x"70",
          3848 => x"05",
          3849 => x"84",
          3850 => x"65",
          3851 => x"5d",
          3852 => x"33",
          3853 => x"83",
          3854 => x"85",
          3855 => x"88",
          3856 => x"7a",
          3857 => x"05",
          3858 => x"84",
          3859 => x"2b",
          3860 => x"14",
          3861 => x"07",
          3862 => x"5c",
          3863 => x"34",
          3864 => x"f4",
          3865 => x"71",
          3866 => x"70",
          3867 => x"75",
          3868 => x"f4",
          3869 => x"33",
          3870 => x"74",
          3871 => x"88",
          3872 => x"f8",
          3873 => x"44",
          3874 => x"74",
          3875 => x"84",
          3876 => x"81",
          3877 => x"2b",
          3878 => x"33",
          3879 => x"06",
          3880 => x"46",
          3881 => x"81",
          3882 => x"5b",
          3883 => x"e5",
          3884 => x"84",
          3885 => x"62",
          3886 => x"51",
          3887 => x"88",
          3888 => x"b7",
          3889 => x"7a",
          3890 => x"58",
          3891 => x"77",
          3892 => x"89",
          3893 => x"3f",
          3894 => x"84",
          3895 => x"80",
          3896 => x"b5",
          3897 => x"89",
          3898 => x"84",
          3899 => x"ba",
          3900 => x"52",
          3901 => x"3f",
          3902 => x"34",
          3903 => x"f4",
          3904 => x"0b",
          3905 => x"56",
          3906 => x"17",
          3907 => x"f0",
          3908 => x"70",
          3909 => x"58",
          3910 => x"73",
          3911 => x"70",
          3912 => x"05",
          3913 => x"34",
          3914 => x"77",
          3915 => x"39",
          3916 => x"51",
          3917 => x"84",
          3918 => x"bb",
          3919 => x"3d",
          3920 => x"53",
          3921 => x"d4",
          3922 => x"ff",
          3923 => x"bb",
          3924 => x"33",
          3925 => x"3d",
          3926 => x"60",
          3927 => x"5c",
          3928 => x"87",
          3929 => x"73",
          3930 => x"38",
          3931 => x"8c",
          3932 => x"d5",
          3933 => x"ff",
          3934 => x"87",
          3935 => x"38",
          3936 => x"80",
          3937 => x"38",
          3938 => x"84",
          3939 => x"16",
          3940 => x"55",
          3941 => x"d5",
          3942 => x"02",
          3943 => x"57",
          3944 => x"38",
          3945 => x"81",
          3946 => x"73",
          3947 => x"0c",
          3948 => x"8e",
          3949 => x"06",
          3950 => x"c0",
          3951 => x"79",
          3952 => x"80",
          3953 => x"81",
          3954 => x"0c",
          3955 => x"81",
          3956 => x"56",
          3957 => x"39",
          3958 => x"9b",
          3959 => x"33",
          3960 => x"26",
          3961 => x"53",
          3962 => x"9b",
          3963 => x"0c",
          3964 => x"72",
          3965 => x"9a",
          3966 => x"0c",
          3967 => x"75",
          3968 => x"3d",
          3969 => x"0b",
          3970 => x"04",
          3971 => x"11",
          3972 => x"70",
          3973 => x"80",
          3974 => x"08",
          3975 => x"8c",
          3976 => x"0c",
          3977 => x"08",
          3978 => x"9b",
          3979 => x"ee",
          3980 => x"7c",
          3981 => x"5b",
          3982 => x"06",
          3983 => x"2e",
          3984 => x"81",
          3985 => x"bb",
          3986 => x"59",
          3987 => x"0d",
          3988 => x"b8",
          3989 => x"5a",
          3990 => x"84",
          3991 => x"38",
          3992 => x"b4",
          3993 => x"a0",
          3994 => x"58",
          3995 => x"38",
          3996 => x"09",
          3997 => x"75",
          3998 => x"51",
          3999 => x"59",
          4000 => x"fb",
          4001 => x"2e",
          4002 => x"18",
          4003 => x"75",
          4004 => x"57",
          4005 => x"b6",
          4006 => x"19",
          4007 => x"0b",
          4008 => x"19",
          4009 => x"80",
          4010 => x"f2",
          4011 => x"0b",
          4012 => x"84",
          4013 => x"74",
          4014 => x"5b",
          4015 => x"2a",
          4016 => x"98",
          4017 => x"90",
          4018 => x"34",
          4019 => x"19",
          4020 => x"a6",
          4021 => x"84",
          4022 => x"05",
          4023 => x"7a",
          4024 => x"fa",
          4025 => x"53",
          4026 => x"d8",
          4027 => x"fd",
          4028 => x"0d",
          4029 => x"81",
          4030 => x"76",
          4031 => x"bb",
          4032 => x"77",
          4033 => x"cc",
          4034 => x"74",
          4035 => x"75",
          4036 => x"19",
          4037 => x"17",
          4038 => x"33",
          4039 => x"83",
          4040 => x"17",
          4041 => x"3f",
          4042 => x"38",
          4043 => x"0c",
          4044 => x"06",
          4045 => x"89",
          4046 => x"5d",
          4047 => x"38",
          4048 => x"56",
          4049 => x"84",
          4050 => x"17",
          4051 => x"3f",
          4052 => x"38",
          4053 => x"0c",
          4054 => x"06",
          4055 => x"7e",
          4056 => x"53",
          4057 => x"38",
          4058 => x"0c",
          4059 => x"a8",
          4060 => x"79",
          4061 => x"33",
          4062 => x"09",
          4063 => x"78",
          4064 => x"51",
          4065 => x"80",
          4066 => x"78",
          4067 => x"75",
          4068 => x"05",
          4069 => x"2b",
          4070 => x"8f",
          4071 => x"81",
          4072 => x"a8",
          4073 => x"79",
          4074 => x"33",
          4075 => x"09",
          4076 => x"78",
          4077 => x"51",
          4078 => x"80",
          4079 => x"78",
          4080 => x"75",
          4081 => x"b8",
          4082 => x"71",
          4083 => x"14",
          4084 => x"33",
          4085 => x"07",
          4086 => x"59",
          4087 => x"54",
          4088 => x"53",
          4089 => x"3f",
          4090 => x"2e",
          4091 => x"bb",
          4092 => x"08",
          4093 => x"08",
          4094 => x"fe",
          4095 => x"82",
          4096 => x"81",
          4097 => x"05",
          4098 => x"f6",
          4099 => x"81",
          4100 => x"70",
          4101 => x"81",
          4102 => x"09",
          4103 => x"84",
          4104 => x"a8",
          4105 => x"08",
          4106 => x"7d",
          4107 => x"84",
          4108 => x"b4",
          4109 => x"81",
          4110 => x"81",
          4111 => x"09",
          4112 => x"84",
          4113 => x"a8",
          4114 => x"5b",
          4115 => x"c5",
          4116 => x"2e",
          4117 => x"54",
          4118 => x"53",
          4119 => x"f1",
          4120 => x"54",
          4121 => x"53",
          4122 => x"3f",
          4123 => x"2e",
          4124 => x"bb",
          4125 => x"08",
          4126 => x"08",
          4127 => x"fb",
          4128 => x"82",
          4129 => x"81",
          4130 => x"05",
          4131 => x"f4",
          4132 => x"81",
          4133 => x"05",
          4134 => x"f3",
          4135 => x"7a",
          4136 => x"3d",
          4137 => x"82",
          4138 => x"9c",
          4139 => x"55",
          4140 => x"24",
          4141 => x"8a",
          4142 => x"3d",
          4143 => x"08",
          4144 => x"58",
          4145 => x"83",
          4146 => x"2e",
          4147 => x"54",
          4148 => x"33",
          4149 => x"08",
          4150 => x"5a",
          4151 => x"ff",
          4152 => x"79",
          4153 => x"5e",
          4154 => x"5a",
          4155 => x"1a",
          4156 => x"3d",
          4157 => x"06",
          4158 => x"1a",
          4159 => x"08",
          4160 => x"38",
          4161 => x"7c",
          4162 => x"81",
          4163 => x"19",
          4164 => x"84",
          4165 => x"81",
          4166 => x"79",
          4167 => x"fc",
          4168 => x"33",
          4169 => x"f0",
          4170 => x"7d",
          4171 => x"b9",
          4172 => x"ba",
          4173 => x"bb",
          4174 => x"fe",
          4175 => x"89",
          4176 => x"08",
          4177 => x"38",
          4178 => x"56",
          4179 => x"82",
          4180 => x"19",
          4181 => x"3f",
          4182 => x"38",
          4183 => x"0c",
          4184 => x"83",
          4185 => x"77",
          4186 => x"7c",
          4187 => x"9f",
          4188 => x"07",
          4189 => x"83",
          4190 => x"08",
          4191 => x"56",
          4192 => x"81",
          4193 => x"81",
          4194 => x"81",
          4195 => x"09",
          4196 => x"84",
          4197 => x"70",
          4198 => x"84",
          4199 => x"74",
          4200 => x"55",
          4201 => x"54",
          4202 => x"51",
          4203 => x"80",
          4204 => x"75",
          4205 => x"7d",
          4206 => x"84",
          4207 => x"88",
          4208 => x"8f",
          4209 => x"81",
          4210 => x"81",
          4211 => x"81",
          4212 => x"81",
          4213 => x"09",
          4214 => x"84",
          4215 => x"70",
          4216 => x"84",
          4217 => x"7e",
          4218 => x"33",
          4219 => x"fb",
          4220 => x"7c",
          4221 => x"3f",
          4222 => x"76",
          4223 => x"33",
          4224 => x"84",
          4225 => x"06",
          4226 => x"83",
          4227 => x"1b",
          4228 => x"84",
          4229 => x"27",
          4230 => x"74",
          4231 => x"38",
          4232 => x"81",
          4233 => x"5c",
          4234 => x"b8",
          4235 => x"57",
          4236 => x"84",
          4237 => x"c5",
          4238 => x"34",
          4239 => x"31",
          4240 => x"5d",
          4241 => x"87",
          4242 => x"2e",
          4243 => x"54",
          4244 => x"33",
          4245 => x"e7",
          4246 => x"52",
          4247 => x"7e",
          4248 => x"83",
          4249 => x"ff",
          4250 => x"34",
          4251 => x"34",
          4252 => x"39",
          4253 => x"7a",
          4254 => x"98",
          4255 => x"06",
          4256 => x"7d",
          4257 => x"1d",
          4258 => x"1d",
          4259 => x"1d",
          4260 => x"7c",
          4261 => x"81",
          4262 => x"80",
          4263 => x"08",
          4264 => x"70",
          4265 => x"38",
          4266 => x"56",
          4267 => x"26",
          4268 => x"82",
          4269 => x"f5",
          4270 => x"81",
          4271 => x"08",
          4272 => x"08",
          4273 => x"25",
          4274 => x"73",
          4275 => x"81",
          4276 => x"84",
          4277 => x"81",
          4278 => x"08",
          4279 => x"f0",
          4280 => x"84",
          4281 => x"08",
          4282 => x"ce",
          4283 => x"08",
          4284 => x"39",
          4285 => x"26",
          4286 => x"51",
          4287 => x"84",
          4288 => x"bb",
          4289 => x"07",
          4290 => x"84",
          4291 => x"ff",
          4292 => x"2e",
          4293 => x"74",
          4294 => x"08",
          4295 => x"57",
          4296 => x"8e",
          4297 => x"f5",
          4298 => x"bb",
          4299 => x"08",
          4300 => x"80",
          4301 => x"90",
          4302 => x"94",
          4303 => x"86",
          4304 => x"19",
          4305 => x"34",
          4306 => x"8c",
          4307 => x"84",
          4308 => x"84",
          4309 => x"2e",
          4310 => x"78",
          4311 => x"08",
          4312 => x"08",
          4313 => x"04",
          4314 => x"38",
          4315 => x"0d",
          4316 => x"73",
          4317 => x"73",
          4318 => x"73",
          4319 => x"74",
          4320 => x"82",
          4321 => x"53",
          4322 => x"72",
          4323 => x"98",
          4324 => x"18",
          4325 => x"94",
          4326 => x"0c",
          4327 => x"9c",
          4328 => x"84",
          4329 => x"84",
          4330 => x"ac",
          4331 => x"ac",
          4332 => x"57",
          4333 => x"17",
          4334 => x"56",
          4335 => x"8a",
          4336 => x"08",
          4337 => x"ff",
          4338 => x"cd",
          4339 => x"bb",
          4340 => x"0b",
          4341 => x"38",
          4342 => x"08",
          4343 => x"31",
          4344 => x"aa",
          4345 => x"8a",
          4346 => x"70",
          4347 => x"5a",
          4348 => x"38",
          4349 => x"08",
          4350 => x"38",
          4351 => x"38",
          4352 => x"75",
          4353 => x"22",
          4354 => x"38",
          4355 => x"0c",
          4356 => x"80",
          4357 => x"3d",
          4358 => x"19",
          4359 => x"5c",
          4360 => x"eb",
          4361 => x"82",
          4362 => x"27",
          4363 => x"08",
          4364 => x"84",
          4365 => x"60",
          4366 => x"08",
          4367 => x"bb",
          4368 => x"84",
          4369 => x"56",
          4370 => x"91",
          4371 => x"ff",
          4372 => x"08",
          4373 => x"ea",
          4374 => x"05",
          4375 => x"8d",
          4376 => x"b0",
          4377 => x"1a",
          4378 => x"57",
          4379 => x"34",
          4380 => x"56",
          4381 => x"81",
          4382 => x"77",
          4383 => x"3f",
          4384 => x"81",
          4385 => x"0c",
          4386 => x"3d",
          4387 => x"53",
          4388 => x"52",
          4389 => x"08",
          4390 => x"83",
          4391 => x"08",
          4392 => x"fe",
          4393 => x"82",
          4394 => x"81",
          4395 => x"05",
          4396 => x"e3",
          4397 => x"22",
          4398 => x"74",
          4399 => x"7c",
          4400 => x"08",
          4401 => x"7d",
          4402 => x"76",
          4403 => x"19",
          4404 => x"84",
          4405 => x"ee",
          4406 => x"7c",
          4407 => x"1e",
          4408 => x"82",
          4409 => x"80",
          4410 => x"d1",
          4411 => x"74",
          4412 => x"38",
          4413 => x"81",
          4414 => x"bb",
          4415 => x"5a",
          4416 => x"5b",
          4417 => x"70",
          4418 => x"81",
          4419 => x"81",
          4420 => x"34",
          4421 => x"ae",
          4422 => x"80",
          4423 => x"74",
          4424 => x"56",
          4425 => x"60",
          4426 => x"80",
          4427 => x"bb",
          4428 => x"81",
          4429 => x"fe",
          4430 => x"94",
          4431 => x"08",
          4432 => x"e1",
          4433 => x"08",
          4434 => x"38",
          4435 => x"b4",
          4436 => x"bb",
          4437 => x"08",
          4438 => x"41",
          4439 => x"a8",
          4440 => x"1a",
          4441 => x"33",
          4442 => x"90",
          4443 => x"81",
          4444 => x"5b",
          4445 => x"33",
          4446 => x"08",
          4447 => x"76",
          4448 => x"74",
          4449 => x"60",
          4450 => x"c1",
          4451 => x"0c",
          4452 => x"0d",
          4453 => x"18",
          4454 => x"06",
          4455 => x"33",
          4456 => x"58",
          4457 => x"33",
          4458 => x"05",
          4459 => x"e7",
          4460 => x"33",
          4461 => x"44",
          4462 => x"79",
          4463 => x"10",
          4464 => x"23",
          4465 => x"77",
          4466 => x"2a",
          4467 => x"90",
          4468 => x"38",
          4469 => x"23",
          4470 => x"41",
          4471 => x"2e",
          4472 => x"39",
          4473 => x"74",
          4474 => x"78",
          4475 => x"05",
          4476 => x"56",
          4477 => x"fd",
          4478 => x"7a",
          4479 => x"04",
          4480 => x"5c",
          4481 => x"84",
          4482 => x"08",
          4483 => x"5d",
          4484 => x"5e",
          4485 => x"1b",
          4486 => x"1b",
          4487 => x"09",
          4488 => x"75",
          4489 => x"51",
          4490 => x"80",
          4491 => x"75",
          4492 => x"b2",
          4493 => x"59",
          4494 => x"19",
          4495 => x"57",
          4496 => x"e5",
          4497 => x"81",
          4498 => x"38",
          4499 => x"81",
          4500 => x"56",
          4501 => x"81",
          4502 => x"5a",
          4503 => x"06",
          4504 => x"38",
          4505 => x"1c",
          4506 => x"8b",
          4507 => x"81",
          4508 => x"5a",
          4509 => x"58",
          4510 => x"38",
          4511 => x"5d",
          4512 => x"7b",
          4513 => x"08",
          4514 => x"fe",
          4515 => x"93",
          4516 => x"08",
          4517 => x"dc",
          4518 => x"08",
          4519 => x"38",
          4520 => x"b4",
          4521 => x"bb",
          4522 => x"08",
          4523 => x"5a",
          4524 => x"dd",
          4525 => x"1c",
          4526 => x"33",
          4527 => x"c5",
          4528 => x"1c",
          4529 => x"55",
          4530 => x"81",
          4531 => x"8d",
          4532 => x"90",
          4533 => x"5e",
          4534 => x"ff",
          4535 => x"f4",
          4536 => x"84",
          4537 => x"38",
          4538 => x"c2",
          4539 => x"1d",
          4540 => x"57",
          4541 => x"38",
          4542 => x"1b",
          4543 => x"40",
          4544 => x"bf",
          4545 => x"81",
          4546 => x"33",
          4547 => x"71",
          4548 => x"80",
          4549 => x"26",
          4550 => x"d1",
          4551 => x"61",
          4552 => x"5b",
          4553 => x"bb",
          4554 => x"de",
          4555 => x"78",
          4556 => x"86",
          4557 => x"2e",
          4558 => x"79",
          4559 => x"7f",
          4560 => x"ff",
          4561 => x"0b",
          4562 => x"04",
          4563 => x"38",
          4564 => x"3d",
          4565 => x"33",
          4566 => x"86",
          4567 => x"1d",
          4568 => x"80",
          4569 => x"17",
          4570 => x"38",
          4571 => x"60",
          4572 => x"05",
          4573 => x"34",
          4574 => x"80",
          4575 => x"56",
          4576 => x"c0",
          4577 => x"3d",
          4578 => x"59",
          4579 => x"70",
          4580 => x"05",
          4581 => x"38",
          4582 => x"79",
          4583 => x"38",
          4584 => x"75",
          4585 => x"2a",
          4586 => x"2a",
          4587 => x"80",
          4588 => x"32",
          4589 => x"d7",
          4590 => x"87",
          4591 => x"58",
          4592 => x"75",
          4593 => x"76",
          4594 => x"2a",
          4595 => x"1f",
          4596 => x"58",
          4597 => x"33",
          4598 => x"16",
          4599 => x"75",
          4600 => x"2e",
          4601 => x"56",
          4602 => x"98",
          4603 => x"71",
          4604 => x"87",
          4605 => x"f8",
          4606 => x"38",
          4607 => x"fe",
          4608 => x"2e",
          4609 => x"56",
          4610 => x"81",
          4611 => x"05",
          4612 => x"84",
          4613 => x"75",
          4614 => x"7e",
          4615 => x"1d",
          4616 => x"84",
          4617 => x"ed",
          4618 => x"84",
          4619 => x"bb",
          4620 => x"1e",
          4621 => x"76",
          4622 => x"40",
          4623 => x"a3",
          4624 => x"52",
          4625 => x"84",
          4626 => x"ff",
          4627 => x"76",
          4628 => x"70",
          4629 => x"81",
          4630 => x"78",
          4631 => x"c9",
          4632 => x"86",
          4633 => x"83",
          4634 => x"bb",
          4635 => x"87",
          4636 => x"75",
          4637 => x"40",
          4638 => x"57",
          4639 => x"83",
          4640 => x"82",
          4641 => x"52",
          4642 => x"84",
          4643 => x"ff",
          4644 => x"75",
          4645 => x"9c",
          4646 => x"81",
          4647 => x"f4",
          4648 => x"58",
          4649 => x"33",
          4650 => x"15",
          4651 => x"ab",
          4652 => x"8c",
          4653 => x"77",
          4654 => x"3d",
          4655 => x"25",
          4656 => x"b9",
          4657 => x"ec",
          4658 => x"84",
          4659 => x"38",
          4660 => x"08",
          4661 => x"d3",
          4662 => x"2e",
          4663 => x"bb",
          4664 => x"08",
          4665 => x"19",
          4666 => x"41",
          4667 => x"bb",
          4668 => x"85",
          4669 => x"58",
          4670 => x"84",
          4671 => x"ef",
          4672 => x"58",
          4673 => x"80",
          4674 => x"33",
          4675 => x"ff",
          4676 => x"74",
          4677 => x"98",
          4678 => x"08",
          4679 => x"5b",
          4680 => x"c9",
          4681 => x"52",
          4682 => x"84",
          4683 => x"ff",
          4684 => x"75",
          4685 => x"08",
          4686 => x"5f",
          4687 => x"0b",
          4688 => x"75",
          4689 => x"7c",
          4690 => x"58",
          4691 => x"38",
          4692 => x"5b",
          4693 => x"7b",
          4694 => x"57",
          4695 => x"34",
          4696 => x"81",
          4697 => x"76",
          4698 => x"78",
          4699 => x"80",
          4700 => x"81",
          4701 => x"51",
          4702 => x"58",
          4703 => x"7f",
          4704 => x"fb",
          4705 => x"53",
          4706 => x"52",
          4707 => x"bb",
          4708 => x"84",
          4709 => x"a8",
          4710 => x"57",
          4711 => x"c9",
          4712 => x"2e",
          4713 => x"54",
          4714 => x"53",
          4715 => x"d1",
          4716 => x"9c",
          4717 => x"74",
          4718 => x"ba",
          4719 => x"57",
          4720 => x"d7",
          4721 => x"d4",
          4722 => x"61",
          4723 => x"3f",
          4724 => x"81",
          4725 => x"83",
          4726 => x"08",
          4727 => x"8a",
          4728 => x"2e",
          4729 => x"fc",
          4730 => x"7f",
          4731 => x"39",
          4732 => x"70",
          4733 => x"38",
          4734 => x"08",
          4735 => x"81",
          4736 => x"c1",
          4737 => x"19",
          4738 => x"33",
          4739 => x"f3",
          4740 => x"5e",
          4741 => x"1c",
          4742 => x"1c",
          4743 => x"70",
          4744 => x"57",
          4745 => x"bc",
          4746 => x"81",
          4747 => x"38",
          4748 => x"ff",
          4749 => x"82",
          4750 => x"70",
          4751 => x"38",
          4752 => x"7a",
          4753 => x"05",
          4754 => x"70",
          4755 => x"08",
          4756 => x"53",
          4757 => x"2e",
          4758 => x"30",
          4759 => x"54",
          4760 => x"2e",
          4761 => x"59",
          4762 => x"81",
          4763 => x"76",
          4764 => x"05",
          4765 => x"1d",
          4766 => x"f3",
          4767 => x"57",
          4768 => x"82",
          4769 => x"33",
          4770 => x"1e",
          4771 => x"33",
          4772 => x"11",
          4773 => x"90",
          4774 => x"33",
          4775 => x"71",
          4776 => x"96",
          4777 => x"41",
          4778 => x"86",
          4779 => x"33",
          4780 => x"84",
          4781 => x"e5",
          4782 => x"11",
          4783 => x"83",
          4784 => x"51",
          4785 => x"08",
          4786 => x"75",
          4787 => x"b3",
          4788 => x"34",
          4789 => x"58",
          4790 => x"78",
          4791 => x"54",
          4792 => x"74",
          4793 => x"25",
          4794 => x"75",
          4795 => x"78",
          4796 => x"56",
          4797 => x"33",
          4798 => x"88",
          4799 => x"54",
          4800 => x"54",
          4801 => x"08",
          4802 => x"27",
          4803 => x"81",
          4804 => x"a0",
          4805 => x"53",
          4806 => x"81",
          4807 => x"13",
          4808 => x"ff",
          4809 => x"2a",
          4810 => x"80",
          4811 => x"5f",
          4812 => x"63",
          4813 => x"65",
          4814 => x"2e",
          4815 => x"2e",
          4816 => x"d9",
          4817 => x"73",
          4818 => x"55",
          4819 => x"42",
          4820 => x"70",
          4821 => x"73",
          4822 => x"ff",
          4823 => x"74",
          4824 => x"80",
          4825 => x"ff",
          4826 => x"9f",
          4827 => x"5b",
          4828 => x"80",
          4829 => x"ff",
          4830 => x"83",
          4831 => x"56",
          4832 => x"38",
          4833 => x"70",
          4834 => x"56",
          4835 => x"5b",
          4836 => x"26",
          4837 => x"74",
          4838 => x"81",
          4839 => x"80",
          4840 => x"81",
          4841 => x"80",
          4842 => x"72",
          4843 => x"46",
          4844 => x"af",
          4845 => x"70",
          4846 => x"54",
          4847 => x"0c",
          4848 => x"42",
          4849 => x"b4",
          4850 => x"8d",
          4851 => x"ff",
          4852 => x"86",
          4853 => x"3d",
          4854 => x"81",
          4855 => x"fe",
          4856 => x"ab",
          4857 => x"8d",
          4858 => x"84",
          4859 => x"80",
          4860 => x"73",
          4861 => x"2e",
          4862 => x"70",
          4863 => x"dd",
          4864 => x"70",
          4865 => x"7d",
          4866 => x"27",
          4867 => x"f8",
          4868 => x"76",
          4869 => x"76",
          4870 => x"70",
          4871 => x"52",
          4872 => x"2e",
          4873 => x"57",
          4874 => x"56",
          4875 => x"c7",
          4876 => x"ff",
          4877 => x"a0",
          4878 => x"ff",
          4879 => x"38",
          4880 => x"fe",
          4881 => x"2e",
          4882 => x"54",
          4883 => x"38",
          4884 => x"ae",
          4885 => x"0b",
          4886 => x"81",
          4887 => x"f4",
          4888 => x"16",
          4889 => x"5d",
          4890 => x"a0",
          4891 => x"70",
          4892 => x"75",
          4893 => x"bb",
          4894 => x"38",
          4895 => x"70",
          4896 => x"51",
          4897 => x"e0",
          4898 => x"75",
          4899 => x"5a",
          4900 => x"88",
          4901 => x"06",
          4902 => x"70",
          4903 => x"ff",
          4904 => x"81",
          4905 => x"2e",
          4906 => x"77",
          4907 => x"06",
          4908 => x"79",
          4909 => x"38",
          4910 => x"85",
          4911 => x"2a",
          4912 => x"38",
          4913 => x"34",
          4914 => x"84",
          4915 => x"bb",
          4916 => x"84",
          4917 => x"06",
          4918 => x"06",
          4919 => x"74",
          4920 => x"98",
          4921 => x"42",
          4922 => x"ce",
          4923 => x"70",
          4924 => x"2e",
          4925 => x"38",
          4926 => x"82",
          4927 => x"81",
          4928 => x"73",
          4929 => x"38",
          4930 => x"80",
          4931 => x"76",
          4932 => x"75",
          4933 => x"53",
          4934 => x"07",
          4935 => x"e3",
          4936 => x"1d",
          4937 => x"fe",
          4938 => x"58",
          4939 => x"70",
          4940 => x"80",
          4941 => x"83",
          4942 => x"33",
          4943 => x"07",
          4944 => x"83",
          4945 => x"0c",
          4946 => x"39",
          4947 => x"f0",
          4948 => x"38",
          4949 => x"17",
          4950 => x"2b",
          4951 => x"5e",
          4952 => x"95",
          4953 => x"39",
          4954 => x"2e",
          4955 => x"39",
          4956 => x"0b",
          4957 => x"04",
          4958 => x"ff",
          4959 => x"59",
          4960 => x"83",
          4961 => x"fc",
          4962 => x"b5",
          4963 => x"84",
          4964 => x"70",
          4965 => x"80",
          4966 => x"83",
          4967 => x"81",
          4968 => x"2e",
          4969 => x"83",
          4970 => x"56",
          4971 => x"38",
          4972 => x"70",
          4973 => x"59",
          4974 => x"59",
          4975 => x"54",
          4976 => x"07",
          4977 => x"9f",
          4978 => x"7d",
          4979 => x"17",
          4980 => x"5f",
          4981 => x"79",
          4982 => x"fa",
          4983 => x"83",
          4984 => x"5a",
          4985 => x"80",
          4986 => x"05",
          4987 => x"1b",
          4988 => x"80",
          4989 => x"90",
          4990 => x"5a",
          4991 => x"05",
          4992 => x"34",
          4993 => x"5b",
          4994 => x"9c",
          4995 => x"58",
          4996 => x"06",
          4997 => x"82",
          4998 => x"38",
          4999 => x"3d",
          5000 => x"02",
          5001 => x"42",
          5002 => x"70",
          5003 => x"d7",
          5004 => x"70",
          5005 => x"85",
          5006 => x"2e",
          5007 => x"56",
          5008 => x"10",
          5009 => x"58",
          5010 => x"96",
          5011 => x"06",
          5012 => x"9b",
          5013 => x"b0",
          5014 => x"06",
          5015 => x"2e",
          5016 => x"16",
          5017 => x"18",
          5018 => x"ff",
          5019 => x"81",
          5020 => x"83",
          5021 => x"2e",
          5022 => x"41",
          5023 => x"5b",
          5024 => x"18",
          5025 => x"7a",
          5026 => x"33",
          5027 => x"bb",
          5028 => x"55",
          5029 => x"56",
          5030 => x"84",
          5031 => x"56",
          5032 => x"2e",
          5033 => x"38",
          5034 => x"85",
          5035 => x"83",
          5036 => x"83",
          5037 => x"c3",
          5038 => x"59",
          5039 => x"83",
          5040 => x"ce",
          5041 => x"5a",
          5042 => x"11",
          5043 => x"71",
          5044 => x"72",
          5045 => x"56",
          5046 => x"a0",
          5047 => x"18",
          5048 => x"70",
          5049 => x"58",
          5050 => x"81",
          5051 => x"19",
          5052 => x"23",
          5053 => x"38",
          5054 => x"bb",
          5055 => x"18",
          5056 => x"74",
          5057 => x"5e",
          5058 => x"80",
          5059 => x"71",
          5060 => x"38",
          5061 => x"12",
          5062 => x"07",
          5063 => x"2b",
          5064 => x"58",
          5065 => x"80",
          5066 => x"5d",
          5067 => x"ce",
          5068 => x"5a",
          5069 => x"52",
          5070 => x"3f",
          5071 => x"84",
          5072 => x"bb",
          5073 => x"26",
          5074 => x"f5",
          5075 => x"f5",
          5076 => x"16",
          5077 => x"0c",
          5078 => x"1d",
          5079 => x"2e",
          5080 => x"8d",
          5081 => x"7d",
          5082 => x"7c",
          5083 => x"70",
          5084 => x"5a",
          5085 => x"58",
          5086 => x"ff",
          5087 => x"18",
          5088 => x"7c",
          5089 => x"34",
          5090 => x"7c",
          5091 => x"23",
          5092 => x"80",
          5093 => x"84",
          5094 => x"8b",
          5095 => x"0d",
          5096 => x"ff",
          5097 => x"91",
          5098 => x"d0",
          5099 => x"fe",
          5100 => x"5f",
          5101 => x"7a",
          5102 => x"81",
          5103 => x"58",
          5104 => x"16",
          5105 => x"9f",
          5106 => x"e0",
          5107 => x"75",
          5108 => x"77",
          5109 => x"ff",
          5110 => x"70",
          5111 => x"58",
          5112 => x"81",
          5113 => x"25",
          5114 => x"39",
          5115 => x"82",
          5116 => x"fe",
          5117 => x"7a",
          5118 => x"2e",
          5119 => x"75",
          5120 => x"25",
          5121 => x"ad",
          5122 => x"38",
          5123 => x"83",
          5124 => x"80",
          5125 => x"84",
          5126 => x"88",
          5127 => x"72",
          5128 => x"71",
          5129 => x"77",
          5130 => x"19",
          5131 => x"ff",
          5132 => x"70",
          5133 => x"9b",
          5134 => x"84",
          5135 => x"42",
          5136 => x"2e",
          5137 => x"34",
          5138 => x"80",
          5139 => x"54",
          5140 => x"33",
          5141 => x"84",
          5142 => x"81",
          5143 => x"75",
          5144 => x"71",
          5145 => x"7b",
          5146 => x"a8",
          5147 => x"58",
          5148 => x"75",
          5149 => x"25",
          5150 => x"38",
          5151 => x"58",
          5152 => x"84",
          5153 => x"78",
          5154 => x"58",
          5155 => x"80",
          5156 => x"1a",
          5157 => x"38",
          5158 => x"18",
          5159 => x"70",
          5160 => x"05",
          5161 => x"5b",
          5162 => x"c5",
          5163 => x"0b",
          5164 => x"5d",
          5165 => x"7e",
          5166 => x"31",
          5167 => x"80",
          5168 => x"e1",
          5169 => x"58",
          5170 => x"84",
          5171 => x"75",
          5172 => x"81",
          5173 => x"58",
          5174 => x"84",
          5175 => x"80",
          5176 => x"58",
          5177 => x"70",
          5178 => x"ff",
          5179 => x"2e",
          5180 => x"38",
          5181 => x"b8",
          5182 => x"5a",
          5183 => x"71",
          5184 => x"40",
          5185 => x"80",
          5186 => x"5a",
          5187 => x"fd",
          5188 => x"e8",
          5189 => x"55",
          5190 => x"d5",
          5191 => x"17",
          5192 => x"33",
          5193 => x"82",
          5194 => x"17",
          5195 => x"d2",
          5196 => x"85",
          5197 => x"18",
          5198 => x"18",
          5199 => x"18",
          5200 => x"75",
          5201 => x"f8",
          5202 => x"82",
          5203 => x"2b",
          5204 => x"88",
          5205 => x"59",
          5206 => x"85",
          5207 => x"cd",
          5208 => x"82",
          5209 => x"2b",
          5210 => x"88",
          5211 => x"40",
          5212 => x"85",
          5213 => x"9d",
          5214 => x"82",
          5215 => x"2b",
          5216 => x"88",
          5217 => x"0c",
          5218 => x"82",
          5219 => x"2b",
          5220 => x"88",
          5221 => x"05",
          5222 => x"40",
          5223 => x"84",
          5224 => x"84",
          5225 => x"84",
          5226 => x"0b",
          5227 => x"83",
          5228 => x"0c",
          5229 => x"17",
          5230 => x"18",
          5231 => x"84",
          5232 => x"06",
          5233 => x"83",
          5234 => x"08",
          5235 => x"8b",
          5236 => x"2e",
          5237 => x"5a",
          5238 => x"2e",
          5239 => x"18",
          5240 => x"ab",
          5241 => x"18",
          5242 => x"8d",
          5243 => x"22",
          5244 => x"17",
          5245 => x"90",
          5246 => x"33",
          5247 => x"71",
          5248 => x"2b",
          5249 => x"d8",
          5250 => x"e8",
          5251 => x"80",
          5252 => x"57",
          5253 => x"5a",
          5254 => x"75",
          5255 => x"05",
          5256 => x"ff",
          5257 => x"3d",
          5258 => x"70",
          5259 => x"76",
          5260 => x"38",
          5261 => x"9f",
          5262 => x"e2",
          5263 => x"80",
          5264 => x"80",
          5265 => x"10",
          5266 => x"55",
          5267 => x"34",
          5268 => x"80",
          5269 => x"7c",
          5270 => x"53",
          5271 => x"ef",
          5272 => x"73",
          5273 => x"04",
          5274 => x"3d",
          5275 => x"81",
          5276 => x"26",
          5277 => x"06",
          5278 => x"80",
          5279 => x"f4",
          5280 => x"5a",
          5281 => x"70",
          5282 => x"59",
          5283 => x"e0",
          5284 => x"ff",
          5285 => x"38",
          5286 => x"54",
          5287 => x"74",
          5288 => x"76",
          5289 => x"30",
          5290 => x"5c",
          5291 => x"81",
          5292 => x"25",
          5293 => x"39",
          5294 => x"60",
          5295 => x"0d",
          5296 => x"33",
          5297 => x"a6",
          5298 => x"3d",
          5299 => x"52",
          5300 => x"08",
          5301 => x"8f",
          5302 => x"84",
          5303 => x"7e",
          5304 => x"5c",
          5305 => x"57",
          5306 => x"ba",
          5307 => x"2e",
          5308 => x"e0",
          5309 => x"78",
          5310 => x"78",
          5311 => x"2e",
          5312 => x"9a",
          5313 => x"70",
          5314 => x"83",
          5315 => x"17",
          5316 => x"0b",
          5317 => x"17",
          5318 => x"34",
          5319 => x"17",
          5320 => x"33",
          5321 => x"66",
          5322 => x"0b",
          5323 => x"34",
          5324 => x"81",
          5325 => x"80",
          5326 => x"7e",
          5327 => x"27",
          5328 => x"83",
          5329 => x"fe",
          5330 => x"70",
          5331 => x"fe",
          5332 => x"57",
          5333 => x"38",
          5334 => x"2a",
          5335 => x"38",
          5336 => x"80",
          5337 => x"77",
          5338 => x"06",
          5339 => x"80",
          5340 => x"a0",
          5341 => x"9b",
          5342 => x"2b",
          5343 => x"5b",
          5344 => x"88",
          5345 => x"82",
          5346 => x"2b",
          5347 => x"88",
          5348 => x"05",
          5349 => x"5e",
          5350 => x"23",
          5351 => x"1b",
          5352 => x"0b",
          5353 => x"80",
          5354 => x"05",
          5355 => x"38",
          5356 => x"80",
          5357 => x"55",
          5358 => x"94",
          5359 => x"2b",
          5360 => x"5b",
          5361 => x"51",
          5362 => x"81",
          5363 => x"2e",
          5364 => x"ff",
          5365 => x"58",
          5366 => x"38",
          5367 => x"2e",
          5368 => x"39",
          5369 => x"5e",
          5370 => x"06",
          5371 => x"88",
          5372 => x"87",
          5373 => x"84",
          5374 => x"7a",
          5375 => x"39",
          5376 => x"98",
          5377 => x"88",
          5378 => x"82",
          5379 => x"2b",
          5380 => x"88",
          5381 => x"05",
          5382 => x"54",
          5383 => x"84",
          5384 => x"0b",
          5385 => x"0c",
          5386 => x"5c",
          5387 => x"39",
          5388 => x"84",
          5389 => x"fa",
          5390 => x"7b",
          5391 => x"84",
          5392 => x"2e",
          5393 => x"81",
          5394 => x"08",
          5395 => x"74",
          5396 => x"84",
          5397 => x"16",
          5398 => x"56",
          5399 => x"17",
          5400 => x"07",
          5401 => x"77",
          5402 => x"7f",
          5403 => x"08",
          5404 => x"58",
          5405 => x"eb",
          5406 => x"52",
          5407 => x"3f",
          5408 => x"38",
          5409 => x"0c",
          5410 => x"0c",
          5411 => x"80",
          5412 => x"94",
          5413 => x"fa",
          5414 => x"33",
          5415 => x"7d",
          5416 => x"17",
          5417 => x"0b",
          5418 => x"17",
          5419 => x"34",
          5420 => x"17",
          5421 => x"33",
          5422 => x"f9",
          5423 => x"1b",
          5424 => x"ff",
          5425 => x"38",
          5426 => x"05",
          5427 => x"ea",
          5428 => x"b0",
          5429 => x"2e",
          5430 => x"70",
          5431 => x"53",
          5432 => x"a1",
          5433 => x"2e",
          5434 => x"0c",
          5435 => x"08",
          5436 => x"33",
          5437 => x"bb",
          5438 => x"80",
          5439 => x"17",
          5440 => x"31",
          5441 => x"a0",
          5442 => x"16",
          5443 => x"06",
          5444 => x"08",
          5445 => x"81",
          5446 => x"7c",
          5447 => x"08",
          5448 => x"81",
          5449 => x"60",
          5450 => x"80",
          5451 => x"9f",
          5452 => x"97",
          5453 => x"8f",
          5454 => x"59",
          5455 => x"80",
          5456 => x"e7",
          5457 => x"df",
          5458 => x"87",
          5459 => x"94",
          5460 => x"56",
          5461 => x"79",
          5462 => x"ff",
          5463 => x"8a",
          5464 => x"06",
          5465 => x"d0",
          5466 => x"27",
          5467 => x"ae",
          5468 => x"98",
          5469 => x"fe",
          5470 => x"a5",
          5471 => x"b0",
          5472 => x"2e",
          5473 => x"2a",
          5474 => x"38",
          5475 => x"38",
          5476 => x"53",
          5477 => x"9f",
          5478 => x"d6",
          5479 => x"59",
          5480 => x"7a",
          5481 => x"08",
          5482 => x"08",
          5483 => x"5a",
          5484 => x"84",
          5485 => x"74",
          5486 => x"04",
          5487 => x"08",
          5488 => x"90",
          5489 => x"52",
          5490 => x"81",
          5491 => x"33",
          5492 => x"84",
          5493 => x"80",
          5494 => x"7e",
          5495 => x"81",
          5496 => x"84",
          5497 => x"9c",
          5498 => x"83",
          5499 => x"55",
          5500 => x"76",
          5501 => x"56",
          5502 => x"70",
          5503 => x"05",
          5504 => x"2e",
          5505 => x"56",
          5506 => x"ff",
          5507 => x"39",
          5508 => x"a3",
          5509 => x"fd",
          5510 => x"9c",
          5511 => x"06",
          5512 => x"08",
          5513 => x"08",
          5514 => x"ef",
          5515 => x"a8",
          5516 => x"05",
          5517 => x"34",
          5518 => x"cf",
          5519 => x"77",
          5520 => x"55",
          5521 => x"0b",
          5522 => x"84",
          5523 => x"91",
          5524 => x"0c",
          5525 => x"61",
          5526 => x"80",
          5527 => x"9f",
          5528 => x"97",
          5529 => x"8f",
          5530 => x"59",
          5531 => x"80",
          5532 => x"cc",
          5533 => x"c4",
          5534 => x"81",
          5535 => x"2e",
          5536 => x"11",
          5537 => x"76",
          5538 => x"38",
          5539 => x"cd",
          5540 => x"78",
          5541 => x"38",
          5542 => x"55",
          5543 => x"81",
          5544 => x"83",
          5545 => x"19",
          5546 => x"7f",
          5547 => x"5b",
          5548 => x"98",
          5549 => x"fe",
          5550 => x"b8",
          5551 => x"b0",
          5552 => x"2e",
          5553 => x"2a",
          5554 => x"38",
          5555 => x"38",
          5556 => x"53",
          5557 => x"9b",
          5558 => x"e9",
          5559 => x"75",
          5560 => x"a8",
          5561 => x"58",
          5562 => x"77",
          5563 => x"55",
          5564 => x"ff",
          5565 => x"89",
          5566 => x"19",
          5567 => x"1a",
          5568 => x"08",
          5569 => x"27",
          5570 => x"0c",
          5571 => x"58",
          5572 => x"1a",
          5573 => x"0c",
          5574 => x"84",
          5575 => x"08",
          5576 => x"57",
          5577 => x"81",
          5578 => x"18",
          5579 => x"bb",
          5580 => x"08",
          5581 => x"ff",
          5582 => x"7a",
          5583 => x"79",
          5584 => x"77",
          5585 => x"05",
          5586 => x"34",
          5587 => x"19",
          5588 => x"1a",
          5589 => x"52",
          5590 => x"bb",
          5591 => x"fc",
          5592 => x"d8",
          5593 => x"d4",
          5594 => x"bb",
          5595 => x"81",
          5596 => x"52",
          5597 => x"3f",
          5598 => x"19",
          5599 => x"1a",
          5600 => x"16",
          5601 => x"bb",
          5602 => x"c7",
          5603 => x"c1",
          5604 => x"0b",
          5605 => x"04",
          5606 => x"84",
          5607 => x"f5",
          5608 => x"80",
          5609 => x"80",
          5610 => x"80",
          5611 => x"19",
          5612 => x"d2",
          5613 => x"76",
          5614 => x"86",
          5615 => x"2e",
          5616 => x"80",
          5617 => x"19",
          5618 => x"2e",
          5619 => x"71",
          5620 => x"81",
          5621 => x"53",
          5622 => x"ff",
          5623 => x"80",
          5624 => x"76",
          5625 => x"90",
          5626 => x"a0",
          5627 => x"77",
          5628 => x"ff",
          5629 => x"34",
          5630 => x"34",
          5631 => x"56",
          5632 => x"8c",
          5633 => x"88",
          5634 => x"90",
          5635 => x"98",
          5636 => x"7a",
          5637 => x"0b",
          5638 => x"18",
          5639 => x"0b",
          5640 => x"83",
          5641 => x"3f",
          5642 => x"81",
          5643 => x"34",
          5644 => x"8d",
          5645 => x"08",
          5646 => x"33",
          5647 => x"59",
          5648 => x"81",
          5649 => x"08",
          5650 => x"17",
          5651 => x"55",
          5652 => x"38",
          5653 => x"09",
          5654 => x"b4",
          5655 => x"7a",
          5656 => x"e9",
          5657 => x"90",
          5658 => x"88",
          5659 => x"18",
          5660 => x"2a",
          5661 => x"2a",
          5662 => x"2a",
          5663 => x"34",
          5664 => x"98",
          5665 => x"34",
          5666 => x"93",
          5667 => x"1c",
          5668 => x"84",
          5669 => x"bf",
          5670 => x"fe",
          5671 => x"92",
          5672 => x"06",
          5673 => x"08",
          5674 => x"9c",
          5675 => x"81",
          5676 => x"3f",
          5677 => x"f2",
          5678 => x"59",
          5679 => x"08",
          5680 => x"09",
          5681 => x"39",
          5682 => x"fb",
          5683 => x"84",
          5684 => x"74",
          5685 => x"72",
          5686 => x"71",
          5687 => x"84",
          5688 => x"96",
          5689 => x"75",
          5690 => x"bb",
          5691 => x"13",
          5692 => x"bb",
          5693 => x"38",
          5694 => x"f6",
          5695 => x"5b",
          5696 => x"81",
          5697 => x"52",
          5698 => x"38",
          5699 => x"e0",
          5700 => x"70",
          5701 => x"bb",
          5702 => x"0b",
          5703 => x"04",
          5704 => x"06",
          5705 => x"38",
          5706 => x"05",
          5707 => x"38",
          5708 => x"79",
          5709 => x"05",
          5710 => x"33",
          5711 => x"99",
          5712 => x"ff",
          5713 => x"70",
          5714 => x"81",
          5715 => x"9f",
          5716 => x"81",
          5717 => x"74",
          5718 => x"9f",
          5719 => x"80",
          5720 => x"5b",
          5721 => x"7a",
          5722 => x"f7",
          5723 => x"39",
          5724 => x"cc",
          5725 => x"3f",
          5726 => x"84",
          5727 => x"bb",
          5728 => x"5c",
          5729 => x"c6",
          5730 => x"84",
          5731 => x"80",
          5732 => x"5a",
          5733 => x"b2",
          5734 => x"57",
          5735 => x"63",
          5736 => x"88",
          5737 => x"57",
          5738 => x"98",
          5739 => x"98",
          5740 => x"84",
          5741 => x"85",
          5742 => x"0d",
          5743 => x"71",
          5744 => x"07",
          5745 => x"7a",
          5746 => x"bb",
          5747 => x"9e",
          5748 => x"e6",
          5749 => x"80",
          5750 => x"52",
          5751 => x"84",
          5752 => x"08",
          5753 => x"0c",
          5754 => x"3d",
          5755 => x"58",
          5756 => x"d8",
          5757 => x"7a",
          5758 => x"84",
          5759 => x"92",
          5760 => x"56",
          5761 => x"84",
          5762 => x"5d",
          5763 => x"53",
          5764 => x"ff",
          5765 => x"80",
          5766 => x"76",
          5767 => x"80",
          5768 => x"12",
          5769 => x"33",
          5770 => x"2e",
          5771 => x"0c",
          5772 => x"3f",
          5773 => x"84",
          5774 => x"51",
          5775 => x"08",
          5776 => x"80",
          5777 => x"12",
          5778 => x"33",
          5779 => x"2e",
          5780 => x"38",
          5781 => x"ff",
          5782 => x"59",
          5783 => x"b4",
          5784 => x"78",
          5785 => x"b8",
          5786 => x"3f",
          5787 => x"79",
          5788 => x"81",
          5789 => x"57",
          5790 => x"78",
          5791 => x"9c",
          5792 => x"18",
          5793 => x"ff",
          5794 => x"75",
          5795 => x"e6",
          5796 => x"34",
          5797 => x"bd",
          5798 => x"80",
          5799 => x"10",
          5800 => x"33",
          5801 => x"2e",
          5802 => x"33",
          5803 => x"1a",
          5804 => x"57",
          5805 => x"5f",
          5806 => x"34",
          5807 => x"38",
          5808 => x"76",
          5809 => x"38",
          5810 => x"bb",
          5811 => x"95",
          5812 => x"2b",
          5813 => x"56",
          5814 => x"94",
          5815 => x"2b",
          5816 => x"5a",
          5817 => x"8d",
          5818 => x"bb",
          5819 => x"ff",
          5820 => x"53",
          5821 => x"52",
          5822 => x"84",
          5823 => x"bb",
          5824 => x"08",
          5825 => x"08",
          5826 => x"fc",
          5827 => x"82",
          5828 => x"81",
          5829 => x"05",
          5830 => x"ff",
          5831 => x"39",
          5832 => x"5c",
          5833 => x"e2",
          5834 => x"f4",
          5835 => x"59",
          5836 => x"06",
          5837 => x"e5",
          5838 => x"79",
          5839 => x"77",
          5840 => x"3d",
          5841 => x"33",
          5842 => x"78",
          5843 => x"59",
          5844 => x"0c",
          5845 => x"0d",
          5846 => x"80",
          5847 => x"80",
          5848 => x"80",
          5849 => x"18",
          5850 => x"ee",
          5851 => x"77",
          5852 => x"74",
          5853 => x"78",
          5854 => x"08",
          5855 => x"85",
          5856 => x"2b",
          5857 => x"fc",
          5858 => x"bb",
          5859 => x"17",
          5860 => x"bb",
          5861 => x"26",
          5862 => x"70",
          5863 => x"19",
          5864 => x"81",
          5865 => x"38",
          5866 => x"94",
          5867 => x"2a",
          5868 => x"2e",
          5869 => x"ff",
          5870 => x"56",
          5871 => x"38",
          5872 => x"76",
          5873 => x"9c",
          5874 => x"98",
          5875 => x"84",
          5876 => x"18",
          5877 => x"80",
          5878 => x"12",
          5879 => x"7a",
          5880 => x"76",
          5881 => x"89",
          5882 => x"2e",
          5883 => x"94",
          5884 => x"38",
          5885 => x"80",
          5886 => x"75",
          5887 => x"81",
          5888 => x"7a",
          5889 => x"70",
          5890 => x"74",
          5891 => x"53",
          5892 => x"56",
          5893 => x"08",
          5894 => x"06",
          5895 => x"79",
          5896 => x"52",
          5897 => x"84",
          5898 => x"0b",
          5899 => x"bb",
          5900 => x"17",
          5901 => x"5a",
          5902 => x"08",
          5903 => x"09",
          5904 => x"18",
          5905 => x"18",
          5906 => x"2e",
          5907 => x"75",
          5908 => x"39",
          5909 => x"bb",
          5910 => x"52",
          5911 => x"bb",
          5912 => x"16",
          5913 => x"bb",
          5914 => x"81",
          5915 => x"fb",
          5916 => x"bc",
          5917 => x"bb",
          5918 => x"bb",
          5919 => x"84",
          5920 => x"98",
          5921 => x"91",
          5922 => x"0c",
          5923 => x"7c",
          5924 => x"38",
          5925 => x"8d",
          5926 => x"84",
          5927 => x"08",
          5928 => x"74",
          5929 => x"3d",
          5930 => x"75",
          5931 => x"84",
          5932 => x"d1",
          5933 => x"59",
          5934 => x"16",
          5935 => x"54",
          5936 => x"16",
          5937 => x"71",
          5938 => x"5d",
          5939 => x"38",
          5940 => x"18",
          5941 => x"51",
          5942 => x"08",
          5943 => x"80",
          5944 => x"fe",
          5945 => x"fe",
          5946 => x"33",
          5947 => x"7a",
          5948 => x"bc",
          5949 => x"54",
          5950 => x"53",
          5951 => x"52",
          5952 => x"22",
          5953 => x"2e",
          5954 => x"84",
          5955 => x"84",
          5956 => x"33",
          5957 => x"84",
          5958 => x"71",
          5959 => x"3d",
          5960 => x"74",
          5961 => x"73",
          5962 => x"72",
          5963 => x"84",
          5964 => x"81",
          5965 => x"53",
          5966 => x"80",
          5967 => x"9e",
          5968 => x"84",
          5969 => x"84",
          5970 => x"74",
          5971 => x"74",
          5972 => x"84",
          5973 => x"07",
          5974 => x"55",
          5975 => x"8a",
          5976 => x"52",
          5977 => x"74",
          5978 => x"84",
          5979 => x"07",
          5980 => x"55",
          5981 => x"51",
          5982 => x"08",
          5983 => x"04",
          5984 => x"3f",
          5985 => x"72",
          5986 => x"56",
          5987 => x"57",
          5988 => x"3d",
          5989 => x"84",
          5990 => x"2e",
          5991 => x"95",
          5992 => x"ff",
          5993 => x"55",
          5994 => x"80",
          5995 => x"58",
          5996 => x"2e",
          5997 => x"b1",
          5998 => x"95",
          5999 => x"84",
          6000 => x"0d",
          6001 => x"3d",
          6002 => x"aa",
          6003 => x"bb",
          6004 => x"74",
          6005 => x"13",
          6006 => x"26",
          6007 => x"bb",
          6008 => x"bb",
          6009 => x"81",
          6010 => x"08",
          6011 => x"77",
          6012 => x"5c",
          6013 => x"82",
          6014 => x"5d",
          6015 => x"53",
          6016 => x"fe",
          6017 => x"80",
          6018 => x"79",
          6019 => x"7d",
          6020 => x"82",
          6021 => x"05",
          6022 => x"90",
          6023 => x"33",
          6024 => x"71",
          6025 => x"70",
          6026 => x"84",
          6027 => x"43",
          6028 => x"40",
          6029 => x"7f",
          6030 => x"33",
          6031 => x"79",
          6032 => x"04",
          6033 => x"17",
          6034 => x"fe",
          6035 => x"84",
          6036 => x"08",
          6037 => x"18",
          6038 => x"55",
          6039 => x"38",
          6040 => x"09",
          6041 => x"b4",
          6042 => x"7c",
          6043 => x"d1",
          6044 => x"77",
          6045 => x"77",
          6046 => x"84",
          6047 => x"bb",
          6048 => x"84",
          6049 => x"84",
          6050 => x"18",
          6051 => x"08",
          6052 => x"7a",
          6053 => x"07",
          6054 => x"39",
          6055 => x"71",
          6056 => x"70",
          6057 => x"06",
          6058 => x"5f",
          6059 => x"39",
          6060 => x"58",
          6061 => x"0c",
          6062 => x"84",
          6063 => x"58",
          6064 => x"58",
          6065 => x"77",
          6066 => x"75",
          6067 => x"86",
          6068 => x"79",
          6069 => x"74",
          6070 => x"33",
          6071 => x"33",
          6072 => x"87",
          6073 => x"94",
          6074 => x"27",
          6075 => x"88",
          6076 => x"75",
          6077 => x"26",
          6078 => x"88",
          6079 => x"0c",
          6080 => x"19",
          6081 => x"5a",
          6082 => x"9c",
          6083 => x"81",
          6084 => x"3f",
          6085 => x"90",
          6086 => x"76",
          6087 => x"3d",
          6088 => x"80",
          6089 => x"ff",
          6090 => x"84",
          6091 => x"38",
          6092 => x"e8",
          6093 => x"82",
          6094 => x"51",
          6095 => x"08",
          6096 => x"11",
          6097 => x"75",
          6098 => x"18",
          6099 => x"74",
          6100 => x"26",
          6101 => x"33",
          6102 => x"84",
          6103 => x"38",
          6104 => x"39",
          6105 => x"74",
          6106 => x"a2",
          6107 => x"fe",
          6108 => x"ff",
          6109 => x"08",
          6110 => x"ae",
          6111 => x"9c",
          6112 => x"bb",
          6113 => x"59",
          6114 => x"08",
          6115 => x"08",
          6116 => x"75",
          6117 => x"52",
          6118 => x"bb",
          6119 => x"80",
          6120 => x"fd",
          6121 => x"84",
          6122 => x"38",
          6123 => x"dc",
          6124 => x"81",
          6125 => x"51",
          6126 => x"08",
          6127 => x"11",
          6128 => x"75",
          6129 => x"0c",
          6130 => x"84",
          6131 => x"ff",
          6132 => x"18",
          6133 => x"fe",
          6134 => x"5a",
          6135 => x"39",
          6136 => x"74",
          6137 => x"39",
          6138 => x"fd",
          6139 => x"19",
          6140 => x"0b",
          6141 => x"39",
          6142 => x"39",
          6143 => x"0d",
          6144 => x"52",
          6145 => x"84",
          6146 => x"08",
          6147 => x"84",
          6148 => x"a8",
          6149 => x"59",
          6150 => x"08",
          6151 => x"02",
          6152 => x"81",
          6153 => x"38",
          6154 => x"c4",
          6155 => x"81",
          6156 => x"b4",
          6157 => x"33",
          6158 => x"73",
          6159 => x"83",
          6160 => x"81",
          6161 => x"38",
          6162 => x"ff",
          6163 => x"bb",
          6164 => x"55",
          6165 => x"08",
          6166 => x"38",
          6167 => x"ff",
          6168 => x"56",
          6169 => x"0b",
          6170 => x"04",
          6171 => x"98",
          6172 => x"5d",
          6173 => x"84",
          6174 => x"84",
          6175 => x"a8",
          6176 => x"2e",
          6177 => x"ff",
          6178 => x"56",
          6179 => x"38",
          6180 => x"56",
          6181 => x"80",
          6182 => x"55",
          6183 => x"08",
          6184 => x"75",
          6185 => x"94",
          6186 => x"84",
          6187 => x"5d",
          6188 => x"17",
          6189 => x"17",
          6190 => x"09",
          6191 => x"75",
          6192 => x"51",
          6193 => x"08",
          6194 => x"58",
          6195 => x"ab",
          6196 => x"34",
          6197 => x"08",
          6198 => x"78",
          6199 => x"84",
          6200 => x"2e",
          6201 => x"81",
          6202 => x"c8",
          6203 => x"7c",
          6204 => x"c9",
          6205 => x"7a",
          6206 => x"84",
          6207 => x"17",
          6208 => x"84",
          6209 => x"27",
          6210 => x"74",
          6211 => x"38",
          6212 => x"08",
          6213 => x"51",
          6214 => x"c5",
          6215 => x"e1",
          6216 => x"9d",
          6217 => x"bb",
          6218 => x"84",
          6219 => x"38",
          6220 => x"cb",
          6221 => x"fe",
          6222 => x"b3",
          6223 => x"19",
          6224 => x"ff",
          6225 => x"84",
          6226 => x"18",
          6227 => x"a1",
          6228 => x"56",
          6229 => x"56",
          6230 => x"39",
          6231 => x"ff",
          6232 => x"b2",
          6233 => x"84",
          6234 => x"75",
          6235 => x"04",
          6236 => x"52",
          6237 => x"84",
          6238 => x"38",
          6239 => x"3d",
          6240 => x"2e",
          6241 => x"f3",
          6242 => x"56",
          6243 => x"7d",
          6244 => x"5d",
          6245 => x"08",
          6246 => x"83",
          6247 => x"81",
          6248 => x"08",
          6249 => x"c9",
          6250 => x"12",
          6251 => x"38",
          6252 => x"5a",
          6253 => x"38",
          6254 => x"19",
          6255 => x"0c",
          6256 => x"55",
          6257 => x"ff",
          6258 => x"8a",
          6259 => x"f9",
          6260 => x"52",
          6261 => x"3f",
          6262 => x"81",
          6263 => x"84",
          6264 => x"b8",
          6265 => x"58",
          6266 => x"bb",
          6267 => x"08",
          6268 => x"18",
          6269 => x"27",
          6270 => x"7a",
          6271 => x"38",
          6272 => x"08",
          6273 => x"51",
          6274 => x"81",
          6275 => x"7c",
          6276 => x"08",
          6277 => x"51",
          6278 => x"08",
          6279 => x"fd",
          6280 => x"2e",
          6281 => x"ff",
          6282 => x"52",
          6283 => x"bb",
          6284 => x"08",
          6285 => x"59",
          6286 => x"94",
          6287 => x"5c",
          6288 => x"7a",
          6289 => x"84",
          6290 => x"22",
          6291 => x"81",
          6292 => x"fe",
          6293 => x"56",
          6294 => x"ff",
          6295 => x"ae",
          6296 => x"0b",
          6297 => x"80",
          6298 => x"34",
          6299 => x"cc",
          6300 => x"83",
          6301 => x"d2",
          6302 => x"80",
          6303 => x"83",
          6304 => x"0b",
          6305 => x"56",
          6306 => x"70",
          6307 => x"75",
          6308 => x"d9",
          6309 => x"ff",
          6310 => x"17",
          6311 => x"f3",
          6312 => x"2e",
          6313 => x"83",
          6314 => x"3f",
          6315 => x"84",
          6316 => x"bb",
          6317 => x"84",
          6318 => x"17",
          6319 => x"7d",
          6320 => x"77",
          6321 => x"7c",
          6322 => x"38",
          6323 => x"7d",
          6324 => x"51",
          6325 => x"08",
          6326 => x"3d",
          6327 => x"80",
          6328 => x"76",
          6329 => x"7b",
          6330 => x"34",
          6331 => x"17",
          6332 => x"1a",
          6333 => x"39",
          6334 => x"34",
          6335 => x"34",
          6336 => x"7d",
          6337 => x"51",
          6338 => x"08",
          6339 => x"b3",
          6340 => x"5f",
          6341 => x"81",
          6342 => x"56",
          6343 => x"ed",
          6344 => x"82",
          6345 => x"b2",
          6346 => x"bb",
          6347 => x"80",
          6348 => x"0c",
          6349 => x"0c",
          6350 => x"52",
          6351 => x"84",
          6352 => x"38",
          6353 => x"06",
          6354 => x"0b",
          6355 => x"55",
          6356 => x"70",
          6357 => x"74",
          6358 => x"7a",
          6359 => x"57",
          6360 => x"ff",
          6361 => x"08",
          6362 => x"84",
          6363 => x"08",
          6364 => x"2e",
          6365 => x"84",
          6366 => x"d0",
          6367 => x"58",
          6368 => x"78",
          6369 => x"78",
          6370 => x"08",
          6371 => x"5e",
          6372 => x"5c",
          6373 => x"ff",
          6374 => x"26",
          6375 => x"06",
          6376 => x"99",
          6377 => x"ff",
          6378 => x"2a",
          6379 => x"06",
          6380 => x"7a",
          6381 => x"2a",
          6382 => x"2e",
          6383 => x"5c",
          6384 => x"08",
          6385 => x"83",
          6386 => x"82",
          6387 => x"b2",
          6388 => x"bb",
          6389 => x"fd",
          6390 => x"3d",
          6391 => x"38",
          6392 => x"bb",
          6393 => x"fd",
          6394 => x"19",
          6395 => x"56",
          6396 => x"75",
          6397 => x"5a",
          6398 => x"33",
          6399 => x"84",
          6400 => x"38",
          6401 => x"34",
          6402 => x"8b",
          6403 => x"57",
          6404 => x"a7",
          6405 => x"7f",
          6406 => x"88",
          6407 => x"57",
          6408 => x"16",
          6409 => x"75",
          6410 => x"22",
          6411 => x"57",
          6412 => x"75",
          6413 => x"2e",
          6414 => x"83",
          6415 => x"17",
          6416 => x"aa",
          6417 => x"85",
          6418 => x"18",
          6419 => x"56",
          6420 => x"33",
          6421 => x"bb",
          6422 => x"5d",
          6423 => x"88",
          6424 => x"76",
          6425 => x"06",
          6426 => x"80",
          6427 => x"75",
          6428 => x"0b",
          6429 => x"08",
          6430 => x"ff",
          6431 => x"fe",
          6432 => x"55",
          6433 => x"b8",
          6434 => x"5a",
          6435 => x"83",
          6436 => x"2e",
          6437 => x"54",
          6438 => x"33",
          6439 => x"84",
          6440 => x"81",
          6441 => x"77",
          6442 => x"7a",
          6443 => x"19",
          6444 => x"78",
          6445 => x"84",
          6446 => x"2e",
          6447 => x"2e",
          6448 => x"db",
          6449 => x"84",
          6450 => x"b1",
          6451 => x"84",
          6452 => x"33",
          6453 => x"90",
          6454 => x"fd",
          6455 => x"2e",
          6456 => x"80",
          6457 => x"84",
          6458 => x"b4",
          6459 => x"33",
          6460 => x"84",
          6461 => x"06",
          6462 => x"83",
          6463 => x"08",
          6464 => x"74",
          6465 => x"82",
          6466 => x"81",
          6467 => x"16",
          6468 => x"52",
          6469 => x"3f",
          6470 => x"b4",
          6471 => x"81",
          6472 => x"3f",
          6473 => x"c9",
          6474 => x"34",
          6475 => x"84",
          6476 => x"18",
          6477 => x"33",
          6478 => x"fc",
          6479 => x"a0",
          6480 => x"17",
          6481 => x"5c",
          6482 => x"80",
          6483 => x"e3",
          6484 => x"3d",
          6485 => x"a3",
          6486 => x"84",
          6487 => x"75",
          6488 => x"04",
          6489 => x"05",
          6490 => x"84",
          6491 => x"38",
          6492 => x"06",
          6493 => x"a7",
          6494 => x"71",
          6495 => x"57",
          6496 => x"81",
          6497 => x"e2",
          6498 => x"bb",
          6499 => x"3d",
          6500 => x"cc",
          6501 => x"92",
          6502 => x"bb",
          6503 => x"84",
          6504 => x"78",
          6505 => x"51",
          6506 => x"08",
          6507 => x"02",
          6508 => x"56",
          6509 => x"18",
          6510 => x"07",
          6511 => x"76",
          6512 => x"76",
          6513 => x"76",
          6514 => x"78",
          6515 => x"51",
          6516 => x"08",
          6517 => x"04",
          6518 => x"80",
          6519 => x"3d",
          6520 => x"84",
          6521 => x"84",
          6522 => x"56",
          6523 => x"70",
          6524 => x"38",
          6525 => x"56",
          6526 => x"81",
          6527 => x"2e",
          6528 => x"58",
          6529 => x"2e",
          6530 => x"5a",
          6531 => x"81",
          6532 => x"16",
          6533 => x"82",
          6534 => x"85",
          6535 => x"17",
          6536 => x"70",
          6537 => x"83",
          6538 => x"84",
          6539 => x"b8",
          6540 => x"71",
          6541 => x"14",
          6542 => x"33",
          6543 => x"57",
          6544 => x"9a",
          6545 => x"80",
          6546 => x"f4",
          6547 => x"84",
          6548 => x"38",
          6549 => x"b8",
          6550 => x"b0",
          6551 => x"b8",
          6552 => x"5b",
          6553 => x"bb",
          6554 => x"fe",
          6555 => x"17",
          6556 => x"31",
          6557 => x"a0",
          6558 => x"16",
          6559 => x"06",
          6560 => x"08",
          6561 => x"81",
          6562 => x"79",
          6563 => x"52",
          6564 => x"3f",
          6565 => x"8d",
          6566 => x"51",
          6567 => x"08",
          6568 => x"38",
          6569 => x"08",
          6570 => x"19",
          6571 => x"75",
          6572 => x"ec",
          6573 => x"76",
          6574 => x"ff",
          6575 => x"58",
          6576 => x"39",
          6577 => x"0d",
          6578 => x"52",
          6579 => x"84",
          6580 => x"08",
          6581 => x"7d",
          6582 => x"58",
          6583 => x"74",
          6584 => x"ff",
          6585 => x"27",
          6586 => x"5c",
          6587 => x"57",
          6588 => x"0c",
          6589 => x"38",
          6590 => x"52",
          6591 => x"3f",
          6592 => x"06",
          6593 => x"83",
          6594 => x"70",
          6595 => x"80",
          6596 => x"77",
          6597 => x"70",
          6598 => x"80",
          6599 => x"81",
          6600 => x"59",
          6601 => x"27",
          6602 => x"96",
          6603 => x"76",
          6604 => x"05",
          6605 => x"70",
          6606 => x"3d",
          6607 => x"5b",
          6608 => x"d1",
          6609 => x"76",
          6610 => x"2e",
          6611 => x"16",
          6612 => x"09",
          6613 => x"79",
          6614 => x"52",
          6615 => x"9d",
          6616 => x"bb",
          6617 => x"56",
          6618 => x"0d",
          6619 => x"e7",
          6620 => x"ff",
          6621 => x"56",
          6622 => x"0d",
          6623 => x"c3",
          6624 => x"a7",
          6625 => x"bb",
          6626 => x"2e",
          6627 => x"57",
          6628 => x"76",
          6629 => x"55",
          6630 => x"83",
          6631 => x"3f",
          6632 => x"ff",
          6633 => x"38",
          6634 => x"84",
          6635 => x"ee",
          6636 => x"e6",
          6637 => x"58",
          6638 => x"08",
          6639 => x"09",
          6640 => x"84",
          6641 => x"08",
          6642 => x"2e",
          6643 => x"79",
          6644 => x"81",
          6645 => x"18",
          6646 => x"bb",
          6647 => x"57",
          6648 => x"57",
          6649 => x"70",
          6650 => x"2e",
          6651 => x"25",
          6652 => x"81",
          6653 => x"2e",
          6654 => x"ef",
          6655 => x"84",
          6656 => x"38",
          6657 => x"38",
          6658 => x"6c",
          6659 => x"58",
          6660 => x"6b",
          6661 => x"6c",
          6662 => x"05",
          6663 => x"34",
          6664 => x"eb",
          6665 => x"76",
          6666 => x"55",
          6667 => x"5a",
          6668 => x"83",
          6669 => x"3f",
          6670 => x"39",
          6671 => x"b4",
          6672 => x"33",
          6673 => x"84",
          6674 => x"c3",
          6675 => x"34",
          6676 => x"5c",
          6677 => x"82",
          6678 => x"38",
          6679 => x"39",
          6680 => x"ee",
          6681 => x"84",
          6682 => x"38",
          6683 => x"78",
          6684 => x"39",
          6685 => x"08",
          6686 => x"51",
          6687 => x"f2",
          6688 => x"80",
          6689 => x"56",
          6690 => x"55",
          6691 => x"54",
          6692 => x"22",
          6693 => x"2e",
          6694 => x"75",
          6695 => x"75",
          6696 => x"a2",
          6697 => x"90",
          6698 => x"56",
          6699 => x"7e",
          6700 => x"55",
          6701 => x"bc",
          6702 => x"70",
          6703 => x"08",
          6704 => x"5f",
          6705 => x"9c",
          6706 => x"58",
          6707 => x"52",
          6708 => x"15",
          6709 => x"26",
          6710 => x"08",
          6711 => x"84",
          6712 => x"bb",
          6713 => x"59",
          6714 => x"2e",
          6715 => x"75",
          6716 => x"3d",
          6717 => x"0c",
          6718 => x"51",
          6719 => x"08",
          6720 => x"73",
          6721 => x"7b",
          6722 => x"56",
          6723 => x"18",
          6724 => x"73",
          6725 => x"96",
          6726 => x"bb",
          6727 => x"19",
          6728 => x"38",
          6729 => x"80",
          6730 => x"0c",
          6731 => x"80",
          6732 => x"9c",
          6733 => x"58",
          6734 => x"76",
          6735 => x"33",
          6736 => x"75",
          6737 => x"97",
          6738 => x"39",
          6739 => x"fe",
          6740 => x"39",
          6741 => x"a3",
          6742 => x"05",
          6743 => x"ff",
          6744 => x"40",
          6745 => x"70",
          6746 => x"56",
          6747 => x"74",
          6748 => x"38",
          6749 => x"24",
          6750 => x"e2",
          6751 => x"80",
          6752 => x"16",
          6753 => x"f9",
          6754 => x"79",
          6755 => x"84",
          6756 => x"5d",
          6757 => x"75",
          6758 => x"7f",
          6759 => x"53",
          6760 => x"3f",
          6761 => x"6d",
          6762 => x"74",
          6763 => x"ff",
          6764 => x"38",
          6765 => x"7f",
          6766 => x"0a",
          6767 => x"06",
          6768 => x"2a",
          6769 => x"2b",
          6770 => x"2e",
          6771 => x"25",
          6772 => x"83",
          6773 => x"38",
          6774 => x"51",
          6775 => x"bb",
          6776 => x"ff",
          6777 => x"71",
          6778 => x"77",
          6779 => x"82",
          6780 => x"83",
          6781 => x"2e",
          6782 => x"11",
          6783 => x"71",
          6784 => x"72",
          6785 => x"83",
          6786 => x"33",
          6787 => x"81",
          6788 => x"75",
          6789 => x"42",
          6790 => x"4e",
          6791 => x"78",
          6792 => x"82",
          6793 => x"26",
          6794 => x"81",
          6795 => x"f9",
          6796 => x"2e",
          6797 => x"83",
          6798 => x"46",
          6799 => x"c2",
          6800 => x"57",
          6801 => x"58",
          6802 => x"26",
          6803 => x"10",
          6804 => x"74",
          6805 => x"ee",
          6806 => x"f4",
          6807 => x"05",
          6808 => x"26",
          6809 => x"08",
          6810 => x"11",
          6811 => x"83",
          6812 => x"a0",
          6813 => x"66",
          6814 => x"31",
          6815 => x"89",
          6816 => x"29",
          6817 => x"79",
          6818 => x"7d",
          6819 => x"56",
          6820 => x"08",
          6821 => x"62",
          6822 => x"38",
          6823 => x"08",
          6824 => x"38",
          6825 => x"89",
          6826 => x"8b",
          6827 => x"3d",
          6828 => x"4e",
          6829 => x"84",
          6830 => x"0c",
          6831 => x"ff",
          6832 => x"91",
          6833 => x"d0",
          6834 => x"b2",
          6835 => x"5c",
          6836 => x"81",
          6837 => x"58",
          6838 => x"62",
          6839 => x"81",
          6840 => x"45",
          6841 => x"70",
          6842 => x"70",
          6843 => x"09",
          6844 => x"38",
          6845 => x"07",
          6846 => x"7a",
          6847 => x"84",
          6848 => x"98",
          6849 => x"3d",
          6850 => x"fe",
          6851 => x"84",
          6852 => x"77",
          6853 => x"75",
          6854 => x"57",
          6855 => x"7f",
          6856 => x"fa",
          6857 => x"38",
          6858 => x"95",
          6859 => x"67",
          6860 => x"70",
          6861 => x"84",
          6862 => x"38",
          6863 => x"80",
          6864 => x"76",
          6865 => x"84",
          6866 => x"81",
          6867 => x"27",
          6868 => x"57",
          6869 => x"57",
          6870 => x"34",
          6871 => x"61",
          6872 => x"70",
          6873 => x"05",
          6874 => x"38",
          6875 => x"82",
          6876 => x"05",
          6877 => x"6a",
          6878 => x"5c",
          6879 => x"90",
          6880 => x"5a",
          6881 => x"9e",
          6882 => x"05",
          6883 => x"26",
          6884 => x"06",
          6885 => x"88",
          6886 => x"f8",
          6887 => x"05",
          6888 => x"61",
          6889 => x"34",
          6890 => x"2a",
          6891 => x"90",
          6892 => x"7e",
          6893 => x"bb",
          6894 => x"83",
          6895 => x"05",
          6896 => x"61",
          6897 => x"05",
          6898 => x"74",
          6899 => x"4b",
          6900 => x"61",
          6901 => x"34",
          6902 => x"59",
          6903 => x"33",
          6904 => x"15",
          6905 => x"05",
          6906 => x"ff",
          6907 => x"54",
          6908 => x"c6",
          6909 => x"08",
          6910 => x"83",
          6911 => x"55",
          6912 => x"ff",
          6913 => x"41",
          6914 => x"87",
          6915 => x"83",
          6916 => x"88",
          6917 => x"81",
          6918 => x"78",
          6919 => x"98",
          6920 => x"65",
          6921 => x"59",
          6922 => x"51",
          6923 => x"08",
          6924 => x"55",
          6925 => x"ff",
          6926 => x"77",
          6927 => x"7f",
          6928 => x"89",
          6929 => x"38",
          6930 => x"83",
          6931 => x"60",
          6932 => x"84",
          6933 => x"1b",
          6934 => x"38",
          6935 => x"86",
          6936 => x"38",
          6937 => x"81",
          6938 => x"2a",
          6939 => x"84",
          6940 => x"81",
          6941 => x"f4",
          6942 => x"6b",
          6943 => x"67",
          6944 => x"67",
          6945 => x"34",
          6946 => x"80",
          6947 => x"f7",
          6948 => x"84",
          6949 => x"57",
          6950 => x"84",
          6951 => x"83",
          6952 => x"05",
          6953 => x"84",
          6954 => x"34",
          6955 => x"88",
          6956 => x"34",
          6957 => x"cc",
          6958 => x"61",
          6959 => x"53",
          6960 => x"3f",
          6961 => x"c9",
          6962 => x"fe",
          6963 => x"84",
          6964 => x"08",
          6965 => x"84",
          6966 => x"e4",
          6967 => x"f6",
          6968 => x"2a",
          6969 => x"56",
          6970 => x"77",
          6971 => x"77",
          6972 => x"58",
          6973 => x"27",
          6974 => x"f5",
          6975 => x"10",
          6976 => x"5c",
          6977 => x"08",
          6978 => x"ff",
          6979 => x"8e",
          6980 => x"08",
          6981 => x"7a",
          6982 => x"7a",
          6983 => x"39",
          6984 => x"f8",
          6985 => x"75",
          6986 => x"49",
          6987 => x"2a",
          6988 => x"98",
          6989 => x"f9",
          6990 => x"34",
          6991 => x"61",
          6992 => x"80",
          6993 => x"34",
          6994 => x"05",
          6995 => x"a6",
          6996 => x"61",
          6997 => x"34",
          6998 => x"ae",
          6999 => x"81",
          7000 => x"05",
          7001 => x"61",
          7002 => x"c0",
          7003 => x"34",
          7004 => x"e0",
          7005 => x"58",
          7006 => x"ff",
          7007 => x"38",
          7008 => x"70",
          7009 => x"74",
          7010 => x"80",
          7011 => x"92",
          7012 => x"f4",
          7013 => x"42",
          7014 => x"54",
          7015 => x"79",
          7016 => x"39",
          7017 => x"3d",
          7018 => x"61",
          7019 => x"05",
          7020 => x"4c",
          7021 => x"05",
          7022 => x"61",
          7023 => x"34",
          7024 => x"89",
          7025 => x"8f",
          7026 => x"76",
          7027 => x"51",
          7028 => x"56",
          7029 => x"34",
          7030 => x"5c",
          7031 => x"34",
          7032 => x"05",
          7033 => x"05",
          7034 => x"f2",
          7035 => x"61",
          7036 => x"83",
          7037 => x"e7",
          7038 => x"61",
          7039 => x"59",
          7040 => x"90",
          7041 => x"34",
          7042 => x"eb",
          7043 => x"34",
          7044 => x"61",
          7045 => x"ef",
          7046 => x"aa",
          7047 => x"60",
          7048 => x"81",
          7049 => x"51",
          7050 => x"55",
          7051 => x"61",
          7052 => x"5a",
          7053 => x"8d",
          7054 => x"81",
          7055 => x"cc",
          7056 => x"9e",
          7057 => x"2e",
          7058 => x"58",
          7059 => x"86",
          7060 => x"76",
          7061 => x"55",
          7062 => x"0d",
          7063 => x"05",
          7064 => x"2e",
          7065 => x"80",
          7066 => x"77",
          7067 => x"34",
          7068 => x"38",
          7069 => x"18",
          7070 => x"fc",
          7071 => x"76",
          7072 => x"7a",
          7073 => x"2a",
          7074 => x"88",
          7075 => x"8d",
          7076 => x"a3",
          7077 => x"05",
          7078 => x"77",
          7079 => x"58",
          7080 => x"a1",
          7081 => x"80",
          7082 => x"80",
          7083 => x"56",
          7084 => x"74",
          7085 => x"0c",
          7086 => x"80",
          7087 => x"ac",
          7088 => x"76",
          7089 => x"bb",
          7090 => x"ba",
          7091 => x"9f",
          7092 => x"11",
          7093 => x"08",
          7094 => x"32",
          7095 => x"70",
          7096 => x"39",
          7097 => x"ff",
          7098 => x"9f",
          7099 => x"02",
          7100 => x"80",
          7101 => x"72",
          7102 => x"bb",
          7103 => x"ff",
          7104 => x"2e",
          7105 => x"2e",
          7106 => x"72",
          7107 => x"83",
          7108 => x"ff",
          7109 => x"c8",
          7110 => x"81",
          7111 => x"bb",
          7112 => x"fe",
          7113 => x"84",
          7114 => x"53",
          7115 => x"53",
          7116 => x"0d",
          7117 => x"06",
          7118 => x"38",
          7119 => x"22",
          7120 => x"0d",
          7121 => x"83",
          7122 => x"83",
          7123 => x"56",
          7124 => x"74",
          7125 => x"30",
          7126 => x"54",
          7127 => x"70",
          7128 => x"2a",
          7129 => x"52",
          7130 => x"cf",
          7131 => x"05",
          7132 => x"25",
          7133 => x"70",
          7134 => x"84",
          7135 => x"83",
          7136 => x"88",
          7137 => x"ca",
          7138 => x"a0",
          7139 => x"51",
          7140 => x"70",
          7141 => x"39",
          7142 => x"57",
          7143 => x"ff",
          7144 => x"16",
          7145 => x"d0",
          7146 => x"06",
          7147 => x"83",
          7148 => x"39",
          7149 => x"31",
          7150 => x"55",
          7151 => x"75",
          7152 => x"39",
          7153 => x"ff",
          7154 => x"ff",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"00",
          7372 => x"00",
          7373 => x"00",
          7374 => x"00",
          7375 => x"00",
          7376 => x"00",
          7377 => x"00",
          7378 => x"00",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"00",
          7383 => x"00",
          7384 => x"00",
          7385 => x"00",
          7386 => x"00",
          7387 => x"00",
          7388 => x"00",
          7389 => x"00",
          7390 => x"00",
          7391 => x"64",
          7392 => x"64",
          7393 => x"66",
          7394 => x"66",
          7395 => x"66",
          7396 => x"6d",
          7397 => x"6d",
          7398 => x"6d",
          7399 => x"6d",
          7400 => x"6d",
          7401 => x"6d",
          7402 => x"68",
          7403 => x"68",
          7404 => x"00",
          7405 => x"72",
          7406 => x"72",
          7407 => x"69",
          7408 => x"74",
          7409 => x"63",
          7410 => x"74",
          7411 => x"6d",
          7412 => x"6b",
          7413 => x"65",
          7414 => x"6f",
          7415 => x"72",
          7416 => x"6d",
          7417 => x"6e",
          7418 => x"2e",
          7419 => x"6d",
          7420 => x"6e",
          7421 => x"00",
          7422 => x"66",
          7423 => x"20",
          7424 => x"00",
          7425 => x"20",
          7426 => x"65",
          7427 => x"6f",
          7428 => x"72",
          7429 => x"61",
          7430 => x"2e",
          7431 => x"61",
          7432 => x"65",
          7433 => x"6f",
          7434 => x"65",
          7435 => x"73",
          7436 => x"6e",
          7437 => x"73",
          7438 => x"20",
          7439 => x"62",
          7440 => x"44",
          7441 => x"6d",
          7442 => x"69",
          7443 => x"00",
          7444 => x"73",
          7445 => x"70",
          7446 => x"64",
          7447 => x"20",
          7448 => x"69",
          7449 => x"00",
          7450 => x"20",
          7451 => x"20",
          7452 => x"00",
          7453 => x"73",
          7454 => x"64",
          7455 => x"6c",
          7456 => x"6e",
          7457 => x"4e",
          7458 => x"66",
          7459 => x"4e",
          7460 => x"66",
          7461 => x"44",
          7462 => x"20",
          7463 => x"49",
          7464 => x"20",
          7465 => x"44",
          7466 => x"6f",
          7467 => x"65",
          7468 => x"0a",
          7469 => x"65",
          7470 => x"20",
          7471 => x"65",
          7472 => x"00",
          7473 => x"00",
          7474 => x"58",
          7475 => x"25",
          7476 => x"20",
          7477 => x"20",
          7478 => x"00",
          7479 => x"20",
          7480 => x"7a",
          7481 => x"73",
          7482 => x"37",
          7483 => x"76",
          7484 => x"20",
          7485 => x"76",
          7486 => x"25",
          7487 => x"0a",
          7488 => x"20",
          7489 => x"20",
          7490 => x"20",
          7491 => x"20",
          7492 => x"30",
          7493 => x"20",
          7494 => x"41",
          7495 => x"20",
          7496 => x"20",
          7497 => x"30",
          7498 => x"5a",
          7499 => x"72",
          7500 => x"6e",
          7501 => x"55",
          7502 => x"20",
          7503 => x"70",
          7504 => x"31",
          7505 => x"65",
          7506 => x"55",
          7507 => x"20",
          7508 => x"70",
          7509 => x"30",
          7510 => x"65",
          7511 => x"49",
          7512 => x"20",
          7513 => x"70",
          7514 => x"4c",
          7515 => x"65",
          7516 => x"50",
          7517 => x"72",
          7518 => x"54",
          7519 => x"74",
          7520 => x"53",
          7521 => x"75",
          7522 => x"2e",
          7523 => x"6c",
          7524 => x"65",
          7525 => x"61",
          7526 => x"2e",
          7527 => x"7a",
          7528 => x"68",
          7529 => x"65",
          7530 => x"69",
          7531 => x"20",
          7532 => x"20",
          7533 => x"73",
          7534 => x"6d",
          7535 => x"2e",
          7536 => x"25",
          7537 => x"30",
          7538 => x"63",
          7539 => x"00",
          7540 => x"62",
          7541 => x"25",
          7542 => x"00",
          7543 => x"20",
          7544 => x"6e",
          7545 => x"52",
          7546 => x"6e",
          7547 => x"63",
          7548 => x"2e",
          7549 => x"69",
          7550 => x"20",
          7551 => x"20",
          7552 => x"43",
          7553 => x"75",
          7554 => x"64",
          7555 => x"0a",
          7556 => x"75",
          7557 => x"64",
          7558 => x"6c",
          7559 => x"25",
          7560 => x"38",
          7561 => x"25",
          7562 => x"34",
          7563 => x"61",
          7564 => x"00",
          7565 => x"78",
          7566 => x"3e",
          7567 => x"30",
          7568 => x"43",
          7569 => x"2e",
          7570 => x"58",
          7571 => x"43",
          7572 => x"2e",
          7573 => x"44",
          7574 => x"6f",
          7575 => x"70",
          7576 => x"25",
          7577 => x"73",
          7578 => x"72",
          7579 => x"73",
          7580 => x"6e",
          7581 => x"63",
          7582 => x"6d",
          7583 => x"3f",
          7584 => x"64",
          7585 => x"25",
          7586 => x"25",
          7587 => x"43",
          7588 => x"61",
          7589 => x"3a",
          7590 => x"73",
          7591 => x"65",
          7592 => x"41",
          7593 => x"73",
          7594 => x"43",
          7595 => x"74",
          7596 => x"20",
          7597 => x"20",
          7598 => x"00",
          7599 => x"43",
          7600 => x"72",
          7601 => x"20",
          7602 => x"20",
          7603 => x"00",
          7604 => x"53",
          7605 => x"61",
          7606 => x"65",
          7607 => x"20",
          7608 => x"00",
          7609 => x"3a",
          7610 => x"5a",
          7611 => x"20",
          7612 => x"20",
          7613 => x"20",
          7614 => x"00",
          7615 => x"53",
          7616 => x"6c",
          7617 => x"71",
          7618 => x"20",
          7619 => x"34",
          7620 => x"20",
          7621 => x"62",
          7622 => x"41",
          7623 => x"20",
          7624 => x"64",
          7625 => x"7a",
          7626 => x"53",
          7627 => x"6f",
          7628 => x"20",
          7629 => x"20",
          7630 => x"34",
          7631 => x"20",
          7632 => x"20",
          7633 => x"20",
          7634 => x"4c",
          7635 => x"57",
          7636 => x"20",
          7637 => x"42",
          7638 => x"00",
          7639 => x"49",
          7640 => x"4c",
          7641 => x"65",
          7642 => x"29",
          7643 => x"54",
          7644 => x"20",
          7645 => x"73",
          7646 => x"29",
          7647 => x"53",
          7648 => x"20",
          7649 => x"65",
          7650 => x"29",
          7651 => x"52",
          7652 => x"20",
          7653 => x"25",
          7654 => x"20",
          7655 => x"20",
          7656 => x"30",
          7657 => x"29",
          7658 => x"49",
          7659 => x"4d",
          7660 => x"25",
          7661 => x"20",
          7662 => x"4d",
          7663 => x"30",
          7664 => x"29",
          7665 => x"57",
          7666 => x"20",
          7667 => x"25",
          7668 => x"20",
          7669 => x"6f",
          7670 => x"67",
          7671 => x"6f",
          7672 => x"00",
          7673 => x"6c",
          7674 => x"75",
          7675 => x"00",
          7676 => x"00",
          7677 => x"00",
          7678 => x"01",
          7679 => x"00",
          7680 => x"00",
          7681 => x"01",
          7682 => x"00",
          7683 => x"00",
          7684 => x"01",
          7685 => x"00",
          7686 => x"00",
          7687 => x"01",
          7688 => x"00",
          7689 => x"00",
          7690 => x"01",
          7691 => x"00",
          7692 => x"00",
          7693 => x"04",
          7694 => x"00",
          7695 => x"00",
          7696 => x"04",
          7697 => x"00",
          7698 => x"00",
          7699 => x"04",
          7700 => x"00",
          7701 => x"00",
          7702 => x"04",
          7703 => x"00",
          7704 => x"00",
          7705 => x"03",
          7706 => x"00",
          7707 => x"00",
          7708 => x"03",
          7709 => x"1b",
          7710 => x"1b",
          7711 => x"1b",
          7712 => x"1b",
          7713 => x"1b",
          7714 => x"1b",
          7715 => x"0e",
          7716 => x"0b",
          7717 => x"06",
          7718 => x"04",
          7719 => x"02",
          7720 => x"48",
          7721 => x"68",
          7722 => x"6c",
          7723 => x"6f",
          7724 => x"63",
          7725 => x"69",
          7726 => x"69",
          7727 => x"61",
          7728 => x"68",
          7729 => x"68",
          7730 => x"21",
          7731 => x"6f",
          7732 => x"65",
          7733 => x"0a",
          7734 => x"75",
          7735 => x"46",
          7736 => x"6f",
          7737 => x"74",
          7738 => x"6f",
          7739 => x"20",
          7740 => x"00",
          7741 => x"00",
          7742 => x"00",
          7743 => x"1b",
          7744 => x"1b",
          7745 => x"7e",
          7746 => x"7e",
          7747 => x"7e",
          7748 => x"7e",
          7749 => x"7e",
          7750 => x"7e",
          7751 => x"7e",
          7752 => x"7e",
          7753 => x"7e",
          7754 => x"7e",
          7755 => x"00",
          7756 => x"00",
          7757 => x"1b",
          7758 => x"1b",
          7759 => x"58",
          7760 => x"25",
          7761 => x"2c",
          7762 => x"00",
          7763 => x"2d",
          7764 => x"63",
          7765 => x"25",
          7766 => x"4b",
          7767 => x"25",
          7768 => x"25",
          7769 => x"52",
          7770 => x"72",
          7771 => x"72",
          7772 => x"30",
          7773 => x"00",
          7774 => x"30",
          7775 => x"00",
          7776 => x"30",
          7777 => x"4e",
          7778 => x"64",
          7779 => x"00",
          7780 => x"22",
          7781 => x"00",
          7782 => x"5b",
          7783 => x"46",
          7784 => x"eb",
          7785 => x"35",
          7786 => x"41",
          7787 => x"41",
          7788 => x"4e",
          7789 => x"20",
          7790 => x"20",
          7791 => x"00",
          7792 => x"00",
          7793 => x"09",
          7794 => x"1e",
          7795 => x"8e",
          7796 => x"49",
          7797 => x"99",
          7798 => x"9c",
          7799 => x"a5",
          7800 => x"ac",
          7801 => x"b4",
          7802 => x"bc",
          7803 => x"c4",
          7804 => x"cc",
          7805 => x"d4",
          7806 => x"dc",
          7807 => x"e4",
          7808 => x"ec",
          7809 => x"f4",
          7810 => x"fc",
          7811 => x"3d",
          7812 => x"3c",
          7813 => x"00",
          7814 => x"01",
          7815 => x"00",
          7816 => x"00",
          7817 => x"00",
          7818 => x"00",
          7819 => x"00",
          7820 => x"00",
          7821 => x"00",
          7822 => x"00",
          7823 => x"00",
          7824 => x"00",
          7825 => x"00",
          7826 => x"00",
          7827 => x"00",
          7828 => x"00",
          7829 => x"25",
          7830 => x"25",
          7831 => x"25",
          7832 => x"25",
          7833 => x"25",
          7834 => x"25",
          7835 => x"25",
          7836 => x"25",
          7837 => x"25",
          7838 => x"25",
          7839 => x"25",
          7840 => x"25",
          7841 => x"03",
          7842 => x"03",
          7843 => x"03",
          7844 => x"22",
          7845 => x"22",
          7846 => x"23",
          7847 => x"00",
          7848 => x"20",
          7849 => x"00",
          7850 => x"00",
          7851 => x"01",
          7852 => x"01",
          7853 => x"01",
          7854 => x"00",
          7855 => x"01",
          7856 => x"01",
          7857 => x"01",
          7858 => x"01",
          7859 => x"01",
          7860 => x"01",
          7861 => x"01",
          7862 => x"01",
          7863 => x"01",
          7864 => x"01",
          7865 => x"01",
          7866 => x"01",
          7867 => x"01",
          7868 => x"01",
          7869 => x"01",
          7870 => x"01",
          7871 => x"01",
          7872 => x"01",
          7873 => x"01",
          7874 => x"01",
          7875 => x"01",
          7876 => x"01",
          7877 => x"02",
          7878 => x"2c",
          7879 => x"2c",
          7880 => x"02",
          7881 => x"00",
          7882 => x"01",
          7883 => x"02",
          7884 => x"02",
          7885 => x"02",
          7886 => x"02",
          7887 => x"02",
          7888 => x"02",
          7889 => x"01",
          7890 => x"02",
          7891 => x"02",
          7892 => x"02",
          7893 => x"02",
          7894 => x"02",
          7895 => x"01",
          7896 => x"02",
          7897 => x"01",
          7898 => x"03",
          7899 => x"03",
          7900 => x"03",
          7901 => x"03",
          7902 => x"03",
          7903 => x"03",
          7904 => x"00",
          7905 => x"03",
          7906 => x"03",
          7907 => x"03",
          7908 => x"01",
          7909 => x"01",
          7910 => x"04",
          7911 => x"00",
          7912 => x"2c",
          7913 => x"01",
          7914 => x"06",
          7915 => x"06",
          7916 => x"00",
          7917 => x"1f",
          7918 => x"1f",
          7919 => x"1f",
          7920 => x"1f",
          7921 => x"1f",
          7922 => x"1f",
          7923 => x"1f",
          7924 => x"1f",
          7925 => x"1f",
          7926 => x"1f",
          7927 => x"06",
          7928 => x"1f",
          7929 => x"00",
          7930 => x"21",
          7931 => x"05",
          7932 => x"01",
          7933 => x"01",
          7934 => x"08",
          7935 => x"00",
          7936 => x"01",
          7937 => x"00",
          7938 => x"01",
          7939 => x"00",
          7940 => x"01",
          7941 => x"00",
          7942 => x"01",
          7943 => x"00",
          7944 => x"01",
          7945 => x"00",
          7946 => x"01",
          7947 => x"00",
          7948 => x"01",
          7949 => x"00",
          7950 => x"01",
          7951 => x"00",
          7952 => x"01",
          7953 => x"00",
          7954 => x"01",
          7955 => x"00",
          7956 => x"01",
          7957 => x"00",
          7958 => x"01",
          7959 => x"00",
          7960 => x"01",
          7961 => x"00",
          7962 => x"01",
          7963 => x"00",
          7964 => x"01",
          7965 => x"00",
          7966 => x"01",
          7967 => x"00",
          7968 => x"01",
          7969 => x"00",
          7970 => x"01",
          7971 => x"00",
          7972 => x"01",
          7973 => x"00",
          7974 => x"01",
          7975 => x"00",
          7976 => x"01",
          7977 => x"00",
          7978 => x"01",
          7979 => x"00",
          7980 => x"01",
          7981 => x"00",
          7982 => x"01",
          7983 => x"00",
          7984 => x"01",
          7985 => x"00",
          7986 => x"01",
          7987 => x"00",
          7988 => x"01",
          7989 => x"00",
          7990 => x"01",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"00",
          7996 => x"01",
          7997 => x"00",
          7998 => x"00",
          7999 => x"05",
          8000 => x"05",
          8001 => x"01",
          8002 => x"01",
          8003 => x"00",
          8004 => x"00",
          8005 => x"00",
          8006 => x"00",
          8007 => x"00",
          8008 => x"00",
          8009 => x"00",
          8010 => x"00",
          8011 => x"00",
          8012 => x"00",
          8013 => x"00",
          8014 => x"00",
          8015 => x"00",
          8016 => x"00",
          8017 => x"00",
          8018 => x"00",
          8019 => x"f0",
          8020 => x"5d",
          8021 => x"75",
          8022 => x"6d",
          8023 => x"65",
          8024 => x"35",
          8025 => x"30",
          8026 => x"f1",
          8027 => x"f0",
          8028 => x"84",
          8029 => x"f0",
          8030 => x"5d",
          8031 => x"55",
          8032 => x"4d",
          8033 => x"45",
          8034 => x"35",
          8035 => x"30",
          8036 => x"f1",
          8037 => x"f0",
          8038 => x"84",
          8039 => x"f0",
          8040 => x"7d",
          8041 => x"55",
          8042 => x"4d",
          8043 => x"45",
          8044 => x"25",
          8045 => x"20",
          8046 => x"f9",
          8047 => x"f0",
          8048 => x"89",
          8049 => x"f0",
          8050 => x"1d",
          8051 => x"15",
          8052 => x"0d",
          8053 => x"05",
          8054 => x"f0",
          8055 => x"f0",
          8056 => x"f0",
          8057 => x"f0",
          8058 => x"84",
          8059 => x"f0",
          8060 => x"b7",
          8061 => x"39",
          8062 => x"1d",
          8063 => x"74",
          8064 => x"7a",
          8065 => x"9d",
          8066 => x"c3",
          8067 => x"f0",
          8068 => x"84",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"f8",
          8083 => x"f3",
          8084 => x"f4",
          8085 => x"f1",
          8086 => x"f2",
          8087 => x"80",
          8088 => x"81",
          8089 => x"82",
          8090 => x"83",
          8091 => x"84",
          8092 => x"85",
          8093 => x"86",
          8094 => x"87",
          8095 => x"88",
          8096 => x"89",
          8097 => x"f6",
          8098 => x"7f",
          8099 => x"f9",
          8100 => x"e0",
          8101 => x"e1",
          8102 => x"71",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"50",
          9104 => x"cc",
          9105 => x"f8",
          9106 => x"e1",
          9107 => x"e3",
          9108 => x"00",
          9109 => x"68",
          9110 => x"20",
          9111 => x"28",
          9112 => x"55",
          9113 => x"08",
          9114 => x"10",
          9115 => x"18",
          9116 => x"c7",
          9117 => x"88",
          9118 => x"90",
          9119 => x"98",
          9120 => x"00",
          9121 => x"00",
          9122 => x"00",
          9123 => x"00",
          9124 => x"00",
          9125 => x"00",
          9126 => x"00",
          9127 => x"00",
          9128 => x"00",
          9129 => x"00",
          9130 => x"00",
          9131 => x"00",
          9132 => x"00",
          9133 => x"00",
          9134 => x"00",
          9135 => x"00",
          9136 => x"01",
        others => X"00"
    );

    shared variable RAM4 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"80",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"09",
             9 => x"83",
            10 => x"00",
            11 => x"00",
            12 => x"73",
            13 => x"83",
            14 => x"ff",
            15 => x"00",
            16 => x"73",
            17 => x"06",
            18 => x"00",
            19 => x"00",
            20 => x"53",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"72",
            26 => x"06",
            27 => x"00",
            28 => x"53",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"00",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"04",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"0b",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"2a",
            49 => x"05",
            50 => x"00",
            51 => x"00",
            52 => x"83",
            53 => x"2b",
            54 => x"51",
            55 => x"00",
            56 => x"70",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"70",
            61 => x"06",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"51",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"06",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"09",
            77 => x"2a",
            78 => x"00",
            79 => x"00",
            80 => x"bf",
            81 => x"08",
            82 => x"00",
            83 => x"00",
            84 => x"75",
            85 => x"50",
            86 => x"88",
            87 => x"00",
            88 => x"75",
            89 => x"50",
            90 => x"88",
            91 => x"00",
            92 => x"0a",
            93 => x"06",
            94 => x"06",
            95 => x"00",
            96 => x"0a",
            97 => x"71",
            98 => x"05",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"52",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"51",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"8c",
           134 => x"04",
           135 => x"0b",
           136 => x"8c",
           137 => x"04",
           138 => x"0b",
           139 => x"8d",
           140 => x"04",
           141 => x"0b",
           142 => x"8d",
           143 => x"04",
           144 => x"0b",
           145 => x"8e",
           146 => x"04",
           147 => x"0b",
           148 => x"8e",
           149 => x"04",
           150 => x"0b",
           151 => x"8f",
           152 => x"04",
           153 => x"0b",
           154 => x"8f",
           155 => x"04",
           156 => x"0b",
           157 => x"90",
           158 => x"04",
           159 => x"0b",
           160 => x"90",
           161 => x"04",
           162 => x"0b",
           163 => x"91",
           164 => x"04",
           165 => x"0b",
           166 => x"91",
           167 => x"04",
           168 => x"0b",
           169 => x"92",
           170 => x"04",
           171 => x"0b",
           172 => x"92",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"90",
           193 => x"90",
           194 => x"bb",
           195 => x"90",
           196 => x"bb",
           197 => x"90",
           198 => x"bb",
           199 => x"90",
           200 => x"bb",
           201 => x"90",
           202 => x"bb",
           203 => x"90",
           204 => x"bb",
           205 => x"90",
           206 => x"bb",
           207 => x"90",
           208 => x"bb",
           209 => x"90",
           210 => x"bb",
           211 => x"90",
           212 => x"bb",
           213 => x"90",
           214 => x"bb",
           215 => x"90",
           216 => x"bb",
           217 => x"bb",
           218 => x"84",
           219 => x"84",
           220 => x"04",
           221 => x"2d",
           222 => x"90",
           223 => x"eb",
           224 => x"80",
           225 => x"ca",
           226 => x"c0",
           227 => x"82",
           228 => x"80",
           229 => x"0c",
           230 => x"08",
           231 => x"90",
           232 => x"90",
           233 => x"bb",
           234 => x"bb",
           235 => x"84",
           236 => x"84",
           237 => x"04",
           238 => x"2d",
           239 => x"90",
           240 => x"95",
           241 => x"80",
           242 => x"f3",
           243 => x"c0",
           244 => x"82",
           245 => x"80",
           246 => x"0c",
           247 => x"08",
           248 => x"90",
           249 => x"90",
           250 => x"bb",
           251 => x"bb",
           252 => x"84",
           253 => x"84",
           254 => x"04",
           255 => x"2d",
           256 => x"90",
           257 => x"97",
           258 => x"80",
           259 => x"e5",
           260 => x"c0",
           261 => x"82",
           262 => x"80",
           263 => x"0c",
           264 => x"08",
           265 => x"90",
           266 => x"90",
           267 => x"bb",
           268 => x"bb",
           269 => x"84",
           270 => x"84",
           271 => x"04",
           272 => x"2d",
           273 => x"90",
           274 => x"c7",
           275 => x"80",
           276 => x"a5",
           277 => x"c0",
           278 => x"83",
           279 => x"80",
           280 => x"0c",
           281 => x"08",
           282 => x"90",
           283 => x"90",
           284 => x"bb",
           285 => x"bb",
           286 => x"84",
           287 => x"84",
           288 => x"04",
           289 => x"2d",
           290 => x"90",
           291 => x"8a",
           292 => x"80",
           293 => x"d7",
           294 => x"c0",
           295 => x"b1",
           296 => x"c0",
           297 => x"81",
           298 => x"80",
           299 => x"0c",
           300 => x"08",
           301 => x"90",
           302 => x"90",
           303 => x"bb",
           304 => x"bb",
           305 => x"3c",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"ff",
           311 => x"83",
           312 => x"fc",
           313 => x"80",
           314 => x"06",
           315 => x"0a",
           316 => x"51",
           317 => x"f0",
           318 => x"05",
           319 => x"04",
           320 => x"00",
           321 => x"84",
           322 => x"84",
           323 => x"86",
           324 => x"7a",
           325 => x"06",
           326 => x"57",
           327 => x"06",
           328 => x"8a",
           329 => x"2a",
           330 => x"25",
           331 => x"75",
           332 => x"08",
           333 => x"ae",
           334 => x"81",
           335 => x"32",
           336 => x"51",
           337 => x"38",
           338 => x"bb",
           339 => x"0b",
           340 => x"04",
           341 => x"84",
           342 => x"0a",
           343 => x"52",
           344 => x"73",
           345 => x"0d",
           346 => x"05",
           347 => x"85",
           348 => x"63",
           349 => x"1f",
           350 => x"81",
           351 => x"54",
           352 => x"d2",
           353 => x"80",
           354 => x"54",
           355 => x"d0",
           356 => x"38",
           357 => x"25",
           358 => x"80",
           359 => x"81",
           360 => x"2e",
           361 => x"7b",
           362 => x"1d",
           363 => x"91",
           364 => x"78",
           365 => x"98",
           366 => x"80",
           367 => x"2c",
           368 => x"24",
           369 => x"72",
           370 => x"58",
           371 => x"76",
           372 => x"81",
           373 => x"33",
           374 => x"9e",
           375 => x"3f",
           376 => x"ff",
           377 => x"06",
           378 => x"74",
           379 => x"17",
           380 => x"72",
           381 => x"73",
           382 => x"80",
           383 => x"76",
           384 => x"58",
           385 => x"39",
           386 => x"5a",
           387 => x"83",
           388 => x"84",
           389 => x"93",
           390 => x"ff",
           391 => x"05",
           392 => x"84",
           393 => x"7e",
           394 => x"75",
           395 => x"08",
           396 => x"7d",
           397 => x"b2",
           398 => x"38",
           399 => x"80",
           400 => x"86",
           401 => x"80",
           402 => x"29",
           403 => x"2e",
           404 => x"fc",
           405 => x"58",
           406 => x"55",
           407 => x"2c",
           408 => x"73",
           409 => x"f7",
           410 => x"41",
           411 => x"80",
           412 => x"90",
           413 => x"06",
           414 => x"96",
           415 => x"73",
           416 => x"06",
           417 => x"2a",
           418 => x"7e",
           419 => x"7a",
           420 => x"2e",
           421 => x"29",
           422 => x"5a",
           423 => x"7c",
           424 => x"78",
           425 => x"05",
           426 => x"80",
           427 => x"72",
           428 => x"80",
           429 => x"98",
           430 => x"9d",
           431 => x"3f",
           432 => x"ff",
           433 => x"55",
           434 => x"2a",
           435 => x"2e",
           436 => x"84",
           437 => x"ca",
           438 => x"38",
           439 => x"7c",
           440 => x"87",
           441 => x"09",
           442 => x"5b",
           443 => x"78",
           444 => x"05",
           445 => x"75",
           446 => x"51",
           447 => x"07",
           448 => x"5b",
           449 => x"7a",
           450 => x"90",
           451 => x"83",
           452 => x"5a",
           453 => x"77",
           454 => x"70",
           455 => x"80",
           456 => x"2c",
           457 => x"7a",
           458 => x"7a",
           459 => x"80",
           460 => x"2c",
           461 => x"b3",
           462 => x"3f",
           463 => x"ff",
           464 => x"2e",
           465 => x"81",
           466 => x"e2",
           467 => x"06",
           468 => x"fe",
           469 => x"05",
           470 => x"39",
           471 => x"07",
           472 => x"80",
           473 => x"80",
           474 => x"5d",
           475 => x"fb",
           476 => x"70",
           477 => x"82",
           478 => x"5b",
           479 => x"7a",
           480 => x"f8",
           481 => x"07",
           482 => x"f7",
           483 => x"84",
           484 => x"58",
           485 => x"51",
           486 => x"83",
           487 => x"2b",
           488 => x"87",
           489 => x"58",
           490 => x"39",
           491 => x"81",
           492 => x"cf",
           493 => x"bb",
           494 => x"71",
           495 => x"7a",
           496 => x"76",
           497 => x"78",
           498 => x"05",
           499 => x"74",
           500 => x"51",
           501 => x"b0",
           502 => x"09",
           503 => x"76",
           504 => x"81",
           505 => x"38",
           506 => x"71",
           507 => x"83",
           508 => x"fa",
           509 => x"ad",
           510 => x"54",
           511 => x"ad",
           512 => x"82",
           513 => x"80",
           514 => x"78",
           515 => x"5a",
           516 => x"51",
           517 => x"a0",
           518 => x"78",
           519 => x"bb",
           520 => x"71",
           521 => x"39",
           522 => x"ff",
           523 => x"39",
           524 => x"53",
           525 => x"84",
           526 => x"55",
           527 => x"11",
           528 => x"81",
           529 => x"56",
           530 => x"d5",
           531 => x"53",
           532 => x"e8",
           533 => x"53",
           534 => x"2e",
           535 => x"05",
           536 => x"38",
           537 => x"84",
           538 => x"08",
           539 => x"74",
           540 => x"83",
           541 => x"bb",
           542 => x"3d",
           543 => x"85",
           544 => x"70",
           545 => x"56",
           546 => x"38",
           547 => x"72",
           548 => x"76",
           549 => x"3d",
           550 => x"33",
           551 => x"52",
           552 => x"2d",
           553 => x"38",
           554 => x"54",
           555 => x"3d",
           556 => x"51",
           557 => x"3d",
           558 => x"81",
           559 => x"56",
           560 => x"82",
           561 => x"ac",
           562 => x"16",
           563 => x"76",
           564 => x"0c",
           565 => x"16",
           566 => x"0c",
           567 => x"81",
           568 => x"73",
           569 => x"e3",
           570 => x"16",
           571 => x"0d",
           572 => x"06",
           573 => x"56",
           574 => x"86",
           575 => x"72",
           576 => x"2e",
           577 => x"53",
           578 => x"81",
           579 => x"05",
           580 => x"54",
           581 => x"0d",
           582 => x"85",
           583 => x"8c",
           584 => x"84",
           585 => x"94",
           586 => x"84",
           587 => x"25",
           588 => x"90",
           589 => x"ff",
           590 => x"72",
           591 => x"bb",
           592 => x"a0",
           593 => x"54",
           594 => x"71",
           595 => x"53",
           596 => x"52",
           597 => x"70",
           598 => x"f0",
           599 => x"3d",
           600 => x"71",
           601 => x"2e",
           602 => x"70",
           603 => x"05",
           604 => x"34",
           605 => x"84",
           606 => x"70",
           607 => x"70",
           608 => x"13",
           609 => x"11",
           610 => x"13",
           611 => x"34",
           612 => x"39",
           613 => x"71",
           614 => x"f7",
           615 => x"bb",
           616 => x"fd",
           617 => x"54",
           618 => x"70",
           619 => x"f0",
           620 => x"3d",
           621 => x"71",
           622 => x"2e",
           623 => x"33",
           624 => x"11",
           625 => x"84",
           626 => x"0d",
           627 => x"80",
           628 => x"81",
           629 => x"2e",
           630 => x"54",
           631 => x"53",
           632 => x"bb",
           633 => x"80",
           634 => x"51",
           635 => x"33",
           636 => x"38",
           637 => x"86",
           638 => x"0c",
           639 => x"77",
           640 => x"3f",
           641 => x"08",
           642 => x"3f",
           643 => x"84",
           644 => x"84",
           645 => x"53",
           646 => x"fe",
           647 => x"73",
           648 => x"04",
           649 => x"54",
           650 => x"38",
           651 => x"70",
           652 => x"71",
           653 => x"ff",
           654 => x"84",
           655 => x"fd",
           656 => x"53",
           657 => x"72",
           658 => x"11",
           659 => x"84",
           660 => x"0d",
           661 => x"80",
           662 => x"3f",
           663 => x"53",
           664 => x"80",
           665 => x"31",
           666 => x"cb",
           667 => x"c3",
           668 => x"72",
           669 => x"55",
           670 => x"72",
           671 => x"77",
           672 => x"2c",
           673 => x"71",
           674 => x"55",
           675 => x"10",
           676 => x"0c",
           677 => x"76",
           678 => x"70",
           679 => x"90",
           680 => x"fe",
           681 => x"83",
           682 => x"70",
           683 => x"25",
           684 => x"2a",
           685 => x"06",
           686 => x"71",
           687 => x"81",
           688 => x"74",
           689 => x"84",
           690 => x"56",
           691 => x"56",
           692 => x"86",
           693 => x"77",
           694 => x"94",
           695 => x"74",
           696 => x"85",
           697 => x"7a",
           698 => x"8b",
           699 => x"bb",
           700 => x"80",
           701 => x"3f",
           702 => x"73",
           703 => x"80",
           704 => x"12",
           705 => x"71",
           706 => x"74",
           707 => x"9f",
           708 => x"72",
           709 => x"06",
           710 => x"1c",
           711 => x"53",
           712 => x"0c",
           713 => x"78",
           714 => x"2c",
           715 => x"73",
           716 => x"75",
           717 => x"fc",
           718 => x"32",
           719 => x"3d",
           720 => x"5b",
           721 => x"70",
           722 => x"09",
           723 => x"78",
           724 => x"2e",
           725 => x"38",
           726 => x"14",
           727 => x"db",
           728 => x"27",
           729 => x"89",
           730 => x"55",
           731 => x"51",
           732 => x"13",
           733 => x"73",
           734 => x"81",
           735 => x"16",
           736 => x"56",
           737 => x"80",
           738 => x"7a",
           739 => x"0c",
           740 => x"70",
           741 => x"73",
           742 => x"38",
           743 => x"55",
           744 => x"90",
           745 => x"81",
           746 => x"14",
           747 => x"27",
           748 => x"0c",
           749 => x"15",
           750 => x"80",
           751 => x"bb",
           752 => x"3d",
           753 => x"7b",
           754 => x"59",
           755 => x"38",
           756 => x"55",
           757 => x"ad",
           758 => x"81",
           759 => x"77",
           760 => x"80",
           761 => x"80",
           762 => x"70",
           763 => x"70",
           764 => x"27",
           765 => x"06",
           766 => x"38",
           767 => x"76",
           768 => x"70",
           769 => x"ff",
           770 => x"75",
           771 => x"75",
           772 => x"04",
           773 => x"33",
           774 => x"81",
           775 => x"78",
           776 => x"e2",
           777 => x"f8",
           778 => x"27",
           779 => x"88",
           780 => x"75",
           781 => x"04",
           782 => x"70",
           783 => x"39",
           784 => x"3d",
           785 => x"bb",
           786 => x"84",
           787 => x"71",
           788 => x"83",
           789 => x"83",
           790 => x"3d",
           791 => x"b3",
           792 => x"d4",
           793 => x"04",
           794 => x"83",
           795 => x"ef",
           796 => x"d0",
           797 => x"0d",
           798 => x"3f",
           799 => x"51",
           800 => x"83",
           801 => x"3d",
           802 => x"db",
           803 => x"9c",
           804 => x"04",
           805 => x"83",
           806 => x"ee",
           807 => x"d1",
           808 => x"0d",
           809 => x"3f",
           810 => x"51",
           811 => x"83",
           812 => x"3d",
           813 => x"83",
           814 => x"b8",
           815 => x"04",
           816 => x"83",
           817 => x"ed",
           818 => x"ec",
           819 => x"84",
           820 => x"80",
           821 => x"70",
           822 => x"59",
           823 => x"38",
           824 => x"ff",
           825 => x"e2",
           826 => x"70",
           827 => x"bb",
           828 => x"80",
           829 => x"af",
           830 => x"80",
           831 => x"06",
           832 => x"aa",
           833 => x"74",
           834 => x"52",
           835 => x"3f",
           836 => x"84",
           837 => x"df",
           838 => x"81",
           839 => x"08",
           840 => x"84",
           841 => x"05",
           842 => x"51",
           843 => x"08",
           844 => x"38",
           845 => x"38",
           846 => x"39",
           847 => x"3f",
           848 => x"f4",
           849 => x"83",
           850 => x"e0",
           851 => x"f8",
           852 => x"05",
           853 => x"7b",
           854 => x"bb",
           855 => x"91",
           856 => x"84",
           857 => x"78",
           858 => x"60",
           859 => x"7e",
           860 => x"84",
           861 => x"f3",
           862 => x"05",
           863 => x"68",
           864 => x"78",
           865 => x"83",
           866 => x"d3",
           867 => x"73",
           868 => x"81",
           869 => x"38",
           870 => x"a7",
           871 => x"51",
           872 => x"e8",
           873 => x"3f",
           874 => x"a0",
           875 => x"79",
           876 => x"33",
           877 => x"83",
           878 => x"27",
           879 => x"70",
           880 => x"2e",
           881 => x"ee",
           882 => x"51",
           883 => x"76",
           884 => x"e9",
           885 => x"58",
           886 => x"84",
           887 => x"54",
           888 => x"9b",
           889 => x"76",
           890 => x"84",
           891 => x"83",
           892 => x"14",
           893 => x"51",
           894 => x"b8",
           895 => x"51",
           896 => x"e8",
           897 => x"3f",
           898 => x"18",
           899 => x"22",
           900 => x"3f",
           901 => x"54",
           902 => x"26",
           903 => x"b4",
           904 => x"e6",
           905 => x"9e",
           906 => x"73",
           907 => x"72",
           908 => x"a0",
           909 => x"53",
           910 => x"74",
           911 => x"e6",
           912 => x"3f",
           913 => x"d0",
           914 => x"ff",
           915 => x"fc",
           916 => x"2e",
           917 => x"59",
           918 => x"3f",
           919 => x"98",
           920 => x"9b",
           921 => x"75",
           922 => x"58",
           923 => x"80",
           924 => x"08",
           925 => x"32",
           926 => x"70",
           927 => x"55",
           928 => x"24",
           929 => x"0b",
           930 => x"04",
           931 => x"08",
           932 => x"8d",
           933 => x"3f",
           934 => x"2a",
           935 => x"b7",
           936 => x"51",
           937 => x"2a",
           938 => x"db",
           939 => x"51",
           940 => x"2a",
           941 => x"ff",
           942 => x"51",
           943 => x"2a",
           944 => x"38",
           945 => x"88",
           946 => x"04",
           947 => x"e8",
           948 => x"8d",
           949 => x"04",
           950 => x"fc",
           951 => x"f5",
           952 => x"72",
           953 => x"51",
           954 => x"9b",
           955 => x"72",
           956 => x"71",
           957 => x"81",
           958 => x"51",
           959 => x"3f",
           960 => x"52",
           961 => x"be",
           962 => x"d5",
           963 => x"9b",
           964 => x"06",
           965 => x"38",
           966 => x"3f",
           967 => x"80",
           968 => x"70",
           969 => x"fe",
           970 => x"9a",
           971 => x"ed",
           972 => x"83",
           973 => x"80",
           974 => x"81",
           975 => x"51",
           976 => x"3f",
           977 => x"52",
           978 => x"bd",
           979 => x"41",
           980 => x"81",
           981 => x"84",
           982 => x"3d",
           983 => x"38",
           984 => x"98",
           985 => x"b8",
           986 => x"52",
           987 => x"83",
           988 => x"5b",
           989 => x"79",
           990 => x"ff",
           991 => x"38",
           992 => x"83",
           993 => x"2e",
           994 => x"70",
           995 => x"38",
           996 => x"7b",
           997 => x"08",
           998 => x"84",
           999 => x"53",
          1000 => x"84",
          1001 => x"33",
          1002 => x"81",
          1003 => x"9b",
          1004 => x"5c",
          1005 => x"f8",
          1006 => x"bb",
          1007 => x"80",
          1008 => x"08",
          1009 => x"91",
          1010 => x"62",
          1011 => x"84",
          1012 => x"80",
          1013 => x"80",
          1014 => x"5b",
          1015 => x"82",
          1016 => x"82",
          1017 => x"d7",
          1018 => x"83",
          1019 => x"7d",
          1020 => x"0a",
          1021 => x"f5",
          1022 => x"bb",
          1023 => x"07",
          1024 => x"5a",
          1025 => x"78",
          1026 => x"38",
          1027 => x"5a",
          1028 => x"61",
          1029 => x"38",
          1030 => x"51",
          1031 => x"51",
          1032 => x"53",
          1033 => x"0b",
          1034 => x"ff",
          1035 => x"81",
          1036 => x"94",
          1037 => x"84",
          1038 => x"0b",
          1039 => x"53",
          1040 => x"cc",
          1041 => x"a0",
          1042 => x"db",
          1043 => x"70",
          1044 => x"2e",
          1045 => x"39",
          1046 => x"3f",
          1047 => x"34",
          1048 => x"53",
          1049 => x"3f",
          1050 => x"38",
          1051 => x"1b",
          1052 => x"fc",
          1053 => x"05",
          1054 => x"d7",
          1055 => x"60",
          1056 => x"82",
          1057 => x"61",
          1058 => x"81",
          1059 => x"aa",
          1060 => x"3f",
          1061 => x"8c",
          1062 => x"83",
          1063 => x"a4",
          1064 => x"8f",
          1065 => x"39",
          1066 => x"52",
          1067 => x"ea",
          1068 => x"39",
          1069 => x"80",
          1070 => x"dd",
          1071 => x"39",
          1072 => x"80",
          1073 => x"84",
          1074 => x"52",
          1075 => x"68",
          1076 => x"80",
          1077 => x"08",
          1078 => x"3f",
          1079 => x"11",
          1080 => x"3f",
          1081 => x"fa",
          1082 => x"d0",
          1083 => x"3d",
          1084 => x"51",
          1085 => x"80",
          1086 => x"f0",
          1087 => x"82",
          1088 => x"38",
          1089 => x"83",
          1090 => x"e6",
          1091 => x"51",
          1092 => x"59",
          1093 => x"9f",
          1094 => x"70",
          1095 => x"f4",
          1096 => x"ba",
          1097 => x"f8",
          1098 => x"53",
          1099 => x"84",
          1100 => x"59",
          1101 => x"c8",
          1102 => x"08",
          1103 => x"a3",
          1104 => x"ae",
          1105 => x"87",
          1106 => x"59",
          1107 => x"53",
          1108 => x"84",
          1109 => x"38",
          1110 => x"80",
          1111 => x"84",
          1112 => x"3d",
          1113 => x"51",
          1114 => x"80",
          1115 => x"51",
          1116 => x"78",
          1117 => x"33",
          1118 => x"2e",
          1119 => x"33",
          1120 => x"cd",
          1121 => x"19",
          1122 => x"3d",
          1123 => x"51",
          1124 => x"80",
          1125 => x"fc",
          1126 => x"ce",
          1127 => x"f7",
          1128 => x"53",
          1129 => x"84",
          1130 => x"38",
          1131 => x"68",
          1132 => x"65",
          1133 => x"7c",
          1134 => x"b8",
          1135 => x"05",
          1136 => x"08",
          1137 => x"fe",
          1138 => x"e7",
          1139 => x"38",
          1140 => x"8c",
          1141 => x"08",
          1142 => x"eb",
          1143 => x"ae",
          1144 => x"84",
          1145 => x"39",
          1146 => x"79",
          1147 => x"fe",
          1148 => x"e7",
          1149 => x"2e",
          1150 => x"db",
          1151 => x"49",
          1152 => x"80",
          1153 => x"84",
          1154 => x"b8",
          1155 => x"05",
          1156 => x"08",
          1157 => x"fe",
          1158 => x"e6",
          1159 => x"2e",
          1160 => x"11",
          1161 => x"3f",
          1162 => x"bb",
          1163 => x"cb",
          1164 => x"7a",
          1165 => x"70",
          1166 => x"f5",
          1167 => x"ca",
          1168 => x"87",
          1169 => x"3d",
          1170 => x"3f",
          1171 => x"78",
          1172 => x"08",
          1173 => x"84",
          1174 => x"39",
          1175 => x"80",
          1176 => x"84",
          1177 => x"5a",
          1178 => x"f3",
          1179 => x"11",
          1180 => x"3f",
          1181 => x"f4",
          1182 => x"8a",
          1183 => x"3d",
          1184 => x"51",
          1185 => x"80",
          1186 => x"7a",
          1187 => x"90",
          1188 => x"2a",
          1189 => x"2e",
          1190 => x"88",
          1191 => x"3f",
          1192 => x"52",
          1193 => x"b4",
          1194 => x"64",
          1195 => x"45",
          1196 => x"80",
          1197 => x"84",
          1198 => x"64",
          1199 => x"b8",
          1200 => x"05",
          1201 => x"08",
          1202 => x"02",
          1203 => x"05",
          1204 => x"f0",
          1205 => x"d2",
          1206 => x"f2",
          1207 => x"05",
          1208 => x"7d",
          1209 => x"ff",
          1210 => x"bb",
          1211 => x"39",
          1212 => x"80",
          1213 => x"84",
          1214 => x"5c",
          1215 => x"68",
          1216 => x"3d",
          1217 => x"51",
          1218 => x"80",
          1219 => x"0c",
          1220 => x"f7",
          1221 => x"06",
          1222 => x"a0",
          1223 => x"7c",
          1224 => x"7b",
          1225 => x"87",
          1226 => x"3f",
          1227 => x"11",
          1228 => x"3f",
          1229 => x"38",
          1230 => x"79",
          1231 => x"f7",
          1232 => x"7b",
          1233 => x"cc",
          1234 => x"89",
          1235 => x"83",
          1236 => x"83",
          1237 => x"59",
          1238 => x"d3",
          1239 => x"83",
          1240 => x"a5",
          1241 => x"8b",
          1242 => x"3f",
          1243 => x"59",
          1244 => x"d4",
          1245 => x"8b",
          1246 => x"83",
          1247 => x"83",
          1248 => x"9b",
          1249 => x"ee",
          1250 => x"80",
          1251 => x"49",
          1252 => x"5d",
          1253 => x"e4",
          1254 => x"f0",
          1255 => x"39",
          1256 => x"fb",
          1257 => x"84",
          1258 => x"70",
          1259 => x"74",
          1260 => x"08",
          1261 => x"84",
          1262 => x"74",
          1263 => x"87",
          1264 => x"87",
          1265 => x"3f",
          1266 => x"08",
          1267 => x"51",
          1268 => x"08",
          1269 => x"87",
          1270 => x"0b",
          1271 => x"ba",
          1272 => x"84",
          1273 => x"e6",
          1274 => x"0c",
          1275 => x"56",
          1276 => x"98",
          1277 => x"83",
          1278 => x"c4",
          1279 => x"52",
          1280 => x"54",
          1281 => x"52",
          1282 => x"8d",
          1283 => x"d3",
          1284 => x"c3",
          1285 => x"d4",
          1286 => x"3f",
          1287 => x"08",
          1288 => x"73",
          1289 => x"81",
          1290 => x"09",
          1291 => x"33",
          1292 => x"70",
          1293 => x"06",
          1294 => x"74",
          1295 => x"80",
          1296 => x"54",
          1297 => x"54",
          1298 => x"2e",
          1299 => x"80",
          1300 => x"a0",
          1301 => x"54",
          1302 => x"25",
          1303 => x"2e",
          1304 => x"54",
          1305 => x"84",
          1306 => x"70",
          1307 => x"ff",
          1308 => x"33",
          1309 => x"70",
          1310 => x"39",
          1311 => x"72",
          1312 => x"38",
          1313 => x"72",
          1314 => x"84",
          1315 => x"fc",
          1316 => x"84",
          1317 => x"74",
          1318 => x"04",
          1319 => x"ff",
          1320 => x"26",
          1321 => x"05",
          1322 => x"8a",
          1323 => x"70",
          1324 => x"33",
          1325 => x"f2",
          1326 => x"74",
          1327 => x"22",
          1328 => x"80",
          1329 => x"52",
          1330 => x"81",
          1331 => x"22",
          1332 => x"33",
          1333 => x"33",
          1334 => x"33",
          1335 => x"33",
          1336 => x"33",
          1337 => x"c0",
          1338 => x"a0",
          1339 => x"0c",
          1340 => x"86",
          1341 => x"5b",
          1342 => x"0c",
          1343 => x"7b",
          1344 => x"7b",
          1345 => x"08",
          1346 => x"98",
          1347 => x"87",
          1348 => x"1c",
          1349 => x"7b",
          1350 => x"08",
          1351 => x"98",
          1352 => x"80",
          1353 => x"59",
          1354 => x"1b",
          1355 => x"1b",
          1356 => x"1b",
          1357 => x"52",
          1358 => x"3f",
          1359 => x"02",
          1360 => x"a8",
          1361 => x"84",
          1362 => x"2c",
          1363 => x"06",
          1364 => x"71",
          1365 => x"04",
          1366 => x"bb",
          1367 => x"51",
          1368 => x"df",
          1369 => x"84",
          1370 => x"2c",
          1371 => x"c7",
          1372 => x"52",
          1373 => x"e8",
          1374 => x"2b",
          1375 => x"2e",
          1376 => x"54",
          1377 => x"84",
          1378 => x"fc",
          1379 => x"f3",
          1380 => x"55",
          1381 => x"87",
          1382 => x"70",
          1383 => x"2e",
          1384 => x"06",
          1385 => x"32",
          1386 => x"38",
          1387 => x"cf",
          1388 => x"c0",
          1389 => x"38",
          1390 => x"0c",
          1391 => x"0d",
          1392 => x"51",
          1393 => x"81",
          1394 => x"71",
          1395 => x"2e",
          1396 => x"70",
          1397 => x"52",
          1398 => x"0d",
          1399 => x"9f",
          1400 => x"bc",
          1401 => x"0d",
          1402 => x"52",
          1403 => x"81",
          1404 => x"ff",
          1405 => x"80",
          1406 => x"70",
          1407 => x"52",
          1408 => x"2a",
          1409 => x"38",
          1410 => x"80",
          1411 => x"06",
          1412 => x"06",
          1413 => x"80",
          1414 => x"52",
          1415 => x"55",
          1416 => x"bb",
          1417 => x"91",
          1418 => x"98",
          1419 => x"72",
          1420 => x"81",
          1421 => x"38",
          1422 => x"2a",
          1423 => x"ce",
          1424 => x"c0",
          1425 => x"06",
          1426 => x"38",
          1427 => x"c0",
          1428 => x"f3",
          1429 => x"83",
          1430 => x"08",
          1431 => x"9c",
          1432 => x"9e",
          1433 => x"c0",
          1434 => x"87",
          1435 => x"0c",
          1436 => x"e0",
          1437 => x"f3",
          1438 => x"83",
          1439 => x"08",
          1440 => x"c4",
          1441 => x"9e",
          1442 => x"23",
          1443 => x"f8",
          1444 => x"f3",
          1445 => x"83",
          1446 => x"84",
          1447 => x"08",
          1448 => x"52",
          1449 => x"85",
          1450 => x"08",
          1451 => x"52",
          1452 => x"71",
          1453 => x"c0",
          1454 => x"06",
          1455 => x"38",
          1456 => x"80",
          1457 => x"88",
          1458 => x"80",
          1459 => x"f4",
          1460 => x"90",
          1461 => x"52",
          1462 => x"52",
          1463 => x"87",
          1464 => x"80",
          1465 => x"83",
          1466 => x"34",
          1467 => x"70",
          1468 => x"70",
          1469 => x"83",
          1470 => x"9e",
          1471 => x"51",
          1472 => x"81",
          1473 => x"0b",
          1474 => x"80",
          1475 => x"2e",
          1476 => x"8d",
          1477 => x"08",
          1478 => x"52",
          1479 => x"71",
          1480 => x"c0",
          1481 => x"51",
          1482 => x"81",
          1483 => x"c0",
          1484 => x"8a",
          1485 => x"34",
          1486 => x"70",
          1487 => x"80",
          1488 => x"f4",
          1489 => x"83",
          1490 => x"71",
          1491 => x"c0",
          1492 => x"52",
          1493 => x"52",
          1494 => x"9e",
          1495 => x"f4",
          1496 => x"52",
          1497 => x"da",
          1498 => x"f4",
          1499 => x"83",
          1500 => x"f4",
          1501 => x"83",
          1502 => x"38",
          1503 => x"9e",
          1504 => x"84",
          1505 => x"73",
          1506 => x"56",
          1507 => x"33",
          1508 => x"91",
          1509 => x"f4",
          1510 => x"83",
          1511 => x"38",
          1512 => x"89",
          1513 => x"82",
          1514 => x"73",
          1515 => x"c2",
          1516 => x"83",
          1517 => x"83",
          1518 => x"51",
          1519 => x"08",
          1520 => x"80",
          1521 => x"3f",
          1522 => x"cc",
          1523 => x"f8",
          1524 => x"51",
          1525 => x"bd",
          1526 => x"54",
          1527 => x"f4",
          1528 => x"8b",
          1529 => x"86",
          1530 => x"0d",
          1531 => x"84",
          1532 => x"84",
          1533 => x"76",
          1534 => x"08",
          1535 => x"88",
          1536 => x"fc",
          1537 => x"51",
          1538 => x"bd",
          1539 => x"54",
          1540 => x"cc",
          1541 => x"86",
          1542 => x"38",
          1543 => x"c0",
          1544 => x"ab",
          1545 => x"da",
          1546 => x"f3",
          1547 => x"ff",
          1548 => x"52",
          1549 => x"3f",
          1550 => x"3f",
          1551 => x"cc",
          1552 => x"f8",
          1553 => x"51",
          1554 => x"bd",
          1555 => x"54",
          1556 => x"f4",
          1557 => x"8b",
          1558 => x"38",
          1559 => x"ff",
          1560 => x"54",
          1561 => x"eb",
          1562 => x"9b",
          1563 => x"80",
          1564 => x"dd",
          1565 => x"f4",
          1566 => x"d1",
          1567 => x"ff",
          1568 => x"54",
          1569 => x"39",
          1570 => x"b4",
          1571 => x"85",
          1572 => x"38",
          1573 => x"83",
          1574 => x"83",
          1575 => x"fb",
          1576 => x"33",
          1577 => x"b8",
          1578 => x"80",
          1579 => x"f3",
          1580 => x"54",
          1581 => x"98",
          1582 => x"80",
          1583 => x"f3",
          1584 => x"54",
          1585 => x"f8",
          1586 => x"80",
          1587 => x"f3",
          1588 => x"54",
          1589 => x"d8",
          1590 => x"80",
          1591 => x"f3",
          1592 => x"54",
          1593 => x"b8",
          1594 => x"80",
          1595 => x"f3",
          1596 => x"54",
          1597 => x"98",
          1598 => x"80",
          1599 => x"df",
          1600 => x"da",
          1601 => x"f4",
          1602 => x"d7",
          1603 => x"8e",
          1604 => x"38",
          1605 => x"52",
          1606 => x"ff",
          1607 => x"83",
          1608 => x"83",
          1609 => x"ff",
          1610 => x"83",
          1611 => x"83",
          1612 => x"ff",
          1613 => x"83",
          1614 => x"83",
          1615 => x"04",
          1616 => x"04",
          1617 => x"84",
          1618 => x"08",
          1619 => x"57",
          1620 => x"51",
          1621 => x"08",
          1622 => x"0b",
          1623 => x"f8",
          1624 => x"84",
          1625 => x"76",
          1626 => x"08",
          1627 => x"bb",
          1628 => x"84",
          1629 => x"80",
          1630 => x"72",
          1631 => x"76",
          1632 => x"83",
          1633 => x"51",
          1634 => x"08",
          1635 => x"77",
          1636 => x"04",
          1637 => x"3f",
          1638 => x"38",
          1639 => x"79",
          1640 => x"08",
          1641 => x"76",
          1642 => x"b0",
          1643 => x"a9",
          1644 => x"3d",
          1645 => x"72",
          1646 => x"2e",
          1647 => x"59",
          1648 => x"f8",
          1649 => x"98",
          1650 => x"52",
          1651 => x"84",
          1652 => x"33",
          1653 => x"73",
          1654 => x"81",
          1655 => x"c1",
          1656 => x"0c",
          1657 => x"aa",
          1658 => x"05",
          1659 => x"08",
          1660 => x"78",
          1661 => x"bb",
          1662 => x"80",
          1663 => x"ff",
          1664 => x"f9",
          1665 => x"05",
          1666 => x"81",
          1667 => x"73",
          1668 => x"38",
          1669 => x"8d",
          1670 => x"84",
          1671 => x"08",
          1672 => x"bb",
          1673 => x"ec",
          1674 => x"82",
          1675 => x"80",
          1676 => x"c0",
          1677 => x"0b",
          1678 => x"84",
          1679 => x"58",
          1680 => x"52",
          1681 => x"ff",
          1682 => x"81",
          1683 => x"bb",
          1684 => x"3d",
          1685 => x"ba",
          1686 => x"08",
          1687 => x"b5",
          1688 => x"75",
          1689 => x"08",
          1690 => x"ff",
          1691 => x"ed",
          1692 => x"81",
          1693 => x"8b",
          1694 => x"94",
          1695 => x"ea",
          1696 => x"2b",
          1697 => x"2e",
          1698 => x"84",
          1699 => x"98",
          1700 => x"2b",
          1701 => x"70",
          1702 => x"08",
          1703 => x"5a",
          1704 => x"74",
          1705 => x"27",
          1706 => x"29",
          1707 => x"57",
          1708 => x"75",
          1709 => x"80",
          1710 => x"57",
          1711 => x"e0",
          1712 => x"78",
          1713 => x"2e",
          1714 => x"81",
          1715 => x"81",
          1716 => x"84",
          1717 => x"97",
          1718 => x"2b",
          1719 => x"5e",
          1720 => x"2e",
          1721 => x"34",
          1722 => x"84",
          1723 => x"57",
          1724 => x"ab",
          1725 => x"7d",
          1726 => x"ff",
          1727 => x"81",
          1728 => x"81",
          1729 => x"26",
          1730 => x"82",
          1731 => x"e4",
          1732 => x"ce",
          1733 => x"70",
          1734 => x"bc",
          1735 => x"fe",
          1736 => x"fe",
          1737 => x"fd",
          1738 => x"38",
          1739 => x"e2",
          1740 => x"0c",
          1741 => x"38",
          1742 => x"57",
          1743 => x"08",
          1744 => x"34",
          1745 => x"39",
          1746 => x"2e",
          1747 => x"52",
          1748 => x"e2",
          1749 => x"e2",
          1750 => x"c8",
          1751 => x"c4",
          1752 => x"fc",
          1753 => x"81",
          1754 => x"7b",
          1755 => x"8e",
          1756 => x"90",
          1757 => x"7c",
          1758 => x"08",
          1759 => x"0b",
          1760 => x"84",
          1761 => x"56",
          1762 => x"e6",
          1763 => x"ce",
          1764 => x"51",
          1765 => x"08",
          1766 => x"84",
          1767 => x"84",
          1768 => x"55",
          1769 => x"b8",
          1770 => x"a5",
          1771 => x"08",
          1772 => x"70",
          1773 => x"26",
          1774 => x"98",
          1775 => x"bc",
          1776 => x"7c",
          1777 => x"08",
          1778 => x"38",
          1779 => x"bb",
          1780 => x"bb",
          1781 => x"53",
          1782 => x"3f",
          1783 => x"33",
          1784 => x"38",
          1785 => x"ff",
          1786 => x"52",
          1787 => x"e6",
          1788 => x"86",
          1789 => x"55",
          1790 => x"ff",
          1791 => x"33",
          1792 => x"33",
          1793 => x"ed",
          1794 => x"15",
          1795 => x"16",
          1796 => x"3f",
          1797 => x"06",
          1798 => x"75",
          1799 => x"e8",
          1800 => x"e2",
          1801 => x"55",
          1802 => x"33",
          1803 => x"33",
          1804 => x"a9",
          1805 => x"33",
          1806 => x"76",
          1807 => x"7a",
          1808 => x"70",
          1809 => x"57",
          1810 => x"84",
          1811 => x"b1",
          1812 => x"98",
          1813 => x"33",
          1814 => x"f8",
          1815 => x"88",
          1816 => x"80",
          1817 => x"98",
          1818 => x"59",
          1819 => x"e6",
          1820 => x"86",
          1821 => x"80",
          1822 => x"c4",
          1823 => x"ff",
          1824 => x"58",
          1825 => x"e8",
          1826 => x"d6",
          1827 => x"80",
          1828 => x"c4",
          1829 => x"fe",
          1830 => x"33",
          1831 => x"77",
          1832 => x"81",
          1833 => x"70",
          1834 => x"57",
          1835 => x"fe",
          1836 => x"74",
          1837 => x"e8",
          1838 => x"3f",
          1839 => x"76",
          1840 => x"06",
          1841 => x"7c",
          1842 => x"e8",
          1843 => x"3f",
          1844 => x"bb",
          1845 => x"06",
          1846 => x"c4",
          1847 => x"38",
          1848 => x"83",
          1849 => x"56",
          1850 => x"87",
          1851 => x"18",
          1852 => x"3f",
          1853 => x"f4",
          1854 => x"9c",
          1855 => x"94",
          1856 => x"f4",
          1857 => x"9c",
          1858 => x"8b",
          1859 => x"75",
          1860 => x"33",
          1861 => x"80",
          1862 => x"84",
          1863 => x"0c",
          1864 => x"33",
          1865 => x"e6",
          1866 => x"96",
          1867 => x"51",
          1868 => x"08",
          1869 => x"84",
          1870 => x"84",
          1871 => x"55",
          1872 => x"ff",
          1873 => x"c8",
          1874 => x"f4",
          1875 => x"81",
          1876 => x"f4",
          1877 => x"05",
          1878 => x"16",
          1879 => x"e6",
          1880 => x"a6",
          1881 => x"2b",
          1882 => x"5a",
          1883 => x"ef",
          1884 => x"51",
          1885 => x"33",
          1886 => x"e2",
          1887 => x"79",
          1888 => x"08",
          1889 => x"74",
          1890 => x"05",
          1891 => x"5c",
          1892 => x"38",
          1893 => x"ff",
          1894 => x"29",
          1895 => x"84",
          1896 => x"75",
          1897 => x"7b",
          1898 => x"84",
          1899 => x"ff",
          1900 => x"29",
          1901 => x"84",
          1902 => x"62",
          1903 => x"81",
          1904 => x"08",
          1905 => x"3f",
          1906 => x"0a",
          1907 => x"33",
          1908 => x"a7",
          1909 => x"80",
          1910 => x"33",
          1911 => x"e6",
          1912 => x"a6",
          1913 => x"51",
          1914 => x"08",
          1915 => x"84",
          1916 => x"84",
          1917 => x"55",
          1918 => x"ff",
          1919 => x"c8",
          1920 => x"7b",
          1921 => x"04",
          1922 => x"06",
          1923 => x"38",
          1924 => x"27",
          1925 => x"2c",
          1926 => x"7b",
          1927 => x"75",
          1928 => x"05",
          1929 => x"52",
          1930 => x"81",
          1931 => x"77",
          1932 => x"3d",
          1933 => x"57",
          1934 => x"56",
          1935 => x"84",
          1936 => x"29",
          1937 => x"79",
          1938 => x"61",
          1939 => x"2b",
          1940 => x"5b",
          1941 => x"38",
          1942 => x"ff",
          1943 => x"29",
          1944 => x"84",
          1945 => x"75",
          1946 => x"08",
          1947 => x"75",
          1948 => x"05",
          1949 => x"57",
          1950 => x"38",
          1951 => x"e2",
          1952 => x"f4",
          1953 => x"83",
          1954 => x"83",
          1955 => x"38",
          1956 => x"cf",
          1957 => x"08",
          1958 => x"ff",
          1959 => x"29",
          1960 => x"84",
          1961 => x"76",
          1962 => x"70",
          1963 => x"ff",
          1964 => x"25",
          1965 => x"f4",
          1966 => x"83",
          1967 => x"55",
          1968 => x"58",
          1969 => x"0b",
          1970 => x"08",
          1971 => x"74",
          1972 => x"ec",
          1973 => x"0b",
          1974 => x"3d",
          1975 => x"80",
          1976 => x"16",
          1977 => x"ff",
          1978 => x"ff",
          1979 => x"84",
          1980 => x"81",
          1981 => x"7b",
          1982 => x"84",
          1983 => x"57",
          1984 => x"38",
          1985 => x"ff",
          1986 => x"52",
          1987 => x"e6",
          1988 => x"c6",
          1989 => x"59",
          1990 => x"ff",
          1991 => x"a9",
          1992 => x"e2",
          1993 => x"ff",
          1994 => x"51",
          1995 => x"c4",
          1996 => x"5d",
          1997 => x"e6",
          1998 => x"f6",
          1999 => x"51",
          2000 => x"08",
          2001 => x"84",
          2002 => x"84",
          2003 => x"55",
          2004 => x"3f",
          2005 => x"34",
          2006 => x"81",
          2007 => x"a9",
          2008 => x"06",
          2009 => x"33",
          2010 => x"f0",
          2011 => x"88",
          2012 => x"e8",
          2013 => x"3f",
          2014 => x"ff",
          2015 => x"ff",
          2016 => x"7a",
          2017 => x"7c",
          2018 => x"80",
          2019 => x"bb",
          2020 => x"f4",
          2021 => x"ce",
          2022 => x"84",
          2023 => x"84",
          2024 => x"05",
          2025 => x"9a",
          2026 => x"c8",
          2027 => x"eb",
          2028 => x"51",
          2029 => x"08",
          2030 => x"84",
          2031 => x"a3",
          2032 => x"05",
          2033 => x"81",
          2034 => x"80",
          2035 => x"70",
          2036 => x"9c",
          2037 => x"56",
          2038 => x"08",
          2039 => x"10",
          2040 => x"54",
          2041 => x"94",
          2042 => x"10",
          2043 => x"57",
          2044 => x"38",
          2045 => x"a6",
          2046 => x"05",
          2047 => x"75",
          2048 => x"f4",
          2049 => x"f8",
          2050 => x"51",
          2051 => x"08",
          2052 => x"83",
          2053 => x"3f",
          2054 => x"0b",
          2055 => x"84",
          2056 => x"77",
          2057 => x"84",
          2058 => x"bb",
          2059 => x"f4",
          2060 => x"51",
          2061 => x"08",
          2062 => x"09",
          2063 => x"84",
          2064 => x"bb",
          2065 => x"84",
          2066 => x"84",
          2067 => x"80",
          2068 => x"f4",
          2069 => x"9c",
          2070 => x"74",
          2071 => x"fc",
          2072 => x"70",
          2073 => x"84",
          2074 => x"f4",
          2075 => x"05",
          2076 => x"52",
          2077 => x"f4",
          2078 => x"05",
          2079 => x"38",
          2080 => x"56",
          2081 => x"76",
          2082 => x"38",
          2083 => x"75",
          2084 => x"c2",
          2085 => x"70",
          2086 => x"27",
          2087 => x"f4",
          2088 => x"d4",
          2089 => x"82",
          2090 => x"05",
          2091 => x"80",
          2092 => x"7f",
          2093 => x"10",
          2094 => x"56",
          2095 => x"88",
          2096 => x"10",
          2097 => x"41",
          2098 => x"ff",
          2099 => x"fe",
          2100 => x"f0",
          2101 => x"9d",
          2102 => x"b6",
          2103 => x"05",
          2104 => x"33",
          2105 => x"38",
          2106 => x"73",
          2107 => x"82",
          2108 => x"86",
          2109 => x"56",
          2110 => x"38",
          2111 => x"fa",
          2112 => x"83",
          2113 => x"90",
          2114 => x"07",
          2115 => x"77",
          2116 => x"05",
          2117 => x"55",
          2118 => x"78",
          2119 => x"84",
          2120 => x"55",
          2121 => x"74",
          2122 => x"13",
          2123 => x"04",
          2124 => x"b4",
          2125 => x"b5",
          2126 => x"5b",
          2127 => x"80",
          2128 => x"ff",
          2129 => x"ff",
          2130 => x"ff",
          2131 => x"5d",
          2132 => x"26",
          2133 => x"56",
          2134 => x"06",
          2135 => x"ff",
          2136 => x"29",
          2137 => x"74",
          2138 => x"33",
          2139 => x"1b",
          2140 => x"80",
          2141 => x"53",
          2142 => x"73",
          2143 => x"b0",
          2144 => x"e8",
          2145 => x"c7",
          2146 => x"70",
          2147 => x"70",
          2148 => x"70",
          2149 => x"56",
          2150 => x"38",
          2151 => x"06",
          2152 => x"79",
          2153 => x"83",
          2154 => x"b5",
          2155 => x"2b",
          2156 => x"07",
          2157 => x"5b",
          2158 => x"be",
          2159 => x"b4",
          2160 => x"10",
          2161 => x"29",
          2162 => x"57",
          2163 => x"80",
          2164 => x"81",
          2165 => x"81",
          2166 => x"83",
          2167 => x"05",
          2168 => x"5e",
          2169 => x"7a",
          2170 => x"53",
          2171 => x"06",
          2172 => x"06",
          2173 => x"58",
          2174 => x"26",
          2175 => x"73",
          2176 => x"79",
          2177 => x"7b",
          2178 => x"78",
          2179 => x"fb",
          2180 => x"ff",
          2181 => x"73",
          2182 => x"9c",
          2183 => x"75",
          2184 => x"76",
          2185 => x"94",
          2186 => x"ff",
          2187 => x"fa",
          2188 => x"08",
          2189 => x"81",
          2190 => x"55",
          2191 => x"ff",
          2192 => x"75",
          2193 => x"77",
          2194 => x"c0",
          2195 => x"06",
          2196 => x"d0",
          2197 => x"84",
          2198 => x"84",
          2199 => x"04",
          2200 => x"02",
          2201 => x"f7",
          2202 => x"79",
          2203 => x"33",
          2204 => x"33",
          2205 => x"80",
          2206 => x"57",
          2207 => x"ff",
          2208 => x"57",
          2209 => x"38",
          2210 => x"74",
          2211 => x"33",
          2212 => x"81",
          2213 => x"26",
          2214 => x"83",
          2215 => x"70",
          2216 => x"33",
          2217 => x"89",
          2218 => x"29",
          2219 => x"26",
          2220 => x"54",
          2221 => x"16",
          2222 => x"75",
          2223 => x"54",
          2224 => x"73",
          2225 => x"b0",
          2226 => x"a0",
          2227 => x"70",
          2228 => x"9f",
          2229 => x"f6",
          2230 => x"b2",
          2231 => x"77",
          2232 => x"73",
          2233 => x"81",
          2234 => x"29",
          2235 => x"a0",
          2236 => x"81",
          2237 => x"71",
          2238 => x"79",
          2239 => x"54",
          2240 => x"80",
          2241 => x"34",
          2242 => x"70",
          2243 => x"b8",
          2244 => x"71",
          2245 => x"75",
          2246 => x"bb",
          2247 => x"83",
          2248 => x"70",
          2249 => x"33",
          2250 => x"f9",
          2251 => x"78",
          2252 => x"b4",
          2253 => x"81",
          2254 => x"81",
          2255 => x"29",
          2256 => x"54",
          2257 => x"fa",
          2258 => x"76",
          2259 => x"e0",
          2260 => x"57",
          2261 => x"fe",
          2262 => x"34",
          2263 => x"ff",
          2264 => x"39",
          2265 => x"56",
          2266 => x"33",
          2267 => x"34",
          2268 => x"39",
          2269 => x"9f",
          2270 => x"9b",
          2271 => x"05",
          2272 => x"33",
          2273 => x"83",
          2274 => x"84",
          2275 => x"83",
          2276 => x"70",
          2277 => x"2e",
          2278 => x"fa",
          2279 => x"0c",
          2280 => x"33",
          2281 => x"2c",
          2282 => x"83",
          2283 => x"b4",
          2284 => x"ff",
          2285 => x"83",
          2286 => x"34",
          2287 => x"3d",
          2288 => x"73",
          2289 => x"06",
          2290 => x"b5",
          2291 => x"86",
          2292 => x"72",
          2293 => x"55",
          2294 => x"70",
          2295 => x"0b",
          2296 => x"04",
          2297 => x"fa",
          2298 => x"05",
          2299 => x"38",
          2300 => x"34",
          2301 => x"8f",
          2302 => x"38",
          2303 => x"51",
          2304 => x"70",
          2305 => x"f0",
          2306 => x"52",
          2307 => x"81",
          2308 => x"fa",
          2309 => x"0c",
          2310 => x"33",
          2311 => x"83",
          2312 => x"84",
          2313 => x"b0",
          2314 => x"fa",
          2315 => x"33",
          2316 => x"83",
          2317 => x"0b",
          2318 => x"bb",
          2319 => x"fa",
          2320 => x"51",
          2321 => x"39",
          2322 => x"70",
          2323 => x"83",
          2324 => x"07",
          2325 => x"93",
          2326 => x"06",
          2327 => x"34",
          2328 => x"81",
          2329 => x"fa",
          2330 => x"b0",
          2331 => x"fa",
          2332 => x"b0",
          2333 => x"51",
          2334 => x"39",
          2335 => x"b0",
          2336 => x"fe",
          2337 => x"ef",
          2338 => x"fa",
          2339 => x"b0",
          2340 => x"51",
          2341 => x"39",
          2342 => x"a0",
          2343 => x"fe",
          2344 => x"8f",
          2345 => x"fd",
          2346 => x"fa",
          2347 => x"b0",
          2348 => x"02",
          2349 => x"c3",
          2350 => x"fa",
          2351 => x"b8",
          2352 => x"59",
          2353 => x"82",
          2354 => x"82",
          2355 => x"0b",
          2356 => x"b4",
          2357 => x"83",
          2358 => x"78",
          2359 => x"80",
          2360 => x"84",
          2361 => x"b4",
          2362 => x"82",
          2363 => x"84",
          2364 => x"33",
          2365 => x"54",
          2366 => x"51",
          2367 => x"fa",
          2368 => x"7a",
          2369 => x"b2",
          2370 => x"3d",
          2371 => x"34",
          2372 => x"0b",
          2373 => x"fa",
          2374 => x"23",
          2375 => x"86",
          2376 => x"79",
          2377 => x"83",
          2378 => x"80",
          2379 => x"79",
          2380 => x"ba",
          2381 => x"e5",
          2382 => x"1a",
          2383 => x"33",
          2384 => x"38",
          2385 => x"3f",
          2386 => x"84",
          2387 => x"34",
          2388 => x"fa",
          2389 => x"0b",
          2390 => x"b8",
          2391 => x"34",
          2392 => x"0b",
          2393 => x"51",
          2394 => x"08",
          2395 => x"a8",
          2396 => x"ff",
          2397 => x"08",
          2398 => x"19",
          2399 => x"fe",
          2400 => x"06",
          2401 => x"7a",
          2402 => x"b8",
          2403 => x"fa",
          2404 => x"c7",
          2405 => x"53",
          2406 => x"70",
          2407 => x"33",
          2408 => x"81",
          2409 => x"81",
          2410 => x"38",
          2411 => x"88",
          2412 => x"33",
          2413 => x"33",
          2414 => x"84",
          2415 => x"80",
          2416 => x"fa",
          2417 => x"71",
          2418 => x"83",
          2419 => x"33",
          2420 => x"fa",
          2421 => x"34",
          2422 => x"06",
          2423 => x"33",
          2424 => x"55",
          2425 => x"d6",
          2426 => x"06",
          2427 => x"38",
          2428 => x"ea",
          2429 => x"b5",
          2430 => x"80",
          2431 => x"57",
          2432 => x"0b",
          2433 => x"04",
          2434 => x"24",
          2435 => x"81",
          2436 => x"51",
          2437 => x"b5",
          2438 => x"15",
          2439 => x"74",
          2440 => x"fe",
          2441 => x"51",
          2442 => x"ff",
          2443 => x"91",
          2444 => x"3f",
          2445 => x"54",
          2446 => x"39",
          2447 => x"39",
          2448 => x"80",
          2449 => x"0d",
          2450 => x"06",
          2451 => x"70",
          2452 => x"73",
          2453 => x"b5",
          2454 => x"3f",
          2455 => x"06",
          2456 => x"38",
          2457 => x"fe",
          2458 => x"34",
          2459 => x"fe",
          2460 => x"d8",
          2461 => x"02",
          2462 => x"08",
          2463 => x"38",
          2464 => x"8a",
          2465 => x"82",
          2466 => x"38",
          2467 => x"b8",
          2468 => x"fa",
          2469 => x"5e",
          2470 => x"c7",
          2471 => x"33",
          2472 => x"22",
          2473 => x"40",
          2474 => x"fa",
          2475 => x"40",
          2476 => x"c7",
          2477 => x"33",
          2478 => x"22",
          2479 => x"11",
          2480 => x"b0",
          2481 => x"1d",
          2482 => x"61",
          2483 => x"33",
          2484 => x"56",
          2485 => x"84",
          2486 => x"78",
          2487 => x"25",
          2488 => x"b3",
          2489 => x"38",
          2490 => x"b8",
          2491 => x"fa",
          2492 => x"40",
          2493 => x"c7",
          2494 => x"33",
          2495 => x"22",
          2496 => x"56",
          2497 => x"fa",
          2498 => x"57",
          2499 => x"80",
          2500 => x"81",
          2501 => x"fa",
          2502 => x"42",
          2503 => x"60",
          2504 => x"58",
          2505 => x"27",
          2506 => x"34",
          2507 => x"3d",
          2508 => x"38",
          2509 => x"8d",
          2510 => x"80",
          2511 => x"84",
          2512 => x"78",
          2513 => x"56",
          2514 => x"ba",
          2515 => x"84",
          2516 => x"18",
          2517 => x"0b",
          2518 => x"84",
          2519 => x"78",
          2520 => x"84",
          2521 => x"83",
          2522 => x"72",
          2523 => x"b9",
          2524 => x"1d",
          2525 => x"b5",
          2526 => x"29",
          2527 => x"fa",
          2528 => x"76",
          2529 => x"b0",
          2530 => x"84",
          2531 => x"83",
          2532 => x"72",
          2533 => x"59",
          2534 => x"d6",
          2535 => x"39",
          2536 => x"80",
          2537 => x"39",
          2538 => x"33",
          2539 => x"33",
          2540 => x"80",
          2541 => x"5d",
          2542 => x"ff",
          2543 => x"59",
          2544 => x"38",
          2545 => x"57",
          2546 => x"83",
          2547 => x"0b",
          2548 => x"ba",
          2549 => x"34",
          2550 => x"0b",
          2551 => x"bb",
          2552 => x"fa",
          2553 => x"fa",
          2554 => x"fa",
          2555 => x"0b",
          2556 => x"bb",
          2557 => x"80",
          2558 => x"38",
          2559 => x"33",
          2560 => x"33",
          2561 => x"11",
          2562 => x"b2",
          2563 => x"70",
          2564 => x"33",
          2565 => x"7d",
          2566 => x"ff",
          2567 => x"38",
          2568 => x"7b",
          2569 => x"78",
          2570 => x"5f",
          2571 => x"c7",
          2572 => x"33",
          2573 => x"22",
          2574 => x"40",
          2575 => x"83",
          2576 => x"05",
          2577 => x"c7",
          2578 => x"33",
          2579 => x"22",
          2580 => x"11",
          2581 => x"b0",
          2582 => x"81",
          2583 => x"7c",
          2584 => x"f9",
          2585 => x"19",
          2586 => x"fa",
          2587 => x"ff",
          2588 => x"2e",
          2589 => x"d7",
          2590 => x"84",
          2591 => x"38",
          2592 => x"84",
          2593 => x"e0",
          2594 => x"83",
          2595 => x"e7",
          2596 => x"0c",
          2597 => x"33",
          2598 => x"06",
          2599 => x"06",
          2600 => x"80",
          2601 => x"72",
          2602 => x"06",
          2603 => x"5c",
          2604 => x"ef",
          2605 => x"7a",
          2606 => x"72",
          2607 => x"b9",
          2608 => x"34",
          2609 => x"33",
          2610 => x"12",
          2611 => x"fa",
          2612 => x"76",
          2613 => x"b0",
          2614 => x"84",
          2615 => x"83",
          2616 => x"72",
          2617 => x"59",
          2618 => x"18",
          2619 => x"06",
          2620 => x"38",
          2621 => x"fb",
          2622 => x"b5",
          2623 => x"5d",
          2624 => x"83",
          2625 => x"83",
          2626 => x"72",
          2627 => x"72",
          2628 => x"5b",
          2629 => x"a0",
          2630 => x"83",
          2631 => x"72",
          2632 => x"a0",
          2633 => x"fa",
          2634 => x"5e",
          2635 => x"80",
          2636 => x"81",
          2637 => x"fa",
          2638 => x"44",
          2639 => x"84",
          2640 => x"70",
          2641 => x"27",
          2642 => x"34",
          2643 => x"80",
          2644 => x"9c",
          2645 => x"33",
          2646 => x"34",
          2647 => x"06",
          2648 => x"81",
          2649 => x"84",
          2650 => x"83",
          2651 => x"80",
          2652 => x"33",
          2653 => x"33",
          2654 => x"39",
          2655 => x"11",
          2656 => x"3f",
          2657 => x"f0",
          2658 => x"57",
          2659 => x"10",
          2660 => x"05",
          2661 => x"fb",
          2662 => x"5c",
          2663 => x"83",
          2664 => x"83",
          2665 => x"e5",
          2666 => x"b4",
          2667 => x"29",
          2668 => x"19",
          2669 => x"34",
          2670 => x"33",
          2671 => x"12",
          2672 => x"b6",
          2673 => x"71",
          2674 => x"33",
          2675 => x"84",
          2676 => x"83",
          2677 => x"72",
          2678 => x"5a",
          2679 => x"1e",
          2680 => x"5c",
          2681 => x"84",
          2682 => x"38",
          2683 => x"34",
          2684 => x"b8",
          2685 => x"bd",
          2686 => x"f3",
          2687 => x"e4",
          2688 => x"9c",
          2689 => x"83",
          2690 => x"83",
          2691 => x"57",
          2692 => x"39",
          2693 => x"34",
          2694 => x"34",
          2695 => x"34",
          2696 => x"5b",
          2697 => x"ba",
          2698 => x"81",
          2699 => x"33",
          2700 => x"81",
          2701 => x"52",
          2702 => x"b0",
          2703 => x"84",
          2704 => x"f9",
          2705 => x"a0",
          2706 => x"f8",
          2707 => x"c0",
          2708 => x"5b",
          2709 => x"7b",
          2710 => x"ba",
          2711 => x"75",
          2712 => x"10",
          2713 => x"04",
          2714 => x"2e",
          2715 => x"84",
          2716 => x"09",
          2717 => x"59",
          2718 => x"fd",
          2719 => x"75",
          2720 => x"d9",
          2721 => x"84",
          2722 => x"7b",
          2723 => x"b5",
          2724 => x"fa",
          2725 => x"81",
          2726 => x"fd",
          2727 => x"fa",
          2728 => x"83",
          2729 => x"84",
          2730 => x"76",
          2731 => x"56",
          2732 => x"39",
          2733 => x"2e",
          2734 => x"84",
          2735 => x"09",
          2736 => x"59",
          2737 => x"fc",
          2738 => x"7a",
          2739 => x"d8",
          2740 => x"06",
          2741 => x"83",
          2742 => x"72",
          2743 => x"11",
          2744 => x"58",
          2745 => x"ff",
          2746 => x"fe",
          2747 => x"84",
          2748 => x"0b",
          2749 => x"84",
          2750 => x"fb",
          2751 => x"77",
          2752 => x"38",
          2753 => x"d0",
          2754 => x"80",
          2755 => x"33",
          2756 => x"84",
          2757 => x"56",
          2758 => x"76",
          2759 => x"84",
          2760 => x"8c",
          2761 => x"fa",
          2762 => x"f7",
          2763 => x"60",
          2764 => x"fa",
          2765 => x"cc",
          2766 => x"84",
          2767 => x"27",
          2768 => x"d8",
          2769 => x"ac",
          2770 => x"70",
          2771 => x"58",
          2772 => x"ba",
          2773 => x"8d",
          2774 => x"83",
          2775 => x"76",
          2776 => x"fa",
          2777 => x"81",
          2778 => x"db",
          2779 => x"84",
          2780 => x"ff",
          2781 => x"ff",
          2782 => x"59",
          2783 => x"77",
          2784 => x"81",
          2785 => x"7f",
          2786 => x"fa",
          2787 => x"11",
          2788 => x"38",
          2789 => x"f9",
          2790 => x"7e",
          2791 => x"d9",
          2792 => x"7a",
          2793 => x"b4",
          2794 => x"ff",
          2795 => x"29",
          2796 => x"fa",
          2797 => x"05",
          2798 => x"8a",
          2799 => x"60",
          2800 => x"ff",
          2801 => x"80",
          2802 => x"f7",
          2803 => x"38",
          2804 => x"23",
          2805 => x"41",
          2806 => x"84",
          2807 => x"8d",
          2808 => x"fa",
          2809 => x"fa",
          2810 => x"76",
          2811 => x"05",
          2812 => x"5c",
          2813 => x"80",
          2814 => x"ff",
          2815 => x"29",
          2816 => x"27",
          2817 => x"57",
          2818 => x"80",
          2819 => x"34",
          2820 => x"70",
          2821 => x"b8",
          2822 => x"71",
          2823 => x"60",
          2824 => x"33",
          2825 => x"70",
          2826 => x"05",
          2827 => x"34",
          2828 => x"b8",
          2829 => x"40",
          2830 => x"38",
          2831 => x"56",
          2832 => x"52",
          2833 => x"3f",
          2834 => x"f8",
          2835 => x"5d",
          2836 => x"38",
          2837 => x"2e",
          2838 => x"fa",
          2839 => x"83",
          2840 => x"76",
          2841 => x"f7",
          2842 => x"38",
          2843 => x"26",
          2844 => x"7d",
          2845 => x"7a",
          2846 => x"05",
          2847 => x"5d",
          2848 => x"83",
          2849 => x"38",
          2850 => x"38",
          2851 => x"71",
          2852 => x"71",
          2853 => x"77",
          2854 => x"84",
          2855 => x"05",
          2856 => x"84",
          2857 => x"41",
          2858 => x"ff",
          2859 => x"29",
          2860 => x"77",
          2861 => x"70",
          2862 => x"76",
          2863 => x"e0",
          2864 => x"d6",
          2865 => x"19",
          2866 => x"34",
          2867 => x"c0",
          2868 => x"79",
          2869 => x"17",
          2870 => x"a8",
          2871 => x"5d",
          2872 => x"33",
          2873 => x"80",
          2874 => x"5d",
          2875 => x"06",
          2876 => x"b0",
          2877 => x"59",
          2878 => x"17",
          2879 => x"7c",
          2880 => x"f8",
          2881 => x"f7",
          2882 => x"39",
          2883 => x"75",
          2884 => x"81",
          2885 => x"83",
          2886 => x"07",
          2887 => x"39",
          2888 => x"83",
          2889 => x"d4",
          2890 => x"06",
          2891 => x"34",
          2892 => x"9f",
          2893 => x"b0",
          2894 => x"83",
          2895 => x"ff",
          2896 => x"fa",
          2897 => x"83",
          2898 => x"fa",
          2899 => x"56",
          2900 => x"39",
          2901 => x"80",
          2902 => x"34",
          2903 => x"81",
          2904 => x"83",
          2905 => x"fa",
          2906 => x"56",
          2907 => x"39",
          2908 => x"86",
          2909 => x"fe",
          2910 => x"fc",
          2911 => x"b0",
          2912 => x"33",
          2913 => x"83",
          2914 => x"fa",
          2915 => x"83",
          2916 => x"fa",
          2917 => x"83",
          2918 => x"fa",
          2919 => x"83",
          2920 => x"fa",
          2921 => x"07",
          2922 => x"cc",
          2923 => x"06",
          2924 => x"34",
          2925 => x"b5",
          2926 => x"3f",
          2927 => x"83",
          2928 => x"83",
          2929 => x"59",
          2930 => x"84",
          2931 => x"0b",
          2932 => x"bb",
          2933 => x"83",
          2934 => x"70",
          2935 => x"e7",
          2936 => x"3d",
          2937 => x"f7",
          2938 => x"38",
          2939 => x"0c",
          2940 => x"0b",
          2941 => x"04",
          2942 => x"39",
          2943 => x"5c",
          2944 => x"83",
          2945 => x"22",
          2946 => x"84",
          2947 => x"83",
          2948 => x"d1",
          2949 => x"81",
          2950 => x"d8",
          2951 => x"80",
          2952 => x"98",
          2953 => x"ef",
          2954 => x"05",
          2955 => x"58",
          2956 => x"81",
          2957 => x"40",
          2958 => x"83",
          2959 => x"fa",
          2960 => x"9f",
          2961 => x"e2",
          2962 => x"84",
          2963 => x"56",
          2964 => x"57",
          2965 => x"70",
          2966 => x"26",
          2967 => x"84",
          2968 => x"83",
          2969 => x"86",
          2970 => x"22",
          2971 => x"83",
          2972 => x"5d",
          2973 => x"2e",
          2974 => x"06",
          2975 => x"84",
          2976 => x"76",
          2977 => x"56",
          2978 => x"ff",
          2979 => x"24",
          2980 => x"56",
          2981 => x"16",
          2982 => x"81",
          2983 => x"57",
          2984 => x"75",
          2985 => x"06",
          2986 => x"58",
          2987 => x"b0",
          2988 => x"ff",
          2989 => x"42",
          2990 => x"84",
          2991 => x"33",
          2992 => x"70",
          2993 => x"05",
          2994 => x"34",
          2995 => x"b8",
          2996 => x"41",
          2997 => x"38",
          2998 => x"80",
          2999 => x"34",
          3000 => x"70",
          3001 => x"b8",
          3002 => x"71",
          3003 => x"78",
          3004 => x"83",
          3005 => x"80",
          3006 => x"33",
          3007 => x"22",
          3008 => x"5d",
          3009 => x"84",
          3010 => x"ff",
          3011 => x"83",
          3012 => x"23",
          3013 => x"5a",
          3014 => x"76",
          3015 => x"33",
          3016 => x"59",
          3017 => x"80",
          3018 => x"88",
          3019 => x"84",
          3020 => x"56",
          3021 => x"57",
          3022 => x"81",
          3023 => x"33",
          3024 => x"33",
          3025 => x"2e",
          3026 => x"a1",
          3027 => x"b4",
          3028 => x"75",
          3029 => x"7c",
          3030 => x"34",
          3031 => x"77",
          3032 => x"70",
          3033 => x"33",
          3034 => x"7a",
          3035 => x"81",
          3036 => x"77",
          3037 => x"27",
          3038 => x"31",
          3039 => x"a8",
          3040 => x"fc",
          3041 => x"fc",
          3042 => x"23",
          3043 => x"b4",
          3044 => x"18",
          3045 => x"77",
          3046 => x"e9",
          3047 => x"05",
          3048 => x"72",
          3049 => x"9c",
          3050 => x"85",
          3051 => x"d7",
          3052 => x"0c",
          3053 => x"02",
          3054 => x"f9",
          3055 => x"f8",
          3056 => x"74",
          3057 => x"56",
          3058 => x"78",
          3059 => x"04",
          3060 => x"73",
          3061 => x"70",
          3062 => x"2a",
          3063 => x"e4",
          3064 => x"2e",
          3065 => x"7b",
          3066 => x"76",
          3067 => x"85",
          3068 => x"fa",
          3069 => x"71",
          3070 => x"83",
          3071 => x"79",
          3072 => x"83",
          3073 => x"74",
          3074 => x"54",
          3075 => x"0b",
          3076 => x"98",
          3077 => x"38",
          3078 => x"83",
          3079 => x"81",
          3080 => x"27",
          3081 => x"14",
          3082 => x"ae",
          3083 => x"2e",
          3084 => x"86",
          3085 => x"34",
          3086 => x"ff",
          3087 => x"c2",
          3088 => x"83",
          3089 => x"81",
          3090 => x"ff",
          3091 => x"98",
          3092 => x"75",
          3093 => x"06",
          3094 => x"06",
          3095 => x"e7",
          3096 => x"73",
          3097 => x"85",
          3098 => x"34",
          3099 => x"f8",
          3100 => x"83",
          3101 => x"5d",
          3102 => x"f8",
          3103 => x"2e",
          3104 => x"54",
          3105 => x"f8",
          3106 => x"2e",
          3107 => x"54",
          3108 => x"06",
          3109 => x"83",
          3110 => x"2e",
          3111 => x"53",
          3112 => x"83",
          3113 => x"27",
          3114 => x"87",
          3115 => x"54",
          3116 => x"81",
          3117 => x"f8",
          3118 => x"ff",
          3119 => x"f6",
          3120 => x"83",
          3121 => x"72",
          3122 => x"10",
          3123 => x"04",
          3124 => x"2e",
          3125 => x"98",
          3126 => x"fc",
          3127 => x"33",
          3128 => x"74",
          3129 => x"c0",
          3130 => x"73",
          3131 => x"94",
          3132 => x"84",
          3133 => x"f0",
          3134 => x"08",
          3135 => x"72",
          3136 => x"76",
          3137 => x"80",
          3138 => x"57",
          3139 => x"79",
          3140 => x"38",
          3141 => x"81",
          3142 => x"06",
          3143 => x"54",
          3144 => x"80",
          3145 => x"ff",
          3146 => x"72",
          3147 => x"58",
          3148 => x"10",
          3149 => x"83",
          3150 => x"70",
          3151 => x"98",
          3152 => x"fd",
          3153 => x"ff",
          3154 => x"ff",
          3155 => x"78",
          3156 => x"84",
          3157 => x"2e",
          3158 => x"30",
          3159 => x"56",
          3160 => x"81",
          3161 => x"f9",
          3162 => x"10",
          3163 => x"54",
          3164 => x"13",
          3165 => x"73",
          3166 => x"53",
          3167 => x"b8",
          3168 => x"78",
          3169 => x"d4",
          3170 => x"3d",
          3171 => x"54",
          3172 => x"92",
          3173 => x"05",
          3174 => x"fa",
          3175 => x"15",
          3176 => x"34",
          3177 => x"fa",
          3178 => x"72",
          3179 => x"f8",
          3180 => x"fc",
          3181 => x"73",
          3182 => x"38",
          3183 => x"87",
          3184 => x"73",
          3185 => x"9c",
          3186 => x"ff",
          3187 => x"83",
          3188 => x"72",
          3189 => x"06",
          3190 => x"f8",
          3191 => x"33",
          3192 => x"33",
          3193 => x"df",
          3194 => x"56",
          3195 => x"81",
          3196 => x"81",
          3197 => x"09",
          3198 => x"39",
          3199 => x"98",
          3200 => x"57",
          3201 => x"84",
          3202 => x"39",
          3203 => x"54",
          3204 => x"b8",
          3205 => x"81",
          3206 => x"f7",
          3207 => x"0c",
          3208 => x"70",
          3209 => x"54",
          3210 => x"74",
          3211 => x"06",
          3212 => x"83",
          3213 => x"34",
          3214 => x"06",
          3215 => x"83",
          3216 => x"34",
          3217 => x"83",
          3218 => x"f6",
          3219 => x"84",
          3220 => x"fe",
          3221 => x"88",
          3222 => x"bb",
          3223 => x"ac",
          3224 => x"0d",
          3225 => x"57",
          3226 => x"83",
          3227 => x"34",
          3228 => x"56",
          3229 => x"87",
          3230 => x"9c",
          3231 => x"ce",
          3232 => x"08",
          3233 => x"70",
          3234 => x"87",
          3235 => x"73",
          3236 => x"db",
          3237 => x"ff",
          3238 => x"71",
          3239 => x"87",
          3240 => x"05",
          3241 => x"87",
          3242 => x"2e",
          3243 => x"98",
          3244 => x"87",
          3245 => x"87",
          3246 => x"26",
          3247 => x"16",
          3248 => x"80",
          3249 => x"52",
          3250 => x"8a",
          3251 => x"3d",
          3252 => x"0c",
          3253 => x"79",
          3254 => x"52",
          3255 => x"88",
          3256 => x"75",
          3257 => x"71",
          3258 => x"70",
          3259 => x"75",
          3260 => x"83",
          3261 => x"34",
          3262 => x"71",
          3263 => x"55",
          3264 => x"0b",
          3265 => x"98",
          3266 => x"80",
          3267 => x"9c",
          3268 => x"51",
          3269 => x"33",
          3270 => x"74",
          3271 => x"2e",
          3272 => x"51",
          3273 => x"38",
          3274 => x"38",
          3275 => x"90",
          3276 => x"52",
          3277 => x"72",
          3278 => x"c0",
          3279 => x"27",
          3280 => x"38",
          3281 => x"75",
          3282 => x"ff",
          3283 => x"75",
          3284 => x"ff",
          3285 => x"51",
          3286 => x"38",
          3287 => x"55",
          3288 => x"71",
          3289 => x"81",
          3290 => x"38",
          3291 => x"0d",
          3292 => x"88",
          3293 => x"fa",
          3294 => x"05",
          3295 => x"90",
          3296 => x"80",
          3297 => x"55",
          3298 => x"90",
          3299 => x"90",
          3300 => x"86",
          3301 => x"80",
          3302 => x"55",
          3303 => x"70",
          3304 => x"05",
          3305 => x"83",
          3306 => x"34",
          3307 => x"75",
          3308 => x"55",
          3309 => x"0b",
          3310 => x"98",
          3311 => x"80",
          3312 => x"9c",
          3313 => x"51",
          3314 => x"33",
          3315 => x"74",
          3316 => x"2e",
          3317 => x"51",
          3318 => x"38",
          3319 => x"38",
          3320 => x"90",
          3321 => x"52",
          3322 => x"72",
          3323 => x"c0",
          3324 => x"27",
          3325 => x"38",
          3326 => x"75",
          3327 => x"ff",
          3328 => x"75",
          3329 => x"06",
          3330 => x"70",
          3331 => x"83",
          3332 => x"0c",
          3333 => x"39",
          3334 => x"51",
          3335 => x"f5",
          3336 => x"16",
          3337 => x"34",
          3338 => x"90",
          3339 => x"87",
          3340 => x"98",
          3341 => x"38",
          3342 => x"08",
          3343 => x"71",
          3344 => x"98",
          3345 => x"27",
          3346 => x"2e",
          3347 => x"08",
          3348 => x"98",
          3349 => x"08",
          3350 => x"15",
          3351 => x"52",
          3352 => x"ff",
          3353 => x"08",
          3354 => x"52",
          3355 => x"06",
          3356 => x"72",
          3357 => x"38",
          3358 => x"88",
          3359 => x"0d",
          3360 => x"08",
          3361 => x"ff",
          3362 => x"70",
          3363 => x"71",
          3364 => x"81",
          3365 => x"2b",
          3366 => x"57",
          3367 => x"24",
          3368 => x"33",
          3369 => x"83",
          3370 => x"12",
          3371 => x"07",
          3372 => x"80",
          3373 => x"33",
          3374 => x"83",
          3375 => x"52",
          3376 => x"73",
          3377 => x"34",
          3378 => x"12",
          3379 => x"07",
          3380 => x"51",
          3381 => x"34",
          3382 => x"0b",
          3383 => x"34",
          3384 => x"14",
          3385 => x"f4",
          3386 => x"71",
          3387 => x"70",
          3388 => x"72",
          3389 => x"0d",
          3390 => x"71",
          3391 => x"11",
          3392 => x"88",
          3393 => x"54",
          3394 => x"34",
          3395 => x"08",
          3396 => x"33",
          3397 => x"56",
          3398 => x"33",
          3399 => x"70",
          3400 => x"86",
          3401 => x"ba",
          3402 => x"33",
          3403 => x"06",
          3404 => x"76",
          3405 => x"ba",
          3406 => x"12",
          3407 => x"07",
          3408 => x"71",
          3409 => x"ff",
          3410 => x"54",
          3411 => x"52",
          3412 => x"34",
          3413 => x"33",
          3414 => x"83",
          3415 => x"12",
          3416 => x"ff",
          3417 => x"55",
          3418 => x"70",
          3419 => x"70",
          3420 => x"71",
          3421 => x"05",
          3422 => x"2b",
          3423 => x"52",
          3424 => x"fc",
          3425 => x"71",
          3426 => x"70",
          3427 => x"34",
          3428 => x"08",
          3429 => x"71",
          3430 => x"05",
          3431 => x"88",
          3432 => x"5c",
          3433 => x"15",
          3434 => x"0d",
          3435 => x"f4",
          3436 => x"38",
          3437 => x"fb",
          3438 => x"ff",
          3439 => x"80",
          3440 => x"80",
          3441 => x"fe",
          3442 => x"55",
          3443 => x"34",
          3444 => x"15",
          3445 => x"ba",
          3446 => x"81",
          3447 => x"08",
          3448 => x"80",
          3449 => x"70",
          3450 => x"88",
          3451 => x"ba",
          3452 => x"ba",
          3453 => x"76",
          3454 => x"34",
          3455 => x"52",
          3456 => x"8e",
          3457 => x"70",
          3458 => x"83",
          3459 => x"84",
          3460 => x"2b",
          3461 => x"81",
          3462 => x"cc",
          3463 => x"33",
          3464 => x"70",
          3465 => x"83",
          3466 => x"53",
          3467 => x"8a",
          3468 => x"73",
          3469 => x"33",
          3470 => x"c1",
          3471 => x"38",
          3472 => x"2b",
          3473 => x"71",
          3474 => x"06",
          3475 => x"79",
          3476 => x"74",
          3477 => x"78",
          3478 => x"2e",
          3479 => x"2b",
          3480 => x"70",
          3481 => x"76",
          3482 => x"ba",
          3483 => x"53",
          3484 => x"34",
          3485 => x"33",
          3486 => x"70",
          3487 => x"05",
          3488 => x"2a",
          3489 => x"75",
          3490 => x"53",
          3491 => x"08",
          3492 => x"15",
          3493 => x"86",
          3494 => x"2b",
          3495 => x"5c",
          3496 => x"72",
          3497 => x"70",
          3498 => x"87",
          3499 => x"88",
          3500 => x"15",
          3501 => x"f4",
          3502 => x"12",
          3503 => x"07",
          3504 => x"75",
          3505 => x"84",
          3506 => x"05",
          3507 => x"88",
          3508 => x"57",
          3509 => x"15",
          3510 => x"05",
          3511 => x"3d",
          3512 => x"33",
          3513 => x"79",
          3514 => x"71",
          3515 => x"5b",
          3516 => x"34",
          3517 => x"08",
          3518 => x"33",
          3519 => x"74",
          3520 => x"71",
          3521 => x"5d",
          3522 => x"86",
          3523 => x"ba",
          3524 => x"33",
          3525 => x"06",
          3526 => x"75",
          3527 => x"ba",
          3528 => x"f1",
          3529 => x"f4",
          3530 => x"38",
          3531 => x"bb",
          3532 => x"51",
          3533 => x"84",
          3534 => x"84",
          3535 => x"a0",
          3536 => x"80",
          3537 => x"51",
          3538 => x"08",
          3539 => x"16",
          3540 => x"84",
          3541 => x"84",
          3542 => x"34",
          3543 => x"f4",
          3544 => x"fe",
          3545 => x"06",
          3546 => x"74",
          3547 => x"84",
          3548 => x"84",
          3549 => x"55",
          3550 => x"15",
          3551 => x"dd",
          3552 => x"65",
          3553 => x"f4",
          3554 => x"84",
          3555 => x"38",
          3556 => x"54",
          3557 => x"05",
          3558 => x"ff",
          3559 => x"06",
          3560 => x"ff",
          3561 => x"70",
          3562 => x"07",
          3563 => x"06",
          3564 => x"83",
          3565 => x"33",
          3566 => x"70",
          3567 => x"53",
          3568 => x"5e",
          3569 => x"38",
          3570 => x"88",
          3571 => x"70",
          3572 => x"71",
          3573 => x"56",
          3574 => x"7a",
          3575 => x"58",
          3576 => x"80",
          3577 => x"77",
          3578 => x"59",
          3579 => x"1e",
          3580 => x"2b",
          3581 => x"33",
          3582 => x"90",
          3583 => x"57",
          3584 => x"38",
          3585 => x"33",
          3586 => x"7a",
          3587 => x"71",
          3588 => x"05",
          3589 => x"88",
          3590 => x"48",
          3591 => x"56",
          3592 => x"34",
          3593 => x"11",
          3594 => x"71",
          3595 => x"33",
          3596 => x"70",
          3597 => x"57",
          3598 => x"87",
          3599 => x"70",
          3600 => x"07",
          3601 => x"5a",
          3602 => x"81",
          3603 => x"1f",
          3604 => x"8b",
          3605 => x"73",
          3606 => x"07",
          3607 => x"5f",
          3608 => x"81",
          3609 => x"1f",
          3610 => x"2b",
          3611 => x"14",
          3612 => x"07",
          3613 => x"5f",
          3614 => x"75",
          3615 => x"70",
          3616 => x"71",
          3617 => x"70",
          3618 => x"05",
          3619 => x"84",
          3620 => x"65",
          3621 => x"5d",
          3622 => x"38",
          3623 => x"95",
          3624 => x"84",
          3625 => x"ba",
          3626 => x"52",
          3627 => x"3f",
          3628 => x"34",
          3629 => x"f4",
          3630 => x"0b",
          3631 => x"5c",
          3632 => x"1d",
          3633 => x"f0",
          3634 => x"70",
          3635 => x"5c",
          3636 => x"77",
          3637 => x"70",
          3638 => x"05",
          3639 => x"34",
          3640 => x"f4",
          3641 => x"80",
          3642 => x"80",
          3643 => x"9b",
          3644 => x"84",
          3645 => x"84",
          3646 => x"11",
          3647 => x"12",
          3648 => x"ff",
          3649 => x"5e",
          3650 => x"34",
          3651 => x"88",
          3652 => x"7b",
          3653 => x"70",
          3654 => x"88",
          3655 => x"f8",
          3656 => x"06",
          3657 => x"5e",
          3658 => x"76",
          3659 => x"05",
          3660 => x"63",
          3661 => x"84",
          3662 => x"ed",
          3663 => x"7b",
          3664 => x"42",
          3665 => x"ff",
          3666 => x"06",
          3667 => x"88",
          3668 => x"70",
          3669 => x"71",
          3670 => x"58",
          3671 => x"f7",
          3672 => x"fa",
          3673 => x"38",
          3674 => x"7b",
          3675 => x"84",
          3676 => x"a0",
          3677 => x"80",
          3678 => x"51",
          3679 => x"08",
          3680 => x"1b",
          3681 => x"84",
          3682 => x"84",
          3683 => x"34",
          3684 => x"f4",
          3685 => x"fe",
          3686 => x"06",
          3687 => x"74",
          3688 => x"05",
          3689 => x"10",
          3690 => x"05",
          3691 => x"81",
          3692 => x"80",
          3693 => x"ff",
          3694 => x"c0",
          3695 => x"82",
          3696 => x"7f",
          3697 => x"3d",
          3698 => x"83",
          3699 => x"2b",
          3700 => x"12",
          3701 => x"07",
          3702 => x"33",
          3703 => x"43",
          3704 => x"5c",
          3705 => x"7a",
          3706 => x"08",
          3707 => x"33",
          3708 => x"74",
          3709 => x"71",
          3710 => x"41",
          3711 => x"64",
          3712 => x"34",
          3713 => x"81",
          3714 => x"ff",
          3715 => x"5a",
          3716 => x"34",
          3717 => x"11",
          3718 => x"71",
          3719 => x"81",
          3720 => x"88",
          3721 => x"45",
          3722 => x"34",
          3723 => x"33",
          3724 => x"83",
          3725 => x"83",
          3726 => x"88",
          3727 => x"55",
          3728 => x"18",
          3729 => x"82",
          3730 => x"2b",
          3731 => x"2b",
          3732 => x"05",
          3733 => x"f4",
          3734 => x"ff",
          3735 => x"ff",
          3736 => x"80",
          3737 => x"80",
          3738 => x"fe",
          3739 => x"56",
          3740 => x"34",
          3741 => x"16",
          3742 => x"ba",
          3743 => x"81",
          3744 => x"08",
          3745 => x"80",
          3746 => x"70",
          3747 => x"88",
          3748 => x"ba",
          3749 => x"ba",
          3750 => x"7f",
          3751 => x"34",
          3752 => x"fc",
          3753 => x"33",
          3754 => x"79",
          3755 => x"71",
          3756 => x"48",
          3757 => x"05",
          3758 => x"ba",
          3759 => x"85",
          3760 => x"2b",
          3761 => x"15",
          3762 => x"2a",
          3763 => x"40",
          3764 => x"87",
          3765 => x"70",
          3766 => x"07",
          3767 => x"59",
          3768 => x"81",
          3769 => x"1f",
          3770 => x"2b",
          3771 => x"33",
          3772 => x"70",
          3773 => x"05",
          3774 => x"5d",
          3775 => x"34",
          3776 => x"08",
          3777 => x"71",
          3778 => x"05",
          3779 => x"2b",
          3780 => x"2a",
          3781 => x"5b",
          3782 => x"34",
          3783 => x"b3",
          3784 => x"71",
          3785 => x"05",
          3786 => x"88",
          3787 => x"5a",
          3788 => x"79",
          3789 => x"70",
          3790 => x"71",
          3791 => x"05",
          3792 => x"88",
          3793 => x"5e",
          3794 => x"86",
          3795 => x"84",
          3796 => x"12",
          3797 => x"ff",
          3798 => x"55",
          3799 => x"84",
          3800 => x"81",
          3801 => x"2b",
          3802 => x"33",
          3803 => x"8f",
          3804 => x"2a",
          3805 => x"5e",
          3806 => x"17",
          3807 => x"70",
          3808 => x"71",
          3809 => x"81",
          3810 => x"ff",
          3811 => x"5e",
          3812 => x"34",
          3813 => x"08",
          3814 => x"33",
          3815 => x"74",
          3816 => x"71",
          3817 => x"05",
          3818 => x"88",
          3819 => x"49",
          3820 => x"57",
          3821 => x"1d",
          3822 => x"84",
          3823 => x"2b",
          3824 => x"14",
          3825 => x"07",
          3826 => x"40",
          3827 => x"7b",
          3828 => x"16",
          3829 => x"2b",
          3830 => x"2a",
          3831 => x"79",
          3832 => x"70",
          3833 => x"71",
          3834 => x"05",
          3835 => x"2b",
          3836 => x"5d",
          3837 => x"75",
          3838 => x"70",
          3839 => x"8b",
          3840 => x"82",
          3841 => x"2b",
          3842 => x"5d",
          3843 => x"34",
          3844 => x"08",
          3845 => x"33",
          3846 => x"56",
          3847 => x"7e",
          3848 => x"3f",
          3849 => x"61",
          3850 => x"06",
          3851 => x"19",
          3852 => x"71",
          3853 => x"33",
          3854 => x"70",
          3855 => x"55",
          3856 => x"85",
          3857 => x"1e",
          3858 => x"8b",
          3859 => x"86",
          3860 => x"2b",
          3861 => x"48",
          3862 => x"05",
          3863 => x"ba",
          3864 => x"33",
          3865 => x"06",
          3866 => x"78",
          3867 => x"ba",
          3868 => x"12",
          3869 => x"07",
          3870 => x"71",
          3871 => x"ff",
          3872 => x"5d",
          3873 => x"40",
          3874 => x"34",
          3875 => x"33",
          3876 => x"83",
          3877 => x"12",
          3878 => x"ff",
          3879 => x"58",
          3880 => x"78",
          3881 => x"06",
          3882 => x"54",
          3883 => x"5f",
          3884 => x"38",
          3885 => x"08",
          3886 => x"df",
          3887 => x"ef",
          3888 => x"0d",
          3889 => x"58",
          3890 => x"54",
          3891 => x"0c",
          3892 => x"d3",
          3893 => x"bb",
          3894 => x"53",
          3895 => x"fe",
          3896 => x"0c",
          3897 => x"0b",
          3898 => x"84",
          3899 => x"76",
          3900 => x"97",
          3901 => x"75",
          3902 => x"ba",
          3903 => x"81",
          3904 => x"08",
          3905 => x"87",
          3906 => x"ba",
          3907 => x"07",
          3908 => x"2a",
          3909 => x"34",
          3910 => x"22",
          3911 => x"08",
          3912 => x"15",
          3913 => x"54",
          3914 => x"cc",
          3915 => x"33",
          3916 => x"38",
          3917 => x"84",
          3918 => x"fe",
          3919 => x"83",
          3920 => x"51",
          3921 => x"81",
          3922 => x"84",
          3923 => x"12",
          3924 => x"84",
          3925 => x"7e",
          3926 => x"5a",
          3927 => x"26",
          3928 => x"54",
          3929 => x"bd",
          3930 => x"98",
          3931 => x"51",
          3932 => x"81",
          3933 => x"38",
          3934 => x"e2",
          3935 => x"fc",
          3936 => x"83",
          3937 => x"bb",
          3938 => x"80",
          3939 => x"5a",
          3940 => x"38",
          3941 => x"60",
          3942 => x"5c",
          3943 => x"87",
          3944 => x"73",
          3945 => x"38",
          3946 => x"8c",
          3947 => x"d7",
          3948 => x"ff",
          3949 => x"87",
          3950 => x"38",
          3951 => x"80",
          3952 => x"38",
          3953 => x"84",
          3954 => x"16",
          3955 => x"55",
          3956 => x"d5",
          3957 => x"05",
          3958 => x"05",
          3959 => x"73",
          3960 => x"33",
          3961 => x"73",
          3962 => x"8c",
          3963 => x"38",
          3964 => x"2e",
          3965 => x"84",
          3966 => x"0a",
          3967 => x"86",
          3968 => x"80",
          3969 => x"0d",
          3970 => x"8c",
          3971 => x"08",
          3972 => x"70",
          3973 => x"8c",
          3974 => x"98",
          3975 => x"72",
          3976 => x"71",
          3977 => x"ff",
          3978 => x"73",
          3979 => x"0d",
          3980 => x"71",
          3981 => x"81",
          3982 => x"83",
          3983 => x"52",
          3984 => x"84",
          3985 => x"81",
          3986 => x"3d",
          3987 => x"53",
          3988 => x"52",
          3989 => x"bb",
          3990 => x"d9",
          3991 => x"34",
          3992 => x"31",
          3993 => x"5c",
          3994 => x"9b",
          3995 => x"2e",
          3996 => x"54",
          3997 => x"33",
          3998 => x"57",
          3999 => x"fe",
          4000 => x"81",
          4001 => x"b8",
          4002 => x"80",
          4003 => x"17",
          4004 => x"84",
          4005 => x"b7",
          4006 => x"d2",
          4007 => x"ba",
          4008 => x"34",
          4009 => x"80",
          4010 => x"c1",
          4011 => x"0b",
          4012 => x"55",
          4013 => x"2a",
          4014 => x"90",
          4015 => x"74",
          4016 => x"34",
          4017 => x"19",
          4018 => x"a5",
          4019 => x"84",
          4020 => x"74",
          4021 => x"81",
          4022 => x"54",
          4023 => x"51",
          4024 => x"80",
          4025 => x"fb",
          4026 => x"2e",
          4027 => x"3d",
          4028 => x"56",
          4029 => x"08",
          4030 => x"84",
          4031 => x"ff",
          4032 => x"81",
          4033 => x"38",
          4034 => x"38",
          4035 => x"a8",
          4036 => x"b4",
          4037 => x"17",
          4038 => x"06",
          4039 => x"b8",
          4040 => x"e3",
          4041 => x"85",
          4042 => x"18",
          4043 => x"ff",
          4044 => x"70",
          4045 => x"5d",
          4046 => x"b5",
          4047 => x"5c",
          4048 => x"06",
          4049 => x"b8",
          4050 => x"93",
          4051 => x"85",
          4052 => x"18",
          4053 => x"ff",
          4054 => x"2b",
          4055 => x"2a",
          4056 => x"ae",
          4057 => x"84",
          4058 => x"2a",
          4059 => x"08",
          4060 => x"18",
          4061 => x"2e",
          4062 => x"54",
          4063 => x"33",
          4064 => x"08",
          4065 => x"5a",
          4066 => x"38",
          4067 => x"b8",
          4068 => x"88",
          4069 => x"5b",
          4070 => x"09",
          4071 => x"2a",
          4072 => x"08",
          4073 => x"18",
          4074 => x"2e",
          4075 => x"54",
          4076 => x"33",
          4077 => x"08",
          4078 => x"5a",
          4079 => x"38",
          4080 => x"05",
          4081 => x"33",
          4082 => x"81",
          4083 => x"75",
          4084 => x"06",
          4085 => x"5e",
          4086 => x"81",
          4087 => x"70",
          4088 => x"e2",
          4089 => x"7b",
          4090 => x"84",
          4091 => x"17",
          4092 => x"84",
          4093 => x"27",
          4094 => x"74",
          4095 => x"38",
          4096 => x"08",
          4097 => x"51",
          4098 => x"39",
          4099 => x"17",
          4100 => x"f6",
          4101 => x"2e",
          4102 => x"bb",
          4103 => x"08",
          4104 => x"18",
          4105 => x"5e",
          4106 => x"bb",
          4107 => x"54",
          4108 => x"53",
          4109 => x"3f",
          4110 => x"2e",
          4111 => x"bb",
          4112 => x"08",
          4113 => x"08",
          4114 => x"fd",
          4115 => x"82",
          4116 => x"81",
          4117 => x"05",
          4118 => x"f4",
          4119 => x"81",
          4120 => x"70",
          4121 => x"da",
          4122 => x"7d",
          4123 => x"84",
          4124 => x"17",
          4125 => x"84",
          4126 => x"27",
          4127 => x"74",
          4128 => x"38",
          4129 => x"08",
          4130 => x"51",
          4131 => x"39",
          4132 => x"08",
          4133 => x"51",
          4134 => x"5b",
          4135 => x"f2",
          4136 => x"59",
          4137 => x"75",
          4138 => x"33",
          4139 => x"78",
          4140 => x"82",
          4141 => x"90",
          4142 => x"1a",
          4143 => x"08",
          4144 => x"38",
          4145 => x"7c",
          4146 => x"81",
          4147 => x"19",
          4148 => x"84",
          4149 => x"81",
          4150 => x"79",
          4151 => x"06",
          4152 => x"58",
          4153 => x"2a",
          4154 => x"83",
          4155 => x"90",
          4156 => x"81",
          4157 => x"a8",
          4158 => x"1a",
          4159 => x"e1",
          4160 => x"7c",
          4161 => x"38",
          4162 => x"81",
          4163 => x"bb",
          4164 => x"58",
          4165 => x"58",
          4166 => x"83",
          4167 => x"11",
          4168 => x"7e",
          4169 => x"5c",
          4170 => x"75",
          4171 => x"79",
          4172 => x"7a",
          4173 => x"34",
          4174 => x"70",
          4175 => x"1b",
          4176 => x"b7",
          4177 => x"5e",
          4178 => x"06",
          4179 => x"b8",
          4180 => x"83",
          4181 => x"85",
          4182 => x"1a",
          4183 => x"79",
          4184 => x"1b",
          4185 => x"55",
          4186 => x"2b",
          4187 => x"71",
          4188 => x"0b",
          4189 => x"1a",
          4190 => x"08",
          4191 => x"38",
          4192 => x"53",
          4193 => x"3f",
          4194 => x"2e",
          4195 => x"bb",
          4196 => x"08",
          4197 => x"08",
          4198 => x"5c",
          4199 => x"33",
          4200 => x"81",
          4201 => x"33",
          4202 => x"08",
          4203 => x"58",
          4204 => x"38",
          4205 => x"7b",
          4206 => x"7a",
          4207 => x"71",
          4208 => x"34",
          4209 => x"39",
          4210 => x"53",
          4211 => x"3f",
          4212 => x"2e",
          4213 => x"bb",
          4214 => x"08",
          4215 => x"08",
          4216 => x"5e",
          4217 => x"19",
          4218 => x"06",
          4219 => x"53",
          4220 => x"c2",
          4221 => x"54",
          4222 => x"1a",
          4223 => x"5c",
          4224 => x"81",
          4225 => x"08",
          4226 => x"a8",
          4227 => x"bb",
          4228 => x"7e",
          4229 => x"55",
          4230 => x"e3",
          4231 => x"52",
          4232 => x"7c",
          4233 => x"53",
          4234 => x"52",
          4235 => x"bb",
          4236 => x"fb",
          4237 => x"1a",
          4238 => x"08",
          4239 => x"08",
          4240 => x"fb",
          4241 => x"82",
          4242 => x"81",
          4243 => x"19",
          4244 => x"fa",
          4245 => x"76",
          4246 => x"3f",
          4247 => x"10",
          4248 => x"ff",
          4249 => x"1f",
          4250 => x"1f",
          4251 => x"88",
          4252 => x"06",
          4253 => x"70",
          4254 => x"0a",
          4255 => x"7d",
          4256 => x"b9",
          4257 => x"ba",
          4258 => x"bb",
          4259 => x"0d",
          4260 => x"7a",
          4261 => x"76",
          4262 => x"1a",
          4263 => x"08",
          4264 => x"d7",
          4265 => x"76",
          4266 => x"76",
          4267 => x"26",
          4268 => x"f0",
          4269 => x"2e",
          4270 => x"84",
          4271 => x"84",
          4272 => x"80",
          4273 => x"55",
          4274 => x"09",
          4275 => x"74",
          4276 => x"04",
          4277 => x"84",
          4278 => x"51",
          4279 => x"bb",
          4280 => x"84",
          4281 => x"2e",
          4282 => x"84",
          4283 => x"dd",
          4284 => x"76",
          4285 => x"79",
          4286 => x"bb",
          4287 => x"84",
          4288 => x"72",
          4289 => x"bb",
          4290 => x"73",
          4291 => x"80",
          4292 => x"81",
          4293 => x"1a",
          4294 => x"57",
          4295 => x"fe",
          4296 => x"51",
          4297 => x"84",
          4298 => x"84",
          4299 => x"7a",
          4300 => x"75",
          4301 => x"05",
          4302 => x"26",
          4303 => x"84",
          4304 => x"1a",
          4305 => x"0c",
          4306 => x"bb",
          4307 => x"bb",
          4308 => x"80",
          4309 => x"52",
          4310 => x"84",
          4311 => x"84",
          4312 => x"0d",
          4313 => x"b9",
          4314 => x"3d",
          4315 => x"58",
          4316 => x"38",
          4317 => x"38",
          4318 => x"55",
          4319 => x"75",
          4320 => x"2a",
          4321 => x"56",
          4322 => x"08",
          4323 => x"98",
          4324 => x"2e",
          4325 => x"19",
          4326 => x"05",
          4327 => x"bb",
          4328 => x"0b",
          4329 => x"04",
          4330 => x"ff",
          4331 => x"2b",
          4332 => x"9c",
          4333 => x"54",
          4334 => x"38",
          4335 => x"19",
          4336 => x"0c",
          4337 => x"ec",
          4338 => x"84",
          4339 => x"81",
          4340 => x"9e",
          4341 => x"84",
          4342 => x"76",
          4343 => x"ff",
          4344 => x"0c",
          4345 => x"7f",
          4346 => x"5c",
          4347 => x"86",
          4348 => x"17",
          4349 => x"b2",
          4350 => x"9d",
          4351 => x"58",
          4352 => x"1a",
          4353 => x"f5",
          4354 => x"18",
          4355 => x"0c",
          4356 => x"8f",
          4357 => x"8a",
          4358 => x"06",
          4359 => x"51",
          4360 => x"5d",
          4361 => x"08",
          4362 => x"84",
          4363 => x"08",
          4364 => x"38",
          4365 => x"17",
          4366 => x"84",
          4367 => x"bb",
          4368 => x"82",
          4369 => x"ff",
          4370 => x"08",
          4371 => x"84",
          4372 => x"80",
          4373 => x"fe",
          4374 => x"27",
          4375 => x"29",
          4376 => x"b4",
          4377 => x"78",
          4378 => x"58",
          4379 => x"74",
          4380 => x"27",
          4381 => x"53",
          4382 => x"b2",
          4383 => x"38",
          4384 => x"18",
          4385 => x"8f",
          4386 => x"08",
          4387 => x"33",
          4388 => x"84",
          4389 => x"08",
          4390 => x"1a",
          4391 => x"27",
          4392 => x"7b",
          4393 => x"38",
          4394 => x"08",
          4395 => x"51",
          4396 => x"19",
          4397 => x"55",
          4398 => x"38",
          4399 => x"1a",
          4400 => x"75",
          4401 => x"22",
          4402 => x"98",
          4403 => x"0b",
          4404 => x"04",
          4405 => x"84",
          4406 => x"98",
          4407 => x"2e",
          4408 => x"5a",
          4409 => x"82",
          4410 => x"55",
          4411 => x"94",
          4412 => x"52",
          4413 => x"84",
          4414 => x"ff",
          4415 => x"76",
          4416 => x"08",
          4417 => x"82",
          4418 => x"70",
          4419 => x"1d",
          4420 => x"78",
          4421 => x"71",
          4422 => x"55",
          4423 => x"43",
          4424 => x"75",
          4425 => x"5d",
          4426 => x"84",
          4427 => x"08",
          4428 => x"75",
          4429 => x"0c",
          4430 => x"19",
          4431 => x"51",
          4432 => x"84",
          4433 => x"ef",
          4434 => x"34",
          4435 => x"84",
          4436 => x"1a",
          4437 => x"33",
          4438 => x"fe",
          4439 => x"a0",
          4440 => x"19",
          4441 => x"fe",
          4442 => x"06",
          4443 => x"06",
          4444 => x"18",
          4445 => x"1f",
          4446 => x"5e",
          4447 => x"55",
          4448 => x"75",
          4449 => x"38",
          4450 => x"1d",
          4451 => x"3d",
          4452 => x"8d",
          4453 => x"81",
          4454 => x"19",
          4455 => x"07",
          4456 => x"77",
          4457 => x"f3",
          4458 => x"83",
          4459 => x"11",
          4460 => x"52",
          4461 => x"38",
          4462 => x"79",
          4463 => x"62",
          4464 => x"8c",
          4465 => x"86",
          4466 => x"2e",
          4467 => x"dd",
          4468 => x"63",
          4469 => x"5e",
          4470 => x"ff",
          4471 => x"c0",
          4472 => x"57",
          4473 => x"05",
          4474 => x"7f",
          4475 => x"59",
          4476 => x"2e",
          4477 => x"0c",
          4478 => x"0d",
          4479 => x"5c",
          4480 => x"3f",
          4481 => x"84",
          4482 => x"40",
          4483 => x"1b",
          4484 => x"b4",
          4485 => x"83",
          4486 => x"2e",
          4487 => x"54",
          4488 => x"33",
          4489 => x"08",
          4490 => x"57",
          4491 => x"81",
          4492 => x"58",
          4493 => x"8b",
          4494 => x"06",
          4495 => x"81",
          4496 => x"2a",
          4497 => x"ef",
          4498 => x"2e",
          4499 => x"7d",
          4500 => x"75",
          4501 => x"05",
          4502 => x"ff",
          4503 => x"e4",
          4504 => x"ab",
          4505 => x"38",
          4506 => x"70",
          4507 => x"05",
          4508 => x"5a",
          4509 => x"dc",
          4510 => x"ff",
          4511 => x"52",
          4512 => x"84",
          4513 => x"2e",
          4514 => x"0c",
          4515 => x"1b",
          4516 => x"51",
          4517 => x"84",
          4518 => x"a4",
          4519 => x"34",
          4520 => x"84",
          4521 => x"1c",
          4522 => x"33",
          4523 => x"fd",
          4524 => x"a0",
          4525 => x"1b",
          4526 => x"fd",
          4527 => x"ab",
          4528 => x"42",
          4529 => x"2a",
          4530 => x"38",
          4531 => x"70",
          4532 => x"59",
          4533 => x"81",
          4534 => x"51",
          4535 => x"5a",
          4536 => x"d9",
          4537 => x"fe",
          4538 => x"ac",
          4539 => x"33",
          4540 => x"c7",
          4541 => x"9a",
          4542 => x"42",
          4543 => x"70",
          4544 => x"55",
          4545 => x"18",
          4546 => x"33",
          4547 => x"75",
          4548 => x"fe",
          4549 => x"a0",
          4550 => x"10",
          4551 => x"1b",
          4552 => x"84",
          4553 => x"fe",
          4554 => x"8c",
          4555 => x"70",
          4556 => x"80",
          4557 => x"38",
          4558 => x"41",
          4559 => x"81",
          4560 => x"84",
          4561 => x"0d",
          4562 => x"bc",
          4563 => x"ea",
          4564 => x"13",
          4565 => x"5e",
          4566 => x"8c",
          4567 => x"74",
          4568 => x"10",
          4569 => x"f4",
          4570 => x"8c",
          4571 => x"81",
          4572 => x"59",
          4573 => x"02",
          4574 => x"58",
          4575 => x"80",
          4576 => x"94",
          4577 => x"58",
          4578 => x"77",
          4579 => x"81",
          4580 => x"ef",
          4581 => x"7a",
          4582 => x"b8",
          4583 => x"58",
          4584 => x"81",
          4585 => x"90",
          4586 => x"60",
          4587 => x"a1",
          4588 => x"25",
          4589 => x"38",
          4590 => x"57",
          4591 => x"b9",
          4592 => x"74",
          4593 => x"84",
          4594 => x"77",
          4595 => x"7a",
          4596 => x"79",
          4597 => x"81",
          4598 => x"38",
          4599 => x"a0",
          4600 => x"16",
          4601 => x"38",
          4602 => x"19",
          4603 => x"34",
          4604 => x"51",
          4605 => x"8b",
          4606 => x"27",
          4607 => x"e4",
          4608 => x"08",
          4609 => x"09",
          4610 => x"db",
          4611 => x"02",
          4612 => x"58",
          4613 => x"5b",
          4614 => x"8c",
          4615 => x"bb",
          4616 => x"51",
          4617 => x"56",
          4618 => x"84",
          4619 => x"98",
          4620 => x"08",
          4621 => x"33",
          4622 => x"82",
          4623 => x"18",
          4624 => x"3f",
          4625 => x"38",
          4626 => x"0c",
          4627 => x"08",
          4628 => x"2e",
          4629 => x"25",
          4630 => x"81",
          4631 => x"2e",
          4632 => x"ee",
          4633 => x"84",
          4634 => x"38",
          4635 => x"38",
          4636 => x"1b",
          4637 => x"08",
          4638 => x"38",
          4639 => x"84",
          4640 => x"1c",
          4641 => x"3f",
          4642 => x"38",
          4643 => x"0c",
          4644 => x"0b",
          4645 => x"70",
          4646 => x"74",
          4647 => x"7b",
          4648 => x"57",
          4649 => x"ff",
          4650 => x"08",
          4651 => x"7c",
          4652 => x"34",
          4653 => x"98",
          4654 => x"80",
          4655 => x"fe",
          4656 => x"51",
          4657 => x"56",
          4658 => x"c7",
          4659 => x"18",
          4660 => x"51",
          4661 => x"77",
          4662 => x"84",
          4663 => x"18",
          4664 => x"a0",
          4665 => x"33",
          4666 => x"84",
          4667 => x"7f",
          4668 => x"53",
          4669 => x"bb",
          4670 => x"fe",
          4671 => x"56",
          4672 => x"81",
          4673 => x"5a",
          4674 => x"06",
          4675 => x"38",
          4676 => x"41",
          4677 => x"1c",
          4678 => x"33",
          4679 => x"82",
          4680 => x"1c",
          4681 => x"3f",
          4682 => x"38",
          4683 => x"0c",
          4684 => x"1c",
          4685 => x"06",
          4686 => x"8f",
          4687 => x"34",
          4688 => x"34",
          4689 => x"5a",
          4690 => x"8b",
          4691 => x"1b",
          4692 => x"33",
          4693 => x"05",
          4694 => x"75",
          4695 => x"57",
          4696 => x"38",
          4697 => x"38",
          4698 => x"76",
          4699 => x"34",
          4700 => x"7d",
          4701 => x"08",
          4702 => x"38",
          4703 => x"38",
          4704 => x"08",
          4705 => x"33",
          4706 => x"84",
          4707 => x"bb",
          4708 => x"08",
          4709 => x"08",
          4710 => x"fb",
          4711 => x"82",
          4712 => x"81",
          4713 => x"05",
          4714 => x"cf",
          4715 => x"76",
          4716 => x"56",
          4717 => x"fa",
          4718 => x"57",
          4719 => x"fa",
          4720 => x"fe",
          4721 => x"53",
          4722 => x"92",
          4723 => x"09",
          4724 => x"08",
          4725 => x"1d",
          4726 => x"27",
          4727 => x"82",
          4728 => x"56",
          4729 => x"58",
          4730 => x"87",
          4731 => x"81",
          4732 => x"fe",
          4733 => x"1c",
          4734 => x"52",
          4735 => x"fc",
          4736 => x"a0",
          4737 => x"18",
          4738 => x"39",
          4739 => x"40",
          4740 => x"98",
          4741 => x"ac",
          4742 => x"80",
          4743 => x"22",
          4744 => x"2e",
          4745 => x"22",
          4746 => x"95",
          4747 => x"ff",
          4748 => x"26",
          4749 => x"11",
          4750 => x"d4",
          4751 => x"30",
          4752 => x"94",
          4753 => x"80",
          4754 => x"1c",
          4755 => x"56",
          4756 => x"85",
          4757 => x"70",
          4758 => x"5b",
          4759 => x"80",
          4760 => x"05",
          4761 => x"70",
          4762 => x"8a",
          4763 => x"88",
          4764 => x"96",
          4765 => x"81",
          4766 => x"81",
          4767 => x"0b",
          4768 => x"11",
          4769 => x"89",
          4770 => x"13",
          4771 => x"9c",
          4772 => x"71",
          4773 => x"14",
          4774 => x"33",
          4775 => x"33",
          4776 => x"5f",
          4777 => x"77",
          4778 => x"16",
          4779 => x"7b",
          4780 => x"81",
          4781 => x"96",
          4782 => x"57",
          4783 => x"07",
          4784 => x"84",
          4785 => x"ff",
          4786 => x"81",
          4787 => x"7a",
          4788 => x"05",
          4789 => x"5b",
          4790 => x"57",
          4791 => x"39",
          4792 => x"80",
          4793 => x"57",
          4794 => x"81",
          4795 => x"08",
          4796 => x"1f",
          4797 => x"fe",
          4798 => x"59",
          4799 => x"5a",
          4800 => x"1c",
          4801 => x"76",
          4802 => x"72",
          4803 => x"38",
          4804 => x"55",
          4805 => x"34",
          4806 => x"89",
          4807 => x"79",
          4808 => x"83",
          4809 => x"70",
          4810 => x"5d",
          4811 => x"0d",
          4812 => x"80",
          4813 => x"af",
          4814 => x"dc",
          4815 => x"81",
          4816 => x"0c",
          4817 => x"42",
          4818 => x"73",
          4819 => x"61",
          4820 => x"53",
          4821 => x"73",
          4822 => x"ff",
          4823 => x"56",
          4824 => x"83",
          4825 => x"30",
          4826 => x"57",
          4827 => x"74",
          4828 => x"80",
          4829 => x"0b",
          4830 => x"06",
          4831 => x"ab",
          4832 => x"16",
          4833 => x"54",
          4834 => x"06",
          4835 => x"fe",
          4836 => x"5d",
          4837 => x"70",
          4838 => x"73",
          4839 => x"39",
          4840 => x"70",
          4841 => x"55",
          4842 => x"70",
          4843 => x"72",
          4844 => x"32",
          4845 => x"51",
          4846 => x"1d",
          4847 => x"41",
          4848 => x"38",
          4849 => x"81",
          4850 => x"83",
          4851 => x"38",
          4852 => x"93",
          4853 => x"70",
          4854 => x"2e",
          4855 => x"0b",
          4856 => x"de",
          4857 => x"bb",
          4858 => x"73",
          4859 => x"25",
          4860 => x"80",
          4861 => x"62",
          4862 => x"2e",
          4863 => x"30",
          4864 => x"59",
          4865 => x"75",
          4866 => x"84",
          4867 => x"38",
          4868 => x"38",
          4869 => x"22",
          4870 => x"2a",
          4871 => x"ae",
          4872 => x"17",
          4873 => x"19",
          4874 => x"fe",
          4875 => x"ff",
          4876 => x"7a",
          4877 => x"ff",
          4878 => x"f1",
          4879 => x"19",
          4880 => x"ae",
          4881 => x"05",
          4882 => x"8f",
          4883 => x"7c",
          4884 => x"8b",
          4885 => x"70",
          4886 => x"72",
          4887 => x"78",
          4888 => x"54",
          4889 => x"74",
          4890 => x"32",
          4891 => x"54",
          4892 => x"83",
          4893 => x"83",
          4894 => x"30",
          4895 => x"07",
          4896 => x"83",
          4897 => x"38",
          4898 => x"07",
          4899 => x"56",
          4900 => x"fc",
          4901 => x"15",
          4902 => x"74",
          4903 => x"76",
          4904 => x"88",
          4905 => x"58",
          4906 => x"83",
          4907 => x"38",
          4908 => x"9d",
          4909 => x"2e",
          4910 => x"82",
          4911 => x"85",
          4912 => x"1d",
          4913 => x"bb",
          4914 => x"84",
          4915 => x"38",
          4916 => x"81",
          4917 => x"81",
          4918 => x"38",
          4919 => x"82",
          4920 => x"73",
          4921 => x"f9",
          4922 => x"11",
          4923 => x"a0",
          4924 => x"85",
          4925 => x"39",
          4926 => x"09",
          4927 => x"54",
          4928 => x"a0",
          4929 => x"23",
          4930 => x"54",
          4931 => x"73",
          4932 => x"13",
          4933 => x"a0",
          4934 => x"51",
          4935 => x"ab",
          4936 => x"08",
          4937 => x"06",
          4938 => x"33",
          4939 => x"74",
          4940 => x"08",
          4941 => x"11",
          4942 => x"2b",
          4943 => x"7d",
          4944 => x"1d",
          4945 => x"b7",
          4946 => x"fe",
          4947 => x"88",
          4948 => x"76",
          4949 => x"82",
          4950 => x"59",
          4951 => x"fd",
          4952 => x"98",
          4953 => x"88",
          4954 => x"d6",
          4955 => x"80",
          4956 => x"0d",
          4957 => x"81",
          4958 => x"1d",
          4959 => x"79",
          4960 => x"5a",
          4961 => x"83",
          4962 => x"3f",
          4963 => x"06",
          4964 => x"78",
          4965 => x"06",
          4966 => x"74",
          4967 => x"80",
          4968 => x"0b",
          4969 => x"06",
          4970 => x"e0",
          4971 => x"19",
          4972 => x"54",
          4973 => x"06",
          4974 => x"15",
          4975 => x"82",
          4976 => x"ff",
          4977 => x"38",
          4978 => x"e0",
          4979 => x"56",
          4980 => x"74",
          4981 => x"55",
          4982 => x"39",
          4983 => x"06",
          4984 => x"38",
          4985 => x"a0",
          4986 => x"81",
          4987 => x"33",
          4988 => x"71",
          4989 => x"0c",
          4990 => x"a0",
          4991 => x"74",
          4992 => x"5a",
          4993 => x"ff",
          4994 => x"33",
          4995 => x"81",
          4996 => x"74",
          4997 => x"f2",
          4998 => x"93",
          4999 => x"69",
          5000 => x"42",
          5001 => x"08",
          5002 => x"85",
          5003 => x"33",
          5004 => x"2e",
          5005 => x"ba",
          5006 => x"33",
          5007 => x"75",
          5008 => x"08",
          5009 => x"85",
          5010 => x"fe",
          5011 => x"2e",
          5012 => x"bb",
          5013 => x"ff",
          5014 => x"80",
          5015 => x"75",
          5016 => x"81",
          5017 => x"51",
          5018 => x"08",
          5019 => x"56",
          5020 => x"80",
          5021 => x"06",
          5022 => x"80",
          5023 => x"b4",
          5024 => x"54",
          5025 => x"18",
          5026 => x"84",
          5027 => x"ff",
          5028 => x"84",
          5029 => x"33",
          5030 => x"07",
          5031 => x"d5",
          5032 => x"8b",
          5033 => x"61",
          5034 => x"2e",
          5035 => x"26",
          5036 => x"80",
          5037 => x"5e",
          5038 => x"06",
          5039 => x"80",
          5040 => x"57",
          5041 => x"83",
          5042 => x"2b",
          5043 => x"70",
          5044 => x"07",
          5045 => x"75",
          5046 => x"82",
          5047 => x"11",
          5048 => x"8d",
          5049 => x"78",
          5050 => x"c5",
          5051 => x"18",
          5052 => x"c4",
          5053 => x"87",
          5054 => x"c9",
          5055 => x"40",
          5056 => x"06",
          5057 => x"38",
          5058 => x"33",
          5059 => x"a4",
          5060 => x"82",
          5061 => x"2b",
          5062 => x"88",
          5063 => x"5a",
          5064 => x"33",
          5065 => x"07",
          5066 => x"81",
          5067 => x"05",
          5068 => x"78",
          5069 => x"b5",
          5070 => x"bb",
          5071 => x"84",
          5072 => x"f5",
          5073 => x"ff",
          5074 => x"9f",
          5075 => x"82",
          5076 => x"19",
          5077 => x"7b",
          5078 => x"83",
          5079 => x"5c",
          5080 => x"38",
          5081 => x"55",
          5082 => x"19",
          5083 => x"56",
          5084 => x"8d",
          5085 => x"38",
          5086 => x"90",
          5087 => x"34",
          5088 => x"77",
          5089 => x"5d",
          5090 => x"18",
          5091 => x"0c",
          5092 => x"77",
          5093 => x"04",
          5094 => x"3d",
          5095 => x"81",
          5096 => x"26",
          5097 => x"06",
          5098 => x"87",
          5099 => x"f4",
          5100 => x"5b",
          5101 => x"70",
          5102 => x"5a",
          5103 => x"e0",
          5104 => x"ff",
          5105 => x"38",
          5106 => x"55",
          5107 => x"75",
          5108 => x"77",
          5109 => x"30",
          5110 => x"5d",
          5111 => x"38",
          5112 => x"7c",
          5113 => x"a9",
          5114 => x"77",
          5115 => x"7d",
          5116 => x"39",
          5117 => x"e9",
          5118 => x"59",
          5119 => x"80",
          5120 => x"83",
          5121 => x"a6",
          5122 => x"59",
          5123 => x"7a",
          5124 => x"33",
          5125 => x"71",
          5126 => x"70",
          5127 => x"33",
          5128 => x"40",
          5129 => x"ff",
          5130 => x"25",
          5131 => x"33",
          5132 => x"31",
          5133 => x"05",
          5134 => x"5b",
          5135 => x"80",
          5136 => x"18",
          5137 => x"55",
          5138 => x"81",
          5139 => x"17",
          5140 => x"bb",
          5141 => x"55",
          5142 => x"58",
          5143 => x"33",
          5144 => x"58",
          5145 => x"06",
          5146 => x"57",
          5147 => x"38",
          5148 => x"80",
          5149 => x"bc",
          5150 => x"82",
          5151 => x"0b",
          5152 => x"7b",
          5153 => x"81",
          5154 => x"77",
          5155 => x"84",
          5156 => x"d1",
          5157 => x"ee",
          5158 => x"7b",
          5159 => x"81",
          5160 => x"1b",
          5161 => x"80",
          5162 => x"85",
          5163 => x"40",
          5164 => x"33",
          5165 => x"71",
          5166 => x"77",
          5167 => x"2e",
          5168 => x"8d",
          5169 => x"bb",
          5170 => x"58",
          5171 => x"0b",
          5172 => x"5d",
          5173 => x"bb",
          5174 => x"0b",
          5175 => x"5a",
          5176 => x"7a",
          5177 => x"31",
          5178 => x"80",
          5179 => x"e1",
          5180 => x"e6",
          5181 => x"05",
          5182 => x"33",
          5183 => x"42",
          5184 => x"75",
          5185 => x"57",
          5186 => x"58",
          5187 => x"80",
          5188 => x"57",
          5189 => x"f9",
          5190 => x"b4",
          5191 => x"17",
          5192 => x"06",
          5193 => x"b8",
          5194 => x"b0",
          5195 => x"2e",
          5196 => x"b4",
          5197 => x"84",
          5198 => x"b6",
          5199 => x"5e",
          5200 => x"06",
          5201 => x"33",
          5202 => x"88",
          5203 => x"07",
          5204 => x"41",
          5205 => x"8b",
          5206 => x"f8",
          5207 => x"33",
          5208 => x"88",
          5209 => x"07",
          5210 => x"44",
          5211 => x"8a",
          5212 => x"f8",
          5213 => x"33",
          5214 => x"88",
          5215 => x"07",
          5216 => x"1e",
          5217 => x"33",
          5218 => x"88",
          5219 => x"07",
          5220 => x"90",
          5221 => x"45",
          5222 => x"34",
          5223 => x"7c",
          5224 => x"23",
          5225 => x"80",
          5226 => x"7b",
          5227 => x"7f",
          5228 => x"b4",
          5229 => x"81",
          5230 => x"3f",
          5231 => x"81",
          5232 => x"08",
          5233 => x"18",
          5234 => x"27",
          5235 => x"82",
          5236 => x"08",
          5237 => x"80",
          5238 => x"8a",
          5239 => x"fc",
          5240 => x"e2",
          5241 => x"5a",
          5242 => x"17",
          5243 => x"e4",
          5244 => x"71",
          5245 => x"14",
          5246 => x"33",
          5247 => x"82",
          5248 => x"f5",
          5249 => x"f9",
          5250 => x"75",
          5251 => x"77",
          5252 => x"75",
          5253 => x"39",
          5254 => x"08",
          5255 => x"51",
          5256 => x"f0",
          5257 => x"64",
          5258 => x"ff",
          5259 => x"e9",
          5260 => x"70",
          5261 => x"80",
          5262 => x"2e",
          5263 => x"54",
          5264 => x"10",
          5265 => x"55",
          5266 => x"74",
          5267 => x"38",
          5268 => x"0c",
          5269 => x"80",
          5270 => x"51",
          5271 => x"54",
          5272 => x"0d",
          5273 => x"92",
          5274 => x"70",
          5275 => x"89",
          5276 => x"ff",
          5277 => x"2e",
          5278 => x"e6",
          5279 => x"59",
          5280 => x"78",
          5281 => x"12",
          5282 => x"38",
          5283 => x"54",
          5284 => x"89",
          5285 => x"57",
          5286 => x"54",
          5287 => x"38",
          5288 => x"70",
          5289 => x"07",
          5290 => x"38",
          5291 => x"7b",
          5292 => x"98",
          5293 => x"79",
          5294 => x"3d",
          5295 => x"05",
          5296 => x"2e",
          5297 => x"9d",
          5298 => x"05",
          5299 => x"84",
          5300 => x"2e",
          5301 => x"75",
          5302 => x"04",
          5303 => x"52",
          5304 => x"08",
          5305 => x"81",
          5306 => x"80",
          5307 => x"83",
          5308 => x"38",
          5309 => x"38",
          5310 => x"80",
          5311 => x"33",
          5312 => x"61",
          5313 => x"7d",
          5314 => x"8e",
          5315 => x"a1",
          5316 => x"91",
          5317 => x"17",
          5318 => x"9a",
          5319 => x"7d",
          5320 => x"38",
          5321 => x"80",
          5322 => x"19",
          5323 => x"55",
          5324 => x"2e",
          5325 => x"7c",
          5326 => x"7b",
          5327 => x"26",
          5328 => x"0c",
          5329 => x"33",
          5330 => x"25",
          5331 => x"5e",
          5332 => x"82",
          5333 => x"84",
          5334 => x"b0",
          5335 => x"7c",
          5336 => x"58",
          5337 => x"81",
          5338 => x"78",
          5339 => x"08",
          5340 => x"67",
          5341 => x"88",
          5342 => x"57",
          5343 => x"77",
          5344 => x"33",
          5345 => x"88",
          5346 => x"07",
          5347 => x"8c",
          5348 => x"58",
          5349 => x"1b",
          5350 => x"91",
          5351 => x"80",
          5352 => x"84",
          5353 => x"81",
          5354 => x"f4",
          5355 => x"78",
          5356 => x"08",
          5357 => x"74",
          5358 => x"89",
          5359 => x"5a",
          5360 => x"25",
          5361 => x"38",
          5362 => x"80",
          5363 => x"51",
          5364 => x"08",
          5365 => x"83",
          5366 => x"ff",
          5367 => x"c1",
          5368 => x"06",
          5369 => x"81",
          5370 => x"38",
          5371 => x"39",
          5372 => x"39",
          5373 => x"39",
          5374 => x"89",
          5375 => x"71",
          5376 => x"07",
          5377 => x"33",
          5378 => x"88",
          5379 => x"07",
          5380 => x"8c",
          5381 => x"5a",
          5382 => x"22",
          5383 => x"80",
          5384 => x"1b",
          5385 => x"1a",
          5386 => x"f4",
          5387 => x"bb",
          5388 => x"76",
          5389 => x"52",
          5390 => x"bb",
          5391 => x"80",
          5392 => x"08",
          5393 => x"84",
          5394 => x"53",
          5395 => x"3f",
          5396 => x"9c",
          5397 => x"59",
          5398 => x"81",
          5399 => x"81",
          5400 => x"55",
          5401 => x"7f",
          5402 => x"16",
          5403 => x"33",
          5404 => x"81",
          5405 => x"16",
          5406 => x"b3",
          5407 => x"85",
          5408 => x"17",
          5409 => x"18",
          5410 => x"38",
          5411 => x"0b",
          5412 => x"34",
          5413 => x"17",
          5414 => x"07",
          5415 => x"8e",
          5416 => x"a1",
          5417 => x"91",
          5418 => x"17",
          5419 => x"9a",
          5420 => x"7d",
          5421 => x"06",
          5422 => x"98",
          5423 => x"83",
          5424 => x"a5",
          5425 => x"fe",
          5426 => x"f9",
          5427 => x"29",
          5428 => x"80",
          5429 => x"15",
          5430 => x"77",
          5431 => x"ff",
          5432 => x"80",
          5433 => x"7a",
          5434 => x"16",
          5435 => x"17",
          5436 => x"84",
          5437 => x"06",
          5438 => x"83",
          5439 => x"08",
          5440 => x"74",
          5441 => x"82",
          5442 => x"81",
          5443 => x"16",
          5444 => x"52",
          5445 => x"3f",
          5446 => x"84",
          5447 => x"39",
          5448 => x"0d",
          5449 => x"59",
          5450 => x"2e",
          5451 => x"2e",
          5452 => x"2e",
          5453 => x"22",
          5454 => x"38",
          5455 => x"81",
          5456 => x"81",
          5457 => x"57",
          5458 => x"38",
          5459 => x"31",
          5460 => x"38",
          5461 => x"83",
          5462 => x"7e",
          5463 => x"2a",
          5464 => x"82",
          5465 => x"75",
          5466 => x"83",
          5467 => x"58",
          5468 => x"08",
          5469 => x"83",
          5470 => x"29",
          5471 => x"80",
          5472 => x"89",
          5473 => x"e6",
          5474 => x"85",
          5475 => x"76",
          5476 => x"ff",
          5477 => x"82",
          5478 => x"2b",
          5479 => x"38",
          5480 => x"7e",
          5481 => x"1b",
          5482 => x"5e",
          5483 => x"75",
          5484 => x"04",
          5485 => x"0d",
          5486 => x"19",
          5487 => x"38",
          5488 => x"1b",
          5489 => x"38",
          5490 => x"18",
          5491 => x"bb",
          5492 => x"33",
          5493 => x"34",
          5494 => x"52",
          5495 => x"3f",
          5496 => x"76",
          5497 => x"75",
          5498 => x"58",
          5499 => x"57",
          5500 => x"59",
          5501 => x"74",
          5502 => x"81",
          5503 => x"80",
          5504 => x"05",
          5505 => x"34",
          5506 => x"ac",
          5507 => x"ff",
          5508 => x"55",
          5509 => x"ff",
          5510 => x"81",
          5511 => x"79",
          5512 => x"19",
          5513 => x"fd",
          5514 => x"1e",
          5515 => x"81",
          5516 => x"59",
          5517 => x"fd",
          5518 => x"33",
          5519 => x"15",
          5520 => x"81",
          5521 => x"bb",
          5522 => x"0b",
          5523 => x"84",
          5524 => x"0d",
          5525 => x"59",
          5526 => x"2e",
          5527 => x"2e",
          5528 => x"2e",
          5529 => x"22",
          5530 => x"38",
          5531 => x"82",
          5532 => x"82",
          5533 => x"2a",
          5534 => x"80",
          5535 => x"7b",
          5536 => x"38",
          5537 => x"89",
          5538 => x"82",
          5539 => x"05",
          5540 => x"aa",
          5541 => x"08",
          5542 => x"74",
          5543 => x"2e",
          5544 => x"88",
          5545 => x"0c",
          5546 => x"2b",
          5547 => x"38",
          5548 => x"08",
          5549 => x"83",
          5550 => x"29",
          5551 => x"80",
          5552 => x"89",
          5553 => x"a6",
          5554 => x"85",
          5555 => x"7b",
          5556 => x"ff",
          5557 => x"82",
          5558 => x"56",
          5559 => x"0b",
          5560 => x"58",
          5561 => x"33",
          5562 => x"15",
          5563 => x"80",
          5564 => x"79",
          5565 => x"08",
          5566 => x"08",
          5567 => x"1d",
          5568 => x"76",
          5569 => x"1a",
          5570 => x"33",
          5571 => x"90",
          5572 => x"84",
          5573 => x"bb",
          5574 => x"19",
          5575 => x"08",
          5576 => x"38",
          5577 => x"81",
          5578 => x"84",
          5579 => x"19",
          5580 => x"83",
          5581 => x"55",
          5582 => x"77",
          5583 => x"56",
          5584 => x"81",
          5585 => x"57",
          5586 => x"90",
          5587 => x"90",
          5588 => x"08",
          5589 => x"84",
          5590 => x"08",
          5591 => x"fe",
          5592 => x"ac",
          5593 => x"84",
          5594 => x"39",
          5595 => x"19",
          5596 => x"c2",
          5597 => x"90",
          5598 => x"90",
          5599 => x"81",
          5600 => x"84",
          5601 => x"fb",
          5602 => x"fb",
          5603 => x"81",
          5604 => x"0d",
          5605 => x"0b",
          5606 => x"04",
          5607 => x"77",
          5608 => x"75",
          5609 => x"74",
          5610 => x"84",
          5611 => x"83",
          5612 => x"56",
          5613 => x"70",
          5614 => x"80",
          5615 => x"56",
          5616 => x"a0",
          5617 => x"77",
          5618 => x"33",
          5619 => x"09",
          5620 => x"76",
          5621 => x"51",
          5622 => x"08",
          5623 => x"59",
          5624 => x"81",
          5625 => x"33",
          5626 => x"34",
          5627 => x"ff",
          5628 => x"18",
          5629 => x"18",
          5630 => x"5c",
          5631 => x"38",
          5632 => x"74",
          5633 => x"74",
          5634 => x"74",
          5635 => x"80",
          5636 => x"a1",
          5637 => x"99",
          5638 => x"80",
          5639 => x"0b",
          5640 => x"95",
          5641 => x"33",
          5642 => x"19",
          5643 => x"0c",
          5644 => x"16",
          5645 => x"17",
          5646 => x"81",
          5647 => x"09",
          5648 => x"84",
          5649 => x"a8",
          5650 => x"5a",
          5651 => x"85",
          5652 => x"2e",
          5653 => x"54",
          5654 => x"53",
          5655 => x"94",
          5656 => x"78",
          5657 => x"74",
          5658 => x"8c",
          5659 => x"88",
          5660 => x"90",
          5661 => x"98",
          5662 => x"7a",
          5663 => x"0b",
          5664 => x"18",
          5665 => x"0b",
          5666 => x"83",
          5667 => x"3f",
          5668 => x"81",
          5669 => x"34",
          5670 => x"ff",
          5671 => x"81",
          5672 => x"78",
          5673 => x"54",
          5674 => x"7b",
          5675 => x"ca",
          5676 => x"fd",
          5677 => x"06",
          5678 => x"19",
          5679 => x"2e",
          5680 => x"c2",
          5681 => x"55",
          5682 => x"54",
          5683 => x"56",
          5684 => x"53",
          5685 => x"52",
          5686 => x"22",
          5687 => x"2e",
          5688 => x"54",
          5689 => x"84",
          5690 => x"81",
          5691 => x"84",
          5692 => x"da",
          5693 => x"39",
          5694 => x"57",
          5695 => x"70",
          5696 => x"52",
          5697 => x"ee",
          5698 => x"e2",
          5699 => x"38",
          5700 => x"84",
          5701 => x"8b",
          5702 => x"0d",
          5703 => x"ff",
          5704 => x"91",
          5705 => x"d0",
          5706 => x"f5",
          5707 => x"58",
          5708 => x"81",
          5709 => x"57",
          5710 => x"70",
          5711 => x"81",
          5712 => x"51",
          5713 => x"70",
          5714 => x"70",
          5715 => x"09",
          5716 => x"38",
          5717 => x"07",
          5718 => x"76",
          5719 => x"1b",
          5720 => x"38",
          5721 => x"24",
          5722 => x"c3",
          5723 => x"3d",
          5724 => x"d3",
          5725 => x"bb",
          5726 => x"84",
          5727 => x"7a",
          5728 => x"51",
          5729 => x"55",
          5730 => x"02",
          5731 => x"58",
          5732 => x"02",
          5733 => x"06",
          5734 => x"7a",
          5735 => x"71",
          5736 => x"5b",
          5737 => x"76",
          5738 => x"0c",
          5739 => x"08",
          5740 => x"38",
          5741 => x"3d",
          5742 => x"33",
          5743 => x"79",
          5744 => x"39",
          5745 => x"84",
          5746 => x"ff",
          5747 => x"80",
          5748 => x"34",
          5749 => x"05",
          5750 => x"3f",
          5751 => x"84",
          5752 => x"3d",
          5753 => x"dd",
          5754 => x"5b",
          5755 => x"80",
          5756 => x"52",
          5757 => x"bb",
          5758 => x"83",
          5759 => x"58",
          5760 => x"38",
          5761 => x"5f",
          5762 => x"76",
          5763 => x"51",
          5764 => x"08",
          5765 => x"59",
          5766 => x"38",
          5767 => x"9a",
          5768 => x"70",
          5769 => x"83",
          5770 => x"3d",
          5771 => x"f6",
          5772 => x"bb",
          5773 => x"7a",
          5774 => x"84",
          5775 => x"38",
          5776 => x"9a",
          5777 => x"70",
          5778 => x"83",
          5779 => x"a4",
          5780 => x"51",
          5781 => x"08",
          5782 => x"ff",
          5783 => x"38",
          5784 => x"fd",
          5785 => x"c8",
          5786 => x"57",
          5787 => x"56",
          5788 => x"57",
          5789 => x"75",
          5790 => x"2e",
          5791 => x"ff",
          5792 => x"19",
          5793 => x"33",
          5794 => x"80",
          5795 => x"7e",
          5796 => x"fd",
          5797 => x"38",
          5798 => x"10",
          5799 => x"70",
          5800 => x"7a",
          5801 => x"70",
          5802 => x"82",
          5803 => x"80",
          5804 => x"16",
          5805 => x"5e",
          5806 => x"ee",
          5807 => x"34",
          5808 => x"df",
          5809 => x"84",
          5810 => x"04",
          5811 => x"98",
          5812 => x"59",
          5813 => x"33",
          5814 => x"90",
          5815 => x"0c",
          5816 => x"a2",
          5817 => x"84",
          5818 => x"38",
          5819 => x"08",
          5820 => x"33",
          5821 => x"59",
          5822 => x"84",
          5823 => x"16",
          5824 => x"84",
          5825 => x"27",
          5826 => x"74",
          5827 => x"38",
          5828 => x"08",
          5829 => x"51",
          5830 => x"dd",
          5831 => x"11",
          5832 => x"84",
          5833 => x"e6",
          5834 => x"59",
          5835 => x"81",
          5836 => x"80",
          5837 => x"5a",
          5838 => x"34",
          5839 => x"e5",
          5840 => x"79",
          5841 => x"7f",
          5842 => x"82",
          5843 => x"84",
          5844 => x"3d",
          5845 => x"76",
          5846 => x"75",
          5847 => x"74",
          5848 => x"84",
          5849 => x"83",
          5850 => x"55",
          5851 => x"55",
          5852 => x"58",
          5853 => x"17",
          5854 => x"83",
          5855 => x"89",
          5856 => x"82",
          5857 => x"fd",
          5858 => x"ff",
          5859 => x"fd",
          5860 => x"75",
          5861 => x"06",
          5862 => x"98",
          5863 => x"2e",
          5864 => x"d3",
          5865 => x"19",
          5866 => x"81",
          5867 => x"80",
          5868 => x"51",
          5869 => x"08",
          5870 => x"9e",
          5871 => x"81",
          5872 => x"75",
          5873 => x"75",
          5874 => x"bb",
          5875 => x"94",
          5876 => x"77",
          5877 => x"9c",
          5878 => x"75",
          5879 => x"22",
          5880 => x"7a",
          5881 => x"80",
          5882 => x"58",
          5883 => x"90",
          5884 => x"33",
          5885 => x"34",
          5886 => x"2e",
          5887 => x"75",
          5888 => x"33",
          5889 => x"59",
          5890 => x"75",
          5891 => x"52",
          5892 => x"84",
          5893 => x"ff",
          5894 => x"54",
          5895 => x"33",
          5896 => x"bb",
          5897 => x"81",
          5898 => x"84",
          5899 => x"90",
          5900 => x"57",
          5901 => x"18",
          5902 => x"2e",
          5903 => x"94",
          5904 => x"94",
          5905 => x"80",
          5906 => x"0c",
          5907 => x"a3",
          5908 => x"84",
          5909 => x"75",
          5910 => x"84",
          5911 => x"81",
          5912 => x"84",
          5913 => x"fc",
          5914 => x"fb",
          5915 => x"98",
          5916 => x"84",
          5917 => x"84",
          5918 => x"38",
          5919 => x"75",
          5920 => x"0b",
          5921 => x"84",
          5922 => x"0d",
          5923 => x"a2",
          5924 => x"52",
          5925 => x"3f",
          5926 => x"84",
          5927 => x"0c",
          5928 => x"8c",
          5929 => x"52",
          5930 => x"bb",
          5931 => x"80",
          5932 => x"2b",
          5933 => x"86",
          5934 => x"5b",
          5935 => x"9c",
          5936 => x"33",
          5937 => x"5d",
          5938 => x"b3",
          5939 => x"86",
          5940 => x"75",
          5941 => x"84",
          5942 => x"74",
          5943 => x"0c",
          5944 => x"0c",
          5945 => x"18",
          5946 => x"07",
          5947 => x"ff",
          5948 => x"89",
          5949 => x"08",
          5950 => x"33",
          5951 => x"13",
          5952 => x"76",
          5953 => x"73",
          5954 => x"bb",
          5955 => x"13",
          5956 => x"bb",
          5957 => x"38",
          5958 => x"f8",
          5959 => x"56",
          5960 => x"54",
          5961 => x"53",
          5962 => x"22",
          5963 => x"2e",
          5964 => x"75",
          5965 => x"2e",
          5966 => x"ff",
          5967 => x"53",
          5968 => x"38",
          5969 => x"52",
          5970 => x"52",
          5971 => x"bb",
          5972 => x"72",
          5973 => x"06",
          5974 => x"0c",
          5975 => x"75",
          5976 => x"52",
          5977 => x"bb",
          5978 => x"72",
          5979 => x"06",
          5980 => x"74",
          5981 => x"84",
          5982 => x"0d",
          5983 => x"d9",
          5984 => x"53",
          5985 => x"54",
          5986 => x"66",
          5987 => x"97",
          5988 => x"bb",
          5989 => x"80",
          5990 => x"0c",
          5991 => x"51",
          5992 => x"08",
          5993 => x"02",
          5994 => x"55",
          5995 => x"80",
          5996 => x"ff",
          5997 => x"0c",
          5998 => x"bb",
          5999 => x"3d",
          6000 => x"95",
          6001 => x"c1",
          6002 => x"84",
          6003 => x"0c",
          6004 => x"94",
          6005 => x"75",
          6006 => x"84",
          6007 => x"84",
          6008 => x"78",
          6009 => x"18",
          6010 => x"59",
          6011 => x"71",
          6012 => x"2e",
          6013 => x"5f",
          6014 => x"75",
          6015 => x"51",
          6016 => x"08",
          6017 => x"5e",
          6018 => x"57",
          6019 => x"7d",
          6020 => x"b8",
          6021 => x"71",
          6022 => x"14",
          6023 => x"33",
          6024 => x"07",
          6025 => x"60",
          6026 => x"05",
          6027 => x"58",
          6028 => x"7a",
          6029 => x"17",
          6030 => x"34",
          6031 => x"0d",
          6032 => x"b8",
          6033 => x"5d",
          6034 => x"bb",
          6035 => x"84",
          6036 => x"a8",
          6037 => x"5f",
          6038 => x"bd",
          6039 => x"2e",
          6040 => x"54",
          6041 => x"53",
          6042 => x"fc",
          6043 => x"82",
          6044 => x"52",
          6045 => x"bb",
          6046 => x"84",
          6047 => x"38",
          6048 => x"bb",
          6049 => x"81",
          6050 => x"17",
          6051 => x"0c",
          6052 => x"81",
          6053 => x"c8",
          6054 => x"33",
          6055 => x"30",
          6056 => x"ff",
          6057 => x"5f",
          6058 => x"8f",
          6059 => x"60",
          6060 => x"18",
          6061 => x"77",
          6062 => x"60",
          6063 => x"7c",
          6064 => x"38",
          6065 => x"38",
          6066 => x"38",
          6067 => x"5a",
          6068 => x"55",
          6069 => x"18",
          6070 => x"18",
          6071 => x"59",
          6072 => x"38",
          6073 => x"08",
          6074 => x"38",
          6075 => x"81",
          6076 => x"75",
          6077 => x"0b",
          6078 => x"19",
          6079 => x"90",
          6080 => x"2b",
          6081 => x"54",
          6082 => x"7a",
          6083 => x"8a",
          6084 => x"83",
          6085 => x"34",
          6086 => x"8c",
          6087 => x"27",
          6088 => x"fe",
          6089 => x"5a",
          6090 => x"e9",
          6091 => x"82",
          6092 => x"2e",
          6093 => x"76",
          6094 => x"84",
          6095 => x"fe",
          6096 => x"75",
          6097 => x"94",
          6098 => x"55",
          6099 => x"7a",
          6100 => x"16",
          6101 => x"bb",
          6102 => x"ee",
          6103 => x"e8",
          6104 => x"55",
          6105 => x"fe",
          6106 => x"51",
          6107 => x"08",
          6108 => x"84",
          6109 => x"81",
          6110 => x"08",
          6111 => x"84",
          6112 => x"08",
          6113 => x"84",
          6114 => x"84",
          6115 => x"38",
          6116 => x"75",
          6117 => x"84",
          6118 => x"08",
          6119 => x"fe",
          6120 => x"5a",
          6121 => x"cb",
          6122 => x"80",
          6123 => x"2e",
          6124 => x"76",
          6125 => x"84",
          6126 => x"fe",
          6127 => x"75",
          6128 => x"18",
          6129 => x"74",
          6130 => x"26",
          6131 => x"90",
          6132 => x"57",
          6133 => x"33",
          6134 => x"e7",
          6135 => x"55",
          6136 => x"ea",
          6137 => x"55",
          6138 => x"90",
          6139 => x"81",
          6140 => x"e0",
          6141 => x"af",
          6142 => x"3d",
          6143 => x"05",
          6144 => x"3f",
          6145 => x"84",
          6146 => x"bb",
          6147 => x"4b",
          6148 => x"52",
          6149 => x"84",
          6150 => x"38",
          6151 => x"2a",
          6152 => x"cd",
          6153 => x"24",
          6154 => x"70",
          6155 => x"ff",
          6156 => x"11",
          6157 => x"07",
          6158 => x"7c",
          6159 => x"2a",
          6160 => x"ed",
          6161 => x"2e",
          6162 => x"84",
          6163 => x"52",
          6164 => x"84",
          6165 => x"e5",
          6166 => x"51",
          6167 => x"08",
          6168 => x"87",
          6169 => x"0d",
          6170 => x"71",
          6171 => x"07",
          6172 => x"bb",
          6173 => x"bb",
          6174 => x"6f",
          6175 => x"ff",
          6176 => x"51",
          6177 => x"08",
          6178 => x"be",
          6179 => x"25",
          6180 => x"74",
          6181 => x"58",
          6182 => x"17",
          6183 => x"56",
          6184 => x"f6",
          6185 => x"bb",
          6186 => x"17",
          6187 => x"b4",
          6188 => x"83",
          6189 => x"2e",
          6190 => x"54",
          6191 => x"33",
          6192 => x"84",
          6193 => x"81",
          6194 => x"77",
          6195 => x"78",
          6196 => x"19",
          6197 => x"52",
          6198 => x"bb",
          6199 => x"80",
          6200 => x"09",
          6201 => x"fe",
          6202 => x"53",
          6203 => x"f2",
          6204 => x"08",
          6205 => x"38",
          6206 => x"b4",
          6207 => x"bb",
          6208 => x"08",
          6209 => x"55",
          6210 => x"de",
          6211 => x"18",
          6212 => x"33",
          6213 => x"fe",
          6214 => x"80",
          6215 => x"f7",
          6216 => x"84",
          6217 => x"38",
          6218 => x"e6",
          6219 => x"80",
          6220 => x"51",
          6221 => x"08",
          6222 => x"94",
          6223 => x"27",
          6224 => x"0c",
          6225 => x"84",
          6226 => x"ff",
          6227 => x"79",
          6228 => x"08",
          6229 => x"90",
          6230 => x"3d",
          6231 => x"ff",
          6232 => x"56",
          6233 => x"38",
          6234 => x"0d",
          6235 => x"70",
          6236 => x"bb",
          6237 => x"8b",
          6238 => x"9f",
          6239 => x"84",
          6240 => x"80",
          6241 => x"06",
          6242 => x"38",
          6243 => x"52",
          6244 => x"84",
          6245 => x"08",
          6246 => x"08",
          6247 => x"84",
          6248 => x"81",
          6249 => x"83",
          6250 => x"e2",
          6251 => x"05",
          6252 => x"8d",
          6253 => x"b0",
          6254 => x"18",
          6255 => x"57",
          6256 => x"34",
          6257 => x"58",
          6258 => x"81",
          6259 => x"78",
          6260 => x"82",
          6261 => x"38",
          6262 => x"ff",
          6263 => x"53",
          6264 => x"52",
          6265 => x"84",
          6266 => x"84",
          6267 => x"a8",
          6268 => x"08",
          6269 => x"5b",
          6270 => x"e1",
          6271 => x"18",
          6272 => x"33",
          6273 => x"39",
          6274 => x"81",
          6275 => x"18",
          6276 => x"7c",
          6277 => x"84",
          6278 => x"2e",
          6279 => x"81",
          6280 => x"08",
          6281 => x"74",
          6282 => x"84",
          6283 => x"17",
          6284 => x"5c",
          6285 => x"18",
          6286 => x"07",
          6287 => x"78",
          6288 => x"bb",
          6289 => x"17",
          6290 => x"57",
          6291 => x"06",
          6292 => x"56",
          6293 => x"34",
          6294 => x"57",
          6295 => x"90",
          6296 => x"75",
          6297 => x"1a",
          6298 => x"80",
          6299 => x"7c",
          6300 => x"80",
          6301 => x"7a",
          6302 => x"74",
          6303 => x"a0",
          6304 => x"58",
          6305 => x"77",
          6306 => x"56",
          6307 => x"80",
          6308 => x"ff",
          6309 => x"f2",
          6310 => x"80",
          6311 => x"83",
          6312 => x"0b",
          6313 => x"cf",
          6314 => x"bb",
          6315 => x"84",
          6316 => x"bb",
          6317 => x"98",
          6318 => x"34",
          6319 => x"34",
          6320 => x"34",
          6321 => x"d9",
          6322 => x"34",
          6323 => x"7d",
          6324 => x"84",
          6325 => x"9f",
          6326 => x"74",
          6327 => x"57",
          6328 => x"39",
          6329 => x"17",
          6330 => x"cd",
          6331 => x"d8",
          6332 => x"a1",
          6333 => x"18",
          6334 => x"18",
          6335 => x"34",
          6336 => x"7d",
          6337 => x"84",
          6338 => x"0d",
          6339 => x"5b",
          6340 => x"70",
          6341 => x"56",
          6342 => x"74",
          6343 => x"38",
          6344 => x"52",
          6345 => x"84",
          6346 => x"08",
          6347 => x"84",
          6348 => x"3d",
          6349 => x"70",
          6350 => x"bb",
          6351 => x"dc",
          6352 => x"a0",
          6353 => x"a0",
          6354 => x"58",
          6355 => x"77",
          6356 => x"55",
          6357 => x"78",
          6358 => x"05",
          6359 => x"34",
          6360 => x"3d",
          6361 => x"3f",
          6362 => x"84",
          6363 => x"08",
          6364 => x"bb",
          6365 => x"33",
          6366 => x"57",
          6367 => x"17",
          6368 => x"59",
          6369 => x"7f",
          6370 => x"5d",
          6371 => x"05",
          6372 => x"33",
          6373 => x"99",
          6374 => x"ff",
          6375 => x"77",
          6376 => x"81",
          6377 => x"9f",
          6378 => x"81",
          6379 => x"78",
          6380 => x"9f",
          6381 => x"80",
          6382 => x"5e",
          6383 => x"7c",
          6384 => x"7b",
          6385 => x"0c",
          6386 => x"52",
          6387 => x"84",
          6388 => x"08",
          6389 => x"aa",
          6390 => x"ac",
          6391 => x"84",
          6392 => x"08",
          6393 => x"8d",
          6394 => x"58",
          6395 => x"33",
          6396 => x"1a",
          6397 => x"05",
          6398 => x"70",
          6399 => x"89",
          6400 => x"19",
          6401 => x"34",
          6402 => x"06",
          6403 => x"38",
          6404 => x"38",
          6405 => x"71",
          6406 => x"5c",
          6407 => x"fe",
          6408 => x"56",
          6409 => x"17",
          6410 => x"05",
          6411 => x"38",
          6412 => x"76",
          6413 => x"7e",
          6414 => x"b8",
          6415 => x"e4",
          6416 => x"2e",
          6417 => x"b4",
          6418 => x"18",
          6419 => x"15",
          6420 => x"06",
          6421 => x"06",
          6422 => x"7b",
          6423 => x"34",
          6424 => x"81",
          6425 => x"7d",
          6426 => x"56",
          6427 => x"81",
          6428 => x"3d",
          6429 => x"74",
          6430 => x"51",
          6431 => x"08",
          6432 => x"38",
          6433 => x"80",
          6434 => x"38",
          6435 => x"7a",
          6436 => x"81",
          6437 => x"16",
          6438 => x"bb",
          6439 => x"57",
          6440 => x"55",
          6441 => x"e5",
          6442 => x"90",
          6443 => x"52",
          6444 => x"bb",
          6445 => x"80",
          6446 => x"84",
          6447 => x"f9",
          6448 => x"3f",
          6449 => x"0c",
          6450 => x"bb",
          6451 => x"18",
          6452 => x"71",
          6453 => x"5c",
          6454 => x"84",
          6455 => x"08",
          6456 => x"bb",
          6457 => x"54",
          6458 => x"16",
          6459 => x"58",
          6460 => x"81",
          6461 => x"08",
          6462 => x"17",
          6463 => x"55",
          6464 => x"38",
          6465 => x"09",
          6466 => x"b4",
          6467 => x"7b",
          6468 => x"82",
          6469 => x"54",
          6470 => x"53",
          6471 => x"ea",
          6472 => x"fc",
          6473 => x"18",
          6474 => x"31",
          6475 => x"a0",
          6476 => x"17",
          6477 => x"06",
          6478 => x"08",
          6479 => x"81",
          6480 => x"79",
          6481 => x"02",
          6482 => x"80",
          6483 => x"96",
          6484 => x"ff",
          6485 => x"56",
          6486 => x"38",
          6487 => x"0d",
          6488 => x"d0",
          6489 => x"bb",
          6490 => x"e0",
          6491 => x"a0",
          6492 => x"74",
          6493 => x"33",
          6494 => x"56",
          6495 => x"55",
          6496 => x"fe",
          6497 => x"84",
          6498 => x"ec",
          6499 => x"3d",
          6500 => x"a2",
          6501 => x"84",
          6502 => x"74",
          6503 => x"04",
          6504 => x"05",
          6505 => x"84",
          6506 => x"38",
          6507 => x"06",
          6508 => x"84",
          6509 => x"2b",
          6510 => x"34",
          6511 => x"34",
          6512 => x"34",
          6513 => x"34",
          6514 => x"78",
          6515 => x"84",
          6516 => x"0d",
          6517 => x"5b",
          6518 => x"9b",
          6519 => x"bb",
          6520 => x"70",
          6521 => x"51",
          6522 => x"81",
          6523 => x"a4",
          6524 => x"25",
          6525 => x"38",
          6526 => x"80",
          6527 => x"08",
          6528 => x"77",
          6529 => x"7a",
          6530 => x"06",
          6531 => x"b8",
          6532 => x"dd",
          6533 => x"2e",
          6534 => x"b4",
          6535 => x"7c",
          6536 => x"74",
          6537 => x"74",
          6538 => x"18",
          6539 => x"33",
          6540 => x"81",
          6541 => x"75",
          6542 => x"5e",
          6543 => x"0c",
          6544 => x"40",
          6545 => x"fe",
          6546 => x"57",
          6547 => x"8d",
          6548 => x"fe",
          6549 => x"fe",
          6550 => x"53",
          6551 => x"52",
          6552 => x"84",
          6553 => x"06",
          6554 => x"83",
          6555 => x"08",
          6556 => x"74",
          6557 => x"82",
          6558 => x"81",
          6559 => x"16",
          6560 => x"52",
          6561 => x"3f",
          6562 => x"16",
          6563 => x"8b",
          6564 => x"fe",
          6565 => x"74",
          6566 => x"84",
          6567 => x"e1",
          6568 => x"84",
          6569 => x"81",
          6570 => x"33",
          6571 => x"27",
          6572 => x"80",
          6573 => x"38",
          6574 => x"57",
          6575 => x"e1",
          6576 => x"3d",
          6577 => x"05",
          6578 => x"3f",
          6579 => x"84",
          6580 => x"8b",
          6581 => x"05",
          6582 => x"38",
          6583 => x"81",
          6584 => x"78",
          6585 => x"3d",
          6586 => x"18",
          6587 => x"7c",
          6588 => x"ff",
          6589 => x"b5",
          6590 => x"dc",
          6591 => x"ff",
          6592 => x"38",
          6593 => x"33",
          6594 => x"78",
          6595 => x"78",
          6596 => x"33",
          6597 => x"74",
          6598 => x"09",
          6599 => x"06",
          6600 => x"77",
          6601 => x"81",
          6602 => x"38",
          6603 => x"81",
          6604 => x"7b",
          6605 => x"a3",
          6606 => x"06",
          6607 => x"fe",
          6608 => x"56",
          6609 => x"80",
          6610 => x"79",
          6611 => x"2e",
          6612 => x"5a",
          6613 => x"80",
          6614 => x"f0",
          6615 => x"84",
          6616 => x"74",
          6617 => x"3d",
          6618 => x"9e",
          6619 => x"ff",
          6620 => x"86",
          6621 => x"3d",
          6622 => x"fe",
          6623 => x"f5",
          6624 => x"84",
          6625 => x"80",
          6626 => x"59",
          6627 => x"33",
          6628 => x"15",
          6629 => x"0b",
          6630 => x"a5",
          6631 => x"56",
          6632 => x"8a",
          6633 => x"bb",
          6634 => x"fe",
          6635 => x"fe",
          6636 => x"52",
          6637 => x"84",
          6638 => x"2e",
          6639 => x"bb",
          6640 => x"16",
          6641 => x"77",
          6642 => x"74",
          6643 => x"38",
          6644 => x"81",
          6645 => x"84",
          6646 => x"ff",
          6647 => x"78",
          6648 => x"08",
          6649 => x"e5",
          6650 => x"80",
          6651 => x"2e",
          6652 => x"81",
          6653 => x"fe",
          6654 => x"57",
          6655 => x"86",
          6656 => x"bf",
          6657 => x"a0",
          6658 => x"05",
          6659 => x"38",
          6660 => x"8b",
          6661 => x"81",
          6662 => x"58",
          6663 => x"fd",
          6664 => x"33",
          6665 => x"15",
          6666 => x"6b",
          6667 => x"0b",
          6668 => x"f5",
          6669 => x"ce",
          6670 => x"54",
          6671 => x"18",
          6672 => x"bb",
          6673 => x"80",
          6674 => x"19",
          6675 => x"31",
          6676 => x"38",
          6677 => x"b1",
          6678 => x"e8",
          6679 => x"fe",
          6680 => x"57",
          6681 => x"b6",
          6682 => x"59",
          6683 => x"a1",
          6684 => x"19",
          6685 => x"33",
          6686 => x"39",
          6687 => x"05",
          6688 => x"89",
          6689 => x"08",
          6690 => x"33",
          6691 => x"15",
          6692 => x"78",
          6693 => x"5f",
          6694 => x"56",
          6695 => x"81",
          6696 => x"38",
          6697 => x"06",
          6698 => x"38",
          6699 => x"70",
          6700 => x"86",
          6701 => x"30",
          6702 => x"84",
          6703 => x"53",
          6704 => x"38",
          6705 => x"82",
          6706 => x"74",
          6707 => x"81",
          6708 => x"75",
          6709 => x"84",
          6710 => x"bb",
          6711 => x"84",
          6712 => x"19",
          6713 => x"78",
          6714 => x"56",
          6715 => x"90",
          6716 => x"84",
          6717 => x"33",
          6718 => x"84",
          6719 => x"38",
          6720 => x"39",
          6721 => x"7d",
          6722 => x"81",
          6723 => x"38",
          6724 => x"de",
          6725 => x"84",
          6726 => x"81",
          6727 => x"d7",
          6728 => x"7b",
          6729 => x"18",
          6730 => x"33",
          6731 => x"34",
          6732 => x"08",
          6733 => x"38",
          6734 => x"15",
          6735 => x"34",
          6736 => x"ff",
          6737 => x"be",
          6738 => x"54",
          6739 => x"a1",
          6740 => x"0d",
          6741 => x"88",
          6742 => x"5f",
          6743 => x"5b",
          6744 => x"79",
          6745 => x"26",
          6746 => x"38",
          6747 => x"92",
          6748 => x"76",
          6749 => x"84",
          6750 => x"74",
          6751 => x"75",
          6752 => x"ba",
          6753 => x"52",
          6754 => x"bb",
          6755 => x"06",
          6756 => x"38",
          6757 => x"57",
          6758 => x"05",
          6759 => x"e9",
          6760 => x"38",
          6761 => x"38",
          6762 => x"38",
          6763 => x"ff",
          6764 => x"80",
          6765 => x"80",
          6766 => x"7f",
          6767 => x"89",
          6768 => x"89",
          6769 => x"80",
          6770 => x"80",
          6771 => x"74",
          6772 => x"df",
          6773 => x"79",
          6774 => x"84",
          6775 => x"83",
          6776 => x"33",
          6777 => x"57",
          6778 => x"06",
          6779 => x"05",
          6780 => x"80",
          6781 => x"83",
          6782 => x"2b",
          6783 => x"70",
          6784 => x"07",
          6785 => x"12",
          6786 => x"07",
          6787 => x"2b",
          6788 => x"0c",
          6789 => x"44",
          6790 => x"4b",
          6791 => x"27",
          6792 => x"80",
          6793 => x"70",
          6794 => x"83",
          6795 => x"82",
          6796 => x"66",
          6797 => x"4a",
          6798 => x"8a",
          6799 => x"2a",
          6800 => x"56",
          6801 => x"77",
          6802 => x"77",
          6803 => x"58",
          6804 => x"27",
          6805 => x"ff",
          6806 => x"84",
          6807 => x"f5",
          6808 => x"84",
          6809 => x"71",
          6810 => x"43",
          6811 => x"5c",
          6812 => x"05",
          6813 => x"72",
          6814 => x"2e",
          6815 => x"90",
          6816 => x"74",
          6817 => x"31",
          6818 => x"52",
          6819 => x"84",
          6820 => x"38",
          6821 => x"dd",
          6822 => x"84",
          6823 => x"f9",
          6824 => x"26",
          6825 => x"39",
          6826 => x"9f",
          6827 => x"81",
          6828 => x"bb",
          6829 => x"90",
          6830 => x"81",
          6831 => x"26",
          6832 => x"06",
          6833 => x"81",
          6834 => x"5f",
          6835 => x"70",
          6836 => x"05",
          6837 => x"57",
          6838 => x"70",
          6839 => x"18",
          6840 => x"18",
          6841 => x"30",
          6842 => x"2e",
          6843 => x"be",
          6844 => x"72",
          6845 => x"4a",
          6846 => x"1c",
          6847 => x"ff",
          6848 => x"9f",
          6849 => x"51",
          6850 => x"bb",
          6851 => x"2a",
          6852 => x"56",
          6853 => x"8e",
          6854 => x"74",
          6855 => x"56",
          6856 => x"ba",
          6857 => x"f9",
          6858 => x"57",
          6859 => x"6e",
          6860 => x"39",
          6861 => x"9d",
          6862 => x"81",
          6863 => x"57",
          6864 => x"0d",
          6865 => x"62",
          6866 => x"60",
          6867 => x"8e",
          6868 => x"61",
          6869 => x"58",
          6870 => x"8b",
          6871 => x"76",
          6872 => x"81",
          6873 => x"ef",
          6874 => x"34",
          6875 => x"8d",
          6876 => x"4b",
          6877 => x"2a",
          6878 => x"61",
          6879 => x"30",
          6880 => x"78",
          6881 => x"92",
          6882 => x"ff",
          6883 => x"ff",
          6884 => x"74",
          6885 => x"34",
          6886 => x"98",
          6887 => x"ff",
          6888 => x"05",
          6889 => x"88",
          6890 => x"7e",
          6891 => x"34",
          6892 => x"84",
          6893 => x"62",
          6894 => x"a7",
          6895 => x"a1",
          6896 => x"aa",
          6897 => x"55",
          6898 => x"2a",
          6899 => x"80",
          6900 => x"05",
          6901 => x"cc",
          6902 => x"58",
          6903 => x"ff",
          6904 => x"fe",
          6905 => x"83",
          6906 => x"81",
          6907 => x"fe",
          6908 => x"84",
          6909 => x"62",
          6910 => x"57",
          6911 => x"34",
          6912 => x"75",
          6913 => x"38",
          6914 => x"2e",
          6915 => x"76",
          6916 => x"70",
          6917 => x"59",
          6918 => x"76",
          6919 => x"57",
          6920 => x"76",
          6921 => x"79",
          6922 => x"84",
          6923 => x"57",
          6924 => x"34",
          6925 => x"1b",
          6926 => x"38",
          6927 => x"ff",
          6928 => x"83",
          6929 => x"26",
          6930 => x"53",
          6931 => x"3f",
          6932 => x"74",
          6933 => x"db",
          6934 => x"38",
          6935 => x"8a",
          6936 => x"38",
          6937 => x"83",
          6938 => x"38",
          6939 => x"70",
          6940 => x"78",
          6941 => x"aa",
          6942 => x"78",
          6943 => x"81",
          6944 => x"05",
          6945 => x"43",
          6946 => x"fc",
          6947 => x"34",
          6948 => x"07",
          6949 => x"bb",
          6950 => x"61",
          6951 => x"c7",
          6952 => x"34",
          6953 => x"05",
          6954 => x"62",
          6955 => x"05",
          6956 => x"83",
          6957 => x"7e",
          6958 => x"78",
          6959 => x"aa",
          6960 => x"f7",
          6961 => x"51",
          6962 => x"bb",
          6963 => x"84",
          6964 => x"0d",
          6965 => x"f9",
          6966 => x"5c",
          6967 => x"91",
          6968 => x"22",
          6969 => x"74",
          6970 => x"56",
          6971 => x"57",
          6972 => x"75",
          6973 => x"fc",
          6974 => x"10",
          6975 => x"5e",
          6976 => x"84",
          6977 => x"fd",
          6978 => x"38",
          6979 => x"84",
          6980 => x"38",
          6981 => x"5b",
          6982 => x"c8",
          6983 => x"2e",
          6984 => x"39",
          6985 => x"2a",
          6986 => x"90",
          6987 => x"75",
          6988 => x"34",
          6989 => x"05",
          6990 => x"a1",
          6991 => x"61",
          6992 => x"05",
          6993 => x"a5",
          6994 => x"61",
          6995 => x"75",
          6996 => x"05",
          6997 => x"61",
          6998 => x"34",
          6999 => x"b1",
          7000 => x"80",
          7001 => x"80",
          7002 => x"05",
          7003 => x"e6",
          7004 => x"05",
          7005 => x"34",
          7006 => x"cd",
          7007 => x"76",
          7008 => x"55",
          7009 => x"54",
          7010 => x"bf",
          7011 => x"08",
          7012 => x"05",
          7013 => x"76",
          7014 => x"52",
          7015 => x"c3",
          7016 => x"9f",
          7017 => x"f8",
          7018 => x"81",
          7019 => x"05",
          7020 => x"84",
          7021 => x"ff",
          7022 => x"05",
          7023 => x"61",
          7024 => x"34",
          7025 => x"39",
          7026 => x"79",
          7027 => x"61",
          7028 => x"57",
          7029 => x"60",
          7030 => x"5e",
          7031 => x"81",
          7032 => x"81",
          7033 => x"80",
          7034 => x"f2",
          7035 => x"61",
          7036 => x"83",
          7037 => x"7a",
          7038 => x"2a",
          7039 => x"7a",
          7040 => x"05",
          7041 => x"83",
          7042 => x"05",
          7043 => x"76",
          7044 => x"83",
          7045 => x"ff",
          7046 => x"53",
          7047 => x"3f",
          7048 => x"79",
          7049 => x"57",
          7050 => x"7e",
          7051 => x"05",
          7052 => x"38",
          7053 => x"54",
          7054 => x"9b",
          7055 => x"06",
          7056 => x"8d",
          7057 => x"05",
          7058 => x"2e",
          7059 => x"80",
          7060 => x"76",
          7061 => x"3d",
          7062 => x"84",
          7063 => x"8a",
          7064 => x"56",
          7065 => x"08",
          7066 => x"75",
          7067 => x"8e",
          7068 => x"88",
          7069 => x"3d",
          7070 => x"52",
          7071 => x"74",
          7072 => x"9f",
          7073 => x"1c",
          7074 => x"39",
          7075 => x"ff",
          7076 => x"ff",
          7077 => x"cc",
          7078 => x"05",
          7079 => x"38",
          7080 => x"2e",
          7081 => x"24",
          7082 => x"05",
          7083 => x"55",
          7084 => x"18",
          7085 => x"55",
          7086 => x"ff",
          7087 => x"52",
          7088 => x"84",
          7089 => x"2e",
          7090 => x"0c",
          7091 => x"b0",
          7092 => x"76",
          7093 => x"7b",
          7094 => x"2a",
          7095 => x"a5",
          7096 => x"3f",
          7097 => x"0c",
          7098 => x"75",
          7099 => x"53",
          7100 => x"38",
          7101 => x"84",
          7102 => x"83",
          7103 => x"b5",
          7104 => x"80",
          7105 => x"51",
          7106 => x"70",
          7107 => x"80",
          7108 => x"e8",
          7109 => x"39",
          7110 => x"84",
          7111 => x"04",
          7112 => x"02",
          7113 => x"80",
          7114 => x"70",
          7115 => x"3d",
          7116 => x"81",
          7117 => x"e9",
          7118 => x"70",
          7119 => x"3d",
          7120 => x"70",
          7121 => x"70",
          7122 => x"56",
          7123 => x"38",
          7124 => x"71",
          7125 => x"07",
          7126 => x"71",
          7127 => x"88",
          7128 => x"14",
          7129 => x"71",
          7130 => x"82",
          7131 => x"80",
          7132 => x"52",
          7133 => x"70",
          7134 => x"04",
          7135 => x"71",
          7136 => x"83",
          7137 => x"c7",
          7138 => x"57",
          7139 => x"16",
          7140 => x"f1",
          7141 => x"06",
          7142 => x"83",
          7143 => x"d0",
          7144 => x"51",
          7145 => x"ff",
          7146 => x"70",
          7147 => x"b9",
          7148 => x"71",
          7149 => x"52",
          7150 => x"10",
          7151 => x"ef",
          7152 => x"ff",
          7153 => x"ff",
          7154 => x"8b",
          7155 => x"75",
          7156 => x"5f",
          7157 => x"49",
          7158 => x"33",
          7159 => x"1d",
          7160 => x"07",
          7161 => x"f1",
          7162 => x"db",
          7163 => x"c5",
          7164 => x"ca",
          7165 => x"64",
          7166 => x"64",
          7167 => x"64",
          7168 => x"64",
          7169 => x"64",
          7170 => x"64",
          7171 => x"64",
          7172 => x"64",
          7173 => x"64",
          7174 => x"64",
          7175 => x"64",
          7176 => x"64",
          7177 => x"64",
          7178 => x"64",
          7179 => x"64",
          7180 => x"64",
          7181 => x"64",
          7182 => x"64",
          7183 => x"64",
          7184 => x"64",
          7185 => x"64",
          7186 => x"64",
          7187 => x"64",
          7188 => x"64",
          7189 => x"64",
          7190 => x"64",
          7191 => x"64",
          7192 => x"64",
          7193 => x"64",
          7194 => x"17",
          7195 => x"64",
          7196 => x"b8",
          7197 => x"3c",
          7198 => x"64",
          7199 => x"64",
          7200 => x"64",
          7201 => x"64",
          7202 => x"64",
          7203 => x"64",
          7204 => x"64",
          7205 => x"64",
          7206 => x"64",
          7207 => x"64",
          7208 => x"64",
          7209 => x"64",
          7210 => x"64",
          7211 => x"64",
          7212 => x"64",
          7213 => x"64",
          7214 => x"64",
          7215 => x"64",
          7216 => x"64",
          7217 => x"64",
          7218 => x"64",
          7219 => x"64",
          7220 => x"64",
          7221 => x"64",
          7222 => x"64",
          7223 => x"64",
          7224 => x"bb",
          7225 => x"64",
          7226 => x"64",
          7227 => x"64",
          7228 => x"64",
          7229 => x"73",
          7230 => x"64",
          7231 => x"64",
          7232 => x"56",
          7233 => x"33",
          7234 => x"57",
          7235 => x"6f",
          7236 => x"10",
          7237 => x"62",
          7238 => x"ac",
          7239 => x"fc",
          7240 => x"44",
          7241 => x"59",
          7242 => x"fd",
          7243 => x"6c",
          7244 => x"fd",
          7245 => x"59",
          7246 => x"b5",
          7247 => x"44",
          7248 => x"82",
          7249 => x"04",
          7250 => x"1d",
          7251 => x"2a",
          7252 => x"2a",
          7253 => x"2a",
          7254 => x"03",
          7255 => x"2a",
          7256 => x"2a",
          7257 => x"2a",
          7258 => x"2a",
          7259 => x"2a",
          7260 => x"2a",
          7261 => x"2a",
          7262 => x"2a",
          7263 => x"2a",
          7264 => x"2a",
          7265 => x"2a",
          7266 => x"30",
          7267 => x"0a",
          7268 => x"f8",
          7269 => x"4d",
          7270 => x"4d",
          7271 => x"52",
          7272 => x"5c",
          7273 => x"b1",
          7274 => x"90",
          7275 => x"34",
          7276 => x"3f",
          7277 => x"68",
          7278 => x"24",
          7279 => x"ca",
          7280 => x"a4",
          7281 => x"51",
          7282 => x"51",
          7283 => x"51",
          7284 => x"6d",
          7285 => x"32",
          7286 => x"51",
          7287 => x"51",
          7288 => x"51",
          7289 => x"51",
          7290 => x"51",
          7291 => x"51",
          7292 => x"51",
          7293 => x"51",
          7294 => x"51",
          7295 => x"ef",
          7296 => x"51",
          7297 => x"92",
          7298 => x"43",
          7299 => x"51",
          7300 => x"51",
          7301 => x"51",
          7302 => x"74",
          7303 => x"e9",
          7304 => x"e9",
          7305 => x"e9",
          7306 => x"e9",
          7307 => x"e9",
          7308 => x"e9",
          7309 => x"e9",
          7310 => x"e9",
          7311 => x"e9",
          7312 => x"e9",
          7313 => x"e9",
          7314 => x"e9",
          7315 => x"e9",
          7316 => x"e9",
          7317 => x"86",
          7318 => x"bb",
          7319 => x"96",
          7320 => x"46",
          7321 => x"e9",
          7322 => x"16",
          7323 => x"f2",
          7324 => x"51",
          7325 => x"2f",
          7326 => x"e9",
          7327 => x"43",
          7328 => x"9f",
          7329 => x"9f",
          7330 => x"9f",
          7331 => x"9f",
          7332 => x"9f",
          7333 => x"9f",
          7334 => x"c1",
          7335 => x"9f",
          7336 => x"9f",
          7337 => x"9f",
          7338 => x"9f",
          7339 => x"18",
          7340 => x"2f",
          7341 => x"01",
          7342 => x"61",
          7343 => x"4a",
          7344 => x"34",
          7345 => x"1d",
          7346 => x"01",
          7347 => x"fd",
          7348 => x"fd",
          7349 => x"fd",
          7350 => x"fd",
          7351 => x"fd",
          7352 => x"fd",
          7353 => x"0d",
          7354 => x"fd",
          7355 => x"fd",
          7356 => x"fd",
          7357 => x"fd",
          7358 => x"fd",
          7359 => x"fd",
          7360 => x"fd",
          7361 => x"fd",
          7362 => x"fd",
          7363 => x"fd",
          7364 => x"fd",
          7365 => x"fd",
          7366 => x"fd",
          7367 => x"fd",
          7368 => x"fd",
          7369 => x"fd",
          7370 => x"fd",
          7371 => x"fd",
          7372 => x"fd",
          7373 => x"fd",
          7374 => x"17",
          7375 => x"fd",
          7376 => x"fd",
          7377 => x"fd",
          7378 => x"fd",
          7379 => x"fd",
          7380 => x"e1",
          7381 => x"b8",
          7382 => x"fd",
          7383 => x"fd",
          7384 => x"ff",
          7385 => x"fd",
          7386 => x"0f",
          7387 => x"fd",
          7388 => x"fd",
          7389 => x"fd",
          7390 => x"17",
          7391 => x"00",
          7392 => x"00",
          7393 => x"00",
          7394 => x"00",
          7395 => x"00",
          7396 => x"00",
          7397 => x"00",
          7398 => x"00",
          7399 => x"00",
          7400 => x"00",
          7401 => x"00",
          7402 => x"00",
          7403 => x"6c",
          7404 => x"00",
          7405 => x"00",
          7406 => x"00",
          7407 => x"00",
          7408 => x"00",
          7409 => x"00",
          7410 => x"00",
          7411 => x"00",
          7412 => x"00",
          7413 => x"6e",
          7414 => x"6f",
          7415 => x"61",
          7416 => x"69",
          7417 => x"74",
          7418 => x"20",
          7419 => x"65",
          7420 => x"2e",
          7421 => x"75",
          7422 => x"74",
          7423 => x"2e",
          7424 => x"65",
          7425 => x"6b",
          7426 => x"65",
          7427 => x"65",
          7428 => x"63",
          7429 => x"64",
          7430 => x"6d",
          7431 => x"74",
          7432 => x"63",
          7433 => x"6c",
          7434 => x"79",
          7435 => x"75",
          7436 => x"69",
          7437 => x"6b",
          7438 => x"61",
          7439 => x"00",
          7440 => x"75",
          7441 => x"20",
          7442 => x"2e",
          7443 => x"69",
          7444 => x"20",
          7445 => x"65",
          7446 => x"65",
          7447 => x"20",
          7448 => x"2e",
          7449 => x"65",
          7450 => x"79",
          7451 => x"2e",
          7452 => x"65",
          7453 => x"65",
          7454 => x"61",
          7455 => x"65",
          7456 => x"00",
          7457 => x"20",
          7458 => x"00",
          7459 => x"20",
          7460 => x"00",
          7461 => x"74",
          7462 => x"00",
          7463 => x"6c",
          7464 => x"00",
          7465 => x"72",
          7466 => x"63",
          7467 => x"00",
          7468 => x"74",
          7469 => x"74",
          7470 => x"74",
          7471 => x"0a",
          7472 => x"64",
          7473 => x"6c",
          7474 => x"00",
          7475 => x"00",
          7476 => x"00",
          7477 => x"58",
          7478 => x"20",
          7479 => x"00",
          7480 => x"25",
          7481 => x"30",
          7482 => x"00",
          7483 => x"00",
          7484 => x"65",
          7485 => x"20",
          7486 => x"2a",
          7487 => x"00",
          7488 => x"65",
          7489 => x"73",
          7490 => x"20",
          7491 => x"25",
          7492 => x"00",
          7493 => x"20",
          7494 => x"20",
          7495 => x"20",
          7496 => x"25",
          7497 => x"00",
          7498 => x"65",
          7499 => x"61",
          7500 => x"00",
          7501 => x"58",
          7502 => x"75",
          7503 => x"54",
          7504 => x"74",
          7505 => x"00",
          7506 => x"58",
          7507 => x"75",
          7508 => x"54",
          7509 => x"74",
          7510 => x"00",
          7511 => x"52",
          7512 => x"75",
          7513 => x"54",
          7514 => x"74",
          7515 => x"00",
          7516 => x"65",
          7517 => x"00",
          7518 => x"6e",
          7519 => x"00",
          7520 => x"20",
          7521 => x"72",
          7522 => x"62",
          7523 => x"6d",
          7524 => x"00",
          7525 => x"63",
          7526 => x"00",
          7527 => x"2e",
          7528 => x"6c",
          7529 => x"6e",
          7530 => x"65",
          7531 => x"64",
          7532 => x"61",
          7533 => x"20",
          7534 => x"79",
          7535 => x"00",
          7536 => x"00",
          7537 => x"20",
          7538 => x"2e",
          7539 => x"00",
          7540 => x"5c",
          7541 => x"73",
          7542 => x"64",
          7543 => x"69",
          7544 => x"00",
          7545 => x"69",
          7546 => x"69",
          7547 => x"2e",
          7548 => x"6c",
          7549 => x"65",
          7550 => x"78",
          7551 => x"00",
          7552 => x"74",
          7553 => x"6f",
          7554 => x"2e",
          7555 => x"63",
          7556 => x"6f",
          7557 => x"38",
          7558 => x"00",
          7559 => x"30",
          7560 => x"00",
          7561 => x"30",
          7562 => x"70",
          7563 => x"2e",
          7564 => x"6c",
          7565 => x"2d",
          7566 => x"25",
          7567 => x"00",
          7568 => x"2e",
          7569 => x"6c",
          7570 => x"00",
          7571 => x"67",
          7572 => x"00",
          7573 => x"6d",
          7574 => x"6d",
          7575 => x"00",
          7576 => x"25",
          7577 => x"6f",
          7578 => x"75",
          7579 => x"61",
          7580 => x"6f",
          7581 => x"6d",
          7582 => x"00",
          7583 => x"25",
          7584 => x"3a",
          7585 => x"64",
          7586 => x"20",
          7587 => x"72",
          7588 => x"00",
          7589 => x"65",
          7590 => x"6d",
          7591 => x"00",
          7592 => x"65",
          7593 => x"20",
          7594 => x"65",
          7595 => x"72",
          7596 => x"73",
          7597 => x"0a",
          7598 => x"20",
          7599 => x"6f",
          7600 => x"74",
          7601 => x"73",
          7602 => x"0a",
          7603 => x"20",
          7604 => x"74",
          7605 => x"72",
          7606 => x"20",
          7607 => x"0a",
          7608 => x"63",
          7609 => x"20",
          7610 => x"20",
          7611 => x"20",
          7612 => x"20",
          7613 => x"0a",
          7614 => x"20",
          7615 => x"43",
          7616 => x"65",
          7617 => x"20",
          7618 => x"30",
          7619 => x"00",
          7620 => x"68",
          7621 => x"52",
          7622 => x"6b",
          7623 => x"25",
          7624 => x"48",
          7625 => x"20",
          7626 => x"6c",
          7627 => x"71",
          7628 => x"20",
          7629 => x"30",
          7630 => x"00",
          7631 => x"00",
          7632 => x"00",
          7633 => x"54",
          7634 => x"20",
          7635 => x"00",
          7636 => x"48",
          7637 => x"53",
          7638 => x"20",
          7639 => x"52",
          7640 => x"6e",
          7641 => x"64",
          7642 => x"20",
          7643 => x"20",
          7644 => x"72",
          7645 => x"64",
          7646 => x"20",
          7647 => x"20",
          7648 => x"63",
          7649 => x"64",
          7650 => x"20",
          7651 => x"20",
          7652 => x"3a",
          7653 => x"00",
          7654 => x"4d",
          7655 => x"25",
          7656 => x"58",
          7657 => x"20",
          7658 => x"41",
          7659 => x"3a",
          7660 => x"00",
          7661 => x"41",
          7662 => x"25",
          7663 => x"58",
          7664 => x"20",
          7665 => x"4d",
          7666 => x"3a",
          7667 => x"00",
          7668 => x"53",
          7669 => x"69",
          7670 => x"6e",
          7671 => x"6d",
          7672 => x"6c",
          7673 => x"69",
          7674 => x"78",
          7675 => x"00",
          7676 => x"00",
          7677 => x"38",
          7678 => x"03",
          7679 => x"00",
          7680 => x"30",
          7681 => x"05",
          7682 => x"00",
          7683 => x"28",
          7684 => x"07",
          7685 => x"00",
          7686 => x"20",
          7687 => x"08",
          7688 => x"00",
          7689 => x"18",
          7690 => x"09",
          7691 => x"00",
          7692 => x"10",
          7693 => x"0d",
          7694 => x"00",
          7695 => x"08",
          7696 => x"0e",
          7697 => x"00",
          7698 => x"00",
          7699 => x"0f",
          7700 => x"00",
          7701 => x"f8",
          7702 => x"11",
          7703 => x"00",
          7704 => x"f0",
          7705 => x"13",
          7706 => x"00",
          7707 => x"e8",
          7708 => x"15",
          7709 => x"00",
          7710 => x"00",
          7711 => x"7e",
          7712 => x"00",
          7713 => x"7e",
          7714 => x"00",
          7715 => x"00",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"20",
          7721 => x"38",
          7722 => x"6e",
          7723 => x"2f",
          7724 => x"68",
          7725 => x"66",
          7726 => x"73",
          7727 => x"00",
          7728 => x"00",
          7729 => x"00",
          7730 => x"74",
          7731 => x"66",
          7732 => x"78",
          7733 => x"6c",
          7734 => x"00",
          7735 => x"74",
          7736 => x"20",
          7737 => x"74",
          7738 => x"65",
          7739 => x"2e",
          7740 => x"0a",
          7741 => x"7e",
          7742 => x"00",
          7743 => x"00",
          7744 => x"30",
          7745 => x"31",
          7746 => x"32",
          7747 => x"33",
          7748 => x"34",
          7749 => x"35",
          7750 => x"37",
          7751 => x"38",
          7752 => x"39",
          7753 => x"30",
          7754 => x"7e",
          7755 => x"7e",
          7756 => x"00",
          7757 => x"00",
          7758 => x"00",
          7759 => x"2c",
          7760 => x"64",
          7761 => x"78",
          7762 => x"64",
          7763 => x"25",
          7764 => x"2c",
          7765 => x"00",
          7766 => x"00",
          7767 => x"00",
          7768 => x"64",
          7769 => x"6f",
          7770 => x"6f",
          7771 => x"25",
          7772 => x"78",
          7773 => x"25",
          7774 => x"78",
          7775 => x"25",
          7776 => x"00",
          7777 => x"20",
          7778 => x"2e",
          7779 => x"00",
          7780 => x"7f",
          7781 => x"3d",
          7782 => x"00",
          7783 => x"00",
          7784 => x"53",
          7785 => x"4e",
          7786 => x"46",
          7787 => x"00",
          7788 => x"20",
          7789 => x"32",
          7790 => x"1c",
          7791 => x"00",
          7792 => x"07",
          7793 => x"1c",
          7794 => x"41",
          7795 => x"49",
          7796 => x"4f",
          7797 => x"9b",
          7798 => x"55",
          7799 => x"ab",
          7800 => x"b3",
          7801 => x"bb",
          7802 => x"c3",
          7803 => x"cb",
          7804 => x"d3",
          7805 => x"db",
          7806 => x"e3",
          7807 => x"eb",
          7808 => x"f3",
          7809 => x"fb",
          7810 => x"3b",
          7811 => x"3a",
          7812 => x"00",
          7813 => x"40",
          7814 => x"00",
          7815 => x"08",
          7816 => x"00",
          7817 => x"e2",
          7818 => x"e7",
          7819 => x"ef",
          7820 => x"c5",
          7821 => x"f4",
          7822 => x"f9",
          7823 => x"a2",
          7824 => x"92",
          7825 => x"fa",
          7826 => x"ba",
          7827 => x"bd",
          7828 => x"bb",
          7829 => x"02",
          7830 => x"56",
          7831 => x"57",
          7832 => x"10",
          7833 => x"1c",
          7834 => x"5f",
          7835 => x"66",
          7836 => x"67",
          7837 => x"59",
          7838 => x"6b",
          7839 => x"88",
          7840 => x"80",
          7841 => x"c0",
          7842 => x"c4",
          7843 => x"b4",
          7844 => x"29",
          7845 => x"64",
          7846 => x"48",
          7847 => x"1a",
          7848 => x"a0",
          7849 => x"17",
          7850 => x"01",
          7851 => x"32",
          7852 => x"4a",
          7853 => x"80",
          7854 => x"82",
          7855 => x"86",
          7856 => x"8a",
          7857 => x"8e",
          7858 => x"91",
          7859 => x"96",
          7860 => x"3d",
          7861 => x"20",
          7862 => x"a2",
          7863 => x"a6",
          7864 => x"aa",
          7865 => x"ae",
          7866 => x"b2",
          7867 => x"b5",
          7868 => x"ba",
          7869 => x"be",
          7870 => x"c2",
          7871 => x"c4",
          7872 => x"ca",
          7873 => x"10",
          7874 => x"de",
          7875 => x"f1",
          7876 => x"28",
          7877 => x"09",
          7878 => x"3d",
          7879 => x"41",
          7880 => x"53",
          7881 => x"55",
          7882 => x"8f",
          7883 => x"5d",
          7884 => x"61",
          7885 => x"65",
          7886 => x"96",
          7887 => x"6d",
          7888 => x"71",
          7889 => x"9f",
          7890 => x"79",
          7891 => x"64",
          7892 => x"81",
          7893 => x"85",
          7894 => x"44",
          7895 => x"8d",
          7896 => x"91",
          7897 => x"fd",
          7898 => x"04",
          7899 => x"8a",
          7900 => x"02",
          7901 => x"08",
          7902 => x"8e",
          7903 => x"f2",
          7904 => x"f4",
          7905 => x"f7",
          7906 => x"30",
          7907 => x"60",
          7908 => x"c1",
          7909 => x"c0",
          7910 => x"26",
          7911 => x"01",
          7912 => x"a0",
          7913 => x"10",
          7914 => x"30",
          7915 => x"51",
          7916 => x"5b",
          7917 => x"5f",
          7918 => x"0e",
          7919 => x"c9",
          7920 => x"db",
          7921 => x"eb",
          7922 => x"08",
          7923 => x"08",
          7924 => x"b9",
          7925 => x"01",
          7926 => x"e0",
          7927 => x"ec",
          7928 => x"4e",
          7929 => x"10",
          7930 => x"d0",
          7931 => x"60",
          7932 => x"75",
          7933 => x"00",
          7934 => x"00",
          7935 => x"f8",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"08",
          7940 => x"00",
          7941 => x"10",
          7942 => x"00",
          7943 => x"18",
          7944 => x"00",
          7945 => x"20",
          7946 => x"00",
          7947 => x"28",
          7948 => x"00",
          7949 => x"30",
          7950 => x"00",
          7951 => x"38",
          7952 => x"00",
          7953 => x"40",
          7954 => x"00",
          7955 => x"44",
          7956 => x"00",
          7957 => x"48",
          7958 => x"00",
          7959 => x"4c",
          7960 => x"00",
          7961 => x"50",
          7962 => x"00",
          7963 => x"54",
          7964 => x"00",
          7965 => x"58",
          7966 => x"00",
          7967 => x"5c",
          7968 => x"00",
          7969 => x"64",
          7970 => x"00",
          7971 => x"68",
          7972 => x"00",
          7973 => x"70",
          7974 => x"00",
          7975 => x"78",
          7976 => x"00",
          7977 => x"80",
          7978 => x"00",
          7979 => x"88",
          7980 => x"00",
          7981 => x"8c",
          7982 => x"00",
          7983 => x"90",
          7984 => x"00",
          7985 => x"98",
          7986 => x"00",
          7987 => x"a0",
          7988 => x"00",
          7989 => x"a8",
          7990 => x"00",
          7991 => x"00",
          7992 => x"ff",
          7993 => x"ff",
          7994 => x"ff",
          7995 => x"00",
          7996 => x"ff",
          7997 => x"00",
          7998 => x"00",
          7999 => x"00",
          8000 => x"00",
          8001 => x"01",
          8002 => x"00",
          8003 => x"00",
          8004 => x"00",
          8005 => x"00",
          8006 => x"00",
          8007 => x"00",
          8008 => x"00",
          8009 => x"00",
          8010 => x"00",
          8011 => x"00",
          8012 => x"00",
          8013 => x"00",
          8014 => x"00",
          8015 => x"00",
          8016 => x"00",
          8017 => x"00",
          8018 => x"fd",
          8019 => x"5b",
          8020 => x"74",
          8021 => x"6c",
          8022 => x"64",
          8023 => x"34",
          8024 => x"20",
          8025 => x"f4",
          8026 => x"f0",
          8027 => x"83",
          8028 => x"fd",
          8029 => x"5b",
          8030 => x"54",
          8031 => x"4c",
          8032 => x"44",
          8033 => x"34",
          8034 => x"20",
          8035 => x"f4",
          8036 => x"f0",
          8037 => x"83",
          8038 => x"fd",
          8039 => x"7b",
          8040 => x"54",
          8041 => x"4c",
          8042 => x"44",
          8043 => x"24",
          8044 => x"20",
          8045 => x"e1",
          8046 => x"f0",
          8047 => x"88",
          8048 => x"fa",
          8049 => x"1b",
          8050 => x"14",
          8051 => x"0c",
          8052 => x"04",
          8053 => x"f0",
          8054 => x"f0",
          8055 => x"f0",
          8056 => x"f0",
          8057 => x"83",
          8058 => x"c9",
          8059 => x"b3",
          8060 => x"31",
          8061 => x"56",
          8062 => x"48",
          8063 => x"3b",
          8064 => x"00",
          8065 => x"c1",
          8066 => x"f0",
          8067 => x"83",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"ec",
          8083 => x"f4",
          8084 => x"f8",
          8085 => x"fc",
          8086 => x"00",
          8087 => x"04",
          8088 => x"0c",
          8089 => x"14",
          8090 => x"1c",
          8091 => x"24",
          8092 => x"2c",
          8093 => x"34",
          8094 => x"3c",
          8095 => x"44",
          8096 => x"4c",
          8097 => x"54",
          8098 => x"5c",
          8099 => x"64",
          8100 => x"68",
          8101 => x"70",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"19",
          9103 => x"00",
          9104 => x"f7",
          9105 => x"ff",
          9106 => x"e2",
          9107 => x"f4",
          9108 => x"67",
          9109 => x"2d",
          9110 => x"27",
          9111 => x"49",
          9112 => x"07",
          9113 => x"0f",
          9114 => x"17",
          9115 => x"3c",
          9116 => x"87",
          9117 => x"8f",
          9118 => x"97",
          9119 => x"c0",
          9120 => x"00",
          9121 => x"00",
          9122 => x"00",
          9123 => x"00",
          9124 => x"00",
          9125 => x"00",
          9126 => x"00",
          9127 => x"00",
          9128 => x"00",
          9129 => x"00",
          9130 => x"00",
          9131 => x"00",
          9132 => x"00",
          9133 => x"00",
          9134 => x"00",
          9135 => x"01",
          9136 => x"01",
        others => X"00"
    );

    shared variable RAM5 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"88",
             5 => x"88",
             6 => x"00",
             7 => x"00",
             8 => x"06",
             9 => x"2a",
            10 => x"00",
            11 => x"00",
            12 => x"ff",
            13 => x"05",
            14 => x"ff",
            15 => x"04",
            16 => x"73",
            17 => x"73",
            18 => x"04",
            19 => x"00",
            20 => x"07",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"81",
            25 => x"0a",
            26 => x"81",
            27 => x"00",
            28 => x"07",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"00",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"51",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"05",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"06",
            49 => x"ff",
            50 => x"00",
            51 => x"00",
            52 => x"73",
            53 => x"83",
            54 => x"0c",
            55 => x"00",
            56 => x"09",
            57 => x"06",
            58 => x"00",
            59 => x"00",
            60 => x"09",
            61 => x"81",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"53",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"09",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"06",
            77 => x"10",
            78 => x"00",
            79 => x"00",
            80 => x"83",
            81 => x"05",
            82 => x"04",
            83 => x"00",
            84 => x"75",
            85 => x"50",
            86 => x"0c",
            87 => x"00",
            88 => x"75",
            89 => x"50",
            90 => x"0c",
            91 => x"00",
            92 => x"06",
            93 => x"71",
            94 => x"05",
            95 => x"00",
            96 => x"06",
            97 => x"54",
            98 => x"ff",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"05",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"53",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"0b",
           134 => x"a6",
           135 => x"0b",
           136 => x"0b",
           137 => x"e6",
           138 => x"0b",
           139 => x"0b",
           140 => x"a6",
           141 => x"0b",
           142 => x"0b",
           143 => x"e8",
           144 => x"0b",
           145 => x"0b",
           146 => x"ac",
           147 => x"0b",
           148 => x"0b",
           149 => x"f0",
           150 => x"0b",
           151 => x"0b",
           152 => x"b4",
           153 => x"0b",
           154 => x"0b",
           155 => x"f8",
           156 => x"0b",
           157 => x"0b",
           158 => x"bc",
           159 => x"0b",
           160 => x"0b",
           161 => x"80",
           162 => x"0b",
           163 => x"0b",
           164 => x"c4",
           165 => x"0b",
           166 => x"0b",
           167 => x"88",
           168 => x"0b",
           169 => x"0b",
           170 => x"cb",
           171 => x"0b",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"bb",
           193 => x"bb",
           194 => x"84",
           195 => x"bb",
           196 => x"84",
           197 => x"bb",
           198 => x"84",
           199 => x"bb",
           200 => x"84",
           201 => x"bb",
           202 => x"84",
           203 => x"bb",
           204 => x"84",
           205 => x"bb",
           206 => x"84",
           207 => x"bb",
           208 => x"84",
           209 => x"bb",
           210 => x"84",
           211 => x"bb",
           212 => x"84",
           213 => x"bb",
           214 => x"84",
           215 => x"bb",
           216 => x"84",
           217 => x"84",
           218 => x"04",
           219 => x"2d",
           220 => x"90",
           221 => x"b8",
           222 => x"80",
           223 => x"d3",
           224 => x"c0",
           225 => x"82",
           226 => x"80",
           227 => x"0c",
           228 => x"08",
           229 => x"90",
           230 => x"90",
           231 => x"bb",
           232 => x"bb",
           233 => x"84",
           234 => x"84",
           235 => x"04",
           236 => x"2d",
           237 => x"90",
           238 => x"b8",
           239 => x"80",
           240 => x"f2",
           241 => x"c0",
           242 => x"82",
           243 => x"80",
           244 => x"0c",
           245 => x"08",
           246 => x"90",
           247 => x"90",
           248 => x"bb",
           249 => x"bb",
           250 => x"84",
           251 => x"84",
           252 => x"04",
           253 => x"2d",
           254 => x"90",
           255 => x"8c",
           256 => x"80",
           257 => x"96",
           258 => x"c0",
           259 => x"82",
           260 => x"80",
           261 => x"0c",
           262 => x"08",
           263 => x"90",
           264 => x"90",
           265 => x"bb",
           266 => x"bb",
           267 => x"84",
           268 => x"84",
           269 => x"04",
           270 => x"2d",
           271 => x"90",
           272 => x"f8",
           273 => x"80",
           274 => x"c8",
           275 => x"c0",
           276 => x"83",
           277 => x"80",
           278 => x"0c",
           279 => x"08",
           280 => x"90",
           281 => x"90",
           282 => x"bb",
           283 => x"bb",
           284 => x"84",
           285 => x"84",
           286 => x"04",
           287 => x"2d",
           288 => x"90",
           289 => x"ba",
           290 => x"80",
           291 => x"d2",
           292 => x"c0",
           293 => x"80",
           294 => x"80",
           295 => x"0c",
           296 => x"80",
           297 => x"0c",
           298 => x"08",
           299 => x"90",
           300 => x"90",
           301 => x"bb",
           302 => x"bb",
           303 => x"84",
           304 => x"84",
           305 => x"04",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"81",
           311 => x"05",
           312 => x"72",
           313 => x"72",
           314 => x"72",
           315 => x"10",
           316 => x"53",
           317 => x"e6",
           318 => x"84",
           319 => x"ec",
           320 => x"04",
           321 => x"70",
           322 => x"52",
           323 => x"3f",
           324 => x"78",
           325 => x"81",
           326 => x"55",
           327 => x"81",
           328 => x"74",
           329 => x"9f",
           330 => x"74",
           331 => x"38",
           332 => x"84",
           333 => x"2e",
           334 => x"70",
           335 => x"8a",
           336 => x"2a",
           337 => x"cb",
           338 => x"84",
           339 => x"80",
           340 => x"0d",
           341 => x"02",
           342 => x"fe",
           343 => x"7e",
           344 => x"3f",
           345 => x"3d",
           346 => x"88",
           347 => x"3f",
           348 => x"61",
           349 => x"8c",
           350 => x"2a",
           351 => x"ff",
           352 => x"80",
           353 => x"2e",
           354 => x"06",
           355 => x"38",
           356 => x"a3",
           357 => x"80",
           358 => x"72",
           359 => x"70",
           360 => x"80",
           361 => x"5b",
           362 => x"8c",
           363 => x"0c",
           364 => x"54",
           365 => x"70",
           366 => x"81",
           367 => x"98",
           368 => x"79",
           369 => x"53",
           370 => x"58",
           371 => x"39",
           372 => x"38",
           373 => x"7c",
           374 => x"ff",
           375 => x"af",
           376 => x"38",
           377 => x"81",
           378 => x"70",
           379 => x"e0",
           380 => x"38",
           381 => x"54",
           382 => x"59",
           383 => x"52",
           384 => x"33",
           385 => x"c7",
           386 => x"88",
           387 => x"7d",
           388 => x"54",
           389 => x"51",
           390 => x"81",
           391 => x"df",
           392 => x"38",
           393 => x"74",
           394 => x"52",
           395 => x"84",
           396 => x"38",
           397 => x"7b",
           398 => x"8f",
           399 => x"80",
           400 => x"7a",
           401 => x"73",
           402 => x"80",
           403 => x"90",
           404 => x"29",
           405 => x"2c",
           406 => x"54",
           407 => x"98",
           408 => x"78",
           409 => x"ff",
           410 => x"2a",
           411 => x"73",
           412 => x"31",
           413 => x"80",
           414 => x"85",
           415 => x"54",
           416 => x"81",
           417 => x"85",
           418 => x"38",
           419 => x"38",
           420 => x"80",
           421 => x"80",
           422 => x"2c",
           423 => x"38",
           424 => x"77",
           425 => x"80",
           426 => x"73",
           427 => x"53",
           428 => x"81",
           429 => x"70",
           430 => x"25",
           431 => x"ef",
           432 => x"81",
           433 => x"55",
           434 => x"87",
           435 => x"80",
           436 => x"2e",
           437 => x"81",
           438 => x"e2",
           439 => x"38",
           440 => x"5e",
           441 => x"2e",
           442 => x"06",
           443 => x"77",
           444 => x"80",
           445 => x"80",
           446 => x"a0",
           447 => x"90",
           448 => x"58",
           449 => x"39",
           450 => x"57",
           451 => x"7e",
           452 => x"55",
           453 => x"05",
           454 => x"33",
           455 => x"80",
           456 => x"90",
           457 => x"5f",
           458 => x"55",
           459 => x"80",
           460 => x"90",
           461 => x"fe",
           462 => x"f7",
           463 => x"ff",
           464 => x"ff",
           465 => x"70",
           466 => x"3f",
           467 => x"ff",
           468 => x"2e",
           469 => x"81",
           470 => x"e2",
           471 => x"0a",
           472 => x"80",
           473 => x"56",
           474 => x"06",
           475 => x"fe",
           476 => x"08",
           477 => x"24",
           478 => x"06",
           479 => x"39",
           480 => x"76",
           481 => x"88",
           482 => x"76",
           483 => x"60",
           484 => x"56",
           485 => x"75",
           486 => x"08",
           487 => x"90",
           488 => x"fe",
           489 => x"33",
           490 => x"ff",
           491 => x"77",
           492 => x"81",
           493 => x"84",
           494 => x"78",
           495 => x"39",
           496 => x"5b",
           497 => x"77",
           498 => x"80",
           499 => x"80",
           500 => x"a0",
           501 => x"52",
           502 => x"2e",
           503 => x"52",
           504 => x"2a",
           505 => x"8c",
           506 => x"78",
           507 => x"7d",
           508 => x"73",
           509 => x"52",
           510 => x"06",
           511 => x"ff",
           512 => x"51",
           513 => x"7a",
           514 => x"39",
           515 => x"2c",
           516 => x"ab",
           517 => x"52",
           518 => x"39",
           519 => x"84",
           520 => x"78",
           521 => x"f3",
           522 => x"83",
           523 => x"99",
           524 => x"08",
           525 => x"3f",
           526 => x"78",
           527 => x"85",
           528 => x"70",
           529 => x"ff",
           530 => x"80",
           531 => x"33",
           532 => x"e6",
           533 => x"08",
           534 => x"80",
           535 => x"81",
           536 => x"88",
           537 => x"39",
           538 => x"e8",
           539 => x"55",
           540 => x"2e",
           541 => x"84",
           542 => x"fa",
           543 => x"0b",
           544 => x"32",
           545 => x"ff",
           546 => x"92",
           547 => x"53",
           548 => x"38",
           549 => x"88",
           550 => x"55",
           551 => x"74",
           552 => x"72",
           553 => x"e3",
           554 => x"33",
           555 => x"ff",
           556 => x"73",
           557 => x"fa",
           558 => x"70",
           559 => x"56",
           560 => x"73",
           561 => x"2e",
           562 => x"88",
           563 => x"56",
           564 => x"75",
           565 => x"8c",
           566 => x"84",
           567 => x"76",
           568 => x"54",
           569 => x"08",
           570 => x"8c",
           571 => x"3d",
           572 => x"ff",
           573 => x"55",
           574 => x"72",
           575 => x"38",
           576 => x"80",
           577 => x"33",
           578 => x"38",
           579 => x"81",
           580 => x"06",
           581 => x"3d",
           582 => x"72",
           583 => x"05",
           584 => x"bb",
           585 => x"51",
           586 => x"bb",
           587 => x"80",
           588 => x"70",
           589 => x"08",
           590 => x"53",
           591 => x"84",
           592 => x"74",
           593 => x"ff",
           594 => x"77",
           595 => x"05",
           596 => x"12",
           597 => x"51",
           598 => x"70",
           599 => x"85",
           600 => x"79",
           601 => x"80",
           602 => x"38",
           603 => x"81",
           604 => x"55",
           605 => x"73",
           606 => x"04",
           607 => x"38",
           608 => x"ff",
           609 => x"ff",
           610 => x"ff",
           611 => x"73",
           612 => x"c7",
           613 => x"53",
           614 => x"70",
           615 => x"84",
           616 => x"04",
           617 => x"54",
           618 => x"51",
           619 => x"70",
           620 => x"85",
           621 => x"78",
           622 => x"80",
           623 => x"53",
           624 => x"ff",
           625 => x"bb",
           626 => x"3d",
           627 => x"72",
           628 => x"70",
           629 => x"71",
           630 => x"14",
           631 => x"13",
           632 => x"84",
           633 => x"72",
           634 => x"ff",
           635 => x"15",
           636 => x"de",
           637 => x"0c",
           638 => x"84",
           639 => x"0d",
           640 => x"c1",
           641 => x"84",
           642 => x"b2",
           643 => x"bb",
           644 => x"bb",
           645 => x"74",
           646 => x"51",
           647 => x"54",
           648 => x"0d",
           649 => x"71",
           650 => x"9f",
           651 => x"51",
           652 => x"52",
           653 => x"38",
           654 => x"70",
           655 => x"04",
           656 => x"55",
           657 => x"38",
           658 => x"ff",
           659 => x"bb",
           660 => x"3d",
           661 => x"76",
           662 => x"f5",
           663 => x"12",
           664 => x"51",
           665 => x"08",
           666 => x"80",
           667 => x"80",
           668 => x"a0",
           669 => x"54",
           670 => x"38",
           671 => x"10",
           672 => x"9f",
           673 => x"75",
           674 => x"52",
           675 => x"73",
           676 => x"84",
           677 => x"0d",
           678 => x"30",
           679 => x"2b",
           680 => x"83",
           681 => x"25",
           682 => x"2a",
           683 => x"80",
           684 => x"71",
           685 => x"8c",
           686 => x"82",
           687 => x"2a",
           688 => x"82",
           689 => x"bb",
           690 => x"54",
           691 => x"56",
           692 => x"52",
           693 => x"75",
           694 => x"81",
           695 => x"29",
           696 => x"53",
           697 => x"78",
           698 => x"2e",
           699 => x"84",
           700 => x"73",
           701 => x"bd",
           702 => x"52",
           703 => x"38",
           704 => x"81",
           705 => x"76",
           706 => x"56",
           707 => x"74",
           708 => x"78",
           709 => x"81",
           710 => x"ff",
           711 => x"55",
           712 => x"84",
           713 => x"0d",
           714 => x"9f",
           715 => x"32",
           716 => x"72",
           717 => x"56",
           718 => x"75",
           719 => x"88",
           720 => x"7d",
           721 => x"08",
           722 => x"2e",
           723 => x"70",
           724 => x"a0",
           725 => x"f5",
           726 => x"d0",
           727 => x"80",
           728 => x"74",
           729 => x"27",
           730 => x"06",
           731 => x"06",
           732 => x"f9",
           733 => x"89",
           734 => x"27",
           735 => x"81",
           736 => x"56",
           737 => x"78",
           738 => x"75",
           739 => x"84",
           740 => x"16",
           741 => x"59",
           742 => x"ff",
           743 => x"33",
           744 => x"38",
           745 => x"38",
           746 => x"d0",
           747 => x"73",
           748 => x"84",
           749 => x"81",
           750 => x"55",
           751 => x"84",
           752 => x"f7",
           753 => x"70",
           754 => x"56",
           755 => x"8f",
           756 => x"33",
           757 => x"73",
           758 => x"2e",
           759 => x"56",
           760 => x"58",
           761 => x"38",
           762 => x"14",
           763 => x"14",
           764 => x"73",
           765 => x"ff",
           766 => x"89",
           767 => x"77",
           768 => x"0c",
           769 => x"26",
           770 => x"38",
           771 => x"56",
           772 => x"0d",
           773 => x"70",
           774 => x"09",
           775 => x"70",
           776 => x"80",
           777 => x"80",
           778 => x"74",
           779 => x"56",
           780 => x"38",
           781 => x"0d",
           782 => x"0c",
           783 => x"ca",
           784 => x"8b",
           785 => x"84",
           786 => x"bb",
           787 => x"52",
           788 => x"10",
           789 => x"04",
           790 => x"83",
           791 => x"ef",
           792 => x"cf",
           793 => x"0d",
           794 => x"3f",
           795 => x"51",
           796 => x"83",
           797 => x"3d",
           798 => x"fc",
           799 => x"c4",
           800 => x"04",
           801 => x"83",
           802 => x"ee",
           803 => x"d1",
           804 => x"0d",
           805 => x"3f",
           806 => x"51",
           807 => x"83",
           808 => x"3d",
           809 => x"a4",
           810 => x"88",
           811 => x"04",
           812 => x"83",
           813 => x"ee",
           814 => x"d2",
           815 => x"0d",
           816 => x"3f",
           817 => x"51",
           818 => x"fe",
           819 => x"02",
           820 => x"58",
           821 => x"30",
           822 => x"57",
           823 => x"83",
           824 => x"81",
           825 => x"80",
           826 => x"3d",
           827 => x"84",
           828 => x"08",
           829 => x"82",
           830 => x"07",
           831 => x"72",
           832 => x"2e",
           833 => x"55",
           834 => x"74",
           835 => x"86",
           836 => x"d3",
           837 => x"51",
           838 => x"0c",
           839 => x"84",
           840 => x"bb",
           841 => x"d4",
           842 => x"77",
           843 => x"84",
           844 => x"85",
           845 => x"fd",
           846 => x"d3",
           847 => x"a6",
           848 => x"51",
           849 => x"54",
           850 => x"d2",
           851 => x"39",
           852 => x"b7",
           853 => x"53",
           854 => x"84",
           855 => x"2e",
           856 => x"77",
           857 => x"04",
           858 => x"55",
           859 => x"52",
           860 => x"08",
           861 => x"04",
           862 => x"8c",
           863 => x"15",
           864 => x"5e",
           865 => x"52",
           866 => x"83",
           867 => x"54",
           868 => x"2e",
           869 => x"a8",
           870 => x"81",
           871 => x"98",
           872 => x"e6",
           873 => x"9f",
           874 => x"d3",
           875 => x"75",
           876 => x"70",
           877 => x"27",
           878 => x"74",
           879 => x"06",
           880 => x"80",
           881 => x"81",
           882 => x"a0",
           883 => x"78",
           884 => x"51",
           885 => x"5c",
           886 => x"bb",
           887 => x"58",
           888 => x"76",
           889 => x"57",
           890 => x"0b",
           891 => x"04",
           892 => x"81",
           893 => x"a0",
           894 => x"fe",
           895 => x"b8",
           896 => x"e6",
           897 => x"df",
           898 => x"73",
           899 => x"72",
           900 => x"e1",
           901 => x"53",
           902 => x"74",
           903 => x"d3",
           904 => x"84",
           905 => x"ea",
           906 => x"38",
           907 => x"38",
           908 => x"db",
           909 => x"08",
           910 => x"78",
           911 => x"84",
           912 => x"e7",
           913 => x"80",
           914 => x"81",
           915 => x"2e",
           916 => x"d0",
           917 => x"90",
           918 => x"c5",
           919 => x"70",
           920 => x"72",
           921 => x"73",
           922 => x"57",
           923 => x"38",
           924 => x"84",
           925 => x"a0",
           926 => x"30",
           927 => x"51",
           928 => x"73",
           929 => x"80",
           930 => x"0d",
           931 => x"80",
           932 => x"9d",
           933 => x"9e",
           934 => x"81",
           935 => x"82",
           936 => x"06",
           937 => x"83",
           938 => x"81",
           939 => x"06",
           940 => x"85",
           941 => x"80",
           942 => x"06",
           943 => x"87",
           944 => x"a9",
           945 => x"72",
           946 => x"0d",
           947 => x"d4",
           948 => x"9c",
           949 => x"0d",
           950 => x"d4",
           951 => x"9b",
           952 => x"53",
           953 => x"81",
           954 => x"51",
           955 => x"3f",
           956 => x"52",
           957 => x"39",
           958 => x"a4",
           959 => x"b6",
           960 => x"51",
           961 => x"ff",
           962 => x"83",
           963 => x"51",
           964 => x"81",
           965 => x"c2",
           966 => x"fe",
           967 => x"3f",
           968 => x"2a",
           969 => x"2e",
           970 => x"51",
           971 => x"9a",
           972 => x"72",
           973 => x"71",
           974 => x"39",
           975 => x"f0",
           976 => x"ae",
           977 => x"51",
           978 => x"ff",
           979 => x"41",
           980 => x"42",
           981 => x"3f",
           982 => x"9b",
           983 => x"b5",
           984 => x"3f",
           985 => x"d6",
           986 => x"80",
           987 => x"0b",
           988 => x"06",
           989 => x"38",
           990 => x"81",
           991 => x"c1",
           992 => x"2e",
           993 => x"a0",
           994 => x"1a",
           995 => x"f6",
           996 => x"38",
           997 => x"70",
           998 => x"bb",
           999 => x"7a",
          1000 => x"3f",
          1001 => x"1b",
          1002 => x"38",
          1003 => x"5b",
          1004 => x"33",
          1005 => x"80",
          1006 => x"84",
          1007 => x"08",
          1008 => x"84",
          1009 => x"51",
          1010 => x"60",
          1011 => x"81",
          1012 => x"e7",
          1013 => x"26",
          1014 => x"5e",
          1015 => x"7a",
          1016 => x"2e",
          1017 => x"83",
          1018 => x"3f",
          1019 => x"57",
          1020 => x"80",
          1021 => x"51",
          1022 => x"84",
          1023 => x"72",
          1024 => x"80",
          1025 => x"5a",
          1026 => x"8d",
          1027 => x"5c",
          1028 => x"32",
          1029 => x"f2",
          1030 => x"7d",
          1031 => x"fc",
          1032 => x"f8",
          1033 => x"3f",
          1034 => x"81",
          1035 => x"38",
          1036 => x"de",
          1037 => x"bb",
          1038 => x"0b",
          1039 => x"94",
          1040 => x"f7",
          1041 => x"2e",
          1042 => x"df",
          1043 => x"33",
          1044 => x"82",
          1045 => x"91",
          1046 => x"d2",
          1047 => x"f8",
          1048 => x"80",
          1049 => x"d7",
          1050 => x"b3",
          1051 => x"85",
          1052 => x"fc",
          1053 => x"e4",
          1054 => x"83",
          1055 => x"3f",
          1056 => x"51",
          1057 => x"08",
          1058 => x"38",
          1059 => x"fb",
          1060 => x"cc",
          1061 => x"fe",
          1062 => x"55",
          1063 => x"d7",
          1064 => x"fd",
          1065 => x"fb",
          1066 => x"81",
          1067 => x"fa",
          1068 => x"e3",
          1069 => x"3f",
          1070 => x"51",
          1071 => x"cb",
          1072 => x"ff",
          1073 => x"bb",
          1074 => x"68",
          1075 => x"3f",
          1076 => x"08",
          1077 => x"84",
          1078 => x"d1",
          1079 => x"84",
          1080 => x"bf",
          1081 => x"f9",
          1082 => x"51",
          1083 => x"b8",
          1084 => x"05",
          1085 => x"08",
          1086 => x"fe",
          1087 => x"e9",
          1088 => x"d0",
          1089 => x"52",
          1090 => x"84",
          1091 => x"7e",
          1092 => x"33",
          1093 => x"78",
          1094 => x"05",
          1095 => x"fe",
          1096 => x"e8",
          1097 => x"2e",
          1098 => x"11",
          1099 => x"3f",
          1100 => x"64",
          1101 => x"d8",
          1102 => x"e4",
          1103 => x"cf",
          1104 => x"78",
          1105 => x"26",
          1106 => x"46",
          1107 => x"11",
          1108 => x"3f",
          1109 => x"9b",
          1110 => x"ff",
          1111 => x"bb",
          1112 => x"b8",
          1113 => x"05",
          1114 => x"08",
          1115 => x"d4",
          1116 => x"59",
          1117 => x"70",
          1118 => x"7d",
          1119 => x"78",
          1120 => x"51",
          1121 => x"81",
          1122 => x"b8",
          1123 => x"05",
          1124 => x"08",
          1125 => x"fe",
          1126 => x"e8",
          1127 => x"2e",
          1128 => x"11",
          1129 => x"3f",
          1130 => x"f3",
          1131 => x"3f",
          1132 => x"38",
          1133 => x"33",
          1134 => x"39",
          1135 => x"80",
          1136 => x"84",
          1137 => x"3d",
          1138 => x"51",
          1139 => x"b1",
          1140 => x"d9",
          1141 => x"e4",
          1142 => x"cc",
          1143 => x"78",
          1144 => x"26",
          1145 => x"d1",
          1146 => x"33",
          1147 => x"3d",
          1148 => x"51",
          1149 => x"80",
          1150 => x"80",
          1151 => x"05",
          1152 => x"ff",
          1153 => x"bb",
          1154 => x"39",
          1155 => x"80",
          1156 => x"84",
          1157 => x"3d",
          1158 => x"51",
          1159 => x"80",
          1160 => x"f8",
          1161 => x"b7",
          1162 => x"84",
          1163 => x"51",
          1164 => x"78",
          1165 => x"79",
          1166 => x"26",
          1167 => x"f4",
          1168 => x"51",
          1169 => x"b9",
          1170 => x"f3",
          1171 => x"52",
          1172 => x"84",
          1173 => x"bb",
          1174 => x"93",
          1175 => x"ff",
          1176 => x"bb",
          1177 => x"33",
          1178 => x"83",
          1179 => x"fc",
          1180 => x"9f",
          1181 => x"83",
          1182 => x"83",
          1183 => x"b8",
          1184 => x"05",
          1185 => x"08",
          1186 => x"5c",
          1187 => x"7a",
          1188 => x"9f",
          1189 => x"80",
          1190 => x"38",
          1191 => x"b4",
          1192 => x"66",
          1193 => x"d9",
          1194 => x"39",
          1195 => x"05",
          1196 => x"ff",
          1197 => x"bb",
          1198 => x"64",
          1199 => x"45",
          1200 => x"80",
          1201 => x"84",
          1202 => x"5e",
          1203 => x"82",
          1204 => x"fe",
          1205 => x"e1",
          1206 => x"2e",
          1207 => x"ce",
          1208 => x"23",
          1209 => x"53",
          1210 => x"84",
          1211 => x"eb",
          1212 => x"ff",
          1213 => x"bb",
          1214 => x"68",
          1215 => x"34",
          1216 => x"b8",
          1217 => x"05",
          1218 => x"08",
          1219 => x"71",
          1220 => x"59",
          1221 => x"81",
          1222 => x"d7",
          1223 => x"52",
          1224 => x"39",
          1225 => x"f3",
          1226 => x"9c",
          1227 => x"f0",
          1228 => x"9b",
          1229 => x"b8",
          1230 => x"22",
          1231 => x"45",
          1232 => x"5c",
          1233 => x"f3",
          1234 => x"f4",
          1235 => x"38",
          1236 => x"39",
          1237 => x"64",
          1238 => x"51",
          1239 => x"39",
          1240 => x"2e",
          1241 => x"fc",
          1242 => x"9c",
          1243 => x"33",
          1244 => x"f3",
          1245 => x"f4",
          1246 => x"38",
          1247 => x"39",
          1248 => x"2e",
          1249 => x"fb",
          1250 => x"7c",
          1251 => x"08",
          1252 => x"33",
          1253 => x"f3",
          1254 => x"f3",
          1255 => x"9c",
          1256 => x"47",
          1257 => x"0b",
          1258 => x"8c",
          1259 => x"52",
          1260 => x"84",
          1261 => x"87",
          1262 => x"3f",
          1263 => x"0c",
          1264 => x"57",
          1265 => x"96",
          1266 => x"77",
          1267 => x"75",
          1268 => x"84",
          1269 => x"0b",
          1270 => x"83",
          1271 => x"be",
          1272 => x"02",
          1273 => x"84",
          1274 => x"13",
          1275 => x"0c",
          1276 => x"95",
          1277 => x"3f",
          1278 => x"51",
          1279 => x"22",
          1280 => x"cc",
          1281 => x"33",
          1282 => x"3f",
          1283 => x"d0",
          1284 => x"51",
          1285 => x"83",
          1286 => x"e2",
          1287 => x"70",
          1288 => x"74",
          1289 => x"70",
          1290 => x"2e",
          1291 => x"70",
          1292 => x"55",
          1293 => x"ff",
          1294 => x"38",
          1295 => x"38",
          1296 => x"53",
          1297 => x"81",
          1298 => x"80",
          1299 => x"39",
          1300 => x"70",
          1301 => x"81",
          1302 => x"80",
          1303 => x"80",
          1304 => x"05",
          1305 => x"70",
          1306 => x"04",
          1307 => x"2e",
          1308 => x"72",
          1309 => x"54",
          1310 => x"e0",
          1311 => x"53",
          1312 => x"f8",
          1313 => x"53",
          1314 => x"bb",
          1315 => x"3d",
          1316 => x"3f",
          1317 => x"38",
          1318 => x"0d",
          1319 => x"33",
          1320 => x"8b",
          1321 => x"ff",
          1322 => x"81",
          1323 => x"52",
          1324 => x"13",
          1325 => x"80",
          1326 => x"52",
          1327 => x"13",
          1328 => x"26",
          1329 => x"87",
          1330 => x"38",
          1331 => x"72",
          1332 => x"13",
          1333 => x"13",
          1334 => x"13",
          1335 => x"13",
          1336 => x"13",
          1337 => x"87",
          1338 => x"98",
          1339 => x"9c",
          1340 => x"0c",
          1341 => x"7f",
          1342 => x"7d",
          1343 => x"7d",
          1344 => x"5c",
          1345 => x"b4",
          1346 => x"c0",
          1347 => x"34",
          1348 => x"85",
          1349 => x"5c",
          1350 => x"a4",
          1351 => x"c0",
          1352 => x"23",
          1353 => x"06",
          1354 => x"86",
          1355 => x"84",
          1356 => x"82",
          1357 => x"06",
          1358 => x"91",
          1359 => x"0d",
          1360 => x"2e",
          1361 => x"3f",
          1362 => x"98",
          1363 => x"81",
          1364 => x"38",
          1365 => x"0d",
          1366 => x"84",
          1367 => x"2c",
          1368 => x"06",
          1369 => x"3f",
          1370 => x"98",
          1371 => x"38",
          1372 => x"54",
          1373 => x"80",
          1374 => x"98",
          1375 => x"ff",
          1376 => x"14",
          1377 => x"71",
          1378 => x"04",
          1379 => x"83",
          1380 => x"53",
          1381 => x"38",
          1382 => x"2a",
          1383 => x"80",
          1384 => x"81",
          1385 => x"81",
          1386 => x"8a",
          1387 => x"71",
          1388 => x"87",
          1389 => x"86",
          1390 => x"72",
          1391 => x"3d",
          1392 => x"06",
          1393 => x"32",
          1394 => x"38",
          1395 => x"80",
          1396 => x"08",
          1397 => x"54",
          1398 => x"3d",
          1399 => x"70",
          1400 => x"f3",
          1401 => x"3d",
          1402 => x"56",
          1403 => x"38",
          1404 => x"81",
          1405 => x"2e",
          1406 => x"08",
          1407 => x"54",
          1408 => x"91",
          1409 => x"e3",
          1410 => x"72",
          1411 => x"81",
          1412 => x"ff",
          1413 => x"70",
          1414 => x"90",
          1415 => x"33",
          1416 => x"84",
          1417 => x"71",
          1418 => x"70",
          1419 => x"53",
          1420 => x"2a",
          1421 => x"b5",
          1422 => x"96",
          1423 => x"70",
          1424 => x"87",
          1425 => x"8a",
          1426 => x"ab",
          1427 => x"f3",
          1428 => x"83",
          1429 => x"08",
          1430 => x"98",
          1431 => x"9e",
          1432 => x"c0",
          1433 => x"87",
          1434 => x"0c",
          1435 => x"dc",
          1436 => x"f3",
          1437 => x"83",
          1438 => x"08",
          1439 => x"c0",
          1440 => x"9e",
          1441 => x"c0",
          1442 => x"f4",
          1443 => x"f3",
          1444 => x"83",
          1445 => x"08",
          1446 => x"f4",
          1447 => x"90",
          1448 => x"52",
          1449 => x"f4",
          1450 => x"90",
          1451 => x"52",
          1452 => x"52",
          1453 => x"87",
          1454 => x"0a",
          1455 => x"83",
          1456 => x"34",
          1457 => x"70",
          1458 => x"70",
          1459 => x"83",
          1460 => x"9e",
          1461 => x"51",
          1462 => x"81",
          1463 => x"0b",
          1464 => x"80",
          1465 => x"2e",
          1466 => x"8a",
          1467 => x"08",
          1468 => x"52",
          1469 => x"71",
          1470 => x"c0",
          1471 => x"06",
          1472 => x"38",
          1473 => x"80",
          1474 => x"81",
          1475 => x"80",
          1476 => x"f4",
          1477 => x"90",
          1478 => x"52",
          1479 => x"52",
          1480 => x"87",
          1481 => x"06",
          1482 => x"38",
          1483 => x"87",
          1484 => x"70",
          1485 => x"90",
          1486 => x"08",
          1487 => x"70",
          1488 => x"83",
          1489 => x"08",
          1490 => x"51",
          1491 => x"87",
          1492 => x"51",
          1493 => x"81",
          1494 => x"c0",
          1495 => x"83",
          1496 => x"81",
          1497 => x"83",
          1498 => x"83",
          1499 => x"38",
          1500 => x"83",
          1501 => x"38",
          1502 => x"c7",
          1503 => x"85",
          1504 => x"74",
          1505 => x"54",
          1506 => x"33",
          1507 => x"93",
          1508 => x"f4",
          1509 => x"83",
          1510 => x"38",
          1511 => x"a7",
          1512 => x"83",
          1513 => x"75",
          1514 => x"54",
          1515 => x"51",
          1516 => x"52",
          1517 => x"3f",
          1518 => x"f4",
          1519 => x"f0",
          1520 => x"b5",
          1521 => x"e4",
          1522 => x"db",
          1523 => x"f3",
          1524 => x"75",
          1525 => x"08",
          1526 => x"54",
          1527 => x"db",
          1528 => x"f4",
          1529 => x"f4",
          1530 => x"3d",
          1531 => x"bd",
          1532 => x"3f",
          1533 => x"29",
          1534 => x"84",
          1535 => x"b4",
          1536 => x"f3",
          1537 => x"75",
          1538 => x"08",
          1539 => x"54",
          1540 => x"dc",
          1541 => x"f4",
          1542 => x"9e",
          1543 => x"51",
          1544 => x"c0",
          1545 => x"83",
          1546 => x"83",
          1547 => x"51",
          1548 => x"08",
          1549 => x"99",
          1550 => x"fc",
          1551 => x"db",
          1552 => x"f3",
          1553 => x"75",
          1554 => x"08",
          1555 => x"54",
          1556 => x"db",
          1557 => x"f4",
          1558 => x"96",
          1559 => x"51",
          1560 => x"33",
          1561 => x"fe",
          1562 => x"bf",
          1563 => x"75",
          1564 => x"83",
          1565 => x"83",
          1566 => x"fc",
          1567 => x"51",
          1568 => x"33",
          1569 => x"d7",
          1570 => x"dd",
          1571 => x"f4",
          1572 => x"90",
          1573 => x"52",
          1574 => x"3f",
          1575 => x"2e",
          1576 => x"90",
          1577 => x"b1",
          1578 => x"73",
          1579 => x"83",
          1580 => x"11",
          1581 => x"b1",
          1582 => x"75",
          1583 => x"83",
          1584 => x"11",
          1585 => x"b0",
          1586 => x"73",
          1587 => x"83",
          1588 => x"11",
          1589 => x"b0",
          1590 => x"74",
          1591 => x"83",
          1592 => x"11",
          1593 => x"b0",
          1594 => x"75",
          1595 => x"83",
          1596 => x"11",
          1597 => x"b0",
          1598 => x"73",
          1599 => x"83",
          1600 => x"83",
          1601 => x"83",
          1602 => x"f9",
          1603 => x"02",
          1604 => x"8c",
          1605 => x"05",
          1606 => x"51",
          1607 => x"04",
          1608 => x"3f",
          1609 => x"51",
          1610 => x"04",
          1611 => x"3f",
          1612 => x"51",
          1613 => x"04",
          1614 => x"3f",
          1615 => x"0c",
          1616 => x"0c",
          1617 => x"96",
          1618 => x"3d",
          1619 => x"70",
          1620 => x"08",
          1621 => x"84",
          1622 => x"ff",
          1623 => x"80",
          1624 => x"3f",
          1625 => x"38",
          1626 => x"84",
          1627 => x"84",
          1628 => x"bb",
          1629 => x"55",
          1630 => x"70",
          1631 => x"78",
          1632 => x"38",
          1633 => x"53",
          1634 => x"84",
          1635 => x"38",
          1636 => x"0d",
          1637 => x"d9",
          1638 => x"e8",
          1639 => x"3f",
          1640 => x"3d",
          1641 => x"34",
          1642 => x"ad",
          1643 => x"0c",
          1644 => x"ab",
          1645 => x"5d",
          1646 => x"a0",
          1647 => x"3d",
          1648 => x"f4",
          1649 => x"bf",
          1650 => x"79",
          1651 => x"3f",
          1652 => x"14",
          1653 => x"38",
          1654 => x"70",
          1655 => x"27",
          1656 => x"84",
          1657 => x"5a",
          1658 => x"80",
          1659 => x"84",
          1660 => x"53",
          1661 => x"84",
          1662 => x"73",
          1663 => x"81",
          1664 => x"fe",
          1665 => x"77",
          1666 => x"38",
          1667 => x"55",
          1668 => x"d4",
          1669 => x"0b",
          1670 => x"73",
          1671 => x"ec",
          1672 => x"84",
          1673 => x"f4",
          1674 => x"51",
          1675 => x"08",
          1676 => x"bd",
          1677 => x"80",
          1678 => x"38",
          1679 => x"19",
          1680 => x"75",
          1681 => x"56",
          1682 => x"09",
          1683 => x"84",
          1684 => x"cd",
          1685 => x"08",
          1686 => x"3d",
          1687 => x"0b",
          1688 => x"5d",
          1689 => x"ec",
          1690 => x"81",
          1691 => x"82",
          1692 => x"38",
          1693 => x"90",
          1694 => x"38",
          1695 => x"51",
          1696 => x"98",
          1697 => x"ff",
          1698 => x"06",
          1699 => x"70",
          1700 => x"98",
          1701 => x"05",
          1702 => x"70",
          1703 => x"5d",
          1704 => x"57",
          1705 => x"75",
          1706 => x"0a",
          1707 => x"2c",
          1708 => x"38",
          1709 => x"57",
          1710 => x"43",
          1711 => x"df",
          1712 => x"42",
          1713 => x"80",
          1714 => x"34",
          1715 => x"38",
          1716 => x"2c",
          1717 => x"70",
          1718 => x"82",
          1719 => x"53",
          1720 => x"78",
          1721 => x"c0",
          1722 => x"bb",
          1723 => x"5b",
          1724 => x"fe",
          1725 => x"38",
          1726 => x"76",
          1727 => x"29",
          1728 => x"70",
          1729 => x"95",
          1730 => x"70",
          1731 => x"df",
          1732 => x"25",
          1733 => x"18",
          1734 => x"ff",
          1735 => x"38",
          1736 => x"2e",
          1737 => x"57",
          1738 => x"c8",
          1739 => x"84",
          1740 => x"60",
          1741 => x"8e",
          1742 => x"05",
          1743 => x"15",
          1744 => x"c0",
          1745 => x"d9",
          1746 => x"80",
          1747 => x"08",
          1748 => x"84",
          1749 => x"84",
          1750 => x"e2",
          1751 => x"e2",
          1752 => x"27",
          1753 => x"52",
          1754 => x"34",
          1755 => x"b5",
          1756 => x"2e",
          1757 => x"38",
          1758 => x"70",
          1759 => x"80",
          1760 => x"34",
          1761 => x"33",
          1762 => x"84",
          1763 => x"b4",
          1764 => x"a0",
          1765 => x"e8",
          1766 => x"3f",
          1767 => x"78",
          1768 => x"06",
          1769 => x"a5",
          1770 => x"fb",
          1771 => x"e8",
          1772 => x"1d",
          1773 => x"92",
          1774 => x"f4",
          1775 => x"8d",
          1776 => x"38",
          1777 => x"70",
          1778 => x"e6",
          1779 => x"84",
          1780 => x"84",
          1781 => x"05",
          1782 => x"b3",
          1783 => x"c8",
          1784 => x"84",
          1785 => x"51",
          1786 => x"08",
          1787 => x"84",
          1788 => x"b3",
          1789 => x"05",
          1790 => x"81",
          1791 => x"c8",
          1792 => x"c4",
          1793 => x"f9",
          1794 => x"81",
          1795 => x"7b",
          1796 => x"c7",
          1797 => x"ff",
          1798 => x"55",
          1799 => x"e6",
          1800 => x"84",
          1801 => x"52",
          1802 => x"c8",
          1803 => x"c4",
          1804 => x"ff",
          1805 => x"c8",
          1806 => x"74",
          1807 => x"5b",
          1808 => x"2b",
          1809 => x"44",
          1810 => x"38",
          1811 => x"ff",
          1812 => x"70",
          1813 => x"c4",
          1814 => x"24",
          1815 => x"52",
          1816 => x"81",
          1817 => x"70",
          1818 => x"56",
          1819 => x"84",
          1820 => x"b1",
          1821 => x"81",
          1822 => x"e2",
          1823 => x"25",
          1824 => x"16",
          1825 => x"e6",
          1826 => x"b0",
          1827 => x"81",
          1828 => x"e2",
          1829 => x"25",
          1830 => x"18",
          1831 => x"52",
          1832 => x"75",
          1833 => x"05",
          1834 => x"5c",
          1835 => x"38",
          1836 => x"55",
          1837 => x"e6",
          1838 => x"f7",
          1839 => x"57",
          1840 => x"ff",
          1841 => x"33",
          1842 => x"e6",
          1843 => x"cf",
          1844 => x"f3",
          1845 => x"ff",
          1846 => x"e2",
          1847 => x"f0",
          1848 => x"10",
          1849 => x"41",
          1850 => x"2b",
          1851 => x"81",
          1852 => x"e2",
          1853 => x"83",
          1854 => x"f4",
          1855 => x"e3",
          1856 => x"83",
          1857 => x"f4",
          1858 => x"74",
          1859 => x"56",
          1860 => x"f0",
          1861 => x"38",
          1862 => x"0b",
          1863 => x"84",
          1864 => x"c8",
          1865 => x"84",
          1866 => x"ae",
          1867 => x"a0",
          1868 => x"e8",
          1869 => x"3f",
          1870 => x"61",
          1871 => x"06",
          1872 => x"51",
          1873 => x"e2",
          1874 => x"34",
          1875 => x"70",
          1876 => x"2e",
          1877 => x"ff",
          1878 => x"ff",
          1879 => x"84",
          1880 => x"ad",
          1881 => x"98",
          1882 => x"33",
          1883 => x"80",
          1884 => x"a0",
          1885 => x"c8",
          1886 => x"84",
          1887 => x"74",
          1888 => x"e8",
          1889 => x"3f",
          1890 => x"0a",
          1891 => x"33",
          1892 => x"d6",
          1893 => x"51",
          1894 => x"0a",
          1895 => x"2c",
          1896 => x"79",
          1897 => x"39",
          1898 => x"34",
          1899 => x"51",
          1900 => x"0a",
          1901 => x"2c",
          1902 => x"75",
          1903 => x"57",
          1904 => x"e8",
          1905 => x"df",
          1906 => x"80",
          1907 => x"c4",
          1908 => x"ff",
          1909 => x"34",
          1910 => x"c8",
          1911 => x"84",
          1912 => x"ab",
          1913 => x"a0",
          1914 => x"e8",
          1915 => x"3f",
          1916 => x"7c",
          1917 => x"06",
          1918 => x"51",
          1919 => x"e2",
          1920 => x"34",
          1921 => x"0d",
          1922 => x"ff",
          1923 => x"de",
          1924 => x"75",
          1925 => x"98",
          1926 => x"38",
          1927 => x"34",
          1928 => x"0a",
          1929 => x"33",
          1930 => x"38",
          1931 => x"34",
          1932 => x"b4",
          1933 => x"33",
          1934 => x"17",
          1935 => x"57",
          1936 => x"0a",
          1937 => x"2c",
          1938 => x"58",
          1939 => x"98",
          1940 => x"06",
          1941 => x"ce",
          1942 => x"51",
          1943 => x"0a",
          1944 => x"2c",
          1945 => x"75",
          1946 => x"e8",
          1947 => x"3f",
          1948 => x"0a",
          1949 => x"33",
          1950 => x"b9",
          1951 => x"80",
          1952 => x"83",
          1953 => x"52",
          1954 => x"3f",
          1955 => x"a6",
          1956 => x"ef",
          1957 => x"e8",
          1958 => x"58",
          1959 => x"0a",
          1960 => x"2c",
          1961 => x"76",
          1962 => x"33",
          1963 => x"81",
          1964 => x"79",
          1965 => x"83",
          1966 => x"38",
          1967 => x"08",
          1968 => x"18",
          1969 => x"80",
          1970 => x"ec",
          1971 => x"38",
          1972 => x"f4",
          1973 => x"80",
          1974 => x"b5",
          1975 => x"51",
          1976 => x"ff",
          1977 => x"25",
          1978 => x"51",
          1979 => x"08",
          1980 => x"08",
          1981 => x"52",
          1982 => x"0b",
          1983 => x"33",
          1984 => x"c4",
          1985 => x"51",
          1986 => x"08",
          1987 => x"84",
          1988 => x"a6",
          1989 => x"05",
          1990 => x"81",
          1991 => x"ff",
          1992 => x"84",
          1993 => x"81",
          1994 => x"7b",
          1995 => x"e2",
          1996 => x"57",
          1997 => x"84",
          1998 => x"a5",
          1999 => x"a0",
          2000 => x"e8",
          2001 => x"3f",
          2002 => x"76",
          2003 => x"06",
          2004 => x"81",
          2005 => x"c4",
          2006 => x"06",
          2007 => x"ff",
          2008 => x"ff",
          2009 => x"c8",
          2010 => x"2e",
          2011 => x"52",
          2012 => x"e6",
          2013 => x"ff",
          2014 => x"51",
          2015 => x"33",
          2016 => x"34",
          2017 => x"80",
          2018 => x"34",
          2019 => x"84",
          2020 => x"83",
          2021 => x"ef",
          2022 => x"3f",
          2023 => x"34",
          2024 => x"81",
          2025 => x"a8",
          2026 => x"e2",
          2027 => x"ef",
          2028 => x"88",
          2029 => x"e8",
          2030 => x"3f",
          2031 => x"ff",
          2032 => x"ff",
          2033 => x"78",
          2034 => x"51",
          2035 => x"33",
          2036 => x"f4",
          2037 => x"5a",
          2038 => x"84",
          2039 => x"70",
          2040 => x"08",
          2041 => x"ff",
          2042 => x"70",
          2043 => x"08",
          2044 => x"b3",
          2045 => x"ff",
          2046 => x"81",
          2047 => x"93",
          2048 => x"f4",
          2049 => x"fe",
          2050 => x"75",
          2051 => x"ec",
          2052 => x"3f",
          2053 => x"89",
          2054 => x"80",
          2055 => x"bb",
          2056 => x"53",
          2057 => x"3f",
          2058 => x"84",
          2059 => x"83",
          2060 => x"7a",
          2061 => x"84",
          2062 => x"2e",
          2063 => x"bb",
          2064 => x"84",
          2065 => x"bb",
          2066 => x"bb",
          2067 => x"57",
          2068 => x"83",
          2069 => x"f4",
          2070 => x"59",
          2071 => x"87",
          2072 => x"1a",
          2073 => x"3f",
          2074 => x"f4",
          2075 => x"9c",
          2076 => x"94",
          2077 => x"f4",
          2078 => x"9c",
          2079 => x"a0",
          2080 => x"5e",
          2081 => x"5d",
          2082 => x"c7",
          2083 => x"39",
          2084 => x"a4",
          2085 => x"05",
          2086 => x"7a",
          2087 => x"f4",
          2088 => x"80",
          2089 => x"70",
          2090 => x"9c",
          2091 => x"56",
          2092 => x"08",
          2093 => x"10",
          2094 => x"54",
          2095 => x"91",
          2096 => x"10",
          2097 => x"57",
          2098 => x"38",
          2099 => x"34",
          2100 => x"34",
          2101 => x"ff",
          2102 => x"f7",
          2103 => x"c3",
          2104 => x"05",
          2105 => x"8d",
          2106 => x"81",
          2107 => x"2e",
          2108 => x"59",
          2109 => x"80",
          2110 => x"90",
          2111 => x"83",
          2112 => x"23",
          2113 => x"71",
          2114 => x"71",
          2115 => x"78",
          2116 => x"84",
          2117 => x"05",
          2118 => x"75",
          2119 => x"33",
          2120 => x"55",
          2121 => x"34",
          2122 => x"ff",
          2123 => x"0d",
          2124 => x"fa",
          2125 => x"fa",
          2126 => x"05",
          2127 => x"b0",
          2128 => x"81",
          2129 => x"81",
          2130 => x"83",
          2131 => x"59",
          2132 => x"73",
          2133 => x"29",
          2134 => x"ff",
          2135 => x"ff",
          2136 => x"75",
          2137 => x"5c",
          2138 => x"b4",
          2139 => x"29",
          2140 => x"7b",
          2141 => x"55",
          2142 => x"80",
          2143 => x"fa",
          2144 => x"34",
          2145 => x"86",
          2146 => x"33",
          2147 => x"33",
          2148 => x"22",
          2149 => x"5e",
          2150 => x"df",
          2151 => x"ff",
          2152 => x"54",
          2153 => x"0b",
          2154 => x"fa",
          2155 => x"98",
          2156 => x"2b",
          2157 => x"56",
          2158 => x"fd",
          2159 => x"fa",
          2160 => x"10",
          2161 => x"90",
          2162 => x"5e",
          2163 => x"b0",
          2164 => x"70",
          2165 => x"70",
          2166 => x"70",
          2167 => x"60",
          2168 => x"40",
          2169 => x"72",
          2170 => x"57",
          2171 => x"ff",
          2172 => x"ff",
          2173 => x"29",
          2174 => x"78",
          2175 => x"79",
          2176 => x"58",
          2177 => x"5c",
          2178 => x"74",
          2179 => x"39",
          2180 => x"53",
          2181 => x"85",
          2182 => x"80",
          2183 => x"b0",
          2184 => x"80",
          2185 => x"80",
          2186 => x"34",
          2187 => x"51",
          2188 => x"70",
          2189 => x"c0",
          2190 => x"54",
          2191 => x"80",
          2192 => x"72",
          2193 => x"70",
          2194 => x"86",
          2195 => x"f7",
          2196 => x"80",
          2197 => x"0b",
          2198 => x"04",
          2199 => x"0c",
          2200 => x"33",
          2201 => x"b8",
          2202 => x"75",
          2203 => x"f8",
          2204 => x"b4",
          2205 => x"a0",
          2206 => x"51",
          2207 => x"83",
          2208 => x"53",
          2209 => x"c4",
          2210 => x"55",
          2211 => x"b4",
          2212 => x"7a",
          2213 => x"7a",
          2214 => x"72",
          2215 => x"22",
          2216 => x"f6",
          2217 => x"82",
          2218 => x"71",
          2219 => x"9f",
          2220 => x"14",
          2221 => x"e0",
          2222 => x"33",
          2223 => x"14",
          2224 => x"38",
          2225 => x"fa",
          2226 => x"55",
          2227 => x"73",
          2228 => x"54",
          2229 => x"b8",
          2230 => x"fa",
          2231 => x"06",
          2232 => x"73",
          2233 => x"31",
          2234 => x"71",
          2235 => x"c7",
          2236 => x"79",
          2237 => x"71",
          2238 => x"75",
          2239 => x"16",
          2240 => x"b9",
          2241 => x"5a",
          2242 => x"77",
          2243 => x"84",
          2244 => x"71",
          2245 => x"72",
          2246 => x"84",
          2247 => x"74",
          2248 => x"22",
          2249 => x"f6",
          2250 => x"fd",
          2251 => x"38",
          2252 => x"fa",
          2253 => x"09",
          2254 => x"31",
          2255 => x"71",
          2256 => x"59",
          2257 => x"83",
          2258 => x"74",
          2259 => x"e0",
          2260 => x"05",
          2261 => x"2e",
          2262 => x"16",
          2263 => x"34",
          2264 => x"f4",
          2265 => x"55",
          2266 => x"15",
          2267 => x"74",
          2268 => x"a9",
          2269 => x"05",
          2270 => x"26",
          2271 => x"fc",
          2272 => x"f8",
          2273 => x"71",
          2274 => x"bb",
          2275 => x"0b",
          2276 => x"33",
          2277 => x"80",
          2278 => x"83",
          2279 => x"84",
          2280 => x"b4",
          2281 => x"9f",
          2282 => x"70",
          2283 => x"fa",
          2284 => x"33",
          2285 => x"25",
          2286 => x"b4",
          2287 => x"86",
          2288 => x"70",
          2289 => x"72",
          2290 => x"fa",
          2291 => x"0c",
          2292 => x"33",
          2293 => x"11",
          2294 => x"38",
          2295 => x"80",
          2296 => x"0d",
          2297 => x"83",
          2298 => x"ff",
          2299 => x"b4",
          2300 => x"b4",
          2301 => x"02",
          2302 => x"b3",
          2303 => x"05",
          2304 => x"33",
          2305 => x"80",
          2306 => x"51",
          2307 => x"09",
          2308 => x"83",
          2309 => x"84",
          2310 => x"b0",
          2311 => x"70",
          2312 => x"bb",
          2313 => x"fa",
          2314 => x"83",
          2315 => x"b0",
          2316 => x"70",
          2317 => x"f1",
          2318 => x"84",
          2319 => x"83",
          2320 => x"07",
          2321 => x"b4",
          2322 => x"51",
          2323 => x"39",
          2324 => x"85",
          2325 => x"ff",
          2326 => x"fb",
          2327 => x"b0",
          2328 => x"33",
          2329 => x"83",
          2330 => x"fa",
          2331 => x"83",
          2332 => x"fa",
          2333 => x"07",
          2334 => x"cc",
          2335 => x"06",
          2336 => x"34",
          2337 => x"81",
          2338 => x"83",
          2339 => x"fa",
          2340 => x"07",
          2341 => x"94",
          2342 => x"06",
          2343 => x"34",
          2344 => x"81",
          2345 => x"34",
          2346 => x"81",
          2347 => x"fa",
          2348 => x"0d",
          2349 => x"80",
          2350 => x"83",
          2351 => x"84",
          2352 => x"5b",
          2353 => x"78",
          2354 => x"81",
          2355 => x"80",
          2356 => x"fa",
          2357 => x"7c",
          2358 => x"04",
          2359 => x"38",
          2360 => x"0b",
          2361 => x"fa",
          2362 => x"34",
          2363 => x"58",
          2364 => x"f7",
          2365 => x"7b",
          2366 => x"f8",
          2367 => x"b8",
          2368 => x"34",
          2369 => x"fa",
          2370 => x"8f",
          2371 => x"fa",
          2372 => x"80",
          2373 => x"83",
          2374 => x"b2",
          2375 => x"ba",
          2376 => x"56",
          2377 => x"52",
          2378 => x"3f",
          2379 => x"5a",
          2380 => x"84",
          2381 => x"83",
          2382 => x"81",
          2383 => x"85",
          2384 => x"dd",
          2385 => x"f9",
          2386 => x"0b",
          2387 => x"b4",
          2388 => x"83",
          2389 => x"80",
          2390 => x"84",
          2391 => x"b4",
          2392 => x"81",
          2393 => x"e8",
          2394 => x"84",
          2395 => x"fe",
          2396 => x"51",
          2397 => x"84",
          2398 => x"e8",
          2399 => x"fe",
          2400 => x"ff",
          2401 => x"0d",
          2402 => x"84",
          2403 => x"83",
          2404 => x"86",
          2405 => x"22",
          2406 => x"05",
          2407 => x"8a",
          2408 => x"72",
          2409 => x"2e",
          2410 => x"b9",
          2411 => x"75",
          2412 => x"f8",
          2413 => x"b5",
          2414 => x"54",
          2415 => x"a0",
          2416 => x"83",
          2417 => x"72",
          2418 => x"75",
          2419 => x"b4",
          2420 => x"83",
          2421 => x"18",
          2422 => x"ff",
          2423 => x"b5",
          2424 => x"57",
          2425 => x"99",
          2426 => x"ff",
          2427 => x"99",
          2428 => x"81",
          2429 => x"fa",
          2430 => x"72",
          2431 => x"33",
          2432 => x"80",
          2433 => x"0d",
          2434 => x"8d",
          2435 => x"09",
          2436 => x"81",
          2437 => x"fa",
          2438 => x"b6",
          2439 => x"33",
          2440 => x"06",
          2441 => x"a0",
          2442 => x"81",
          2443 => x"ff",
          2444 => x"a5",
          2445 => x"54",
          2446 => x"fa",
          2447 => x"f2",
          2448 => x"3f",
          2449 => x"3d",
          2450 => x"81",
          2451 => x"33",
          2452 => x"53",
          2453 => x"fa",
          2454 => x"d5",
          2455 => x"ff",
          2456 => x"a5",
          2457 => x"34",
          2458 => x"b5",
          2459 => x"3f",
          2460 => x"ef",
          2461 => x"0d",
          2462 => x"80",
          2463 => x"b8",
          2464 => x"78",
          2465 => x"24",
          2466 => x"b9",
          2467 => x"84",
          2468 => x"83",
          2469 => x"58",
          2470 => x"86",
          2471 => x"f8",
          2472 => x"b2",
          2473 => x"42",
          2474 => x"83",
          2475 => x"05",
          2476 => x"86",
          2477 => x"f8",
          2478 => x"b2",
          2479 => x"29",
          2480 => x"fa",
          2481 => x"81",
          2482 => x"76",
          2483 => x"f9",
          2484 => x"19",
          2485 => x"0b",
          2486 => x"04",
          2487 => x"79",
          2488 => x"9b",
          2489 => x"cc",
          2490 => x"84",
          2491 => x"83",
          2492 => x"5e",
          2493 => x"86",
          2494 => x"f8",
          2495 => x"b2",
          2496 => x"59",
          2497 => x"83",
          2498 => x"5b",
          2499 => x"b0",
          2500 => x"70",
          2501 => x"83",
          2502 => x"44",
          2503 => x"33",
          2504 => x"1f",
          2505 => x"77",
          2506 => x"b5",
          2507 => x"9c",
          2508 => x"b7",
          2509 => x"78",
          2510 => x"38",
          2511 => x"0b",
          2512 => x"04",
          2513 => x"19",
          2514 => x"84",
          2515 => x"77",
          2516 => x"88",
          2517 => x"80",
          2518 => x"0b",
          2519 => x"04",
          2520 => x"0b",
          2521 => x"33",
          2522 => x"33",
          2523 => x"84",
          2524 => x"80",
          2525 => x"fa",
          2526 => x"71",
          2527 => x"83",
          2528 => x"33",
          2529 => x"fa",
          2530 => x"34",
          2531 => x"06",
          2532 => x"33",
          2533 => x"58",
          2534 => x"99",
          2535 => x"89",
          2536 => x"3f",
          2537 => x"ae",
          2538 => x"b5",
          2539 => x"b4",
          2540 => x"a0",
          2541 => x"51",
          2542 => x"ff",
          2543 => x"51",
          2544 => x"a4",
          2545 => x"57",
          2546 => x"75",
          2547 => x"80",
          2548 => x"84",
          2549 => x"86",
          2550 => x"81",
          2551 => x"84",
          2552 => x"83",
          2553 => x"83",
          2554 => x"83",
          2555 => x"80",
          2556 => x"84",
          2557 => x"78",
          2558 => x"a7",
          2559 => x"f8",
          2560 => x"b5",
          2561 => x"29",
          2562 => x"fa",
          2563 => x"05",
          2564 => x"8a",
          2565 => x"5c",
          2566 => x"81",
          2567 => x"83",
          2568 => x"34",
          2569 => x"06",
          2570 => x"05",
          2571 => x"86",
          2572 => x"f8",
          2573 => x"b2",
          2574 => x"42",
          2575 => x"34",
          2576 => x"62",
          2577 => x"86",
          2578 => x"f8",
          2579 => x"b2",
          2580 => x"29",
          2581 => x"fa",
          2582 => x"34",
          2583 => x"58",
          2584 => x"b8",
          2585 => x"ff",
          2586 => x"83",
          2587 => x"58",
          2588 => x"bb",
          2589 => x"83",
          2590 => x"38",
          2591 => x"f9",
          2592 => x"26",
          2593 => x"c6",
          2594 => x"0b",
          2595 => x"51",
          2596 => x"84",
          2597 => x"b4",
          2598 => x"ff",
          2599 => x"ff",
          2600 => x"a0",
          2601 => x"41",
          2602 => x"ff",
          2603 => x"45",
          2604 => x"82",
          2605 => x"06",
          2606 => x"06",
          2607 => x"84",
          2608 => x"1b",
          2609 => x"b5",
          2610 => x"29",
          2611 => x"83",
          2612 => x"33",
          2613 => x"fa",
          2614 => x"34",
          2615 => x"06",
          2616 => x"33",
          2617 => x"40",
          2618 => x"d6",
          2619 => x"ff",
          2620 => x"ac",
          2621 => x"92",
          2622 => x"fa",
          2623 => x"06",
          2624 => x"38",
          2625 => x"33",
          2626 => x"06",
          2627 => x"06",
          2628 => x"5b",
          2629 => x"c7",
          2630 => x"33",
          2631 => x"22",
          2632 => x"56",
          2633 => x"83",
          2634 => x"5a",
          2635 => x"b0",
          2636 => x"70",
          2637 => x"83",
          2638 => x"5b",
          2639 => x"33",
          2640 => x"05",
          2641 => x"7f",
          2642 => x"b5",
          2643 => x"ba",
          2644 => x"0c",
          2645 => x"17",
          2646 => x"7a",
          2647 => x"ff",
          2648 => x"39",
          2649 => x"0b",
          2650 => x"04",
          2651 => x"b9",
          2652 => x"b4",
          2653 => x"b5",
          2654 => x"f4",
          2655 => x"dc",
          2656 => x"ff",
          2657 => x"fb",
          2658 => x"11",
          2659 => x"79",
          2660 => x"ca",
          2661 => x"23",
          2662 => x"33",
          2663 => x"34",
          2664 => x"33",
          2665 => x"f9",
          2666 => x"fa",
          2667 => x"72",
          2668 => x"80",
          2669 => x"05",
          2670 => x"b5",
          2671 => x"29",
          2672 => x"fa",
          2673 => x"76",
          2674 => x"b0",
          2675 => x"34",
          2676 => x"06",
          2677 => x"33",
          2678 => x"42",
          2679 => x"d6",
          2680 => x"06",
          2681 => x"38",
          2682 => x"e2",
          2683 => x"b5",
          2684 => x"84",
          2685 => x"f3",
          2686 => x"75",
          2687 => x"ea",
          2688 => x"0c",
          2689 => x"33",
          2690 => x"33",
          2691 => x"33",
          2692 => x"b9",
          2693 => x"ec",
          2694 => x"ed",
          2695 => x"ee",
          2696 => x"33",
          2697 => x"84",
          2698 => x"09",
          2699 => x"b5",
          2700 => x"33",
          2701 => x"c0",
          2702 => x"ec",
          2703 => x"3f",
          2704 => x"83",
          2705 => x"60",
          2706 => x"83",
          2707 => x"fe",
          2708 => x"33",
          2709 => x"77",
          2710 => x"84",
          2711 => x"41",
          2712 => x"10",
          2713 => x"08",
          2714 => x"80",
          2715 => x"33",
          2716 => x"70",
          2717 => x"42",
          2718 => x"34",
          2719 => x"56",
          2720 => x"ba",
          2721 => x"06",
          2722 => x"75",
          2723 => x"fa",
          2724 => x"83",
          2725 => x"70",
          2726 => x"2e",
          2727 => x"83",
          2728 => x"0b",
          2729 => x"33",
          2730 => x"57",
          2731 => x"17",
          2732 => x"f9",
          2733 => x"80",
          2734 => x"33",
          2735 => x"70",
          2736 => x"41",
          2737 => x"34",
          2738 => x"5b",
          2739 => x"ba",
          2740 => x"81",
          2741 => x"33",
          2742 => x"33",
          2743 => x"80",
          2744 => x"5a",
          2745 => x"ff",
          2746 => x"ff",
          2747 => x"7e",
          2748 => x"80",
          2749 => x"39",
          2750 => x"2e",
          2751 => x"58",
          2752 => x"d9",
          2753 => x"fb",
          2754 => x"75",
          2755 => x"d9",
          2756 => x"05",
          2757 => x"5e",
          2758 => x"57",
          2759 => x"39",
          2760 => x"2e",
          2761 => x"83",
          2762 => x"b8",
          2763 => x"75",
          2764 => x"83",
          2765 => x"e5",
          2766 => x"0b",
          2767 => x"76",
          2768 => x"ba",
          2769 => x"e5",
          2770 => x"17",
          2771 => x"33",
          2772 => x"84",
          2773 => x"2e",
          2774 => x"75",
          2775 => x"52",
          2776 => x"3f",
          2777 => x"57",
          2778 => x"ba",
          2779 => x"06",
          2780 => x"81",
          2781 => x"81",
          2782 => x"5b",
          2783 => x"38",
          2784 => x"76",
          2785 => x"77",
          2786 => x"83",
          2787 => x"ff",
          2788 => x"b4",
          2789 => x"34",
          2790 => x"5f",
          2791 => x"ba",
          2792 => x"5b",
          2793 => x"fa",
          2794 => x"81",
          2795 => x"74",
          2796 => x"83",
          2797 => x"29",
          2798 => x"f9",
          2799 => x"5d",
          2800 => x"83",
          2801 => x"57",
          2802 => x"b8",
          2803 => x"d6",
          2804 => x"b2",
          2805 => x"31",
          2806 => x"38",
          2807 => x"27",
          2808 => x"83",
          2809 => x"83",
          2810 => x"76",
          2811 => x"81",
          2812 => x"29",
          2813 => x"a0",
          2814 => x"81",
          2815 => x"71",
          2816 => x"7f",
          2817 => x"1a",
          2818 => x"b9",
          2819 => x"5d",
          2820 => x"7c",
          2821 => x"84",
          2822 => x"71",
          2823 => x"77",
          2824 => x"17",
          2825 => x"7b",
          2826 => x"81",
          2827 => x"5e",
          2828 => x"84",
          2829 => x"43",
          2830 => x"99",
          2831 => x"33",
          2832 => x"80",
          2833 => x"b1",
          2834 => x"b8",
          2835 => x"33",
          2836 => x"94",
          2837 => x"78",
          2838 => x"83",
          2839 => x"06",
          2840 => x"5c",
          2841 => x"b8",
          2842 => x"89",
          2843 => x"76",
          2844 => x"61",
          2845 => x"38",
          2846 => x"62",
          2847 => x"1f",
          2848 => x"79",
          2849 => x"ac",
          2850 => x"a4",
          2851 => x"2b",
          2852 => x"07",
          2853 => x"57",
          2854 => x"70",
          2855 => x"84",
          2856 => x"38",
          2857 => x"33",
          2858 => x"81",
          2859 => x"73",
          2860 => x"77",
          2861 => x"1b",
          2862 => x"75",
          2863 => x"f4",
          2864 => x"99",
          2865 => x"e0",
          2866 => x"5a",
          2867 => x"f4",
          2868 => x"34",
          2869 => x"81",
          2870 => x"f4",
          2871 => x"06",
          2872 => x"b0",
          2873 => x"2b",
          2874 => x"58",
          2875 => x"81",
          2876 => x"fa",
          2877 => x"06",
          2878 => x"b6",
          2879 => x"33",
          2880 => x"b8",
          2881 => x"b8",
          2882 => x"ee",
          2883 => x"56",
          2884 => x"70",
          2885 => x"39",
          2886 => x"85",
          2887 => x"e5",
          2888 => x"06",
          2889 => x"34",
          2890 => x"f9",
          2891 => x"b0",
          2892 => x"81",
          2893 => x"fa",
          2894 => x"0b",
          2895 => x"81",
          2896 => x"83",
          2897 => x"75",
          2898 => x"83",
          2899 => x"07",
          2900 => x"fd",
          2901 => x"06",
          2902 => x"b0",
          2903 => x"33",
          2904 => x"75",
          2905 => x"83",
          2906 => x"07",
          2907 => x"c5",
          2908 => x"06",
          2909 => x"34",
          2910 => x"81",
          2911 => x"fa",
          2912 => x"b0",
          2913 => x"75",
          2914 => x"83",
          2915 => x"75",
          2916 => x"83",
          2917 => x"75",
          2918 => x"83",
          2919 => x"75",
          2920 => x"83",
          2921 => x"d0",
          2922 => x"fd",
          2923 => x"bf",
          2924 => x"b0",
          2925 => x"fa",
          2926 => x"c9",
          2927 => x"33",
          2928 => x"33",
          2929 => x"33",
          2930 => x"0b",
          2931 => x"81",
          2932 => x"84",
          2933 => x"77",
          2934 => x"33",
          2935 => x"56",
          2936 => x"9c",
          2937 => x"fe",
          2938 => x"a1",
          2939 => x"80",
          2940 => x"80",
          2941 => x"0d",
          2942 => x"e9",
          2943 => x"5c",
          2944 => x"10",
          2945 => x"05",
          2946 => x"0b",
          2947 => x"0b",
          2948 => x"51",
          2949 => x"70",
          2950 => x"e6",
          2951 => x"34",
          2952 => x"ef",
          2953 => x"3f",
          2954 => x"ff",
          2955 => x"06",
          2956 => x"52",
          2957 => x"33",
          2958 => x"75",
          2959 => x"83",
          2960 => x"70",
          2961 => x"f0",
          2962 => x"05",
          2963 => x"59",
          2964 => x"75",
          2965 => x"33",
          2966 => x"77",
          2967 => x"33",
          2968 => x"06",
          2969 => x"11",
          2970 => x"b2",
          2971 => x"70",
          2972 => x"33",
          2973 => x"81",
          2974 => x"ff",
          2975 => x"24",
          2976 => x"56",
          2977 => x"16",
          2978 => x"81",
          2979 => x"76",
          2980 => x"33",
          2981 => x"ff",
          2982 => x"7b",
          2983 => x"57",
          2984 => x"38",
          2985 => x"ff",
          2986 => x"79",
          2987 => x"c7",
          2988 => x"81",
          2989 => x"42",
          2990 => x"38",
          2991 => x"17",
          2992 => x"7b",
          2993 => x"81",
          2994 => x"5f",
          2995 => x"84",
          2996 => x"59",
          2997 => x"b1",
          2998 => x"b9",
          2999 => x"5d",
          3000 => x"7d",
          3001 => x"84",
          3002 => x"71",
          3003 => x"75",
          3004 => x"39",
          3005 => x"b9",
          3006 => x"b4",
          3007 => x"b2",
          3008 => x"5f",
          3009 => x"38",
          3010 => x"06",
          3011 => x"27",
          3012 => x"b2",
          3013 => x"58",
          3014 => x"57",
          3015 => x"f8",
          3016 => x"52",
          3017 => x"38",
          3018 => x"eb",
          3019 => x"05",
          3020 => x"40",
          3021 => x"75",
          3022 => x"09",
          3023 => x"b5",
          3024 => x"b4",
          3025 => x"ff",
          3026 => x"f6",
          3027 => x"fa",
          3028 => x"56",
          3029 => x"39",
          3030 => x"b4",
          3031 => x"56",
          3032 => x"76",
          3033 => x"b0",
          3034 => x"75",
          3035 => x"70",
          3036 => x"33",
          3037 => x"76",
          3038 => x"7b",
          3039 => x"f1",
          3040 => x"34",
          3041 => x"23",
          3042 => x"b2",
          3043 => x"fa",
          3044 => x"b6",
          3045 => x"33",
          3046 => x"34",
          3047 => x"97",
          3048 => x"54",
          3049 => x"db",
          3050 => x"0c",
          3051 => x"51",
          3052 => x"84",
          3053 => x"0d",
          3054 => x"83",
          3055 => x"83",
          3056 => x"59",
          3057 => x"14",
          3058 => x"59",
          3059 => x"0d",
          3060 => x"53",
          3061 => x"32",
          3062 => x"9f",
          3063 => x"f8",
          3064 => x"81",
          3065 => x"54",
          3066 => x"25",
          3067 => x"2e",
          3068 => x"83",
          3069 => x"72",
          3070 => x"05",
          3071 => x"71",
          3072 => x"06",
          3073 => x"58",
          3074 => x"f0",
          3075 => x"80",
          3076 => x"c0",
          3077 => x"f6",
          3078 => x"76",
          3079 => x"70",
          3080 => x"74",
          3081 => x"a4",
          3082 => x"f8",
          3083 => x"76",
          3084 => x"2e",
          3085 => x"15",
          3086 => x"81",
          3087 => x"f8",
          3088 => x"33",
          3089 => x"70",
          3090 => x"27",
          3091 => x"70",
          3092 => x"54",
          3093 => x"ff",
          3094 => x"81",
          3095 => x"85",
          3096 => x"34",
          3097 => x"2e",
          3098 => x"de",
          3099 => x"83",
          3100 => x"70",
          3101 => x"33",
          3102 => x"83",
          3103 => x"ff",
          3104 => x"33",
          3105 => x"83",
          3106 => x"ff",
          3107 => x"33",
          3108 => x"ff",
          3109 => x"38",
          3110 => x"81",
          3111 => x"06",
          3112 => x"38",
          3113 => x"74",
          3114 => x"08",
          3115 => x"08",
          3116 => x"38",
          3117 => x"83",
          3118 => x"81",
          3119 => x"fe",
          3120 => x"77",
          3121 => x"53",
          3122 => x"10",
          3123 => x"08",
          3124 => x"80",
          3125 => x"c0",
          3126 => x"27",
          3127 => x"8a",
          3128 => x"38",
          3129 => x"87",
          3130 => x"0c",
          3131 => x"2e",
          3132 => x"54",
          3133 => x"81",
          3134 => x"e4",
          3135 => x"38",
          3136 => x"c3",
          3137 => x"39",
          3138 => x"56",
          3139 => x"38",
          3140 => x"b4",
          3141 => x"79",
          3142 => x"ff",
          3143 => x"2b",
          3144 => x"73",
          3145 => x"81",
          3146 => x"87",
          3147 => x"57",
          3148 => x"78",
          3149 => x"11",
          3150 => x"05",
          3151 => x"c0",
          3152 => x"57",
          3153 => x"2e",
          3154 => x"59",
          3155 => x"39",
          3156 => x"0b",
          3157 => x"81",
          3158 => x"70",
          3159 => x"59",
          3160 => x"09",
          3161 => x"2e",
          3162 => x"10",
          3163 => x"5d",
          3164 => x"81",
          3165 => x"93",
          3166 => x"33",
          3167 => x"84",
          3168 => x"38",
          3169 => x"cc",
          3170 => x"8f",
          3171 => x"f0",
          3172 => x"2e",
          3173 => x"81",
          3174 => x"34",
          3175 => x"cc",
          3176 => x"15",
          3177 => x"34",
          3178 => x"53",
          3179 => x"83",
          3180 => x"27",
          3181 => x"54",
          3182 => x"fc",
          3183 => x"05",
          3184 => x"74",
          3185 => x"98",
          3186 => x"81",
          3187 => x"0b",
          3188 => x"39",
          3189 => x"81",
          3190 => x"83",
          3191 => x"dd",
          3192 => x"de",
          3193 => x"f8",
          3194 => x"5e",
          3195 => x"09",
          3196 => x"7a",
          3197 => x"2e",
          3198 => x"93",
          3199 => x"f8",
          3200 => x"33",
          3201 => x"73",
          3202 => x"ac",
          3203 => x"58",
          3204 => x"84",
          3205 => x"39",
          3206 => x"2e",
          3207 => x"e4",
          3208 => x"33",
          3209 => x"5a",
          3210 => x"55",
          3211 => x"ff",
          3212 => x"27",
          3213 => x"b4",
          3214 => x"ff",
          3215 => x"27",
          3216 => x"b5",
          3217 => x"52",
          3218 => x"59",
          3219 => x"39",
          3220 => x"51",
          3221 => x"f9",
          3222 => x"fc",
          3223 => x"f5",
          3224 => x"3d",
          3225 => x"53",
          3226 => x"34",
          3227 => x"71",
          3228 => x"55",
          3229 => x"0b",
          3230 => x"98",
          3231 => x"80",
          3232 => x"9c",
          3233 => x"51",
          3234 => x"33",
          3235 => x"74",
          3236 => x"2e",
          3237 => x"51",
          3238 => x"38",
          3239 => x"38",
          3240 => x"90",
          3241 => x"52",
          3242 => x"72",
          3243 => x"c0",
          3244 => x"27",
          3245 => x"38",
          3246 => x"75",
          3247 => x"ff",
          3248 => x"75",
          3249 => x"06",
          3250 => x"2e",
          3251 => x"88",
          3252 => x"84",
          3253 => x"0d",
          3254 => x"56",
          3255 => x"73",
          3256 => x"70",
          3257 => x"57",
          3258 => x"51",
          3259 => x"56",
          3260 => x"34",
          3261 => x"13",
          3262 => x"e1",
          3263 => x"08",
          3264 => x"80",
          3265 => x"c0",
          3266 => x"55",
          3267 => x"98",
          3268 => x"08",
          3269 => x"14",
          3270 => x"52",
          3271 => x"fe",
          3272 => x"08",
          3273 => x"c8",
          3274 => x"c0",
          3275 => x"ce",
          3276 => x"08",
          3277 => x"74",
          3278 => x"87",
          3279 => x"73",
          3280 => x"db",
          3281 => x"72",
          3282 => x"55",
          3283 => x"53",
          3284 => x"81",
          3285 => x"74",
          3286 => x"aa",
          3287 => x"11",
          3288 => x"38",
          3289 => x"70",
          3290 => x"f0",
          3291 => x"3d",
          3292 => x"0c",
          3293 => x"39",
          3294 => x"a3",
          3295 => x"f5",
          3296 => x"80",
          3297 => x"51",
          3298 => x"72",
          3299 => x"75",
          3300 => x"72",
          3301 => x"08",
          3302 => x"54",
          3303 => x"70",
          3304 => x"81",
          3305 => x"38",
          3306 => x"15",
          3307 => x"e2",
          3308 => x"08",
          3309 => x"80",
          3310 => x"c0",
          3311 => x"55",
          3312 => x"98",
          3313 => x"08",
          3314 => x"14",
          3315 => x"52",
          3316 => x"fe",
          3317 => x"08",
          3318 => x"c8",
          3319 => x"c0",
          3320 => x"ce",
          3321 => x"08",
          3322 => x"74",
          3323 => x"87",
          3324 => x"73",
          3325 => x"db",
          3326 => x"72",
          3327 => x"55",
          3328 => x"53",
          3329 => x"ff",
          3330 => x"51",
          3331 => x"2e",
          3332 => x"84",
          3333 => x"e8",
          3334 => x"08",
          3335 => x"83",
          3336 => x"81",
          3337 => x"e8",
          3338 => x"f5",
          3339 => x"54",
          3340 => x"c0",
          3341 => x"f6",
          3342 => x"9c",
          3343 => x"38",
          3344 => x"c0",
          3345 => x"74",
          3346 => x"ff",
          3347 => x"9c",
          3348 => x"c0",
          3349 => x"9c",
          3350 => x"81",
          3351 => x"55",
          3352 => x"81",
          3353 => x"a4",
          3354 => x"ff",
          3355 => x"ff",
          3356 => x"38",
          3357 => x"d5",
          3358 => x"e6",
          3359 => x"3d",
          3360 => x"f4",
          3361 => x"83",
          3362 => x"11",
          3363 => x"2b",
          3364 => x"33",
          3365 => x"90",
          3366 => x"5d",
          3367 => x"71",
          3368 => x"11",
          3369 => x"71",
          3370 => x"81",
          3371 => x"2b",
          3372 => x"52",
          3373 => x"13",
          3374 => x"71",
          3375 => x"2a",
          3376 => x"34",
          3377 => x"13",
          3378 => x"84",
          3379 => x"2b",
          3380 => x"54",
          3381 => x"14",
          3382 => x"80",
          3383 => x"13",
          3384 => x"84",
          3385 => x"ba",
          3386 => x"33",
          3387 => x"07",
          3388 => x"74",
          3389 => x"3d",
          3390 => x"33",
          3391 => x"75",
          3392 => x"71",
          3393 => x"58",
          3394 => x"12",
          3395 => x"f4",
          3396 => x"12",
          3397 => x"07",
          3398 => x"12",
          3399 => x"07",
          3400 => x"77",
          3401 => x"84",
          3402 => x"12",
          3403 => x"ff",
          3404 => x"52",
          3405 => x"84",
          3406 => x"81",
          3407 => x"2b",
          3408 => x"33",
          3409 => x"8f",
          3410 => x"2a",
          3411 => x"54",
          3412 => x"14",
          3413 => x"70",
          3414 => x"71",
          3415 => x"81",
          3416 => x"ff",
          3417 => x"53",
          3418 => x"34",
          3419 => x"08",
          3420 => x"33",
          3421 => x"74",
          3422 => x"98",
          3423 => x"5d",
          3424 => x"25",
          3425 => x"33",
          3426 => x"07",
          3427 => x"75",
          3428 => x"f4",
          3429 => x"33",
          3430 => x"74",
          3431 => x"71",
          3432 => x"5c",
          3433 => x"82",
          3434 => x"3d",
          3435 => x"ba",
          3436 => x"8f",
          3437 => x"51",
          3438 => x"84",
          3439 => x"a0",
          3440 => x"80",
          3441 => x"51",
          3442 => x"08",
          3443 => x"16",
          3444 => x"84",
          3445 => x"84",
          3446 => x"34",
          3447 => x"f4",
          3448 => x"fe",
          3449 => x"06",
          3450 => x"74",
          3451 => x"84",
          3452 => x"84",
          3453 => x"55",
          3454 => x"15",
          3455 => x"7b",
          3456 => x"27",
          3457 => x"05",
          3458 => x"70",
          3459 => x"08",
          3460 => x"88",
          3461 => x"55",
          3462 => x"80",
          3463 => x"70",
          3464 => x"07",
          3465 => x"70",
          3466 => x"56",
          3467 => x"27",
          3468 => x"75",
          3469 => x"13",
          3470 => x"75",
          3471 => x"85",
          3472 => x"83",
          3473 => x"33",
          3474 => x"ff",
          3475 => x"70",
          3476 => x"51",
          3477 => x"51",
          3478 => x"75",
          3479 => x"83",
          3480 => x"07",
          3481 => x"5a",
          3482 => x"84",
          3483 => x"53",
          3484 => x"14",
          3485 => x"70",
          3486 => x"07",
          3487 => x"74",
          3488 => x"88",
          3489 => x"52",
          3490 => x"06",
          3491 => x"f4",
          3492 => x"81",
          3493 => x"19",
          3494 => x"8b",
          3495 => x"58",
          3496 => x"34",
          3497 => x"08",
          3498 => x"33",
          3499 => x"70",
          3500 => x"86",
          3501 => x"ba",
          3502 => x"85",
          3503 => x"2b",
          3504 => x"52",
          3505 => x"34",
          3506 => x"78",
          3507 => x"71",
          3508 => x"5c",
          3509 => x"85",
          3510 => x"84",
          3511 => x"8b",
          3512 => x"15",
          3513 => x"07",
          3514 => x"33",
          3515 => x"5a",
          3516 => x"12",
          3517 => x"f4",
          3518 => x"12",
          3519 => x"07",
          3520 => x"33",
          3521 => x"58",
          3522 => x"70",
          3523 => x"84",
          3524 => x"12",
          3525 => x"ff",
          3526 => x"57",
          3527 => x"84",
          3528 => x"fe",
          3529 => x"ba",
          3530 => x"a0",
          3531 => x"84",
          3532 => x"77",
          3533 => x"08",
          3534 => x"04",
          3535 => x"0c",
          3536 => x"82",
          3537 => x"f4",
          3538 => x"f4",
          3539 => x"81",
          3540 => x"76",
          3541 => x"34",
          3542 => x"17",
          3543 => x"ba",
          3544 => x"05",
          3545 => x"ff",
          3546 => x"56",
          3547 => x"34",
          3548 => x"10",
          3549 => x"55",
          3550 => x"83",
          3551 => x"fe",
          3552 => x"0d",
          3553 => x"ba",
          3554 => x"2e",
          3555 => x"af",
          3556 => x"81",
          3557 => x"fb",
          3558 => x"ff",
          3559 => x"ff",
          3560 => x"83",
          3561 => x"11",
          3562 => x"2b",
          3563 => x"ff",
          3564 => x"73",
          3565 => x"12",
          3566 => x"2b",
          3567 => x"44",
          3568 => x"52",
          3569 => x"fd",
          3570 => x"71",
          3571 => x"19",
          3572 => x"2b",
          3573 => x"56",
          3574 => x"38",
          3575 => x"1b",
          3576 => x"60",
          3577 => x"58",
          3578 => x"18",
          3579 => x"76",
          3580 => x"8b",
          3581 => x"70",
          3582 => x"71",
          3583 => x"53",
          3584 => x"ba",
          3585 => x"12",
          3586 => x"07",
          3587 => x"33",
          3588 => x"7e",
          3589 => x"71",
          3590 => x"57",
          3591 => x"59",
          3592 => x"1d",
          3593 => x"84",
          3594 => x"2b",
          3595 => x"14",
          3596 => x"07",
          3597 => x"40",
          3598 => x"7b",
          3599 => x"16",
          3600 => x"2b",
          3601 => x"2a",
          3602 => x"79",
          3603 => x"70",
          3604 => x"71",
          3605 => x"05",
          3606 => x"2b",
          3607 => x"5d",
          3608 => x"75",
          3609 => x"70",
          3610 => x"8b",
          3611 => x"82",
          3612 => x"2b",
          3613 => x"5d",
          3614 => x"34",
          3615 => x"08",
          3616 => x"33",
          3617 => x"56",
          3618 => x"7e",
          3619 => x"3f",
          3620 => x"61",
          3621 => x"06",
          3622 => x"b6",
          3623 => x"0c",
          3624 => x"0b",
          3625 => x"84",
          3626 => x"60",
          3627 => x"a0",
          3628 => x"7e",
          3629 => x"ba",
          3630 => x"81",
          3631 => x"08",
          3632 => x"87",
          3633 => x"ba",
          3634 => x"07",
          3635 => x"2a",
          3636 => x"34",
          3637 => x"22",
          3638 => x"08",
          3639 => x"15",
          3640 => x"ba",
          3641 => x"76",
          3642 => x"7f",
          3643 => x"f4",
          3644 => x"bb",
          3645 => x"1c",
          3646 => x"71",
          3647 => x"81",
          3648 => x"ff",
          3649 => x"5b",
          3650 => x"1c",
          3651 => x"7c",
          3652 => x"34",
          3653 => x"08",
          3654 => x"71",
          3655 => x"ff",
          3656 => x"ff",
          3657 => x"57",
          3658 => x"34",
          3659 => x"83",
          3660 => x"5b",
          3661 => x"61",
          3662 => x"51",
          3663 => x"39",
          3664 => x"06",
          3665 => x"ff",
          3666 => x"ff",
          3667 => x"71",
          3668 => x"1b",
          3669 => x"2b",
          3670 => x"54",
          3671 => x"f9",
          3672 => x"24",
          3673 => x"8f",
          3674 => x"61",
          3675 => x"39",
          3676 => x"0c",
          3677 => x"82",
          3678 => x"f4",
          3679 => x"f4",
          3680 => x"81",
          3681 => x"7e",
          3682 => x"34",
          3683 => x"19",
          3684 => x"ba",
          3685 => x"05",
          3686 => x"ff",
          3687 => x"44",
          3688 => x"89",
          3689 => x"10",
          3690 => x"f8",
          3691 => x"34",
          3692 => x"39",
          3693 => x"83",
          3694 => x"fb",
          3695 => x"2e",
          3696 => x"3f",
          3697 => x"95",
          3698 => x"33",
          3699 => x"83",
          3700 => x"87",
          3701 => x"2b",
          3702 => x"15",
          3703 => x"2a",
          3704 => x"53",
          3705 => x"34",
          3706 => x"f4",
          3707 => x"12",
          3708 => x"07",
          3709 => x"33",
          3710 => x"5b",
          3711 => x"73",
          3712 => x"05",
          3713 => x"33",
          3714 => x"81",
          3715 => x"5c",
          3716 => x"1e",
          3717 => x"82",
          3718 => x"2b",
          3719 => x"33",
          3720 => x"70",
          3721 => x"57",
          3722 => x"1d",
          3723 => x"70",
          3724 => x"71",
          3725 => x"33",
          3726 => x"70",
          3727 => x"5c",
          3728 => x"83",
          3729 => x"1f",
          3730 => x"88",
          3731 => x"83",
          3732 => x"84",
          3733 => x"ba",
          3734 => x"ff",
          3735 => x"84",
          3736 => x"a0",
          3737 => x"80",
          3738 => x"51",
          3739 => x"08",
          3740 => x"17",
          3741 => x"84",
          3742 => x"84",
          3743 => x"34",
          3744 => x"f4",
          3745 => x"fe",
          3746 => x"06",
          3747 => x"61",
          3748 => x"84",
          3749 => x"84",
          3750 => x"5d",
          3751 => x"1c",
          3752 => x"54",
          3753 => x"1a",
          3754 => x"07",
          3755 => x"33",
          3756 => x"5c",
          3757 => x"84",
          3758 => x"84",
          3759 => x"33",
          3760 => x"83",
          3761 => x"87",
          3762 => x"88",
          3763 => x"59",
          3764 => x"64",
          3765 => x"1d",
          3766 => x"2b",
          3767 => x"2a",
          3768 => x"7f",
          3769 => x"70",
          3770 => x"8b",
          3771 => x"70",
          3772 => x"07",
          3773 => x"77",
          3774 => x"5a",
          3775 => x"17",
          3776 => x"f4",
          3777 => x"33",
          3778 => x"74",
          3779 => x"88",
          3780 => x"88",
          3781 => x"41",
          3782 => x"05",
          3783 => x"fa",
          3784 => x"33",
          3785 => x"79",
          3786 => x"71",
          3787 => x"5e",
          3788 => x"34",
          3789 => x"08",
          3790 => x"33",
          3791 => x"74",
          3792 => x"71",
          3793 => x"56",
          3794 => x"60",
          3795 => x"34",
          3796 => x"81",
          3797 => x"ff",
          3798 => x"58",
          3799 => x"34",
          3800 => x"33",
          3801 => x"83",
          3802 => x"12",
          3803 => x"2b",
          3804 => x"88",
          3805 => x"42",
          3806 => x"83",
          3807 => x"1f",
          3808 => x"2b",
          3809 => x"33",
          3810 => x"81",
          3811 => x"54",
          3812 => x"7c",
          3813 => x"f4",
          3814 => x"12",
          3815 => x"07",
          3816 => x"33",
          3817 => x"78",
          3818 => x"71",
          3819 => x"57",
          3820 => x"5a",
          3821 => x"85",
          3822 => x"17",
          3823 => x"8b",
          3824 => x"86",
          3825 => x"2b",
          3826 => x"52",
          3827 => x"34",
          3828 => x"08",
          3829 => x"88",
          3830 => x"88",
          3831 => x"34",
          3832 => x"08",
          3833 => x"33",
          3834 => x"74",
          3835 => x"88",
          3836 => x"45",
          3837 => x"34",
          3838 => x"08",
          3839 => x"71",
          3840 => x"05",
          3841 => x"88",
          3842 => x"45",
          3843 => x"1a",
          3844 => x"f4",
          3845 => x"12",
          3846 => x"62",
          3847 => x"5d",
          3848 => x"fb",
          3849 => x"05",
          3850 => x"ff",
          3851 => x"86",
          3852 => x"2b",
          3853 => x"1c",
          3854 => x"07",
          3855 => x"41",
          3856 => x"61",
          3857 => x"70",
          3858 => x"71",
          3859 => x"05",
          3860 => x"88",
          3861 => x"5f",
          3862 => x"86",
          3863 => x"84",
          3864 => x"12",
          3865 => x"ff",
          3866 => x"55",
          3867 => x"84",
          3868 => x"81",
          3869 => x"2b",
          3870 => x"33",
          3871 => x"8f",
          3872 => x"2a",
          3873 => x"58",
          3874 => x"1e",
          3875 => x"70",
          3876 => x"71",
          3877 => x"81",
          3878 => x"ff",
          3879 => x"49",
          3880 => x"34",
          3881 => x"ff",
          3882 => x"52",
          3883 => x"08",
          3884 => x"93",
          3885 => x"84",
          3886 => x"51",
          3887 => x"27",
          3888 => x"3d",
          3889 => x"08",
          3890 => x"77",
          3891 => x"84",
          3892 => x"e4",
          3893 => x"84",
          3894 => x"77",
          3895 => x"51",
          3896 => x"84",
          3897 => x"f4",
          3898 => x"0b",
          3899 => x"53",
          3900 => x"b5",
          3901 => x"76",
          3902 => x"84",
          3903 => x"34",
          3904 => x"f4",
          3905 => x"0b",
          3906 => x"84",
          3907 => x"80",
          3908 => x"88",
          3909 => x"17",
          3910 => x"f0",
          3911 => x"f4",
          3912 => x"82",
          3913 => x"77",
          3914 => x"fe",
          3915 => x"05",
          3916 => x"87",
          3917 => x"71",
          3918 => x"04",
          3919 => x"52",
          3920 => x"71",
          3921 => x"08",
          3922 => x"72",
          3923 => x"80",
          3924 => x"0c",
          3925 => x"7c",
          3926 => x"33",
          3927 => x"74",
          3928 => x"33",
          3929 => x"73",
          3930 => x"c0",
          3931 => x"76",
          3932 => x"08",
          3933 => x"a7",
          3934 => x"73",
          3935 => x"74",
          3936 => x"2e",
          3937 => x"84",
          3938 => x"84",
          3939 => x"06",
          3940 => x"ac",
          3941 => x"7e",
          3942 => x"5a",
          3943 => x"26",
          3944 => x"54",
          3945 => x"bd",
          3946 => x"98",
          3947 => x"51",
          3948 => x"81",
          3949 => x"38",
          3950 => x"e2",
          3951 => x"fc",
          3952 => x"83",
          3953 => x"bb",
          3954 => x"80",
          3955 => x"5a",
          3956 => x"38",
          3957 => x"84",
          3958 => x"9f",
          3959 => x"71",
          3960 => x"12",
          3961 => x"53",
          3962 => x"98",
          3963 => x"96",
          3964 => x"83",
          3965 => x"bb",
          3966 => x"80",
          3967 => x"0c",
          3968 => x"0c",
          3969 => x"3d",
          3970 => x"92",
          3971 => x"71",
          3972 => x"51",
          3973 => x"98",
          3974 => x"c0",
          3975 => x"81",
          3976 => x"52",
          3977 => x"2e",
          3978 => x"54",
          3979 => x"3d",
          3980 => x"33",
          3981 => x"09",
          3982 => x"75",
          3983 => x"80",
          3984 => x"3f",
          3985 => x"38",
          3986 => x"8c",
          3987 => x"08",
          3988 => x"33",
          3989 => x"84",
          3990 => x"06",
          3991 => x"19",
          3992 => x"08",
          3993 => x"08",
          3994 => x"ff",
          3995 => x"82",
          3996 => x"81",
          3997 => x"18",
          3998 => x"33",
          3999 => x"06",
          4000 => x"76",
          4001 => x"38",
          4002 => x"57",
          4003 => x"ff",
          4004 => x"0b",
          4005 => x"84",
          4006 => x"80",
          4007 => x"0b",
          4008 => x"19",
          4009 => x"34",
          4010 => x"80",
          4011 => x"e1",
          4012 => x"08",
          4013 => x"88",
          4014 => x"74",
          4015 => x"34",
          4016 => x"19",
          4017 => x"a4",
          4018 => x"84",
          4019 => x"75",
          4020 => x"55",
          4021 => x"08",
          4022 => x"81",
          4023 => x"33",
          4024 => x"34",
          4025 => x"51",
          4026 => x"80",
          4027 => x"f3",
          4028 => x"56",
          4029 => x"17",
          4030 => x"77",
          4031 => x"04",
          4032 => x"2e",
          4033 => x"a5",
          4034 => x"dd",
          4035 => x"2a",
          4036 => x"5b",
          4037 => x"83",
          4038 => x"81",
          4039 => x"53",
          4040 => x"f8",
          4041 => x"2e",
          4042 => x"b4",
          4043 => x"83",
          4044 => x"1c",
          4045 => x"53",
          4046 => x"2e",
          4047 => x"71",
          4048 => x"81",
          4049 => x"53",
          4050 => x"f8",
          4051 => x"2e",
          4052 => x"b4",
          4053 => x"83",
          4054 => x"88",
          4055 => x"84",
          4056 => x"fe",
          4057 => x"bb",
          4058 => x"88",
          4059 => x"17",
          4060 => x"83",
          4061 => x"7b",
          4062 => x"81",
          4063 => x"17",
          4064 => x"84",
          4065 => x"81",
          4066 => x"df",
          4067 => x"05",
          4068 => x"71",
          4069 => x"57",
          4070 => x"2e",
          4071 => x"87",
          4072 => x"17",
          4073 => x"83",
          4074 => x"7b",
          4075 => x"81",
          4076 => x"17",
          4077 => x"84",
          4078 => x"81",
          4079 => x"f7",
          4080 => x"77",
          4081 => x"12",
          4082 => x"07",
          4083 => x"2b",
          4084 => x"80",
          4085 => x"5c",
          4086 => x"04",
          4087 => x"17",
          4088 => x"f6",
          4089 => x"08",
          4090 => x"38",
          4091 => x"b4",
          4092 => x"bb",
          4093 => x"08",
          4094 => x"55",
          4095 => x"f7",
          4096 => x"18",
          4097 => x"33",
          4098 => x"df",
          4099 => x"b8",
          4100 => x"5c",
          4101 => x"7b",
          4102 => x"84",
          4103 => x"17",
          4104 => x"a0",
          4105 => x"33",
          4106 => x"84",
          4107 => x"81",
          4108 => x"70",
          4109 => x"bb",
          4110 => x"7b",
          4111 => x"84",
          4112 => x"17",
          4113 => x"84",
          4114 => x"27",
          4115 => x"74",
          4116 => x"38",
          4117 => x"08",
          4118 => x"51",
          4119 => x"39",
          4120 => x"17",
          4121 => x"f4",
          4122 => x"08",
          4123 => x"38",
          4124 => x"b4",
          4125 => x"bb",
          4126 => x"08",
          4127 => x"55",
          4128 => x"84",
          4129 => x"18",
          4130 => x"33",
          4131 => x"ec",
          4132 => x"18",
          4133 => x"33",
          4134 => x"81",
          4135 => x"39",
          4136 => x"57",
          4137 => x"38",
          4138 => x"78",
          4139 => x"74",
          4140 => x"2e",
          4141 => x"0c",
          4142 => x"a8",
          4143 => x"1a",
          4144 => x"b6",
          4145 => x"7c",
          4146 => x"38",
          4147 => x"81",
          4148 => x"bb",
          4149 => x"58",
          4150 => x"58",
          4151 => x"fe",
          4152 => x"06",
          4153 => x"88",
          4154 => x"0b",
          4155 => x"0c",
          4156 => x"09",
          4157 => x"2a",
          4158 => x"b4",
          4159 => x"85",
          4160 => x"5d",
          4161 => x"bd",
          4162 => x"52",
          4163 => x"84",
          4164 => x"ff",
          4165 => x"79",
          4166 => x"2b",
          4167 => x"83",
          4168 => x"06",
          4169 => x"5e",
          4170 => x"56",
          4171 => x"5a",
          4172 => x"5b",
          4173 => x"1a",
          4174 => x"16",
          4175 => x"b4",
          4176 => x"2e",
          4177 => x"71",
          4178 => x"81",
          4179 => x"53",
          4180 => x"f0",
          4181 => x"2e",
          4182 => x"b4",
          4183 => x"38",
          4184 => x"81",
          4185 => x"7a",
          4186 => x"84",
          4187 => x"06",
          4188 => x"81",
          4189 => x"a8",
          4190 => x"1a",
          4191 => x"dd",
          4192 => x"70",
          4193 => x"9b",
          4194 => x"7f",
          4195 => x"84",
          4196 => x"19",
          4197 => x"1b",
          4198 => x"56",
          4199 => x"19",
          4200 => x"38",
          4201 => x"19",
          4202 => x"84",
          4203 => x"81",
          4204 => x"83",
          4205 => x"05",
          4206 => x"38",
          4207 => x"06",
          4208 => x"76",
          4209 => x"cb",
          4210 => x"70",
          4211 => x"8b",
          4212 => x"7c",
          4213 => x"84",
          4214 => x"19",
          4215 => x"1b",
          4216 => x"40",
          4217 => x"82",
          4218 => x"81",
          4219 => x"1e",
          4220 => x"ee",
          4221 => x"81",
          4222 => x"81",
          4223 => x"81",
          4224 => x"09",
          4225 => x"84",
          4226 => x"70",
          4227 => x"84",
          4228 => x"74",
          4229 => x"33",
          4230 => x"fc",
          4231 => x"76",
          4232 => x"3f",
          4233 => x"76",
          4234 => x"33",
          4235 => x"84",
          4236 => x"06",
          4237 => x"83",
          4238 => x"1b",
          4239 => x"84",
          4240 => x"27",
          4241 => x"74",
          4242 => x"38",
          4243 => x"81",
          4244 => x"5a",
          4245 => x"53",
          4246 => x"f3",
          4247 => x"76",
          4248 => x"83",
          4249 => x"b8",
          4250 => x"b9",
          4251 => x"fd",
          4252 => x"fc",
          4253 => x"33",
          4254 => x"f0",
          4255 => x"58",
          4256 => x"75",
          4257 => x"79",
          4258 => x"7a",
          4259 => x"3d",
          4260 => x"5a",
          4261 => x"57",
          4262 => x"9c",
          4263 => x"19",
          4264 => x"80",
          4265 => x"38",
          4266 => x"08",
          4267 => x"77",
          4268 => x"51",
          4269 => x"80",
          4270 => x"bb",
          4271 => x"bb",
          4272 => x"07",
          4273 => x"55",
          4274 => x"2e",
          4275 => x"55",
          4276 => x"0d",
          4277 => x"bb",
          4278 => x"79",
          4279 => x"84",
          4280 => x"bb",
          4281 => x"ff",
          4282 => x"bb",
          4283 => x"fe",
          4284 => x"08",
          4285 => x"52",
          4286 => x"84",
          4287 => x"38",
          4288 => x"70",
          4289 => x"84",
          4290 => x"55",
          4291 => x"08",
          4292 => x"54",
          4293 => x"9c",
          4294 => x"70",
          4295 => x"2e",
          4296 => x"78",
          4297 => x"08",
          4298 => x"bb",
          4299 => x"55",
          4300 => x"38",
          4301 => x"fe",
          4302 => x"78",
          4303 => x"0c",
          4304 => x"84",
          4305 => x"84",
          4306 => x"84",
          4307 => x"84",
          4308 => x"73",
          4309 => x"7a",
          4310 => x"bb",
          4311 => x"bb",
          4312 => x"3d",
          4313 => x"ff",
          4314 => x"f8",
          4315 => x"55",
          4316 => x"df",
          4317 => x"d7",
          4318 => x"08",
          4319 => x"56",
          4320 => x"85",
          4321 => x"5a",
          4322 => x"17",
          4323 => x"0c",
          4324 => x"80",
          4325 => x"98",
          4326 => x"b8",
          4327 => x"84",
          4328 => x"82",
          4329 => x"0d",
          4330 => x"2e",
          4331 => x"89",
          4332 => x"38",
          4333 => x"14",
          4334 => x"8d",
          4335 => x"b0",
          4336 => x"19",
          4337 => x"51",
          4338 => x"55",
          4339 => x"38",
          4340 => x"ff",
          4341 => x"bb",
          4342 => x"73",
          4343 => x"38",
          4344 => x"84",
          4345 => x"0d",
          4346 => x"05",
          4347 => x"27",
          4348 => x"98",
          4349 => x"2e",
          4350 => x"7a",
          4351 => x"57",
          4352 => x"88",
          4353 => x"81",
          4354 => x"90",
          4355 => x"18",
          4356 => x"0c",
          4357 => x"0c",
          4358 => x"2a",
          4359 => x"76",
          4360 => x"08",
          4361 => x"84",
          4362 => x"bb",
          4363 => x"19",
          4364 => x"91",
          4365 => x"94",
          4366 => x"3f",
          4367 => x"84",
          4368 => x"38",
          4369 => x"2e",
          4370 => x"84",
          4371 => x"bb",
          4372 => x"7d",
          4373 => x"08",
          4374 => x"78",
          4375 => x"71",
          4376 => x"7b",
          4377 => x"80",
          4378 => x"05",
          4379 => x"38",
          4380 => x"75",
          4381 => x"1c",
          4382 => x"e4",
          4383 => x"e7",
          4384 => x"98",
          4385 => x"0c",
          4386 => x"19",
          4387 => x"1a",
          4388 => x"bb",
          4389 => x"84",
          4390 => x"a8",
          4391 => x"08",
          4392 => x"5c",
          4393 => x"db",
          4394 => x"1a",
          4395 => x"33",
          4396 => x"8a",
          4397 => x"06",
          4398 => x"a7",
          4399 => x"9c",
          4400 => x"58",
          4401 => x"19",
          4402 => x"05",
          4403 => x"81",
          4404 => x"0d",
          4405 => x"5c",
          4406 => x"70",
          4407 => x"80",
          4408 => x"75",
          4409 => x"2e",
          4410 => x"58",
          4411 => x"81",
          4412 => x"19",
          4413 => x"3f",
          4414 => x"38",
          4415 => x"0c",
          4416 => x"1c",
          4417 => x"2e",
          4418 => x"06",
          4419 => x"86",
          4420 => x"30",
          4421 => x"25",
          4422 => x"57",
          4423 => x"06",
          4424 => x"38",
          4425 => x"ff",
          4426 => x"3f",
          4427 => x"84",
          4428 => x"56",
          4429 => x"84",
          4430 => x"b4",
          4431 => x"33",
          4432 => x"bb",
          4433 => x"fe",
          4434 => x"1a",
          4435 => x"31",
          4436 => x"a0",
          4437 => x"19",
          4438 => x"06",
          4439 => x"08",
          4440 => x"81",
          4441 => x"57",
          4442 => x"81",
          4443 => x"81",
          4444 => x"8d",
          4445 => x"90",
          4446 => x"5e",
          4447 => x"ff",
          4448 => x"56",
          4449 => x"be",
          4450 => x"98",
          4451 => x"94",
          4452 => x"39",
          4453 => x"09",
          4454 => x"9b",
          4455 => x"2b",
          4456 => x"38",
          4457 => x"29",
          4458 => x"5b",
          4459 => x"81",
          4460 => x"07",
          4461 => x"c5",
          4462 => x"38",
          4463 => x"75",
          4464 => x"57",
          4465 => x"70",
          4466 => x"80",
          4467 => x"fe",
          4468 => x"80",
          4469 => x"06",
          4470 => x"ff",
          4471 => x"fe",
          4472 => x"8b",
          4473 => x"29",
          4474 => x"40",
          4475 => x"19",
          4476 => x"7e",
          4477 => x"1d",
          4478 => x"3d",
          4479 => x"08",
          4480 => x"cf",
          4481 => x"bb",
          4482 => x"70",
          4483 => x"b8",
          4484 => x"58",
          4485 => x"38",
          4486 => x"78",
          4487 => x"81",
          4488 => x"1b",
          4489 => x"84",
          4490 => x"81",
          4491 => x"76",
          4492 => x"33",
          4493 => x"38",
          4494 => x"ff",
          4495 => x"76",
          4496 => x"83",
          4497 => x"81",
          4498 => x"8f",
          4499 => x"78",
          4500 => x"2a",
          4501 => x"81",
          4502 => x"81",
          4503 => x"76",
          4504 => x"38",
          4505 => x"a7",
          4506 => x"78",
          4507 => x"81",
          4508 => x"1a",
          4509 => x"81",
          4510 => x"81",
          4511 => x"80",
          4512 => x"bb",
          4513 => x"80",
          4514 => x"84",
          4515 => x"b4",
          4516 => x"33",
          4517 => x"bb",
          4518 => x"fe",
          4519 => x"1c",
          4520 => x"31",
          4521 => x"a0",
          4522 => x"1b",
          4523 => x"06",
          4524 => x"08",
          4525 => x"81",
          4526 => x"57",
          4527 => x"39",
          4528 => x"06",
          4529 => x"86",
          4530 => x"93",
          4531 => x"06",
          4532 => x"0c",
          4533 => x"38",
          4534 => x"7b",
          4535 => x"08",
          4536 => x"fc",
          4537 => x"2e",
          4538 => x"0b",
          4539 => x"19",
          4540 => x"06",
          4541 => x"33",
          4542 => x"59",
          4543 => x"33",
          4544 => x"5b",
          4545 => x"84",
          4546 => x"71",
          4547 => x"57",
          4548 => x"81",
          4549 => x"81",
          4550 => x"7a",
          4551 => x"81",
          4552 => x"75",
          4553 => x"06",
          4554 => x"58",
          4555 => x"33",
          4556 => x"75",
          4557 => x"8d",
          4558 => x"41",
          4559 => x"70",
          4560 => x"39",
          4561 => x"3d",
          4562 => x"ff",
          4563 => x"39",
          4564 => x"ab",
          4565 => x"5d",
          4566 => x"74",
          4567 => x"5d",
          4568 => x"70",
          4569 => x"74",
          4570 => x"40",
          4571 => x"70",
          4572 => x"05",
          4573 => x"38",
          4574 => x"06",
          4575 => x"38",
          4576 => x"0b",
          4577 => x"7b",
          4578 => x"55",
          4579 => x"70",
          4580 => x"74",
          4581 => x"38",
          4582 => x"2e",
          4583 => x"8f",
          4584 => x"76",
          4585 => x"72",
          4586 => x"57",
          4587 => x"a0",
          4588 => x"80",
          4589 => x"ca",
          4590 => x"05",
          4591 => x"55",
          4592 => x"55",
          4593 => x"78",
          4594 => x"38",
          4595 => x"76",
          4596 => x"38",
          4597 => x"38",
          4598 => x"a2",
          4599 => x"74",
          4600 => x"81",
          4601 => x"8e",
          4602 => x"81",
          4603 => x"77",
          4604 => x"7d",
          4605 => x"08",
          4606 => x"7b",
          4607 => x"80",
          4608 => x"84",
          4609 => x"2e",
          4610 => x"80",
          4611 => x"08",
          4612 => x"57",
          4613 => x"81",
          4614 => x"52",
          4615 => x"84",
          4616 => x"7d",
          4617 => x"08",
          4618 => x"38",
          4619 => x"59",
          4620 => x"18",
          4621 => x"18",
          4622 => x"06",
          4623 => x"b8",
          4624 => x"a4",
          4625 => x"85",
          4626 => x"19",
          4627 => x"1e",
          4628 => x"e5",
          4629 => x"80",
          4630 => x"2e",
          4631 => x"7b",
          4632 => x"51",
          4633 => x"56",
          4634 => x"88",
          4635 => x"89",
          4636 => x"ff",
          4637 => x"1e",
          4638 => x"af",
          4639 => x"7f",
          4640 => x"b8",
          4641 => x"9c",
          4642 => x"85",
          4643 => x"1d",
          4644 => x"a0",
          4645 => x"76",
          4646 => x"55",
          4647 => x"08",
          4648 => x"05",
          4649 => x"34",
          4650 => x"1e",
          4651 => x"5a",
          4652 => x"1d",
          4653 => x"0c",
          4654 => x"70",
          4655 => x"74",
          4656 => x"7d",
          4657 => x"08",
          4658 => x"fd",
          4659 => x"b4",
          4660 => x"33",
          4661 => x"08",
          4662 => x"38",
          4663 => x"b4",
          4664 => x"74",
          4665 => x"18",
          4666 => x"38",
          4667 => x"39",
          4668 => x"31",
          4669 => x"84",
          4670 => x"08",
          4671 => x"08",
          4672 => x"75",
          4673 => x"05",
          4674 => x"ff",
          4675 => x"e4",
          4676 => x"43",
          4677 => x"b4",
          4678 => x"1c",
          4679 => x"06",
          4680 => x"b8",
          4681 => x"dc",
          4682 => x"85",
          4683 => x"1d",
          4684 => x"8c",
          4685 => x"ff",
          4686 => x"34",
          4687 => x"1c",
          4688 => x"1c",
          4689 => x"77",
          4690 => x"2e",
          4691 => x"81",
          4692 => x"18",
          4693 => x"81",
          4694 => x"75",
          4695 => x"ff",
          4696 => x"cb",
          4697 => x"b3",
          4698 => x"58",
          4699 => x"7b",
          4700 => x"52",
          4701 => x"84",
          4702 => x"f1",
          4703 => x"a9",
          4704 => x"1c",
          4705 => x"1d",
          4706 => x"56",
          4707 => x"84",
          4708 => x"1c",
          4709 => x"84",
          4710 => x"27",
          4711 => x"61",
          4712 => x"38",
          4713 => x"08",
          4714 => x"51",
          4715 => x"39",
          4716 => x"43",
          4717 => x"06",
          4718 => x"70",
          4719 => x"38",
          4720 => x"5d",
          4721 => x"08",
          4722 => x"cf",
          4723 => x"2e",
          4724 => x"84",
          4725 => x"a8",
          4726 => x"08",
          4727 => x"7e",
          4728 => x"08",
          4729 => x"41",
          4730 => x"fc",
          4731 => x"39",
          4732 => x"fc",
          4733 => x"b4",
          4734 => x"61",
          4735 => x"3f",
          4736 => x"08",
          4737 => x"81",
          4738 => x"e3",
          4739 => x"08",
          4740 => x"34",
          4741 => x"38",
          4742 => x"38",
          4743 => x"70",
          4744 => x"78",
          4745 => x"70",
          4746 => x"82",
          4747 => x"83",
          4748 => x"ff",
          4749 => x"76",
          4750 => x"79",
          4751 => x"70",
          4752 => x"18",
          4753 => x"34",
          4754 => x"9c",
          4755 => x"58",
          4756 => x"74",
          4757 => x"32",
          4758 => x"55",
          4759 => x"72",
          4760 => x"81",
          4761 => x"77",
          4762 => x"58",
          4763 => x"18",
          4764 => x"34",
          4765 => x"77",
          4766 => x"34",
          4767 => x"80",
          4768 => x"8c",
          4769 => x"73",
          4770 => x"8b",
          4771 => x"08",
          4772 => x"33",
          4773 => x"81",
          4774 => x"75",
          4775 => x"16",
          4776 => x"07",
          4777 => x"55",
          4778 => x"98",
          4779 => x"54",
          4780 => x"04",
          4781 => x"1d",
          4782 => x"5b",
          4783 => x"74",
          4784 => x"bb",
          4785 => x"81",
          4786 => x"27",
          4787 => x"73",
          4788 => x"78",
          4789 => x"56",
          4790 => x"5c",
          4791 => x"ba",
          4792 => x"07",
          4793 => x"55",
          4794 => x"34",
          4795 => x"1f",
          4796 => x"89",
          4797 => x"2e",
          4798 => x"57",
          4799 => x"11",
          4800 => x"9c",
          4801 => x"88",
          4802 => x"53",
          4803 => x"8a",
          4804 => x"06",
          4805 => x"5a",
          4806 => x"71",
          4807 => x"56",
          4808 => x"72",
          4809 => x"30",
          4810 => x"53",
          4811 => x"3d",
          4812 => x"5c",
          4813 => x"74",
          4814 => x"80",
          4815 => x"2e",
          4816 => x"1d",
          4817 => x"41",
          4818 => x"38",
          4819 => x"57",
          4820 => x"55",
          4821 => x"0c",
          4822 => x"ff",
          4823 => x"18",
          4824 => x"73",
          4825 => x"70",
          4826 => x"07",
          4827 => x"38",
          4828 => x"74",
          4829 => x"a0",
          4830 => x"ff",
          4831 => x"81",
          4832 => x"81",
          4833 => x"56",
          4834 => x"ff",
          4835 => x"81",
          4836 => x"18",
          4837 => x"70",
          4838 => x"57",
          4839 => x"cb",
          4840 => x"30",
          4841 => x"58",
          4842 => x"14",
          4843 => x"55",
          4844 => x"dc",
          4845 => x"07",
          4846 => x"88",
          4847 => x"3d",
          4848 => x"90",
          4849 => x"51",
          4850 => x"08",
          4851 => x"8d",
          4852 => x"0c",
          4853 => x"33",
          4854 => x"80",
          4855 => x"80",
          4856 => x"51",
          4857 => x"84",
          4858 => x"81",
          4859 => x"80",
          4860 => x"7d",
          4861 => x"80",
          4862 => x"af",
          4863 => x"70",
          4864 => x"54",
          4865 => x"9f",
          4866 => x"2e",
          4867 => x"d1",
          4868 => x"a7",
          4869 => x"70",
          4870 => x"9f",
          4871 => x"7c",
          4872 => x"ff",
          4873 => x"77",
          4874 => x"2e",
          4875 => x"83",
          4876 => x"56",
          4877 => x"83",
          4878 => x"82",
          4879 => x"77",
          4880 => x"78",
          4881 => x"fe",
          4882 => x"2e",
          4883 => x"54",
          4884 => x"38",
          4885 => x"74",
          4886 => x"53",
          4887 => x"88",
          4888 => x"57",
          4889 => x"38",
          4890 => x"ae",
          4891 => x"5a",
          4892 => x"72",
          4893 => x"26",
          4894 => x"70",
          4895 => x"7c",
          4896 => x"2e",
          4897 => x"83",
          4898 => x"83",
          4899 => x"76",
          4900 => x"81",
          4901 => x"77",
          4902 => x"53",
          4903 => x"57",
          4904 => x"7c",
          4905 => x"06",
          4906 => x"7d",
          4907 => x"e3",
          4908 => x"75",
          4909 => x"80",
          4910 => x"7d",
          4911 => x"2e",
          4912 => x"ab",
          4913 => x"84",
          4914 => x"54",
          4915 => x"ac",
          4916 => x"09",
          4917 => x"2a",
          4918 => x"f0",
          4919 => x"78",
          4920 => x"56",
          4921 => x"57",
          4922 => x"79",
          4923 => x"7c",
          4924 => x"fd",
          4925 => x"8a",
          4926 => x"2e",
          4927 => x"22",
          4928 => x"fc",
          4929 => x"7b",
          4930 => x"ae",
          4931 => x"54",
          4932 => x"81",
          4933 => x"79",
          4934 => x"7b",
          4935 => x"08",
          4936 => x"84",
          4937 => x"81",
          4938 => x"1c",
          4939 => x"5d",
          4940 => x"1c",
          4941 => x"d3",
          4942 => x"88",
          4943 => x"54",
          4944 => x"88",
          4945 => x"fe",
          4946 => x"2e",
          4947 => x"fb",
          4948 => x"07",
          4949 => x"7d",
          4950 => x"06",
          4951 => x"06",
          4952 => x"fd",
          4953 => x"7c",
          4954 => x"38",
          4955 => x"34",
          4956 => x"3d",
          4957 => x"38",
          4958 => x"ff",
          4959 => x"38",
          4960 => x"5c",
          4961 => x"5a",
          4962 => x"bd",
          4963 => x"ff",
          4964 => x"55",
          4965 => x"ff",
          4966 => x"54",
          4967 => x"74",
          4968 => x"ac",
          4969 => x"ff",
          4970 => x"80",
          4971 => x"81",
          4972 => x"56",
          4973 => x"ff",
          4974 => x"bf",
          4975 => x"7d",
          4976 => x"53",
          4977 => x"93",
          4978 => x"06",
          4979 => x"58",
          4980 => x"59",
          4981 => x"16",
          4982 => x"b3",
          4983 => x"ff",
          4984 => x"ae",
          4985 => x"1d",
          4986 => x"34",
          4987 => x"14",
          4988 => x"2b",
          4989 => x"1f",
          4990 => x"1b",
          4991 => x"72",
          4992 => x"05",
          4993 => x"5b",
          4994 => x"1d",
          4995 => x"09",
          4996 => x"39",
          4997 => x"f6",
          4998 => x"0c",
          4999 => x"67",
          5000 => x"33",
          5001 => x"7e",
          5002 => x"2e",
          5003 => x"5b",
          5004 => x"ba",
          5005 => x"75",
          5006 => x"e0",
          5007 => x"38",
          5008 => x"70",
          5009 => x"2e",
          5010 => x"81",
          5011 => x"80",
          5012 => x"ff",
          5013 => x"81",
          5014 => x"7c",
          5015 => x"34",
          5016 => x"33",
          5017 => x"33",
          5018 => x"84",
          5019 => x"41",
          5020 => x"78",
          5021 => x"81",
          5022 => x"38",
          5023 => x"0b",
          5024 => x"81",
          5025 => x"81",
          5026 => x"3f",
          5027 => x"38",
          5028 => x"0c",
          5029 => x"17",
          5030 => x"2b",
          5031 => x"d4",
          5032 => x"26",
          5033 => x"42",
          5034 => x"84",
          5035 => x"81",
          5036 => x"33",
          5037 => x"07",
          5038 => x"81",
          5039 => x"33",
          5040 => x"07",
          5041 => x"17",
          5042 => x"90",
          5043 => x"33",
          5044 => x"71",
          5045 => x"56",
          5046 => x"33",
          5047 => x"ff",
          5048 => x"59",
          5049 => x"38",
          5050 => x"80",
          5051 => x"8a",
          5052 => x"87",
          5053 => x"61",
          5054 => x"80",
          5055 => x"56",
          5056 => x"8f",
          5057 => x"98",
          5058 => x"18",
          5059 => x"74",
          5060 => x"33",
          5061 => x"88",
          5062 => x"07",
          5063 => x"44",
          5064 => x"17",
          5065 => x"2b",
          5066 => x"2e",
          5067 => x"2a",
          5068 => x"38",
          5069 => x"ec",
          5070 => x"84",
          5071 => x"38",
          5072 => x"ff",
          5073 => x"83",
          5074 => x"75",
          5075 => x"5d",
          5076 => x"a4",
          5077 => x"0c",
          5078 => x"7c",
          5079 => x"22",
          5080 => x"e0",
          5081 => x"19",
          5082 => x"10",
          5083 => x"05",
          5084 => x"59",
          5085 => x"b8",
          5086 => x"0b",
          5087 => x"18",
          5088 => x"7c",
          5089 => x"05",
          5090 => x"86",
          5091 => x"18",
          5092 => x"58",
          5093 => x"0d",
          5094 => x"97",
          5095 => x"70",
          5096 => x"89",
          5097 => x"ff",
          5098 => x"2e",
          5099 => x"e6",
          5100 => x"5a",
          5101 => x"79",
          5102 => x"12",
          5103 => x"38",
          5104 => x"55",
          5105 => x"89",
          5106 => x"58",
          5107 => x"55",
          5108 => x"38",
          5109 => x"70",
          5110 => x"07",
          5111 => x"98",
          5112 => x"83",
          5113 => x"f9",
          5114 => x"38",
          5115 => x"58",
          5116 => x"c0",
          5117 => x"81",
          5118 => x"81",
          5119 => x"70",
          5120 => x"77",
          5121 => x"83",
          5122 => x"83",
          5123 => x"5b",
          5124 => x"16",
          5125 => x"2b",
          5126 => x"33",
          5127 => x"1b",
          5128 => x"40",
          5129 => x"0c",
          5130 => x"80",
          5131 => x"1d",
          5132 => x"71",
          5133 => x"f0",
          5134 => x"43",
          5135 => x"7a",
          5136 => x"83",
          5137 => x"7a",
          5138 => x"38",
          5139 => x"81",
          5140 => x"84",
          5141 => x"ff",
          5142 => x"84",
          5143 => x"7f",
          5144 => x"83",
          5145 => x"81",
          5146 => x"33",
          5147 => x"b7",
          5148 => x"70",
          5149 => x"7f",
          5150 => x"38",
          5151 => x"80",
          5152 => x"58",
          5153 => x"38",
          5154 => x"38",
          5155 => x"1a",
          5156 => x"fe",
          5157 => x"80",
          5158 => x"58",
          5159 => x"70",
          5160 => x"ff",
          5161 => x"2e",
          5162 => x"38",
          5163 => x"b8",
          5164 => x"5d",
          5165 => x"71",
          5166 => x"40",
          5167 => x"80",
          5168 => x"39",
          5169 => x"84",
          5170 => x"75",
          5171 => x"85",
          5172 => x"40",
          5173 => x"84",
          5174 => x"83",
          5175 => x"5c",
          5176 => x"33",
          5177 => x"71",
          5178 => x"77",
          5179 => x"2e",
          5180 => x"83",
          5181 => x"81",
          5182 => x"5c",
          5183 => x"58",
          5184 => x"38",
          5185 => x"77",
          5186 => x"81",
          5187 => x"33",
          5188 => x"07",
          5189 => x"06",
          5190 => x"5a",
          5191 => x"83",
          5192 => x"81",
          5193 => x"53",
          5194 => x"ff",
          5195 => x"80",
          5196 => x"77",
          5197 => x"79",
          5198 => x"84",
          5199 => x"57",
          5200 => x"81",
          5201 => x"11",
          5202 => x"71",
          5203 => x"72",
          5204 => x"5e",
          5205 => x"84",
          5206 => x"06",
          5207 => x"11",
          5208 => x"71",
          5209 => x"72",
          5210 => x"47",
          5211 => x"86",
          5212 => x"06",
          5213 => x"11",
          5214 => x"71",
          5215 => x"72",
          5216 => x"94",
          5217 => x"11",
          5218 => x"71",
          5219 => x"72",
          5220 => x"62",
          5221 => x"5c",
          5222 => x"77",
          5223 => x"5d",
          5224 => x"18",
          5225 => x"0c",
          5226 => x"39",
          5227 => x"7a",
          5228 => x"54",
          5229 => x"53",
          5230 => x"b3",
          5231 => x"09",
          5232 => x"84",
          5233 => x"a8",
          5234 => x"08",
          5235 => x"60",
          5236 => x"84",
          5237 => x"74",
          5238 => x"81",
          5239 => x"58",
          5240 => x"80",
          5241 => x"5f",
          5242 => x"88",
          5243 => x"80",
          5244 => x"33",
          5245 => x"81",
          5246 => x"75",
          5247 => x"7d",
          5248 => x"40",
          5249 => x"2e",
          5250 => x"39",
          5251 => x"3d",
          5252 => x"39",
          5253 => x"bf",
          5254 => x"18",
          5255 => x"33",
          5256 => x"39",
          5257 => x"33",
          5258 => x"5d",
          5259 => x"80",
          5260 => x"33",
          5261 => x"2e",
          5262 => x"ba",
          5263 => x"33",
          5264 => x"73",
          5265 => x"08",
          5266 => x"80",
          5267 => x"86",
          5268 => x"75",
          5269 => x"38",
          5270 => x"05",
          5271 => x"08",
          5272 => x"3d",
          5273 => x"0c",
          5274 => x"11",
          5275 => x"73",
          5276 => x"81",
          5277 => x"79",
          5278 => x"83",
          5279 => x"7e",
          5280 => x"33",
          5281 => x"9f",
          5282 => x"89",
          5283 => x"56",
          5284 => x"26",
          5285 => x"06",
          5286 => x"58",
          5287 => x"85",
          5288 => x"32",
          5289 => x"79",
          5290 => x"92",
          5291 => x"83",
          5292 => x"fe",
          5293 => x"7a",
          5294 => x"e6",
          5295 => x"fb",
          5296 => x"80",
          5297 => x"54",
          5298 => x"84",
          5299 => x"bb",
          5300 => x"80",
          5301 => x"56",
          5302 => x"0d",
          5303 => x"70",
          5304 => x"84",
          5305 => x"2e",
          5306 => x"7c",
          5307 => x"2e",
          5308 => x"f2",
          5309 => x"bb",
          5310 => x"77",
          5311 => x"11",
          5312 => x"07",
          5313 => x"56",
          5314 => x"0b",
          5315 => x"34",
          5316 => x"0b",
          5317 => x"8b",
          5318 => x"0b",
          5319 => x"34",
          5320 => x"d7",
          5321 => x"34",
          5322 => x"9e",
          5323 => x"7e",
          5324 => x"80",
          5325 => x"08",
          5326 => x"81",
          5327 => x"7b",
          5328 => x"7a",
          5329 => x"05",
          5330 => x"80",
          5331 => x"06",
          5332 => x"fe",
          5333 => x"70",
          5334 => x"82",
          5335 => x"5d",
          5336 => x"06",
          5337 => x"2a",
          5338 => x"38",
          5339 => x"11",
          5340 => x"0c",
          5341 => x"71",
          5342 => x"40",
          5343 => x"38",
          5344 => x"11",
          5345 => x"71",
          5346 => x"72",
          5347 => x"60",
          5348 => x"41",
          5349 => x"84",
          5350 => x"0b",
          5351 => x"0c",
          5352 => x"5c",
          5353 => x"70",
          5354 => x"74",
          5355 => x"59",
          5356 => x"1a",
          5357 => x"38",
          5358 => x"70",
          5359 => x"5a",
          5360 => x"80",
          5361 => x"e7",
          5362 => x"7c",
          5363 => x"79",
          5364 => x"84",
          5365 => x"26",
          5366 => x"08",
          5367 => x"56",
          5368 => x"91",
          5369 => x"2a",
          5370 => x"99",
          5371 => x"ce",
          5372 => x"c6",
          5373 => x"be",
          5374 => x"ff",
          5375 => x"33",
          5376 => x"7a",
          5377 => x"11",
          5378 => x"71",
          5379 => x"72",
          5380 => x"62",
          5381 => x"55",
          5382 => x"1b",
          5383 => x"34",
          5384 => x"9c",
          5385 => x"a8",
          5386 => x"fd",
          5387 => x"84",
          5388 => x"57",
          5389 => x"74",
          5390 => x"84",
          5391 => x"08",
          5392 => x"84",
          5393 => x"bb",
          5394 => x"80",
          5395 => x"a0",
          5396 => x"38",
          5397 => x"08",
          5398 => x"38",
          5399 => x"33",
          5400 => x"7c",
          5401 => x"80",
          5402 => x"b4",
          5403 => x"16",
          5404 => x"06",
          5405 => x"b8",
          5406 => x"a3",
          5407 => x"2e",
          5408 => x"b4",
          5409 => x"90",
          5410 => x"b5",
          5411 => x"80",
          5412 => x"17",
          5413 => x"94",
          5414 => x"2b",
          5415 => x"0b",
          5416 => x"34",
          5417 => x"0b",
          5418 => x"8b",
          5419 => x"0b",
          5420 => x"34",
          5421 => x"81",
          5422 => x"77",
          5423 => x"75",
          5424 => x"f8",
          5425 => x"08",
          5426 => x"27",
          5427 => x"71",
          5428 => x"74",
          5429 => x"2a",
          5430 => x"54",
          5431 => x"51",
          5432 => x"08",
          5433 => x"80",
          5434 => x"b4",
          5435 => x"81",
          5436 => x"3f",
          5437 => x"81",
          5438 => x"08",
          5439 => x"17",
          5440 => x"55",
          5441 => x"38",
          5442 => x"09",
          5443 => x"b4",
          5444 => x"77",
          5445 => x"fb",
          5446 => x"bb",
          5447 => x"ee",
          5448 => x"3d",
          5449 => x"5b",
          5450 => x"80",
          5451 => x"80",
          5452 => x"80",
          5453 => x"1a",
          5454 => x"b4",
          5455 => x"76",
          5456 => x"74",
          5457 => x"06",
          5458 => x"c8",
          5459 => x"71",
          5460 => x"ca",
          5461 => x"75",
          5462 => x"38",
          5463 => x"89",
          5464 => x"75",
          5465 => x"81",
          5466 => x"2e",
          5467 => x"7e",
          5468 => x"19",
          5469 => x"27",
          5470 => x"78",
          5471 => x"74",
          5472 => x"7a",
          5473 => x"80",
          5474 => x"27",
          5475 => x"54",
          5476 => x"51",
          5477 => x"08",
          5478 => x"98",
          5479 => x"87",
          5480 => x"31",
          5481 => x"94",
          5482 => x"0c",
          5483 => x"56",
          5484 => x"0d",
          5485 => x"3d",
          5486 => x"9c",
          5487 => x"c8",
          5488 => x"a8",
          5489 => x"a3",
          5490 => x"81",
          5491 => x"84",
          5492 => x"19",
          5493 => x"1a",
          5494 => x"7a",
          5495 => x"ec",
          5496 => x"38",
          5497 => x"56",
          5498 => x"31",
          5499 => x"79",
          5500 => x"57",
          5501 => x"38",
          5502 => x"70",
          5503 => x"75",
          5504 => x"81",
          5505 => x"5a",
          5506 => x"fe",
          5507 => x"51",
          5508 => x"08",
          5509 => x"51",
          5510 => x"08",
          5511 => x"74",
          5512 => x"9c",
          5513 => x"27",
          5514 => x"29",
          5515 => x"70",
          5516 => x"05",
          5517 => x"2e",
          5518 => x"57",
          5519 => x"ff",
          5520 => x"39",
          5521 => x"84",
          5522 => x"82",
          5523 => x"bb",
          5524 => x"3d",
          5525 => x"5c",
          5526 => x"80",
          5527 => x"80",
          5528 => x"80",
          5529 => x"1a",
          5530 => x"a8",
          5531 => x"76",
          5532 => x"74",
          5533 => x"81",
          5534 => x"76",
          5535 => x"08",
          5536 => x"84",
          5537 => x"82",
          5538 => x"7c",
          5539 => x"ff",
          5540 => x"7c",
          5541 => x"19",
          5542 => x"38",
          5543 => x"ff",
          5544 => x"0c",
          5545 => x"1a",
          5546 => x"98",
          5547 => x"f9",
          5548 => x"19",
          5549 => x"27",
          5550 => x"78",
          5551 => x"74",
          5552 => x"7b",
          5553 => x"81",
          5554 => x"27",
          5555 => x"54",
          5556 => x"51",
          5557 => x"08",
          5558 => x"31",
          5559 => x"80",
          5560 => x"05",
          5561 => x"57",
          5562 => x"ff",
          5563 => x"33",
          5564 => x"34",
          5565 => x"7f",
          5566 => x"1b",
          5567 => x"8c",
          5568 => x"74",
          5569 => x"8c",
          5570 => x"19",
          5571 => x"7a",
          5572 => x"bb",
          5573 => x"84",
          5574 => x"9c",
          5575 => x"19",
          5576 => x"9b",
          5577 => x"52",
          5578 => x"3f",
          5579 => x"94",
          5580 => x"76",
          5581 => x"59",
          5582 => x"58",
          5583 => x"56",
          5584 => x"70",
          5585 => x"05",
          5586 => x"38",
          5587 => x"79",
          5588 => x"19",
          5589 => x"3f",
          5590 => x"84",
          5591 => x"58",
          5592 => x"ff",
          5593 => x"55",
          5594 => x"e4",
          5595 => x"a8",
          5596 => x"98",
          5597 => x"38",
          5598 => x"75",
          5599 => x"39",
          5600 => x"3f",
          5601 => x"74",
          5602 => x"57",
          5603 => x"34",
          5604 => x"3d",
          5605 => x"82",
          5606 => x"0d",
          5607 => x"57",
          5608 => x"56",
          5609 => x"55",
          5610 => x"22",
          5611 => x"2e",
          5612 => x"76",
          5613 => x"33",
          5614 => x"7a",
          5615 => x"2b",
          5616 => x"7b",
          5617 => x"08",
          5618 => x"17",
          5619 => x"2e",
          5620 => x"54",
          5621 => x"33",
          5622 => x"84",
          5623 => x"81",
          5624 => x"78",
          5625 => x"11",
          5626 => x"18",
          5627 => x"83",
          5628 => x"9a",
          5629 => x"9b",
          5630 => x"19",
          5631 => x"c8",
          5632 => x"34",
          5633 => x"34",
          5634 => x"34",
          5635 => x"34",
          5636 => x"34",
          5637 => x"0b",
          5638 => x"34",
          5639 => x"81",
          5640 => x"98",
          5641 => x"19",
          5642 => x"90",
          5643 => x"84",
          5644 => x"b4",
          5645 => x"81",
          5646 => x"3f",
          5647 => x"2e",
          5648 => x"bb",
          5649 => x"08",
          5650 => x"08",
          5651 => x"fe",
          5652 => x"82",
          5653 => x"81",
          5654 => x"05",
          5655 => x"ff",
          5656 => x"39",
          5657 => x"34",
          5658 => x"34",
          5659 => x"74",
          5660 => x"74",
          5661 => x"74",
          5662 => x"80",
          5663 => x"a1",
          5664 => x"99",
          5665 => x"80",
          5666 => x"0b",
          5667 => x"be",
          5668 => x"33",
          5669 => x"19",
          5670 => x"51",
          5671 => x"08",
          5672 => x"74",
          5673 => x"81",
          5674 => x"52",
          5675 => x"93",
          5676 => x"08",
          5677 => x"ff",
          5678 => x"a0",
          5679 => x"77",
          5680 => x"fc",
          5681 => x"52",
          5682 => x"08",
          5683 => x"89",
          5684 => x"08",
          5685 => x"33",
          5686 => x"13",
          5687 => x"77",
          5688 => x"75",
          5689 => x"73",
          5690 => x"04",
          5691 => x"3f",
          5692 => x"72",
          5693 => x"d5",
          5694 => x"5b",
          5695 => x"75",
          5696 => x"26",
          5697 => x"70",
          5698 => x"84",
          5699 => x"90",
          5700 => x"0b",
          5701 => x"04",
          5702 => x"3d",
          5703 => x"81",
          5704 => x"26",
          5705 => x"06",
          5706 => x"80",
          5707 => x"5b",
          5708 => x"70",
          5709 => x"05",
          5710 => x"52",
          5711 => x"70",
          5712 => x"13",
          5713 => x"13",
          5714 => x"30",
          5715 => x"2e",
          5716 => x"be",
          5717 => x"72",
          5718 => x"52",
          5719 => x"84",
          5720 => x"99",
          5721 => x"83",
          5722 => x"fe",
          5723 => x"98",
          5724 => x"d2",
          5725 => x"84",
          5726 => x"74",
          5727 => x"04",
          5728 => x"05",
          5729 => x"08",
          5730 => x"38",
          5731 => x"2b",
          5732 => x"38",
          5733 => x"81",
          5734 => x"38",
          5735 => x"33",
          5736 => x"5a",
          5737 => x"38",
          5738 => x"84",
          5739 => x"84",
          5740 => x"8f",
          5741 => x"98",
          5742 => x"17",
          5743 => x"07",
          5744 => x"cc",
          5745 => x"74",
          5746 => x"04",
          5747 => x"08",
          5748 => x"7c",
          5749 => x"b4",
          5750 => x"84",
          5751 => x"bb",
          5752 => x"d9",
          5753 => x"80",
          5754 => x"08",
          5755 => x"38",
          5756 => x"a0",
          5757 => x"84",
          5758 => x"08",
          5759 => x"08",
          5760 => x"b1",
          5761 => x"33",
          5762 => x"54",
          5763 => x"33",
          5764 => x"84",
          5765 => x"81",
          5766 => x"d4",
          5767 => x"33",
          5768 => x"63",
          5769 => x"78",
          5770 => x"db",
          5771 => x"a4",
          5772 => x"84",
          5773 => x"52",
          5774 => x"bb",
          5775 => x"bb",
          5776 => x"33",
          5777 => x"63",
          5778 => x"7d",
          5779 => x"2e",
          5780 => x"7a",
          5781 => x"84",
          5782 => x"2e",
          5783 => x"d8",
          5784 => x"3d",
          5785 => x"be",
          5786 => x"5b",
          5787 => x"1f",
          5788 => x"5f",
          5789 => x"56",
          5790 => x"80",
          5791 => x"56",
          5792 => x"ff",
          5793 => x"75",
          5794 => x"18",
          5795 => x"af",
          5796 => x"79",
          5797 => x"8a",
          5798 => x"70",
          5799 => x"08",
          5800 => x"7e",
          5801 => x"17",
          5802 => x"38",
          5803 => x"38",
          5804 => x"76",
          5805 => x"05",
          5806 => x"26",
          5807 => x"5e",
          5808 => x"81",
          5809 => x"78",
          5810 => x"0d",
          5811 => x"71",
          5812 => x"07",
          5813 => x"16",
          5814 => x"71",
          5815 => x"3d",
          5816 => x"ff",
          5817 => x"59",
          5818 => x"96",
          5819 => x"16",
          5820 => x"17",
          5821 => x"81",
          5822 => x"38",
          5823 => x"b4",
          5824 => x"bb",
          5825 => x"08",
          5826 => x"55",
          5827 => x"f6",
          5828 => x"17",
          5829 => x"33",
          5830 => x"fb",
          5831 => x"08",
          5832 => x"0b",
          5833 => x"83",
          5834 => x"43",
          5835 => x"09",
          5836 => x"39",
          5837 => x"59",
          5838 => x"5e",
          5839 => x"80",
          5840 => x"5a",
          5841 => x"34",
          5842 => x"39",
          5843 => x"bb",
          5844 => x"f5",
          5845 => x"58",
          5846 => x"56",
          5847 => x"55",
          5848 => x"22",
          5849 => x"2e",
          5850 => x"77",
          5851 => x"33",
          5852 => x"08",
          5853 => x"94",
          5854 => x"2e",
          5855 => x"70",
          5856 => x"2e",
          5857 => x"51",
          5858 => x"08",
          5859 => x"55",
          5860 => x"08",
          5861 => x"76",
          5862 => x"31",
          5863 => x"80",
          5864 => x"80",
          5865 => x"08",
          5866 => x"70",
          5867 => x"7a",
          5868 => x"76",
          5869 => x"84",
          5870 => x"2e",
          5871 => x"38",
          5872 => x"55",
          5873 => x"38",
          5874 => x"84",
          5875 => x"19",
          5876 => x"58",
          5877 => x"17",
          5878 => x"58",
          5879 => x"18",
          5880 => x"05",
          5881 => x"7a",
          5882 => x"08",
          5883 => x"27",
          5884 => x"17",
          5885 => x"18",
          5886 => x"80",
          5887 => x"56",
          5888 => x"17",
          5889 => x"56",
          5890 => x"54",
          5891 => x"33",
          5892 => x"bb",
          5893 => x"80",
          5894 => x"81",
          5895 => x"11",
          5896 => x"84",
          5897 => x"38",
          5898 => x"74",
          5899 => x"04",
          5900 => x"06",
          5901 => x"94",
          5902 => x"7a",
          5903 => x"79",
          5904 => x"0b",
          5905 => x"75",
          5906 => x"18",
          5907 => x"fd",
          5908 => x"0b",
          5909 => x"04",
          5910 => x"3f",
          5911 => x"39",
          5912 => x"3f",
          5913 => x"74",
          5914 => x"58",
          5915 => x"ff",
          5916 => x"56",
          5917 => x"38",
          5918 => x"d8",
          5919 => x"0c",
          5920 => x"82",
          5921 => x"bb",
          5922 => x"3d",
          5923 => x"2e",
          5924 => x"05",
          5925 => x"8c",
          5926 => x"bb",
          5927 => x"76",
          5928 => x"0c",
          5929 => x"7d",
          5930 => x"84",
          5931 => x"08",
          5932 => x"98",
          5933 => x"38",
          5934 => x"06",
          5935 => x"38",
          5936 => x"12",
          5937 => x"33",
          5938 => x"2e",
          5939 => x"58",
          5940 => x"52",
          5941 => x"bb",
          5942 => x"38",
          5943 => x"76",
          5944 => x"76",
          5945 => x"94",
          5946 => x"2b",
          5947 => x"5a",
          5948 => x"55",
          5949 => x"74",
          5950 => x"72",
          5951 => x"86",
          5952 => x"71",
          5953 => x"57",
          5954 => x"84",
          5955 => x"81",
          5956 => x"84",
          5957 => x"dc",
          5958 => x"39",
          5959 => x"89",
          5960 => x"08",
          5961 => x"33",
          5962 => x"14",
          5963 => x"78",
          5964 => x"59",
          5965 => x"80",
          5966 => x"51",
          5967 => x"08",
          5968 => x"b5",
          5969 => x"76",
          5970 => x"72",
          5971 => x"84",
          5972 => x"70",
          5973 => x"08",
          5974 => x"84",
          5975 => x"53",
          5976 => x"72",
          5977 => x"84",
          5978 => x"70",
          5979 => x"08",
          5980 => x"52",
          5981 => x"bb",
          5982 => x"3d",
          5983 => x"fe",
          5984 => x"06",
          5985 => x"08",
          5986 => x"0d",
          5987 => x"53",
          5988 => x"84",
          5989 => x"08",
          5990 => x"84",
          5991 => x"75",
          5992 => x"84",
          5993 => x"38",
          5994 => x"2b",
          5995 => x"76",
          5996 => x"51",
          5997 => x"84",
          5998 => x"84",
          5999 => x"ed",
          6000 => x"53",
          6001 => x"51",
          6002 => x"5a",
          6003 => x"75",
          6004 => x"11",
          6005 => x"75",
          6006 => x"79",
          6007 => x"04",
          6008 => x"5b",
          6009 => x"a8",
          6010 => x"5d",
          6011 => x"1d",
          6012 => x"76",
          6013 => x"78",
          6014 => x"54",
          6015 => x"33",
          6016 => x"84",
          6017 => x"81",
          6018 => x"5b",
          6019 => x"5e",
          6020 => x"17",
          6021 => x"33",
          6022 => x"81",
          6023 => x"75",
          6024 => x"06",
          6025 => x"05",
          6026 => x"ff",
          6027 => x"53",
          6028 => x"38",
          6029 => x"84",
          6030 => x"18",
          6031 => x"3d",
          6032 => x"53",
          6033 => x"52",
          6034 => x"84",
          6035 => x"bb",
          6036 => x"08",
          6037 => x"08",
          6038 => x"fe",
          6039 => x"82",
          6040 => x"81",
          6041 => x"05",
          6042 => x"fe",
          6043 => x"39",
          6044 => x"75",
          6045 => x"84",
          6046 => x"38",
          6047 => x"f7",
          6048 => x"84",
          6049 => x"05",
          6050 => x"9c",
          6051 => x"7f",
          6052 => x"33",
          6053 => x"fe",
          6054 => x"11",
          6055 => x"70",
          6056 => x"83",
          6057 => x"59",
          6058 => x"fe",
          6059 => x"81",
          6060 => x"94",
          6061 => x"58",
          6062 => x"82",
          6063 => x"0d",
          6064 => x"9f",
          6065 => x"97",
          6066 => x"8f",
          6067 => x"5a",
          6068 => x"80",
          6069 => x"91",
          6070 => x"90",
          6071 => x"56",
          6072 => x"eb",
          6073 => x"19",
          6074 => x"fb",
          6075 => x"55",
          6076 => x"08",
          6077 => x"80",
          6078 => x"8c",
          6079 => x"74",
          6080 => x"98",
          6081 => x"81",
          6082 => x"52",
          6083 => x"fa",
          6084 => x"2e",
          6085 => x"19",
          6086 => x"0c",
          6087 => x"79",
          6088 => x"51",
          6089 => x"08",
          6090 => x"80",
          6091 => x"2e",
          6092 => x"ff",
          6093 => x"52",
          6094 => x"bb",
          6095 => x"08",
          6096 => x"59",
          6097 => x"16",
          6098 => x"07",
          6099 => x"78",
          6100 => x"81",
          6101 => x"84",
          6102 => x"fd",
          6103 => x"fd",
          6104 => x"5a",
          6105 => x"0c",
          6106 => x"77",
          6107 => x"84",
          6108 => x"bb",
          6109 => x"76",
          6110 => x"84",
          6111 => x"38",
          6112 => x"79",
          6113 => x"bb",
          6114 => x"bb",
          6115 => x"96",
          6116 => x"53",
          6117 => x"3f",
          6118 => x"84",
          6119 => x"51",
          6120 => x"08",
          6121 => x"80",
          6122 => x"2e",
          6123 => x"ff",
          6124 => x"52",
          6125 => x"bb",
          6126 => x"08",
          6127 => x"59",
          6128 => x"94",
          6129 => x"55",
          6130 => x"7a",
          6131 => x"57",
          6132 => x"81",
          6133 => x"19",
          6134 => x"57",
          6135 => x"06",
          6136 => x"fc",
          6137 => x"5a",
          6138 => x"08",
          6139 => x"39",
          6140 => x"fd",
          6141 => x"ff",
          6142 => x"db",
          6143 => x"9c",
          6144 => x"b4",
          6145 => x"bb",
          6146 => x"84",
          6147 => x"7d",
          6148 => x"70",
          6149 => x"bb",
          6150 => x"de",
          6151 => x"85",
          6152 => x"77",
          6153 => x"7b",
          6154 => x"33",
          6155 => x"7b",
          6156 => x"9b",
          6157 => x"2b",
          6158 => x"58",
          6159 => x"84",
          6160 => x"80",
          6161 => x"7b",
          6162 => x"41",
          6163 => x"70",
          6164 => x"bb",
          6165 => x"fe",
          6166 => x"74",
          6167 => x"84",
          6168 => x"38",
          6169 => x"3d",
          6170 => x"33",
          6171 => x"7d",
          6172 => x"84",
          6173 => x"84",
          6174 => x"08",
          6175 => x"74",
          6176 => x"78",
          6177 => x"84",
          6178 => x"2e",
          6179 => x"80",
          6180 => x"38",
          6181 => x"08",
          6182 => x"9c",
          6183 => x"82",
          6184 => x"fe",
          6185 => x"84",
          6186 => x"b8",
          6187 => x"5a",
          6188 => x"38",
          6189 => x"7a",
          6190 => x"81",
          6191 => x"17",
          6192 => x"bb",
          6193 => x"56",
          6194 => x"56",
          6195 => x"e5",
          6196 => x"90",
          6197 => x"80",
          6198 => x"84",
          6199 => x"08",
          6200 => x"2e",
          6201 => x"56",
          6202 => x"08",
          6203 => x"fe",
          6204 => x"84",
          6205 => x"a6",
          6206 => x"34",
          6207 => x"84",
          6208 => x"18",
          6209 => x"33",
          6210 => x"fe",
          6211 => x"a0",
          6212 => x"17",
          6213 => x"58",
          6214 => x"27",
          6215 => x"fe",
          6216 => x"5a",
          6217 => x"cb",
          6218 => x"fd",
          6219 => x"2e",
          6220 => x"76",
          6221 => x"84",
          6222 => x"11",
          6223 => x"7b",
          6224 => x"18",
          6225 => x"7b",
          6226 => x"26",
          6227 => x"39",
          6228 => x"84",
          6229 => x"fd",
          6230 => x"9f",
          6231 => x"51",
          6232 => x"08",
          6233 => x"8a",
          6234 => x"3d",
          6235 => x"3d",
          6236 => x"84",
          6237 => x"08",
          6238 => x"0c",
          6239 => x"08",
          6240 => x"02",
          6241 => x"81",
          6242 => x"b9",
          6243 => x"70",
          6244 => x"bb",
          6245 => x"84",
          6246 => x"84",
          6247 => x"bb",
          6248 => x"75",
          6249 => x"08",
          6250 => x"80",
          6251 => x"fe",
          6252 => x"27",
          6253 => x"29",
          6254 => x"b4",
          6255 => x"79",
          6256 => x"58",
          6257 => x"74",
          6258 => x"27",
          6259 => x"53",
          6260 => x"ef",
          6261 => x"df",
          6262 => x"56",
          6263 => x"08",
          6264 => x"33",
          6265 => x"56",
          6266 => x"bb",
          6267 => x"08",
          6268 => x"18",
          6269 => x"33",
          6270 => x"fe",
          6271 => x"a0",
          6272 => x"17",
          6273 => x"ca",
          6274 => x"55",
          6275 => x"9c",
          6276 => x"52",
          6277 => x"bb",
          6278 => x"80",
          6279 => x"08",
          6280 => x"84",
          6281 => x"53",
          6282 => x"3f",
          6283 => x"9c",
          6284 => x"5a",
          6285 => x"81",
          6286 => x"81",
          6287 => x"55",
          6288 => x"84",
          6289 => x"8a",
          6290 => x"06",
          6291 => x"81",
          6292 => x"1f",
          6293 => x"57",
          6294 => x"7d",
          6295 => x"58",
          6296 => x"59",
          6297 => x"cf",
          6298 => x"34",
          6299 => x"7d",
          6300 => x"77",
          6301 => x"5b",
          6302 => x"55",
          6303 => x"59",
          6304 => x"57",
          6305 => x"33",
          6306 => x"16",
          6307 => x"0b",
          6308 => x"83",
          6309 => x"80",
          6310 => x"7a",
          6311 => x"74",
          6312 => x"81",
          6313 => x"92",
          6314 => x"84",
          6315 => x"56",
          6316 => x"84",
          6317 => x"0b",
          6318 => x"17",
          6319 => x"18",
          6320 => x"18",
          6321 => x"80",
          6322 => x"16",
          6323 => x"34",
          6324 => x"bb",
          6325 => x"0c",
          6326 => x"55",
          6327 => x"2a",
          6328 => x"fd",
          6329 => x"cc",
          6330 => x"80",
          6331 => x"80",
          6332 => x"fe",
          6333 => x"94",
          6334 => x"95",
          6335 => x"16",
          6336 => x"34",
          6337 => x"bb",
          6338 => x"3d",
          6339 => x"59",
          6340 => x"79",
          6341 => x"26",
          6342 => x"38",
          6343 => x"af",
          6344 => x"05",
          6345 => x"3f",
          6346 => x"84",
          6347 => x"bb",
          6348 => x"a6",
          6349 => x"3d",
          6350 => x"84",
          6351 => x"08",
          6352 => x"81",
          6353 => x"38",
          6354 => x"58",
          6355 => x"33",
          6356 => x"15",
          6357 => x"b0",
          6358 => x"81",
          6359 => x"59",
          6360 => x"b3",
          6361 => x"8e",
          6362 => x"bb",
          6363 => x"3d",
          6364 => x"84",
          6365 => x"76",
          6366 => x"57",
          6367 => x"82",
          6368 => x"5d",
          6369 => x"80",
          6370 => x"72",
          6371 => x"81",
          6372 => x"5b",
          6373 => x"77",
          6374 => x"81",
          6375 => x"58",
          6376 => x"70",
          6377 => x"70",
          6378 => x"09",
          6379 => x"38",
          6380 => x"07",
          6381 => x"7a",
          6382 => x"1e",
          6383 => x"38",
          6384 => x"39",
          6385 => x"7f",
          6386 => x"05",
          6387 => x"3f",
          6388 => x"84",
          6389 => x"6c",
          6390 => x"fe",
          6391 => x"3f",
          6392 => x"84",
          6393 => x"0b",
          6394 => x"05",
          6395 => x"57",
          6396 => x"ff",
          6397 => x"cb",
          6398 => x"33",
          6399 => x"7e",
          6400 => x"8b",
          6401 => x"1e",
          6402 => x"81",
          6403 => x"c5",
          6404 => x"bd",
          6405 => x"33",
          6406 => x"58",
          6407 => x"38",
          6408 => x"5e",
          6409 => x"8a",
          6410 => x"08",
          6411 => x"b5",
          6412 => x"08",
          6413 => x"5f",
          6414 => x"53",
          6415 => x"fe",
          6416 => x"80",
          6417 => x"77",
          6418 => x"d8",
          6419 => x"81",
          6420 => x"81",
          6421 => x"ff",
          6422 => x"34",
          6423 => x"18",
          6424 => x"09",
          6425 => x"5e",
          6426 => x"2a",
          6427 => x"57",
          6428 => x"aa",
          6429 => x"56",
          6430 => x"78",
          6431 => x"84",
          6432 => x"f5",
          6433 => x"57",
          6434 => x"b4",
          6435 => x"7e",
          6436 => x"38",
          6437 => x"81",
          6438 => x"84",
          6439 => x"ff",
          6440 => x"77",
          6441 => x"5a",
          6442 => x"34",
          6443 => x"80",
          6444 => x"84",
          6445 => x"08",
          6446 => x"74",
          6447 => x"74",
          6448 => x"d6",
          6449 => x"84",
          6450 => x"84",
          6451 => x"95",
          6452 => x"2b",
          6453 => x"56",
          6454 => x"08",
          6455 => x"84",
          6456 => x"84",
          6457 => x"81",
          6458 => x"81",
          6459 => x"81",
          6460 => x"09",
          6461 => x"84",
          6462 => x"a8",
          6463 => x"59",
          6464 => x"a0",
          6465 => x"2e",
          6466 => x"54",
          6467 => x"53",
          6468 => x"e2",
          6469 => x"81",
          6470 => x"70",
          6471 => x"e1",
          6472 => x"08",
          6473 => x"83",
          6474 => x"08",
          6475 => x"74",
          6476 => x"82",
          6477 => x"81",
          6478 => x"17",
          6479 => x"52",
          6480 => x"3f",
          6481 => x"0d",
          6482 => x"05",
          6483 => x"53",
          6484 => x"51",
          6485 => x"08",
          6486 => x"8a",
          6487 => x"3d",
          6488 => x"3d",
          6489 => x"84",
          6490 => x"08",
          6491 => x"81",
          6492 => x"38",
          6493 => x"12",
          6494 => x"51",
          6495 => x"78",
          6496 => x"51",
          6497 => x"08",
          6498 => x"04",
          6499 => x"96",
          6500 => x"ff",
          6501 => x"55",
          6502 => x"38",
          6503 => x"0d",
          6504 => x"d0",
          6505 => x"bb",
          6506 => x"e0",
          6507 => x"a0",
          6508 => x"60",
          6509 => x"90",
          6510 => x"17",
          6511 => x"17",
          6512 => x"17",
          6513 => x"17",
          6514 => x"34",
          6515 => x"bb",
          6516 => x"3d",
          6517 => x"5d",
          6518 => x"52",
          6519 => x"84",
          6520 => x"30",
          6521 => x"25",
          6522 => x"38",
          6523 => x"81",
          6524 => x"80",
          6525 => x"8c",
          6526 => x"78",
          6527 => x"11",
          6528 => x"08",
          6529 => x"33",
          6530 => x"81",
          6531 => x"53",
          6532 => x"fe",
          6533 => x"80",
          6534 => x"76",
          6535 => x"38",
          6536 => x"56",
          6537 => x"56",
          6538 => x"75",
          6539 => x"12",
          6540 => x"07",
          6541 => x"2b",
          6542 => x"5d",
          6543 => x"84",
          6544 => x"80",
          6545 => x"55",
          6546 => x"08",
          6547 => x"81",
          6548 => x"06",
          6549 => x"57",
          6550 => x"08",
          6551 => x"33",
          6552 => x"59",
          6553 => x"81",
          6554 => x"08",
          6555 => x"17",
          6556 => x"55",
          6557 => x"38",
          6558 => x"09",
          6559 => x"b4",
          6560 => x"7a",
          6561 => x"9b",
          6562 => x"b8",
          6563 => x"db",
          6564 => x"2e",
          6565 => x"52",
          6566 => x"bb",
          6567 => x"fe",
          6568 => x"bb",
          6569 => x"18",
          6570 => x"75",
          6571 => x"78",
          6572 => x"58",
          6573 => x"f2",
          6574 => x"5c",
          6575 => x"fc",
          6576 => x"e1",
          6577 => x"b4",
          6578 => x"a4",
          6579 => x"bb",
          6580 => x"5d",
          6581 => x"81",
          6582 => x"f4",
          6583 => x"70",
          6584 => x"9f",
          6585 => x"90",
          6586 => x"81",
          6587 => x"75",
          6588 => x"81",
          6589 => x"83",
          6590 => x"9f",
          6591 => x"ff",
          6592 => x"e0",
          6593 => x"94",
          6594 => x"58",
          6595 => x"56",
          6596 => x"70",
          6597 => x"58",
          6598 => x"2e",
          6599 => x"ff",
          6600 => x"ff",
          6601 => x"26",
          6602 => x"8f",
          6603 => x"70",
          6604 => x"76",
          6605 => x"1a",
          6606 => x"ff",
          6607 => x"26",
          6608 => x"86",
          6609 => x"79",
          6610 => x"56",
          6611 => x"a0",
          6612 => x"1a",
          6613 => x"47",
          6614 => x"fe",
          6615 => x"55",
          6616 => x"38",
          6617 => x"a1",
          6618 => x"51",
          6619 => x"83",
          6620 => x"38",
          6621 => x"a1",
          6622 => x"56",
          6623 => x"fe",
          6624 => x"55",
          6625 => x"79",
          6626 => x"7e",
          6627 => x"58",
          6628 => x"ff",
          6629 => x"81",
          6630 => x"da",
          6631 => x"74",
          6632 => x"fe",
          6633 => x"84",
          6634 => x"06",
          6635 => x"2e",
          6636 => x"76",
          6637 => x"bb",
          6638 => x"75",
          6639 => x"84",
          6640 => x"98",
          6641 => x"08",
          6642 => x"55",
          6643 => x"d7",
          6644 => x"52",
          6645 => x"3f",
          6646 => x"38",
          6647 => x"0c",
          6648 => x"17",
          6649 => x"81",
          6650 => x"70",
          6651 => x"80",
          6652 => x"79",
          6653 => x"51",
          6654 => x"08",
          6655 => x"ff",
          6656 => x"fd",
          6657 => x"38",
          6658 => x"81",
          6659 => x"f4",
          6660 => x"34",
          6661 => x"70",
          6662 => x"05",
          6663 => x"2e",
          6664 => x"58",
          6665 => x"ff",
          6666 => x"39",
          6667 => x"81",
          6668 => x"d7",
          6669 => x"fd",
          6670 => x"81",
          6671 => x"81",
          6672 => x"84",
          6673 => x"06",
          6674 => x"83",
          6675 => x"08",
          6676 => x"8a",
          6677 => x"2e",
          6678 => x"fd",
          6679 => x"51",
          6680 => x"08",
          6681 => x"fd",
          6682 => x"58",
          6683 => x"fe",
          6684 => x"a0",
          6685 => x"18",
          6686 => x"a9",
          6687 => x"88",
          6688 => x"57",
          6689 => x"76",
          6690 => x"74",
          6691 => x"86",
          6692 => x"78",
          6693 => x"73",
          6694 => x"33",
          6695 => x"2e",
          6696 => x"9c",
          6697 => x"81",
          6698 => x"8c",
          6699 => x"2b",
          6700 => x"fd",
          6701 => x"70",
          6702 => x"bb",
          6703 => x"42",
          6704 => x"88",
          6705 => x"38",
          6706 => x"59",
          6707 => x"3f",
          6708 => x"08",
          6709 => x"bb",
          6710 => x"84",
          6711 => x"38",
          6712 => x"81",
          6713 => x"74",
          6714 => x"87",
          6715 => x"0c",
          6716 => x"bb",
          6717 => x"15",
          6718 => x"bb",
          6719 => x"ad",
          6720 => x"a7",
          6721 => x"7a",
          6722 => x"38",
          6723 => x"e6",
          6724 => x"fe",
          6725 => x"56",
          6726 => x"77",
          6727 => x"74",
          6728 => x"55",
          6729 => x"88",
          6730 => x"17",
          6731 => x"18",
          6732 => x"16",
          6733 => x"e9",
          6734 => x"84",
          6735 => x"16",
          6736 => x"54",
          6737 => x"fe",
          6738 => x"81",
          6739 => x"ff",
          6740 => x"3d",
          6741 => x"02",
          6742 => x"42",
          6743 => x"5f",
          6744 => x"38",
          6745 => x"9f",
          6746 => x"9b",
          6747 => x"85",
          6748 => x"80",
          6749 => x"10",
          6750 => x"5a",
          6751 => x"34",
          6752 => x"84",
          6753 => x"81",
          6754 => x"84",
          6755 => x"81",
          6756 => x"ab",
          6757 => x"8a",
          6758 => x"fc",
          6759 => x"d0",
          6760 => x"98",
          6761 => x"90",
          6762 => x"88",
          6763 => x"83",
          6764 => x"84",
          6765 => x"81",
          6766 => x"1f",
          6767 => x"7e",
          6768 => x"70",
          6769 => x"60",
          6770 => x"70",
          6771 => x"57",
          6772 => x"84",
          6773 => x"52",
          6774 => x"57",
          6775 => x"60",
          6776 => x"05",
          6777 => x"8e",
          6778 => x"81",
          6779 => x"61",
          6780 => x"62",
          6781 => x"18",
          6782 => x"90",
          6783 => x"33",
          6784 => x"71",
          6785 => x"82",
          6786 => x"2b",
          6787 => x"88",
          6788 => x"3d",
          6789 => x"0c",
          6790 => x"5a",
          6791 => x"79",
          6792 => x"81",
          6793 => x"2a",
          6794 => x"2e",
          6795 => x"64",
          6796 => x"47",
          6797 => x"30",
          6798 => x"2e",
          6799 => x"8c",
          6800 => x"22",
          6801 => x"74",
          6802 => x"56",
          6803 => x"57",
          6804 => x"75",
          6805 => x"fc",
          6806 => x"10",
          6807 => x"9f",
          6808 => x"bb",
          6809 => x"05",
          6810 => x"4c",
          6811 => x"81",
          6812 => x"68",
          6813 => x"06",
          6814 => x"83",
          6815 => x"77",
          6816 => x"57",
          6817 => x"7c",
          6818 => x"31",
          6819 => x"bb",
          6820 => x"f6",
          6821 => x"82",
          6822 => x"bb",
          6823 => x"89",
          6824 => x"c0",
          6825 => x"a3",
          6826 => x"0c",
          6827 => x"04",
          6828 => x"84",
          6829 => x"bb",
          6830 => x"70",
          6831 => x"89",
          6832 => x"ff",
          6833 => x"2e",
          6834 => x"f4",
          6835 => x"7a",
          6836 => x"81",
          6837 => x"59",
          6838 => x"17",
          6839 => x"9f",
          6840 => x"e0",
          6841 => x"76",
          6842 => x"78",
          6843 => x"ff",
          6844 => x"70",
          6845 => x"4a",
          6846 => x"81",
          6847 => x"25",
          6848 => x"39",
          6849 => x"79",
          6850 => x"84",
          6851 => x"83",
          6852 => x"40",
          6853 => x"55",
          6854 => x"38",
          6855 => x"81",
          6856 => x"ff",
          6857 => x"56",
          6858 => x"93",
          6859 => x"82",
          6860 => x"8b",
          6861 => x"26",
          6862 => x"5b",
          6863 => x"8e",
          6864 => x"3d",
          6865 => x"55",
          6866 => x"f5",
          6867 => x"5b",
          6868 => x"80",
          6869 => x"05",
          6870 => x"38",
          6871 => x"55",
          6872 => x"70",
          6873 => x"74",
          6874 => x"65",
          6875 => x"61",
          6876 => x"06",
          6877 => x"88",
          6878 => x"81",
          6879 => x"70",
          6880 => x"34",
          6881 => x"61",
          6882 => x"ff",
          6883 => x"ff",
          6884 => x"34",
          6885 => x"05",
          6886 => x"61",
          6887 => x"34",
          6888 => x"9b",
          6889 => x"7e",
          6890 => x"34",
          6891 => x"05",
          6892 => x"0c",
          6893 => x"34",
          6894 => x"61",
          6895 => x"34",
          6896 => x"61",
          6897 => x"06",
          6898 => x"88",
          6899 => x"ff",
          6900 => x"a6",
          6901 => x"e6",
          6902 => x"05",
          6903 => x"34",
          6904 => x"83",
          6905 => x"60",
          6906 => x"34",
          6907 => x"51",
          6908 => x"bb",
          6909 => x"5c",
          6910 => x"61",
          6911 => x"58",
          6912 => x"63",
          6913 => x"c0",
          6914 => x"81",
          6915 => x"34",
          6916 => x"64",
          6917 => x"2a",
          6918 => x"34",
          6919 => x"7c",
          6920 => x"38",
          6921 => x"52",
          6922 => x"bb",
          6923 => x"61",
          6924 => x"58",
          6925 => x"78",
          6926 => x"c9",
          6927 => x"2e",
          6928 => x"2e",
          6929 => x"66",
          6930 => x"7a",
          6931 => x"8b",
          6932 => x"38",
          6933 => x"75",
          6934 => x"93",
          6935 => x"26",
          6936 => x"83",
          6937 => x"61",
          6938 => x"b3",
          6939 => x"75",
          6940 => x"59",
          6941 => x"ff",
          6942 => x"47",
          6943 => x"34",
          6944 => x"83",
          6945 => x"6c",
          6946 => x"51",
          6947 => x"05",
          6948 => x"bf",
          6949 => x"84",
          6950 => x"7e",
          6951 => x"83",
          6952 => x"05",
          6953 => x"c9",
          6954 => x"34",
          6955 => x"cb",
          6956 => x"61",
          6957 => x"5f",
          6958 => x"54",
          6959 => x"c3",
          6960 => x"08",
          6961 => x"79",
          6962 => x"84",
          6963 => x"bb",
          6964 => x"3d",
          6965 => x"55",
          6966 => x"45",
          6967 => x"78",
          6968 => x"b8",
          6969 => x"38",
          6970 => x"b8",
          6971 => x"57",
          6972 => x"76",
          6973 => x"51",
          6974 => x"08",
          6975 => x"2a",
          6976 => x"bb",
          6977 => x"47",
          6978 => x"cb",
          6979 => x"bb",
          6980 => x"e6",
          6981 => x"2a",
          6982 => x"f8",
          6983 => x"80",
          6984 => x"ab",
          6985 => x"88",
          6986 => x"75",
          6987 => x"34",
          6988 => x"05",
          6989 => x"c3",
          6990 => x"34",
          6991 => x"cc",
          6992 => x"a4",
          6993 => x"61",
          6994 => x"78",
          6995 => x"56",
          6996 => x"ac",
          6997 => x"80",
          6998 => x"05",
          6999 => x"61",
          7000 => x"34",
          7001 => x"61",
          7002 => x"c2",
          7003 => x"83",
          7004 => x"81",
          7005 => x"58",
          7006 => x"f9",
          7007 => x"33",
          7008 => x"15",
          7009 => x"81",
          7010 => x"fe",
          7011 => x"84",
          7012 => x"61",
          7013 => x"34",
          7014 => x"60",
          7015 => x"fc",
          7016 => x"0c",
          7017 => x"04",
          7018 => x"70",
          7019 => x"81",
          7020 => x"61",
          7021 => x"34",
          7022 => x"87",
          7023 => x"ff",
          7024 => x"05",
          7025 => x"b1",
          7026 => x"52",
          7027 => x"80",
          7028 => x"05",
          7029 => x"38",
          7030 => x"05",
          7031 => x"70",
          7032 => x"70",
          7033 => x"34",
          7034 => x"80",
          7035 => x"c1",
          7036 => x"61",
          7037 => x"5b",
          7038 => x"88",
          7039 => x"34",
          7040 => x"ea",
          7041 => x"61",
          7042 => x"ec",
          7043 => x"34",
          7044 => x"61",
          7045 => x"34",
          7046 => x"1f",
          7047 => x"eb",
          7048 => x"52",
          7049 => x"61",
          7050 => x"0d",
          7051 => x"ff",
          7052 => x"b8",
          7053 => x"05",
          7054 => x"ff",
          7055 => x"81",
          7056 => x"74",
          7057 => x"81",
          7058 => x"8a",
          7059 => x"38",
          7060 => x"38",
          7061 => x"8e",
          7062 => x"02",
          7063 => x"77",
          7064 => x"08",
          7065 => x"17",
          7066 => x"77",
          7067 => x"24",
          7068 => x"19",
          7069 => x"8b",
          7070 => x"17",
          7071 => x"3f",
          7072 => x"07",
          7073 => x"81",
          7074 => x"d3",
          7075 => x"3f",
          7076 => x"80",
          7077 => x"80",
          7078 => x"81",
          7079 => x"f4",
          7080 => x"8a",
          7081 => x"76",
          7082 => x"8c",
          7083 => x"16",
          7084 => x"84",
          7085 => x"7c",
          7086 => x"3d",
          7087 => x"05",
          7088 => x"3f",
          7089 => x"7a",
          7090 => x"84",
          7091 => x"ff",
          7092 => x"52",
          7093 => x"74",
          7094 => x"9f",
          7095 => x"ff",
          7096 => x"eb",
          7097 => x"84",
          7098 => x"0d",
          7099 => x"52",
          7100 => x"90",
          7101 => x"71",
          7102 => x"04",
          7103 => x"83",
          7104 => x"73",
          7105 => x"22",
          7106 => x"12",
          7107 => x"71",
          7108 => x"83",
          7109 => x"e1",
          7110 => x"06",
          7111 => x"0d",
          7112 => x"22",
          7113 => x"51",
          7114 => x"38",
          7115 => x"84",
          7116 => x"09",
          7117 => x"26",
          7118 => x"05",
          7119 => x"84",
          7120 => x"51",
          7121 => x"38",
          7122 => x"c8",
          7123 => x"d9",
          7124 => x"75",
          7125 => x"26",
          7126 => x"38",
          7127 => x"71",
          7128 => x"70",
          7129 => x"38",
          7130 => x"70",
          7131 => x"70",
          7132 => x"55",
          7133 => x"51",
          7134 => x"0d",
          7135 => x"39",
          7136 => x"10",
          7137 => x"04",
          7138 => x"06",
          7139 => x"b0",
          7140 => x"51",
          7141 => x"ff",
          7142 => x"70",
          7143 => x"39",
          7144 => x"57",
          7145 => x"ff",
          7146 => x"16",
          7147 => x"ff",
          7148 => x"76",
          7149 => x"58",
          7150 => x"31",
          7151 => x"fe",
          7152 => x"ff",
          7153 => x"00",
          7154 => x"19",
          7155 => x"19",
          7156 => x"19",
          7157 => x"19",
          7158 => x"19",
          7159 => x"19",
          7160 => x"19",
          7161 => x"18",
          7162 => x"18",
          7163 => x"18",
          7164 => x"1e",
          7165 => x"1f",
          7166 => x"1f",
          7167 => x"1f",
          7168 => x"1f",
          7169 => x"1f",
          7170 => x"1f",
          7171 => x"1f",
          7172 => x"1f",
          7173 => x"1f",
          7174 => x"1f",
          7175 => x"1f",
          7176 => x"1f",
          7177 => x"1f",
          7178 => x"1f",
          7179 => x"1f",
          7180 => x"1f",
          7181 => x"1f",
          7182 => x"1f",
          7183 => x"1f",
          7184 => x"1f",
          7185 => x"1f",
          7186 => x"1f",
          7187 => x"1f",
          7188 => x"1f",
          7189 => x"1f",
          7190 => x"1f",
          7191 => x"1f",
          7192 => x"1f",
          7193 => x"1f",
          7194 => x"24",
          7195 => x"1f",
          7196 => x"24",
          7197 => x"22",
          7198 => x"1f",
          7199 => x"1f",
          7200 => x"1f",
          7201 => x"1f",
          7202 => x"1f",
          7203 => x"1f",
          7204 => x"1f",
          7205 => x"1f",
          7206 => x"1f",
          7207 => x"1f",
          7208 => x"1f",
          7209 => x"1f",
          7210 => x"1f",
          7211 => x"1f",
          7212 => x"1f",
          7213 => x"1f",
          7214 => x"1f",
          7215 => x"1f",
          7216 => x"1f",
          7217 => x"1f",
          7218 => x"1f",
          7219 => x"1f",
          7220 => x"1f",
          7221 => x"1f",
          7222 => x"1f",
          7223 => x"1f",
          7224 => x"21",
          7225 => x"1f",
          7226 => x"1f",
          7227 => x"1f",
          7228 => x"1f",
          7229 => x"21",
          7230 => x"1f",
          7231 => x"1f",
          7232 => x"21",
          7233 => x"32",
          7234 => x"32",
          7235 => x"32",
          7236 => x"3c",
          7237 => x"39",
          7238 => x"3b",
          7239 => x"37",
          7240 => x"3a",
          7241 => x"37",
          7242 => x"34",
          7243 => x"38",
          7244 => x"34",
          7245 => x"37",
          7246 => x"36",
          7247 => x"47",
          7248 => x"47",
          7249 => x"47",
          7250 => x"47",
          7251 => x"48",
          7252 => x"48",
          7253 => x"48",
          7254 => x"48",
          7255 => x"48",
          7256 => x"48",
          7257 => x"48",
          7258 => x"48",
          7259 => x"48",
          7260 => x"48",
          7261 => x"48",
          7262 => x"48",
          7263 => x"48",
          7264 => x"48",
          7265 => x"48",
          7266 => x"49",
          7267 => x"49",
          7268 => x"48",
          7269 => x"48",
          7270 => x"48",
          7271 => x"49",
          7272 => x"48",
          7273 => x"48",
          7274 => x"48",
          7275 => x"48",
          7276 => x"56",
          7277 => x"55",
          7278 => x"55",
          7279 => x"56",
          7280 => x"56",
          7281 => x"53",
          7282 => x"53",
          7283 => x"53",
          7284 => x"56",
          7285 => x"57",
          7286 => x"53",
          7287 => x"53",
          7288 => x"53",
          7289 => x"53",
          7290 => x"53",
          7291 => x"53",
          7292 => x"53",
          7293 => x"53",
          7294 => x"53",
          7295 => x"55",
          7296 => x"53",
          7297 => x"55",
          7298 => x"54",
          7299 => x"53",
          7300 => x"53",
          7301 => x"53",
          7302 => x"5a",
          7303 => x"59",
          7304 => x"59",
          7305 => x"59",
          7306 => x"59",
          7307 => x"59",
          7308 => x"59",
          7309 => x"59",
          7310 => x"59",
          7311 => x"59",
          7312 => x"59",
          7313 => x"59",
          7314 => x"59",
          7315 => x"59",
          7316 => x"59",
          7317 => x"5a",
          7318 => x"5a",
          7319 => x"5a",
          7320 => x"5b",
          7321 => x"59",
          7322 => x"5b",
          7323 => x"5a",
          7324 => x"5a",
          7325 => x"5a",
          7326 => x"59",
          7327 => x"64",
          7328 => x"62",
          7329 => x"62",
          7330 => x"62",
          7331 => x"62",
          7332 => x"62",
          7333 => x"62",
          7334 => x"5f",
          7335 => x"62",
          7336 => x"62",
          7337 => x"62",
          7338 => x"62",
          7339 => x"64",
          7340 => x"64",
          7341 => x"64",
          7342 => x"df",
          7343 => x"df",
          7344 => x"df",
          7345 => x"df",
          7346 => x"0e",
          7347 => x"0b",
          7348 => x"0b",
          7349 => x"0b",
          7350 => x"0b",
          7351 => x"0b",
          7352 => x"0b",
          7353 => x"0f",
          7354 => x"0b",
          7355 => x"0b",
          7356 => x"0b",
          7357 => x"0b",
          7358 => x"0b",
          7359 => x"0b",
          7360 => x"0b",
          7361 => x"0b",
          7362 => x"0b",
          7363 => x"0b",
          7364 => x"0b",
          7365 => x"0b",
          7366 => x"0b",
          7367 => x"0b",
          7368 => x"0b",
          7369 => x"0b",
          7370 => x"0b",
          7371 => x"0b",
          7372 => x"0b",
          7373 => x"0b",
          7374 => x"0e",
          7375 => x"0b",
          7376 => x"0b",
          7377 => x"0b",
          7378 => x"0b",
          7379 => x"0b",
          7380 => x"0e",
          7381 => x"0e",
          7382 => x"0b",
          7383 => x"0b",
          7384 => x"0e",
          7385 => x"0b",
          7386 => x"0e",
          7387 => x"0b",
          7388 => x"0b",
          7389 => x"0b",
          7390 => x"0e",
          7391 => x"00",
          7392 => x"00",
          7393 => x"00",
          7394 => x"00",
          7395 => x"00",
          7396 => x"00",
          7397 => x"00",
          7398 => x"00",
          7399 => x"00",
          7400 => x"68",
          7401 => x"64",
          7402 => x"64",
          7403 => x"6c",
          7404 => x"70",
          7405 => x"74",
          7406 => x"00",
          7407 => x"00",
          7408 => x"00",
          7409 => x"30",
          7410 => x"00",
          7411 => x"00",
          7412 => x"00",
          7413 => x"6b",
          7414 => x"72",
          7415 => x"72",
          7416 => x"20",
          7417 => x"63",
          7418 => x"6f",
          7419 => x"70",
          7420 => x"73",
          7421 => x"73",
          7422 => x"6e",
          7423 => x"79",
          7424 => x"6c",
          7425 => x"63",
          7426 => x"6d",
          7427 => x"70",
          7428 => x"20",
          7429 => x"65",
          7430 => x"72",
          7431 => x"72",
          7432 => x"20",
          7433 => x"62",
          7434 => x"73",
          7435 => x"6f",
          7436 => x"64",
          7437 => x"73",
          7438 => x"6e",
          7439 => x"00",
          7440 => x"6e",
          7441 => x"73",
          7442 => x"64",
          7443 => x"20",
          7444 => x"65",
          7445 => x"74",
          7446 => x"6c",
          7447 => x"65",
          7448 => x"64",
          7449 => x"6c",
          7450 => x"64",
          7451 => x"73",
          7452 => x"63",
          7453 => x"69",
          7454 => x"76",
          7455 => x"6c",
          7456 => x"00",
          7457 => x"68",
          7458 => x"00",
          7459 => x"65",
          7460 => x"00",
          7461 => x"6f",
          7462 => x"2e",
          7463 => x"61",
          7464 => x"2e",
          7465 => x"72",
          7466 => x"63",
          7467 => x"00",
          7468 => x"79",
          7469 => x"61",
          7470 => x"79",
          7471 => x"2e",
          7472 => x"61",
          7473 => x"38",
          7474 => x"20",
          7475 => x"00",
          7476 => x"00",
          7477 => x"34",
          7478 => x"20",
          7479 => x"00",
          7480 => x"20",
          7481 => x"2f",
          7482 => x"00",
          7483 => x"00",
          7484 => x"72",
          7485 => x"29",
          7486 => x"2a",
          7487 => x"3a",
          7488 => x"73",
          7489 => x"73",
          7490 => x"20",
          7491 => x"20",
          7492 => x"00",
          7493 => x"70",
          7494 => x"73",
          7495 => x"20",
          7496 => x"20",
          7497 => x"00",
          7498 => x"74",
          7499 => x"48",
          7500 => x"00",
          7501 => x"54",
          7502 => x"72",
          7503 => x"52",
          7504 => x"6e",
          7505 => x"00",
          7506 => x"54",
          7507 => x"72",
          7508 => x"52",
          7509 => x"6e",
          7510 => x"00",
          7511 => x"57",
          7512 => x"72",
          7513 => x"43",
          7514 => x"6e",
          7515 => x"00",
          7516 => x"74",
          7517 => x"00",
          7518 => x"69",
          7519 => x"74",
          7520 => x"67",
          7521 => x"65",
          7522 => x"61",
          7523 => x"69",
          7524 => x"00",
          7525 => x"65",
          7526 => x"00",
          7527 => x"75",
          7528 => x"69",
          7529 => x"69",
          7530 => x"73",
          7531 => x"72",
          7532 => x"65",
          7533 => x"74",
          7534 => x"6c",
          7535 => x"00",
          7536 => x"00",
          7537 => x"64",
          7538 => x"64",
          7539 => x"55",
          7540 => x"3a",
          7541 => x"25",
          7542 => x"6c",
          7543 => x"74",
          7544 => x"00",
          7545 => x"74",
          7546 => x"6c",
          7547 => x"2e",
          7548 => x"6c",
          7549 => x"64",
          7550 => x"6c",
          7551 => x"00",
          7552 => x"65",
          7553 => x"63",
          7554 => x"29",
          7555 => x"65",
          7556 => x"63",
          7557 => x"30",
          7558 => x"0a",
          7559 => x"25",
          7560 => x"00",
          7561 => x"25",
          7562 => x"6d",
          7563 => x"2e",
          7564 => x"38",
          7565 => x"29",
          7566 => x"28",
          7567 => x"00",
          7568 => x"67",
          7569 => x"38",
          7570 => x"2d",
          7571 => x"6e",
          7572 => x"00",
          7573 => x"65",
          7574 => x"6f",
          7575 => x"00",
          7576 => x"5c",
          7577 => x"6d",
          7578 => x"61",
          7579 => x"63",
          7580 => x"72",
          7581 => x"6f",
          7582 => x"00",
          7583 => x"2f",
          7584 => x"64",
          7585 => x"25",
          7586 => x"43",
          7587 => x"75",
          7588 => x"00",
          7589 => x"63",
          7590 => x"65",
          7591 => x"00",
          7592 => x"73",
          7593 => x"20",
          7594 => x"73",
          7595 => x"6f",
          7596 => x"73",
          7597 => x"58",
          7598 => x"20",
          7599 => x"6d",
          7600 => x"72",
          7601 => x"73",
          7602 => x"58",
          7603 => x"20",
          7604 => x"53",
          7605 => x"64",
          7606 => x"20",
          7607 => x"58",
          7608 => x"73",
          7609 => x"20",
          7610 => x"20",
          7611 => x"20",
          7612 => x"20",
          7613 => x"58",
          7614 => x"20",
          7615 => x"20",
          7616 => x"72",
          7617 => x"20",
          7618 => x"25",
          7619 => x"00",
          7620 => x"73",
          7621 => x"44",
          7622 => x"63",
          7623 => x"20",
          7624 => x"4d",
          7625 => x"20",
          7626 => x"43",
          7627 => x"65",
          7628 => x"20",
          7629 => x"25",
          7630 => x"00",
          7631 => x"49",
          7632 => x"32",
          7633 => x"43",
          7634 => x"20",
          7635 => x"00",
          7636 => x"53",
          7637 => x"55",
          7638 => x"20",
          7639 => x"54",
          7640 => x"6e",
          7641 => x"32",
          7642 => x"20",
          7643 => x"20",
          7644 => x"65",
          7645 => x"32",
          7646 => x"20",
          7647 => x"44",
          7648 => x"69",
          7649 => x"32",
          7650 => x"20",
          7651 => x"20",
          7652 => x"58",
          7653 => x"0a",
          7654 => x"41",
          7655 => x"28",
          7656 => x"38",
          7657 => x"20",
          7658 => x"52",
          7659 => x"58",
          7660 => x"0a",
          7661 => x"52",
          7662 => x"28",
          7663 => x"38",
          7664 => x"20",
          7665 => x"41",
          7666 => x"58",
          7667 => x"0a",
          7668 => x"20",
          7669 => x"66",
          7670 => x"6b",
          7671 => x"4f",
          7672 => x"61",
          7673 => x"64",
          7674 => x"65",
          7675 => x"4f",
          7676 => x"00",
          7677 => x"f1",
          7678 => x"00",
          7679 => x"00",
          7680 => x"f1",
          7681 => x"00",
          7682 => x"00",
          7683 => x"f1",
          7684 => x"00",
          7685 => x"00",
          7686 => x"f1",
          7687 => x"00",
          7688 => x"00",
          7689 => x"f1",
          7690 => x"00",
          7691 => x"00",
          7692 => x"f1",
          7693 => x"00",
          7694 => x"00",
          7695 => x"f1",
          7696 => x"00",
          7697 => x"00",
          7698 => x"f1",
          7699 => x"00",
          7700 => x"00",
          7701 => x"f0",
          7702 => x"00",
          7703 => x"00",
          7704 => x"f0",
          7705 => x"00",
          7706 => x"00",
          7707 => x"f0",
          7708 => x"00",
          7709 => x"43",
          7710 => x"41",
          7711 => x"35",
          7712 => x"46",
          7713 => x"32",
          7714 => x"00",
          7715 => x"00",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"79",
          7721 => x"30",
          7722 => x"6e",
          7723 => x"6e",
          7724 => x"20",
          7725 => x"20",
          7726 => x"69",
          7727 => x"2e",
          7728 => x"79",
          7729 => x"00",
          7730 => x"73",
          7731 => x"66",
          7732 => x"6c",
          7733 => x"36",
          7734 => x"00",
          7735 => x"20",
          7736 => x"74",
          7737 => x"73",
          7738 => x"6c",
          7739 => x"46",
          7740 => x"73",
          7741 => x"31",
          7742 => x"41",
          7743 => x"43",
          7744 => x"31",
          7745 => x"31",
          7746 => x"31",
          7747 => x"31",
          7748 => x"31",
          7749 => x"31",
          7750 => x"31",
          7751 => x"31",
          7752 => x"31",
          7753 => x"32",
          7754 => x"32",
          7755 => x"33",
          7756 => x"46",
          7757 => x"00",
          7758 => x"00",
          7759 => x"64",
          7760 => x"25",
          7761 => x"32",
          7762 => x"25",
          7763 => x"3a",
          7764 => x"64",
          7765 => x"2c",
          7766 => x"00",
          7767 => x"00",
          7768 => x"25",
          7769 => x"70",
          7770 => x"73",
          7771 => x"3a",
          7772 => x"32",
          7773 => x"3a",
          7774 => x"32",
          7775 => x"3a",
          7776 => x"00",
          7777 => x"74",
          7778 => x"64",
          7779 => x"00",
          7780 => x"7c",
          7781 => x"3b",
          7782 => x"54",
          7783 => x"00",
          7784 => x"4f",
          7785 => x"20",
          7786 => x"20",
          7787 => x"20",
          7788 => x"45",
          7789 => x"33",
          7790 => x"f3",
          7791 => x"00",
          7792 => x"05",
          7793 => x"18",
          7794 => x"45",
          7795 => x"45",
          7796 => x"92",
          7797 => x"9a",
          7798 => x"4f",
          7799 => x"aa",
          7800 => x"b2",
          7801 => x"ba",
          7802 => x"c2",
          7803 => x"ca",
          7804 => x"d2",
          7805 => x"da",
          7806 => x"e2",
          7807 => x"ea",
          7808 => x"f2",
          7809 => x"fa",
          7810 => x"2c",
          7811 => x"2a",
          7812 => x"00",
          7813 => x"00",
          7814 => x"00",
          7815 => x"00",
          7816 => x"00",
          7817 => x"00",
          7818 => x"00",
          7819 => x"00",
          7820 => x"00",
          7821 => x"00",
          7822 => x"00",
          7823 => x"00",
          7824 => x"01",
          7825 => x"00",
          7826 => x"00",
          7827 => x"00",
          7828 => x"00",
          7829 => x"25",
          7830 => x"25",
          7831 => x"25",
          7832 => x"25",
          7833 => x"25",
          7834 => x"25",
          7835 => x"25",
          7836 => x"25",
          7837 => x"25",
          7838 => x"25",
          7839 => x"25",
          7840 => x"25",
          7841 => x"03",
          7842 => x"03",
          7843 => x"03",
          7844 => x"22",
          7845 => x"22",
          7846 => x"22",
          7847 => x"22",
          7848 => x"00",
          7849 => x"03",
          7850 => x"00",
          7851 => x"01",
          7852 => x"01",
          7853 => x"01",
          7854 => x"01",
          7855 => x"01",
          7856 => x"01",
          7857 => x"01",
          7858 => x"01",
          7859 => x"01",
          7860 => x"02",
          7861 => x"02",
          7862 => x"01",
          7863 => x"01",
          7864 => x"01",
          7865 => x"01",
          7866 => x"01",
          7867 => x"01",
          7868 => x"01",
          7869 => x"01",
          7870 => x"01",
          7871 => x"01",
          7872 => x"01",
          7873 => x"01",
          7874 => x"01",
          7875 => x"01",
          7876 => x"01",
          7877 => x"00",
          7878 => x"02",
          7879 => x"02",
          7880 => x"02",
          7881 => x"02",
          7882 => x"01",
          7883 => x"02",
          7884 => x"02",
          7885 => x"02",
          7886 => x"01",
          7887 => x"02",
          7888 => x"02",
          7889 => x"01",
          7890 => x"02",
          7891 => x"2c",
          7892 => x"02",
          7893 => x"02",
          7894 => x"02",
          7895 => x"02",
          7896 => x"02",
          7897 => x"03",
          7898 => x"00",
          7899 => x"03",
          7900 => x"00",
          7901 => x"03",
          7902 => x"03",
          7903 => x"03",
          7904 => x"03",
          7905 => x"03",
          7906 => x"04",
          7907 => x"04",
          7908 => x"04",
          7909 => x"04",
          7910 => x"04",
          7911 => x"00",
          7912 => x"1e",
          7913 => x"1f",
          7914 => x"1f",
          7915 => x"1f",
          7916 => x"1f",
          7917 => x"1f",
          7918 => x"00",
          7919 => x"1f",
          7920 => x"1f",
          7921 => x"1f",
          7922 => x"06",
          7923 => x"06",
          7924 => x"1f",
          7925 => x"00",
          7926 => x"1f",
          7927 => x"1f",
          7928 => x"21",
          7929 => x"02",
          7930 => x"24",
          7931 => x"2c",
          7932 => x"2c",
          7933 => x"2d",
          7934 => x"00",
          7935 => x"e6",
          7936 => x"00",
          7937 => x"e7",
          7938 => x"00",
          7939 => x"e7",
          7940 => x"00",
          7941 => x"e7",
          7942 => x"00",
          7943 => x"e7",
          7944 => x"00",
          7945 => x"e7",
          7946 => x"00",
          7947 => x"e7",
          7948 => x"00",
          7949 => x"e7",
          7950 => x"00",
          7951 => x"e7",
          7952 => x"00",
          7953 => x"e7",
          7954 => x"00",
          7955 => x"e7",
          7956 => x"00",
          7957 => x"e7",
          7958 => x"00",
          7959 => x"e7",
          7960 => x"00",
          7961 => x"e7",
          7962 => x"00",
          7963 => x"e7",
          7964 => x"00",
          7965 => x"e7",
          7966 => x"00",
          7967 => x"e7",
          7968 => x"00",
          7969 => x"e7",
          7970 => x"00",
          7971 => x"e7",
          7972 => x"00",
          7973 => x"e7",
          7974 => x"00",
          7975 => x"e7",
          7976 => x"00",
          7977 => x"e7",
          7978 => x"00",
          7979 => x"e7",
          7980 => x"00",
          7981 => x"e7",
          7982 => x"00",
          7983 => x"e7",
          7984 => x"00",
          7985 => x"e7",
          7986 => x"00",
          7987 => x"e7",
          7988 => x"00",
          7989 => x"e7",
          7990 => x"00",
          7991 => x"00",
          7992 => x"7f",
          7993 => x"7f",
          7994 => x"7f",
          7995 => x"00",
          7996 => x"ff",
          7997 => x"00",
          7998 => x"00",
          7999 => x"e1",
          8000 => x"00",
          8001 => x"01",
          8002 => x"00",
          8003 => x"00",
          8004 => x"00",
          8005 => x"00",
          8006 => x"00",
          8007 => x"00",
          8008 => x"00",
          8009 => x"00",
          8010 => x"00",
          8011 => x"00",
          8012 => x"00",
          8013 => x"00",
          8014 => x"00",
          8015 => x"00",
          8016 => x"00",
          8017 => x"00",
          8018 => x"5f",
          8019 => x"40",
          8020 => x"73",
          8021 => x"6b",
          8022 => x"63",
          8023 => x"33",
          8024 => x"2d",
          8025 => x"f3",
          8026 => x"f0",
          8027 => x"82",
          8028 => x"58",
          8029 => x"40",
          8030 => x"53",
          8031 => x"4b",
          8032 => x"43",
          8033 => x"33",
          8034 => x"2d",
          8035 => x"f3",
          8036 => x"f0",
          8037 => x"82",
          8038 => x"58",
          8039 => x"60",
          8040 => x"53",
          8041 => x"4b",
          8042 => x"43",
          8043 => x"23",
          8044 => x"3d",
          8045 => x"e0",
          8046 => x"f0",
          8047 => x"87",
          8048 => x"1e",
          8049 => x"00",
          8050 => x"13",
          8051 => x"0b",
          8052 => x"03",
          8053 => x"f0",
          8054 => x"f0",
          8055 => x"f0",
          8056 => x"f0",
          8057 => x"82",
          8058 => x"cf",
          8059 => x"d7",
          8060 => x"41",
          8061 => x"6c",
          8062 => x"d9",
          8063 => x"7e",
          8064 => x"d1",
          8065 => x"c2",
          8066 => x"f0",
          8067 => x"82",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"f1",
          8083 => x"f1",
          8084 => x"f1",
          8085 => x"f1",
          8086 => x"f2",
          8087 => x"f2",
          8088 => x"f2",
          8089 => x"f2",
          8090 => x"f2",
          8091 => x"f2",
          8092 => x"f2",
          8093 => x"f2",
          8094 => x"f2",
          8095 => x"f2",
          8096 => x"f2",
          8097 => x"f2",
          8098 => x"f2",
          8099 => x"f2",
          8100 => x"f2",
          8101 => x"f2",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"32",
          9103 => x"00",
          9104 => x"f6",
          9105 => x"fe",
          9106 => x"c6",
          9107 => x"ef",
          9108 => x"66",
          9109 => x"2e",
          9110 => x"26",
          9111 => x"57",
          9112 => x"06",
          9113 => x"0e",
          9114 => x"16",
          9115 => x"be",
          9116 => x"86",
          9117 => x"8e",
          9118 => x"96",
          9119 => x"a5",
          9120 => x"00",
          9121 => x"00",
          9122 => x"00",
          9123 => x"00",
          9124 => x"00",
          9125 => x"00",
          9126 => x"00",
          9127 => x"00",
          9128 => x"00",
          9129 => x"00",
          9130 => x"00",
          9131 => x"00",
          9132 => x"00",
          9133 => x"00",
          9134 => x"00",
          9135 => x"01",
          9136 => x"01",
        others => X"00"
    );

    shared variable RAM6 : ramArray :=
    (
             0 => x"0d",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"83",
             9 => x"2b",
            10 => x"00",
            11 => x"00",
            12 => x"ff",
            13 => x"82",
            14 => x"83",
            15 => x"a5",
            16 => x"05",
            17 => x"09",
            18 => x"51",
            19 => x"00",
            20 => x"2e",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"10",
            26 => x"0a",
            27 => x"00",
            28 => x"2e",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"04",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"53",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"81",
            45 => x"04",
            46 => x"00",
            47 => x"00",
            48 => x"9f",
            49 => x"06",
            50 => x"00",
            51 => x"00",
            52 => x"06",
            53 => x"05",
            54 => x"06",
            55 => x"00",
            56 => x"05",
            57 => x"81",
            58 => x"00",
            59 => x"00",
            60 => x"05",
            61 => x"09",
            62 => x"00",
            63 => x"00",
            64 => x"04",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"05",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"73",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"83",
            77 => x"10",
            78 => x"00",
            79 => x"00",
            80 => x"0b",
            81 => x"10",
            82 => x"b5",
            83 => x"00",
            84 => x"08",
            85 => x"2d",
            86 => x"8c",
            87 => x"00",
            88 => x"08",
            89 => x"2d",
            90 => x"8c",
            91 => x"00",
            92 => x"09",
            93 => x"54",
            94 => x"ff",
            95 => x"00",
            96 => x"09",
            97 => x"70",
            98 => x"05",
            99 => x"04",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"10",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"04",
           133 => x"0b",
           134 => x"8c",
           135 => x"04",
           136 => x"0b",
           137 => x"8c",
           138 => x"04",
           139 => x"0b",
           140 => x"8d",
           141 => x"04",
           142 => x"0b",
           143 => x"8d",
           144 => x"04",
           145 => x"0b",
           146 => x"8e",
           147 => x"04",
           148 => x"0b",
           149 => x"8e",
           150 => x"04",
           151 => x"0b",
           152 => x"8f",
           153 => x"04",
           154 => x"0b",
           155 => x"8f",
           156 => x"04",
           157 => x"0b",
           158 => x"90",
           159 => x"04",
           160 => x"0b",
           161 => x"91",
           162 => x"04",
           163 => x"0b",
           164 => x"91",
           165 => x"04",
           166 => x"0b",
           167 => x"92",
           168 => x"04",
           169 => x"0b",
           170 => x"92",
           171 => x"04",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"84",
           193 => x"84",
           194 => x"04",
           195 => x"84",
           196 => x"04",
           197 => x"84",
           198 => x"04",
           199 => x"84",
           200 => x"04",
           201 => x"84",
           202 => x"04",
           203 => x"84",
           204 => x"04",
           205 => x"84",
           206 => x"04",
           207 => x"84",
           208 => x"04",
           209 => x"84",
           210 => x"04",
           211 => x"84",
           212 => x"04",
           213 => x"84",
           214 => x"04",
           215 => x"84",
           216 => x"04",
           217 => x"2d",
           218 => x"90",
           219 => x"e1",
           220 => x"80",
           221 => x"d2",
           222 => x"c0",
           223 => x"80",
           224 => x"80",
           225 => x"0c",
           226 => x"08",
           227 => x"90",
           228 => x"90",
           229 => x"bb",
           230 => x"bb",
           231 => x"84",
           232 => x"84",
           233 => x"04",
           234 => x"2d",
           235 => x"90",
           236 => x"fc",
           237 => x"80",
           238 => x"de",
           239 => x"c0",
           240 => x"82",
           241 => x"80",
           242 => x"0c",
           243 => x"08",
           244 => x"90",
           245 => x"90",
           246 => x"bb",
           247 => x"bb",
           248 => x"84",
           249 => x"84",
           250 => x"04",
           251 => x"2d",
           252 => x"90",
           253 => x"94",
           254 => x"80",
           255 => x"95",
           256 => x"c0",
           257 => x"83",
           258 => x"80",
           259 => x"0c",
           260 => x"08",
           261 => x"90",
           262 => x"90",
           263 => x"bb",
           264 => x"bb",
           265 => x"84",
           266 => x"84",
           267 => x"04",
           268 => x"2d",
           269 => x"90",
           270 => x"86",
           271 => x"80",
           272 => x"a1",
           273 => x"c0",
           274 => x"82",
           275 => x"80",
           276 => x"0c",
           277 => x"08",
           278 => x"90",
           279 => x"90",
           280 => x"bb",
           281 => x"bb",
           282 => x"84",
           283 => x"84",
           284 => x"04",
           285 => x"2d",
           286 => x"90",
           287 => x"a9",
           288 => x"80",
           289 => x"d0",
           290 => x"c0",
           291 => x"80",
           292 => x"80",
           293 => x"0c",
           294 => x"08",
           295 => x"90",
           296 => x"08",
           297 => x"90",
           298 => x"90",
           299 => x"bb",
           300 => x"bb",
           301 => x"84",
           302 => x"84",
           303 => x"04",
           304 => x"2d",
           305 => x"90",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"73",
           311 => x"81",
           312 => x"07",
           313 => x"72",
           314 => x"09",
           315 => x"0a",
           316 => x"51",
           317 => x"84",
           318 => x"70",
           319 => x"93",
           320 => x"ca",
           321 => x"70",
           322 => x"74",
           323 => x"c5",
           324 => x"0d",
           325 => x"32",
           326 => x"58",
           327 => x"09",
           328 => x"77",
           329 => x"07",
           330 => x"80",
           331 => x"b2",
           332 => x"bb",
           333 => x"ff",
           334 => x"75",
           335 => x"73",
           336 => x"9f",
           337 => x"24",
           338 => x"71",
           339 => x"04",
           340 => x"3d",
           341 => x"86",
           342 => x"56",
           343 => x"53",
           344 => x"9d",
           345 => x"8d",
           346 => x"3d",
           347 => x"85",
           348 => x"0d",
           349 => x"70",
           350 => x"81",
           351 => x"5b",
           352 => x"06",
           353 => x"7b",
           354 => x"81",
           355 => x"81",
           356 => x"81",
           357 => x"70",
           358 => x"38",
           359 => x"2a",
           360 => x"7e",
           361 => x"07",
           362 => x"38",
           363 => x"84",
           364 => x"2a",
           365 => x"05",
           366 => x"70",
           367 => x"70",
           368 => x"80",
           369 => x"06",
           370 => x"33",
           371 => x"b8",
           372 => x"93",
           373 => x"8a",
           374 => x"38",
           375 => x"8b",
           376 => x"cc",
           377 => x"70",
           378 => x"81",
           379 => x"38",
           380 => x"97",
           381 => x"05",
           382 => x"54",
           383 => x"7c",
           384 => x"7c",
           385 => x"fe",
           386 => x"39",
           387 => x"08",
           388 => x"41",
           389 => x"75",
           390 => x"08",
           391 => x"18",
           392 => x"88",
           393 => x"55",
           394 => x"79",
           395 => x"bb",
           396 => x"c5",
           397 => x"2b",
           398 => x"2e",
           399 => x"fc",
           400 => x"55",
           401 => x"5f",
           402 => x"80",
           403 => x"79",
           404 => x"80",
           405 => x"90",
           406 => x"06",
           407 => x"75",
           408 => x"54",
           409 => x"83",
           410 => x"86",
           411 => x"54",
           412 => x"79",
           413 => x"83",
           414 => x"2e",
           415 => x"06",
           416 => x"2a",
           417 => x"7a",
           418 => x"97",
           419 => x"8f",
           420 => x"7e",
           421 => x"80",
           422 => x"90",
           423 => x"9d",
           424 => x"3f",
           425 => x"80",
           426 => x"54",
           427 => x"06",
           428 => x"79",
           429 => x"05",
           430 => x"75",
           431 => x"87",
           432 => x"29",
           433 => x"5b",
           434 => x"7a",
           435 => x"7a",
           436 => x"e3",
           437 => x"2e",
           438 => x"81",
           439 => x"96",
           440 => x"52",
           441 => x"94",
           442 => x"81",
           443 => x"38",
           444 => x"80",
           445 => x"55",
           446 => x"52",
           447 => x"7a",
           448 => x"33",
           449 => x"c8",
           450 => x"f8",
           451 => x"08",
           452 => x"42",
           453 => x"84",
           454 => x"13",
           455 => x"84",
           456 => x"70",
           457 => x"41",
           458 => x"5c",
           459 => x"84",
           460 => x"70",
           461 => x"25",
           462 => x"85",
           463 => x"83",
           464 => x"ff",
           465 => x"75",
           466 => x"d8",
           467 => x"ff",
           468 => x"ff",
           469 => x"70",
           470 => x"3f",
           471 => x"fc",
           472 => x"fc",
           473 => x"58",
           474 => x"81",
           475 => x"38",
           476 => x"71",
           477 => x"7e",
           478 => x"bf",
           479 => x"ad",
           480 => x"5b",
           481 => x"7a",
           482 => x"59",
           483 => x"7f",
           484 => x"06",
           485 => x"38",
           486 => x"84",
           487 => x"31",
           488 => x"58",
           489 => x"7c",
           490 => x"f7",
           491 => x"08",
           492 => x"79",
           493 => x"3f",
           494 => x"06",
           495 => x"c4",
           496 => x"58",
           497 => x"39",
           498 => x"80",
           499 => x"54",
           500 => x"52",
           501 => x"7c",
           502 => x"90",
           503 => x"7c",
           504 => x"88",
           505 => x"fb",
           506 => x"2c",
           507 => x"2c",
           508 => x"53",
           509 => x"7c",
           510 => x"81",
           511 => x"38",
           512 => x"2a",
           513 => x"5b",
           514 => x"c8",
           515 => x"98",
           516 => x"52",
           517 => x"7c",
           518 => x"be",
           519 => x"3f",
           520 => x"06",
           521 => x"fd",
           522 => x"71",
           523 => x"fd",
           524 => x"e4",
           525 => x"b5",
           526 => x"0d",
           527 => x"08",
           528 => x"32",
           529 => x"57",
           530 => x"06",
           531 => x"56",
           532 => x"84",
           533 => x"14",
           534 => x"08",
           535 => x"70",
           536 => x"2e",
           537 => x"d7",
           538 => x"e6",
           539 => x"08",
           540 => x"80",
           541 => x"75",
           542 => x"04",
           543 => x"80",
           544 => x"81",
           545 => x"57",
           546 => x"06",
           547 => x"33",
           548 => x"98",
           549 => x"0c",
           550 => x"05",
           551 => x"38",
           552 => x"53",
           553 => x"2e",
           554 => x"56",
           555 => x"39",
           556 => x"52",
           557 => x"04",
           558 => x"33",
           559 => x"56",
           560 => x"38",
           561 => x"80",
           562 => x"72",
           563 => x"08",
           564 => x"05",
           565 => x"13",
           566 => x"bb",
           567 => x"52",
           568 => x"08",
           569 => x"84",
           570 => x"05",
           571 => x"fb",
           572 => x"81",
           573 => x"55",
           574 => x"38",
           575 => x"b3",
           576 => x"71",
           577 => x"70",
           578 => x"f0",
           579 => x"08",
           580 => x"ff",
           581 => x"87",
           582 => x"53",
           583 => x"81",
           584 => x"84",
           585 => x"75",
           586 => x"84",
           587 => x"08",
           588 => x"33",
           589 => x"84",
           590 => x"07",
           591 => x"73",
           592 => x"04",
           593 => x"34",
           594 => x"75",
           595 => x"81",
           596 => x"ff",
           597 => x"33",
           598 => x"34",
           599 => x"0c",
           600 => x"76",
           601 => x"70",
           602 => x"a1",
           603 => x"70",
           604 => x"05",
           605 => x"38",
           606 => x"0d",
           607 => x"d9",
           608 => x"13",
           609 => x"34",
           610 => x"38",
           611 => x"33",
           612 => x"38",
           613 => x"53",
           614 => x"51",
           615 => x"31",
           616 => x"0d",
           617 => x"54",
           618 => x"33",
           619 => x"34",
           620 => x"0c",
           621 => x"75",
           622 => x"70",
           623 => x"05",
           624 => x"34",
           625 => x"84",
           626 => x"fc",
           627 => x"54",
           628 => x"75",
           629 => x"71",
           630 => x"81",
           631 => x"ff",
           632 => x"70",
           633 => x"04",
           634 => x"53",
           635 => x"ff",
           636 => x"2e",
           637 => x"84",
           638 => x"bb",
           639 => x"3d",
           640 => x"80",
           641 => x"bb",
           642 => x"b4",
           643 => x"84",
           644 => x"84",
           645 => x"34",
           646 => x"08",
           647 => x"08",
           648 => x"3d",
           649 => x"71",
           650 => x"2e",
           651 => x"33",
           652 => x"12",
           653 => x"ea",
           654 => x"52",
           655 => x"0d",
           656 => x"72",
           657 => x"8e",
           658 => x"34",
           659 => x"84",
           660 => x"fa",
           661 => x"52",
           662 => x"80",
           663 => x"e0",
           664 => x"73",
           665 => x"84",
           666 => x"26",
           667 => x"2e",
           668 => x"2a",
           669 => x"54",
           670 => x"a8",
           671 => x"74",
           672 => x"11",
           673 => x"06",
           674 => x"52",
           675 => x"38",
           676 => x"bb",
           677 => x"3d",
           678 => x"70",
           679 => x"84",
           680 => x"70",
           681 => x"80",
           682 => x"71",
           683 => x"70",
           684 => x"74",
           685 => x"73",
           686 => x"10",
           687 => x"81",
           688 => x"30",
           689 => x"84",
           690 => x"51",
           691 => x"51",
           692 => x"54",
           693 => x"0d",
           694 => x"54",
           695 => x"73",
           696 => x"0c",
           697 => x"0d",
           698 => x"80",
           699 => x"3f",
           700 => x"52",
           701 => x"fe",
           702 => x"31",
           703 => x"c5",
           704 => x"38",
           705 => x"31",
           706 => x"80",
           707 => x"10",
           708 => x"07",
           709 => x"70",
           710 => x"31",
           711 => x"58",
           712 => x"bb",
           713 => x"3d",
           714 => x"7a",
           715 => x"7d",
           716 => x"57",
           717 => x"55",
           718 => x"08",
           719 => x"0c",
           720 => x"7b",
           721 => x"77",
           722 => x"a0",
           723 => x"15",
           724 => x"73",
           725 => x"80",
           726 => x"38",
           727 => x"26",
           728 => x"a0",
           729 => x"74",
           730 => x"ff",
           731 => x"ff",
           732 => x"38",
           733 => x"54",
           734 => x"78",
           735 => x"13",
           736 => x"56",
           737 => x"38",
           738 => x"56",
           739 => x"bb",
           740 => x"70",
           741 => x"56",
           742 => x"fe",
           743 => x"70",
           744 => x"a6",
           745 => x"a0",
           746 => x"38",
           747 => x"89",
           748 => x"bb",
           749 => x"58",
           750 => x"55",
           751 => x"0b",
           752 => x"04",
           753 => x"80",
           754 => x"56",
           755 => x"06",
           756 => x"70",
           757 => x"38",
           758 => x"b0",
           759 => x"80",
           760 => x"8a",
           761 => x"c4",
           762 => x"e0",
           763 => x"d0",
           764 => x"90",
           765 => x"81",
           766 => x"81",
           767 => x"38",
           768 => x"79",
           769 => x"a0",
           770 => x"84",
           771 => x"81",
           772 => x"3d",
           773 => x"0c",
           774 => x"2e",
           775 => x"15",
           776 => x"73",
           777 => x"73",
           778 => x"a0",
           779 => x"80",
           780 => x"e1",
           781 => x"3d",
           782 => x"78",
           783 => x"fe",
           784 => x"0c",
           785 => x"3f",
           786 => x"84",
           787 => x"73",
           788 => x"10",
           789 => x"08",
           790 => x"3f",
           791 => x"51",
           792 => x"83",
           793 => x"3d",
           794 => x"9d",
           795 => x"84",
           796 => x"04",
           797 => x"83",
           798 => x"ee",
           799 => x"d0",
           800 => x"0d",
           801 => x"3f",
           802 => x"51",
           803 => x"83",
           804 => x"3d",
           805 => x"c5",
           806 => x"cc",
           807 => x"04",
           808 => x"83",
           809 => x"ee",
           810 => x"d2",
           811 => x"0d",
           812 => x"3f",
           813 => x"51",
           814 => x"83",
           815 => x"3d",
           816 => x"ed",
           817 => x"d4",
           818 => x"04",
           819 => x"08",
           820 => x"5b",
           821 => x"79",
           822 => x"57",
           823 => x"26",
           824 => x"70",
           825 => x"74",
           826 => x"8c",
           827 => x"3f",
           828 => x"84",
           829 => x"51",
           830 => x"78",
           831 => x"2a",
           832 => x"80",
           833 => x"08",
           834 => x"38",
           835 => x"f5",
           836 => x"83",
           837 => x"e0",
           838 => x"84",
           839 => x"bb",
           840 => x"84",
           841 => x"fb",
           842 => x"52",
           843 => x"bb",
           844 => x"ff",
           845 => x"fe",
           846 => x"59",
           847 => x"f4",
           848 => x"78",
           849 => x"08",
           850 => x"83",
           851 => x"94",
           852 => x"05",
           853 => x"80",
           854 => x"3f",
           855 => x"80",
           856 => x"38",
           857 => x"0d",
           858 => x"61",
           859 => x"7f",
           860 => x"84",
           861 => x"0d",
           862 => x"02",
           863 => x"73",
           864 => x"5d",
           865 => x"7a",
           866 => x"3f",
           867 => x"80",
           868 => x"90",
           869 => x"82",
           870 => x"27",
           871 => x"d3",
           872 => x"84",
           873 => x"ec",
           874 => x"83",
           875 => x"56",
           876 => x"18",
           877 => x"7a",
           878 => x"9f",
           879 => x"73",
           880 => x"74",
           881 => x"27",
           882 => x"52",
           883 => x"56",
           884 => x"a4",
           885 => x"1c",
           886 => x"84",
           887 => x"2c",
           888 => x"38",
           889 => x"1e",
           890 => x"ff",
           891 => x"0d",
           892 => x"3f",
           893 => x"54",
           894 => x"26",
           895 => x"d3",
           896 => x"84",
           897 => x"ea",
           898 => x"38",
           899 => x"38",
           900 => x"db",
           901 => x"08",
           902 => x"78",
           903 => x"83",
           904 => x"14",
           905 => x"51",
           906 => x"ff",
           907 => x"df",
           908 => x"51",
           909 => x"e8",
           910 => x"3f",
           911 => x"39",
           912 => x"e9",
           913 => x"39",
           914 => x"08",
           915 => x"a8",
           916 => x"80",
           917 => x"38",
           918 => x"9b",
           919 => x"2b",
           920 => x"30",
           921 => x"07",
           922 => x"59",
           923 => x"e8",
           924 => x"bb",
           925 => x"70",
           926 => x"70",
           927 => x"06",
           928 => x"80",
           929 => x"39",
           930 => x"3d",
           931 => x"96",
           932 => x"51",
           933 => x"9d",
           934 => x"72",
           935 => x"71",
           936 => x"81",
           937 => x"72",
           938 => x"71",
           939 => x"81",
           940 => x"72",
           941 => x"71",
           942 => x"81",
           943 => x"72",
           944 => x"71",
           945 => x"53",
           946 => x"3d",
           947 => x"83",
           948 => x"51",
           949 => x"3d",
           950 => x"83",
           951 => x"51",
           952 => x"06",
           953 => x"39",
           954 => x"90",
           955 => x"d7",
           956 => x"51",
           957 => x"c2",
           958 => x"d5",
           959 => x"9b",
           960 => x"06",
           961 => x"38",
           962 => x"3f",
           963 => x"80",
           964 => x"70",
           965 => x"fe",
           966 => x"9a",
           967 => x"8f",
           968 => x"84",
           969 => x"80",
           970 => x"81",
           971 => x"51",
           972 => x"3f",
           973 => x"52",
           974 => x"bd",
           975 => x"d5",
           976 => x"9a",
           977 => x"06",
           978 => x"38",
           979 => x"70",
           980 => x"0c",
           981 => x"c9",
           982 => x"06",
           983 => x"84",
           984 => x"ad",
           985 => x"51",
           986 => x"53",
           987 => x"0b",
           988 => x"ff",
           989 => x"f1",
           990 => x"78",
           991 => x"83",
           992 => x"80",
           993 => x"7b",
           994 => x"81",
           995 => x"2e",
           996 => x"be",
           997 => x"05",
           998 => x"84",
           999 => x"54",
          1000 => x"cf",
          1001 => x"84",
          1002 => x"84",
          1003 => x"5d",
          1004 => x"3d",
          1005 => x"38",
          1006 => x"3f",
          1007 => x"84",
          1008 => x"bb",
          1009 => x"05",
          1010 => x"08",
          1011 => x"2e",
          1012 => x"51",
          1013 => x"8f",
          1014 => x"3d",
          1015 => x"38",
          1016 => x"81",
          1017 => x"53",
          1018 => x"d2",
          1019 => x"b4",
          1020 => x"90",
          1021 => x"7c",
          1022 => x"08",
          1023 => x"70",
          1024 => x"42",
          1025 => x"81",
          1026 => x"2e",
          1027 => x"06",
          1028 => x"81",
          1029 => x"81",
          1030 => x"38",
          1031 => x"d6",
          1032 => x"80",
          1033 => x"b1",
          1034 => x"70",
          1035 => x"91",
          1036 => x"84",
          1037 => x"84",
          1038 => x"0b",
          1039 => x"de",
          1040 => x"82",
          1041 => x"80",
          1042 => x"51",
          1043 => x"f8",
          1044 => x"7d",
          1045 => x"38",
          1046 => x"a1",
          1047 => x"ef",
          1048 => x"54",
          1049 => x"a7",
          1050 => x"fc",
          1051 => x"0c",
          1052 => x"26",
          1053 => x"bf",
          1054 => x"53",
          1055 => x"ec",
          1056 => x"b0",
          1057 => x"84",
          1058 => x"aa",
          1059 => x"41",
          1060 => x"de",
          1061 => x"3f",
          1062 => x"7b",
          1063 => x"83",
          1064 => x"3f",
          1065 => x"fa",
          1066 => x"39",
          1067 => x"3f",
          1068 => x"fa",
          1069 => x"85",
          1070 => x"c8",
          1071 => x"fa",
          1072 => x"53",
          1073 => x"84",
          1074 => x"38",
          1075 => x"ea",
          1076 => x"84",
          1077 => x"bb",
          1078 => x"d0",
          1079 => x"ff",
          1080 => x"eb",
          1081 => x"2e",
          1082 => x"9c",
          1083 => x"04",
          1084 => x"80",
          1085 => x"84",
          1086 => x"3d",
          1087 => x"51",
          1088 => x"86",
          1089 => x"78",
          1090 => x"3f",
          1091 => x"52",
          1092 => x"7e",
          1093 => x"38",
          1094 => x"84",
          1095 => x"3d",
          1096 => x"51",
          1097 => x"80",
          1098 => x"f0",
          1099 => x"a4",
          1100 => x"38",
          1101 => x"83",
          1102 => x"e6",
          1103 => x"51",
          1104 => x"59",
          1105 => x"9f",
          1106 => x"70",
          1107 => x"84",
          1108 => x"e0",
          1109 => x"f8",
          1110 => x"53",
          1111 => x"84",
          1112 => x"38",
          1113 => x"80",
          1114 => x"84",
          1115 => x"d8",
          1116 => x"5d",
          1117 => x"65",
          1118 => x"7a",
          1119 => x"54",
          1120 => x"e4",
          1121 => x"5c",
          1122 => x"39",
          1123 => x"80",
          1124 => x"84",
          1125 => x"3d",
          1126 => x"51",
          1127 => x"80",
          1128 => x"f8",
          1129 => x"b8",
          1130 => x"f6",
          1131 => x"aa",
          1132 => x"93",
          1133 => x"5b",
          1134 => x"eb",
          1135 => x"ff",
          1136 => x"bb",
          1137 => x"b8",
          1138 => x"05",
          1139 => x"08",
          1140 => x"83",
          1141 => x"e6",
          1142 => x"51",
          1143 => x"59",
          1144 => x"9f",
          1145 => x"49",
          1146 => x"05",
          1147 => x"b8",
          1148 => x"05",
          1149 => x"08",
          1150 => x"02",
          1151 => x"81",
          1152 => x"53",
          1153 => x"84",
          1154 => x"b4",
          1155 => x"ff",
          1156 => x"bb",
          1157 => x"b8",
          1158 => x"05",
          1159 => x"08",
          1160 => x"fe",
          1161 => x"e6",
          1162 => x"38",
          1163 => x"98",
          1164 => x"59",
          1165 => x"7a",
          1166 => x"79",
          1167 => x"3f",
          1168 => x"05",
          1169 => x"08",
          1170 => x"88",
          1171 => x"08",
          1172 => x"bb",
          1173 => x"84",
          1174 => x"f4",
          1175 => x"53",
          1176 => x"84",
          1177 => x"88",
          1178 => x"38",
          1179 => x"fe",
          1180 => x"e5",
          1181 => x"38",
          1182 => x"2e",
          1183 => x"47",
          1184 => x"80",
          1185 => x"84",
          1186 => x"5c",
          1187 => x"5c",
          1188 => x"07",
          1189 => x"79",
          1190 => x"83",
          1191 => x"d6",
          1192 => x"53",
          1193 => x"83",
          1194 => x"f4",
          1195 => x"84",
          1196 => x"53",
          1197 => x"84",
          1198 => x"38",
          1199 => x"05",
          1200 => x"ff",
          1201 => x"bb",
          1202 => x"64",
          1203 => x"70",
          1204 => x"3d",
          1205 => x"51",
          1206 => x"80",
          1207 => x"80",
          1208 => x"40",
          1209 => x"11",
          1210 => x"3f",
          1211 => x"f1",
          1212 => x"53",
          1213 => x"84",
          1214 => x"38",
          1215 => x"7c",
          1216 => x"39",
          1217 => x"80",
          1218 => x"84",
          1219 => x"64",
          1220 => x"46",
          1221 => x"09",
          1222 => x"83",
          1223 => x"c0",
          1224 => x"91",
          1225 => x"3f",
          1226 => x"d4",
          1227 => x"fe",
          1228 => x"e0",
          1229 => x"2e",
          1230 => x"05",
          1231 => x"78",
          1232 => x"33",
          1233 => x"83",
          1234 => x"83",
          1235 => x"a1",
          1236 => x"b5",
          1237 => x"3f",
          1238 => x"f8",
          1239 => x"cc",
          1240 => x"80",
          1241 => x"49",
          1242 => x"d3",
          1243 => x"8a",
          1244 => x"83",
          1245 => x"83",
          1246 => x"9b",
          1247 => x"dd",
          1248 => x"80",
          1249 => x"47",
          1250 => x"5d",
          1251 => x"e0",
          1252 => x"86",
          1253 => x"83",
          1254 => x"83",
          1255 => x"fb",
          1256 => x"05",
          1257 => x"80",
          1258 => x"94",
          1259 => x"80",
          1260 => x"bb",
          1261 => x"55",
          1262 => x"af",
          1263 => x"77",
          1264 => x"56",
          1265 => x"da",
          1266 => x"2b",
          1267 => x"52",
          1268 => x"bb",
          1269 => x"83",
          1270 => x"80",
          1271 => x"81",
          1272 => x"83",
          1273 => x"5e",
          1274 => x"88",
          1275 => x"e8",
          1276 => x"3f",
          1277 => x"8d",
          1278 => x"c4",
          1279 => x"70",
          1280 => x"d3",
          1281 => x"15",
          1282 => x"f2",
          1283 => x"51",
          1284 => x"80",
          1285 => x"52",
          1286 => x"ec",
          1287 => x"77",
          1288 => x"53",
          1289 => x"33",
          1290 => x"a0",
          1291 => x"15",
          1292 => x"53",
          1293 => x"81",
          1294 => x"82",
          1295 => x"e7",
          1296 => x"06",
          1297 => x"38",
          1298 => x"73",
          1299 => x"e1",
          1300 => x"54",
          1301 => x"38",
          1302 => x"70",
          1303 => x"72",
          1304 => x"81",
          1305 => x"51",
          1306 => x"0d",
          1307 => x"80",
          1308 => x"80",
          1309 => x"54",
          1310 => x"54",
          1311 => x"53",
          1312 => x"fe",
          1313 => x"76",
          1314 => x"84",
          1315 => x"86",
          1316 => x"dc",
          1317 => x"e5",
          1318 => x"3d",
          1319 => x"11",
          1320 => x"70",
          1321 => x"33",
          1322 => x"26",
          1323 => x"83",
          1324 => x"85",
          1325 => x"26",
          1326 => x"85",
          1327 => x"88",
          1328 => x"e7",
          1329 => x"54",
          1330 => x"cc",
          1331 => x"0c",
          1332 => x"82",
          1333 => x"83",
          1334 => x"84",
          1335 => x"85",
          1336 => x"86",
          1337 => x"74",
          1338 => x"c0",
          1339 => x"98",
          1340 => x"84",
          1341 => x"0d",
          1342 => x"81",
          1343 => x"5e",
          1344 => x"08",
          1345 => x"98",
          1346 => x"87",
          1347 => x"1c",
          1348 => x"79",
          1349 => x"08",
          1350 => x"98",
          1351 => x"87",
          1352 => x"1c",
          1353 => x"ff",
          1354 => x"58",
          1355 => x"56",
          1356 => x"54",
          1357 => x"ff",
          1358 => x"bf",
          1359 => x"3d",
          1360 => x"81",
          1361 => x"de",
          1362 => x"70",
          1363 => x"09",
          1364 => x"e3",
          1365 => x"3d",
          1366 => x"3f",
          1367 => x"98",
          1368 => x"81",
          1369 => x"9e",
          1370 => x"70",
          1371 => x"d2",
          1372 => x"70",
          1373 => x"51",
          1374 => x"08",
          1375 => x"71",
          1376 => x"81",
          1377 => x"38",
          1378 => x"0d",
          1379 => x"33",
          1380 => x"06",
          1381 => x"f4",
          1382 => x"96",
          1383 => x"70",
          1384 => x"70",
          1385 => x"72",
          1386 => x"2e",
          1387 => x"52",
          1388 => x"51",
          1389 => x"2e",
          1390 => x"74",
          1391 => x"86",
          1392 => x"81",
          1393 => x"81",
          1394 => x"cb",
          1395 => x"71",
          1396 => x"84",
          1397 => x"53",
          1398 => x"ff",
          1399 => x"30",
          1400 => x"83",
          1401 => x"fa",
          1402 => x"70",
          1403 => x"e7",
          1404 => x"70",
          1405 => x"80",
          1406 => x"94",
          1407 => x"53",
          1408 => x"71",
          1409 => x"70",
          1410 => x"53",
          1411 => x"2a",
          1412 => x"81",
          1413 => x"52",
          1414 => x"94",
          1415 => x"75",
          1416 => x"76",
          1417 => x"04",
          1418 => x"51",
          1419 => x"06",
          1420 => x"93",
          1421 => x"ff",
          1422 => x"70",
          1423 => x"52",
          1424 => x"0d",
          1425 => x"2a",
          1426 => x"84",
          1427 => x"83",
          1428 => x"08",
          1429 => x"94",
          1430 => x"9e",
          1431 => x"c0",
          1432 => x"87",
          1433 => x"0c",
          1434 => x"d8",
          1435 => x"f3",
          1436 => x"83",
          1437 => x"08",
          1438 => x"bc",
          1439 => x"9e",
          1440 => x"c0",
          1441 => x"87",
          1442 => x"f3",
          1443 => x"83",
          1444 => x"08",
          1445 => x"8c",
          1446 => x"83",
          1447 => x"9e",
          1448 => x"51",
          1449 => x"83",
          1450 => x"9e",
          1451 => x"51",
          1452 => x"81",
          1453 => x"0b",
          1454 => x"80",
          1455 => x"2e",
          1456 => x"87",
          1457 => x"08",
          1458 => x"52",
          1459 => x"71",
          1460 => x"c0",
          1461 => x"06",
          1462 => x"38",
          1463 => x"80",
          1464 => x"90",
          1465 => x"80",
          1466 => x"f4",
          1467 => x"90",
          1468 => x"52",
          1469 => x"52",
          1470 => x"87",
          1471 => x"80",
          1472 => x"83",
          1473 => x"34",
          1474 => x"70",
          1475 => x"70",
          1476 => x"83",
          1477 => x"9e",
          1478 => x"51",
          1479 => x"81",
          1480 => x"0b",
          1481 => x"80",
          1482 => x"83",
          1483 => x"34",
          1484 => x"06",
          1485 => x"f4",
          1486 => x"90",
          1487 => x"52",
          1488 => x"71",
          1489 => x"90",
          1490 => x"53",
          1491 => x"0b",
          1492 => x"06",
          1493 => x"38",
          1494 => x"87",
          1495 => x"70",
          1496 => x"04",
          1497 => x"0d",
          1498 => x"3f",
          1499 => x"a0",
          1500 => x"3f",
          1501 => x"f0",
          1502 => x"85",
          1503 => x"75",
          1504 => x"55",
          1505 => x"33",
          1506 => x"8f",
          1507 => x"f4",
          1508 => x"83",
          1509 => x"38",
          1510 => x"c5",
          1511 => x"83",
          1512 => x"74",
          1513 => x"56",
          1514 => x"33",
          1515 => x"c0",
          1516 => x"08",
          1517 => x"9a",
          1518 => x"da",
          1519 => x"f3",
          1520 => x"ff",
          1521 => x"c1",
          1522 => x"83",
          1523 => x"83",
          1524 => x"52",
          1525 => x"84",
          1526 => x"31",
          1527 => x"83",
          1528 => x"83",
          1529 => x"83",
          1530 => x"87",
          1531 => x"56",
          1532 => x"bf",
          1533 => x"c0",
          1534 => x"bb",
          1535 => x"ff",
          1536 => x"83",
          1537 => x"52",
          1538 => x"84",
          1539 => x"31",
          1540 => x"83",
          1541 => x"83",
          1542 => x"ff",
          1543 => x"f8",
          1544 => x"51",
          1545 => x"52",
          1546 => x"3f",
          1547 => x"f4",
          1548 => x"f0",
          1549 => x"b3",
          1550 => x"bf",
          1551 => x"83",
          1552 => x"83",
          1553 => x"52",
          1554 => x"84",
          1555 => x"31",
          1556 => x"83",
          1557 => x"83",
          1558 => x"fe",
          1559 => x"80",
          1560 => x"8e",
          1561 => x"38",
          1562 => x"ff",
          1563 => x"56",
          1564 => x"39",
          1565 => x"3f",
          1566 => x"2e",
          1567 => x"a0",
          1568 => x"87",
          1569 => x"38",
          1570 => x"83",
          1571 => x"83",
          1572 => x"fc",
          1573 => x"33",
          1574 => x"d2",
          1575 => x"80",
          1576 => x"f4",
          1577 => x"ff",
          1578 => x"54",
          1579 => x"39",
          1580 => x"08",
          1581 => x"ff",
          1582 => x"56",
          1583 => x"39",
          1584 => x"08",
          1585 => x"ff",
          1586 => x"54",
          1587 => x"39",
          1588 => x"08",
          1589 => x"ff",
          1590 => x"55",
          1591 => x"39",
          1592 => x"08",
          1593 => x"ff",
          1594 => x"56",
          1595 => x"39",
          1596 => x"08",
          1597 => x"ff",
          1598 => x"54",
          1599 => x"39",
          1600 => x"3f",
          1601 => x"3f",
          1602 => x"2e",
          1603 => x"0d",
          1604 => x"26",
          1605 => x"8c",
          1606 => x"b4",
          1607 => x"0d",
          1608 => x"c2",
          1609 => x"c4",
          1610 => x"0d",
          1611 => x"aa",
          1612 => x"d4",
          1613 => x"0d",
          1614 => x"92",
          1615 => x"80",
          1616 => x"84",
          1617 => x"c0",
          1618 => x"aa",
          1619 => x"81",
          1620 => x"ec",
          1621 => x"bb",
          1622 => x"57",
          1623 => x"55",
          1624 => x"8e",
          1625 => x"a4",
          1626 => x"bb",
          1627 => x"0b",
          1628 => x"84",
          1629 => x"55",
          1630 => x"30",
          1631 => x"55",
          1632 => x"b0",
          1633 => x"08",
          1634 => x"bb",
          1635 => x"9a",
          1636 => x"3d",
          1637 => x"ad",
          1638 => x"06",
          1639 => x"89",
          1640 => x"ab",
          1641 => x"76",
          1642 => x"ff",
          1643 => x"84",
          1644 => x"0d",
          1645 => x"72",
          1646 => x"73",
          1647 => x"8d",
          1648 => x"83",
          1649 => x"ff",
          1650 => x"53",
          1651 => x"f7",
          1652 => x"84",
          1653 => x"88",
          1654 => x"16",
          1655 => x"76",
          1656 => x"bb",
          1657 => x"1a",
          1658 => x"ff",
          1659 => x"bb",
          1660 => x"1b",
          1661 => x"3f",
          1662 => x"54",
          1663 => x"70",
          1664 => x"27",
          1665 => x"33",
          1666 => x"e5",
          1667 => x"55",
          1668 => x"fe",
          1669 => x"80",
          1670 => x"39",
          1671 => x"f4",
          1672 => x"3f",
          1673 => x"83",
          1674 => x"77",
          1675 => x"84",
          1676 => x"ff",
          1677 => x"55",
          1678 => x"9d",
          1679 => x"70",
          1680 => x"53",
          1681 => x"52",
          1682 => x"2e",
          1683 => x"0b",
          1684 => x"04",
          1685 => x"3d",
          1686 => x"be",
          1687 => x"80",
          1688 => x"33",
          1689 => x"f4",
          1690 => x"76",
          1691 => x"2e",
          1692 => x"88",
          1693 => x"78",
          1694 => x"f8",
          1695 => x"80",
          1696 => x"08",
          1697 => x"79",
          1698 => x"ff",
          1699 => x"2b",
          1700 => x"70",
          1701 => x"2c",
          1702 => x"05",
          1703 => x"49",
          1704 => x"81",
          1705 => x"78",
          1706 => x"80",
          1707 => x"98",
          1708 => x"ec",
          1709 => x"56",
          1710 => x"33",
          1711 => x"83",
          1712 => x"56",
          1713 => x"76",
          1714 => x"bc",
          1715 => x"ba",
          1716 => x"98",
          1717 => x"2b",
          1718 => x"70",
          1719 => x"5f",
          1720 => x"7a",
          1721 => x"e2",
          1722 => x"84",
          1723 => x"2c",
          1724 => x"06",
          1725 => x"8f",
          1726 => x"57",
          1727 => x"0a",
          1728 => x"2c",
          1729 => x"76",
          1730 => x"16",
          1731 => x"83",
          1732 => x"62",
          1733 => x"08",
          1734 => x"2e",
          1735 => x"bc",
          1736 => x"80",
          1737 => x"81",
          1738 => x"fe",
          1739 => x"76",
          1740 => x"76",
          1741 => x"fd",
          1742 => x"a4",
          1743 => x"e8",
          1744 => x"e2",
          1745 => x"34",
          1746 => x"75",
          1747 => x"e8",
          1748 => x"3f",
          1749 => x"7a",
          1750 => x"84",
          1751 => x"84",
          1752 => x"78",
          1753 => x"08",
          1754 => x"c8",
          1755 => x"ff",
          1756 => x"93",
          1757 => x"90",
          1758 => x"05",
          1759 => x"38",
          1760 => x"7c",
          1761 => x"c8",
          1762 => x"38",
          1763 => x"ff",
          1764 => x"52",
          1765 => x"e6",
          1766 => x"b8",
          1767 => x"59",
          1768 => x"ff",
          1769 => x"ff",
          1770 => x"34",
          1771 => x"f4",
          1772 => x"ff",
          1773 => x"76",
          1774 => x"83",
          1775 => x"75",
          1776 => x"f7",
          1777 => x"05",
          1778 => x"fa",
          1779 => x"3f",
          1780 => x"34",
          1781 => x"81",
          1782 => x"b7",
          1783 => x"e2",
          1784 => x"ff",
          1785 => x"88",
          1786 => x"e8",
          1787 => x"3f",
          1788 => x"ff",
          1789 => x"ff",
          1790 => x"74",
          1791 => x"e2",
          1792 => x"e2",
          1793 => x"27",
          1794 => x"52",
          1795 => x"34",
          1796 => x"b2",
          1797 => x"81",
          1798 => x"57",
          1799 => x"84",
          1800 => x"76",
          1801 => x"33",
          1802 => x"e2",
          1803 => x"e2",
          1804 => x"26",
          1805 => x"e2",
          1806 => x"56",
          1807 => x"15",
          1808 => x"98",
          1809 => x"06",
          1810 => x"ef",
          1811 => x"51",
          1812 => x"33",
          1813 => x"e2",
          1814 => x"77",
          1815 => x"08",
          1816 => x"74",
          1817 => x"05",
          1818 => x"5d",
          1819 => x"38",
          1820 => x"ff",
          1821 => x"29",
          1822 => x"84",
          1823 => x"75",
          1824 => x"7b",
          1825 => x"84",
          1826 => x"ff",
          1827 => x"29",
          1828 => x"84",
          1829 => x"7a",
          1830 => x"81",
          1831 => x"08",
          1832 => x"3f",
          1833 => x"0a",
          1834 => x"33",
          1835 => x"a7",
          1836 => x"33",
          1837 => x"84",
          1838 => x"af",
          1839 => x"05",
          1840 => x"81",
          1841 => x"c4",
          1842 => x"84",
          1843 => x"af",
          1844 => x"51",
          1845 => x"81",
          1846 => x"84",
          1847 => x"80",
          1848 => x"10",
          1849 => x"57",
          1850 => x"82",
          1851 => x"05",
          1852 => x"e8",
          1853 => x"0c",
          1854 => x"83",
          1855 => x"83",
          1856 => x"3f",
          1857 => x"83",
          1858 => x"5e",
          1859 => x"08",
          1860 => x"f4",
          1861 => x"de",
          1862 => x"80",
          1863 => x"bb",
          1864 => x"e2",
          1865 => x"38",
          1866 => x"ff",
          1867 => x"52",
          1868 => x"e6",
          1869 => x"80",
          1870 => x"42",
          1871 => x"ff",
          1872 => x"80",
          1873 => x"84",
          1874 => x"c4",
          1875 => x"33",
          1876 => x"80",
          1877 => x"33",
          1878 => x"34",
          1879 => x"34",
          1880 => x"ff",
          1881 => x"70",
          1882 => x"c4",
          1883 => x"24",
          1884 => x"52",
          1885 => x"e2",
          1886 => x"2c",
          1887 => x"56",
          1888 => x"e6",
          1889 => x"e0",
          1890 => x"80",
          1891 => x"c4",
          1892 => x"f3",
          1893 => x"88",
          1894 => x"80",
          1895 => x"98",
          1896 => x"55",
          1897 => x"af",
          1898 => x"77",
          1899 => x"33",
          1900 => x"80",
          1901 => x"98",
          1902 => x"5b",
          1903 => x"16",
          1904 => x"e6",
          1905 => x"ab",
          1906 => x"81",
          1907 => x"e2",
          1908 => x"24",
          1909 => x"7c",
          1910 => x"e2",
          1911 => x"38",
          1912 => x"ff",
          1913 => x"52",
          1914 => x"e6",
          1915 => x"90",
          1916 => x"5d",
          1917 => x"ff",
          1918 => x"80",
          1919 => x"84",
          1920 => x"c4",
          1921 => x"3d",
          1922 => x"81",
          1923 => x"f1",
          1924 => x"76",
          1925 => x"70",
          1926 => x"a1",
          1927 => x"1c",
          1928 => x"ff",
          1929 => x"c8",
          1930 => x"e1",
          1931 => x"c8",
          1932 => x"59",
          1933 => x"c4",
          1934 => x"81",
          1935 => x"75",
          1936 => x"80",
          1937 => x"98",
          1938 => x"5c",
          1939 => x"77",
          1940 => x"ff",
          1941 => x"f0",
          1942 => x"88",
          1943 => x"80",
          1944 => x"98",
          1945 => x"42",
          1946 => x"e6",
          1947 => x"90",
          1948 => x"80",
          1949 => x"c4",
          1950 => x"ff",
          1951 => x"51",
          1952 => x"08",
          1953 => x"08",
          1954 => x"f2",
          1955 => x"86",
          1956 => x"77",
          1957 => x"e6",
          1958 => x"52",
          1959 => x"80",
          1960 => x"98",
          1961 => x"57",
          1962 => x"c8",
          1963 => x"79",
          1964 => x"75",
          1965 => x"39",
          1966 => x"81",
          1967 => x"76",
          1968 => x"84",
          1969 => x"38",
          1970 => x"f4",
          1971 => x"d9",
          1972 => x"83",
          1973 => x"3f",
          1974 => x"3d",
          1975 => x"74",
          1976 => x"0c",
          1977 => x"80",
          1978 => x"75",
          1979 => x"84",
          1980 => x"84",
          1981 => x"75",
          1982 => x"93",
          1983 => x"c8",
          1984 => x"f2",
          1985 => x"88",
          1986 => x"e8",
          1987 => x"3f",
          1988 => x"ff",
          1989 => x"ff",
          1990 => x"78",
          1991 => x"51",
          1992 => x"08",
          1993 => x"08",
          1994 => x"52",
          1995 => x"84",
          1996 => x"57",
          1997 => x"38",
          1998 => x"ff",
          1999 => x"52",
          2000 => x"e6",
          2001 => x"e0",
          2002 => x"57",
          2003 => x"ff",
          2004 => x"a9",
          2005 => x"e2",
          2006 => x"ff",
          2007 => x"51",
          2008 => x"81",
          2009 => x"e2",
          2010 => x"80",
          2011 => x"08",
          2012 => x"84",
          2013 => x"a4",
          2014 => x"88",
          2015 => x"c8",
          2016 => x"c8",
          2017 => x"39",
          2018 => x"c8",
          2019 => x"7b",
          2020 => x"04",
          2021 => x"2e",
          2022 => x"f2",
          2023 => x"c4",
          2024 => x"06",
          2025 => x"ff",
          2026 => x"84",
          2027 => x"2e",
          2028 => x"52",
          2029 => x"e6",
          2030 => x"f8",
          2031 => x"51",
          2032 => x"33",
          2033 => x"34",
          2034 => x"74",
          2035 => x"f4",
          2036 => x"83",
          2037 => x"52",
          2038 => x"bb",
          2039 => x"33",
          2040 => x"70",
          2041 => x"5b",
          2042 => x"33",
          2043 => x"70",
          2044 => x"f4",
          2045 => x"51",
          2046 => x"33",
          2047 => x"56",
          2048 => x"83",
          2049 => x"3d",
          2050 => x"52",
          2051 => x"f4",
          2052 => x"fc",
          2053 => x"de",
          2054 => x"34",
          2055 => x"84",
          2056 => x"93",
          2057 => x"a8",
          2058 => x"38",
          2059 => x"5d",
          2060 => x"52",
          2061 => x"bb",
          2062 => x"7b",
          2063 => x"84",
          2064 => x"3f",
          2065 => x"84",
          2066 => x"84",
          2067 => x"57",
          2068 => x"06",
          2069 => x"83",
          2070 => x"57",
          2071 => x"2b",
          2072 => x"81",
          2073 => x"fb",
          2074 => x"83",
          2075 => x"f4",
          2076 => x"e3",
          2077 => x"83",
          2078 => x"f4",
          2079 => x"74",
          2080 => x"06",
          2081 => x"80",
          2082 => x"fe",
          2083 => x"d0",
          2084 => x"ff",
          2085 => x"81",
          2086 => x"93",
          2087 => x"83",
          2088 => x"51",
          2089 => x"33",
          2090 => x"f4",
          2091 => x"40",
          2092 => x"84",
          2093 => x"70",
          2094 => x"08",
          2095 => x"ff",
          2096 => x"70",
          2097 => x"08",
          2098 => x"ea",
          2099 => x"f4",
          2100 => x"f4",
          2101 => x"51",
          2102 => x"38",
          2103 => x"80",
          2104 => x"c7",
          2105 => x"81",
          2106 => x"38",
          2107 => x"82",
          2108 => x"80",
          2109 => x"57",
          2110 => x"2e",
          2111 => x"75",
          2112 => x"b2",
          2113 => x"2b",
          2114 => x"07",
          2115 => x"5b",
          2116 => x"70",
          2117 => x"84",
          2118 => x"38",
          2119 => x"b0",
          2120 => x"31",
          2121 => x"15",
          2122 => x"34",
          2123 => x"3d",
          2124 => x"83",
          2125 => x"83",
          2126 => x"74",
          2127 => x"c7",
          2128 => x"70",
          2129 => x"70",
          2130 => x"70",
          2131 => x"5d",
          2132 => x"73",
          2133 => x"75",
          2134 => x"81",
          2135 => x"83",
          2136 => x"70",
          2137 => x"5b",
          2138 => x"fa",
          2139 => x"7d",
          2140 => x"5c",
          2141 => x"7d",
          2142 => x"38",
          2143 => x"83",
          2144 => x"56",
          2145 => x"59",
          2146 => x"f8",
          2147 => x"f7",
          2148 => x"b2",
          2149 => x"57",
          2150 => x"81",
          2151 => x"81",
          2152 => x"54",
          2153 => x"80",
          2154 => x"83",
          2155 => x"70",
          2156 => x"88",
          2157 => x"56",
          2158 => x"38",
          2159 => x"83",
          2160 => x"70",
          2161 => x"71",
          2162 => x"11",
          2163 => x"c7",
          2164 => x"33",
          2165 => x"33",
          2166 => x"22",
          2167 => x"29",
          2168 => x"5f",
          2169 => x"38",
          2170 => x"19",
          2171 => x"81",
          2172 => x"ff",
          2173 => x"75",
          2174 => x"7b",
          2175 => x"53",
          2176 => x"5b",
          2177 => x"06",
          2178 => x"39",
          2179 => x"9a",
          2180 => x"8c",
          2181 => x"34",
          2182 => x"8e",
          2183 => x"ff",
          2184 => x"56",
          2185 => x"8e",
          2186 => x"74",
          2187 => x"83",
          2188 => x"e0",
          2189 => x"86",
          2190 => x"07",
          2191 => x"70",
          2192 => x"53",
          2193 => x"08",
          2194 => x"72",
          2195 => x"81",
          2196 => x"34",
          2197 => x"80",
          2198 => x"0d",
          2199 => x"84",
          2200 => x"05",
          2201 => x"84",
          2202 => x"53",
          2203 => x"b8",
          2204 => x"fa",
          2205 => x"c7",
          2206 => x"5f",
          2207 => x"70",
          2208 => x"33",
          2209 => x"83",
          2210 => x"05",
          2211 => x"fa",
          2212 => x"06",
          2213 => x"72",
          2214 => x"53",
          2215 => x"b2",
          2216 => x"b8",
          2217 => x"26",
          2218 => x"76",
          2219 => x"9f",
          2220 => x"70",
          2221 => x"e0",
          2222 => x"54",
          2223 => x"81",
          2224 => x"e3",
          2225 => x"83",
          2226 => x"54",
          2227 => x"74",
          2228 => x"14",
          2229 => x"84",
          2230 => x"83",
          2231 => x"ff",
          2232 => x"54",
          2233 => x"74",
          2234 => x"71",
          2235 => x"86",
          2236 => x"80",
          2237 => x"06",
          2238 => x"57",
          2239 => x"d6",
          2240 => x"84",
          2241 => x"05",
          2242 => x"33",
          2243 => x"15",
          2244 => x"33",
          2245 => x"55",
          2246 => x"72",
          2247 => x"04",
          2248 => x"b2",
          2249 => x"b8",
          2250 => x"27",
          2251 => x"dd",
          2252 => x"83",
          2253 => x"2e",
          2254 => x"76",
          2255 => x"71",
          2256 => x"52",
          2257 => x"38",
          2258 => x"15",
          2259 => x"0b",
          2260 => x"81",
          2261 => x"80",
          2262 => x"e0",
          2263 => x"57",
          2264 => x"fd",
          2265 => x"33",
          2266 => x"b6",
          2267 => x"33",
          2268 => x"fc",
          2269 => x"84",
          2270 => x"86",
          2271 => x"c4",
          2272 => x"b8",
          2273 => x"38",
          2274 => x"84",
          2275 => x"80",
          2276 => x"b4",
          2277 => x"72",
          2278 => x"70",
          2279 => x"bb",
          2280 => x"fa",
          2281 => x"70",
          2282 => x"54",
          2283 => x"83",
          2284 => x"f7",
          2285 => x"75",
          2286 => x"fa",
          2287 => x"0c",
          2288 => x"33",
          2289 => x"2c",
          2290 => x"83",
          2291 => x"84",
          2292 => x"b5",
          2293 => x"ff",
          2294 => x"83",
          2295 => x"34",
          2296 => x"3d",
          2297 => x"34",
          2298 => x"33",
          2299 => x"fe",
          2300 => x"fa",
          2301 => x"0d",
          2302 => x"26",
          2303 => x"98",
          2304 => x"b0",
          2305 => x"2b",
          2306 => x"07",
          2307 => x"2e",
          2308 => x"0b",
          2309 => x"bb",
          2310 => x"fa",
          2311 => x"51",
          2312 => x"84",
          2313 => x"83",
          2314 => x"70",
          2315 => x"fa",
          2316 => x"51",
          2317 => x"80",
          2318 => x"0b",
          2319 => x"04",
          2320 => x"84",
          2321 => x"ff",
          2322 => x"07",
          2323 => x"a5",
          2324 => x"06",
          2325 => x"34",
          2326 => x"81",
          2327 => x"fa",
          2328 => x"b0",
          2329 => x"70",
          2330 => x"83",
          2331 => x"70",
          2332 => x"83",
          2333 => x"d0",
          2334 => x"fe",
          2335 => x"bf",
          2336 => x"b0",
          2337 => x"33",
          2338 => x"70",
          2339 => x"83",
          2340 => x"c0",
          2341 => x"fe",
          2342 => x"af",
          2343 => x"b0",
          2344 => x"33",
          2345 => x"b0",
          2346 => x"33",
          2347 => x"83",
          2348 => x"3d",
          2349 => x"05",
          2350 => x"33",
          2351 => x"33",
          2352 => x"5d",
          2353 => x"38",
          2354 => x"2e",
          2355 => x"34",
          2356 => x"83",
          2357 => x"23",
          2358 => x"0d",
          2359 => x"db",
          2360 => x"81",
          2361 => x"83",
          2362 => x"b5",
          2363 => x"79",
          2364 => x"b8",
          2365 => x"55",
          2366 => x"e4",
          2367 => x"84",
          2368 => x"fc",
          2369 => x"83",
          2370 => x"34",
          2371 => x"b8",
          2372 => x"34",
          2373 => x"0b",
          2374 => x"fa",
          2375 => x"84",
          2376 => x"33",
          2377 => x"7a",
          2378 => x"b2",
          2379 => x"5a",
          2380 => x"10",
          2381 => x"59",
          2382 => x"3f",
          2383 => x"ba",
          2384 => x"26",
          2385 => x"fe",
          2386 => x"80",
          2387 => x"fa",
          2388 => x"7c",
          2389 => x"04",
          2390 => x"0b",
          2391 => x"fa",
          2392 => x"34",
          2393 => x"f8",
          2394 => x"bb",
          2395 => x"fe",
          2396 => x"e8",
          2397 => x"bb",
          2398 => x"f8",
          2399 => x"51",
          2400 => x"81",
          2401 => x"3d",
          2402 => x"33",
          2403 => x"33",
          2404 => x"12",
          2405 => x"b2",
          2406 => x"29",
          2407 => x"f9",
          2408 => x"57",
          2409 => x"89",
          2410 => x"81",
          2411 => x"38",
          2412 => x"b8",
          2413 => x"fa",
          2414 => x"56",
          2415 => x"c7",
          2416 => x"33",
          2417 => x"22",
          2418 => x"53",
          2419 => x"fa",
          2420 => x"54",
          2421 => x"80",
          2422 => x"81",
          2423 => x"fa",
          2424 => x"5b",
          2425 => x"84",
          2426 => x"81",
          2427 => x"81",
          2428 => x"77",
          2429 => x"83",
          2430 => x"53",
          2431 => x"fc",
          2432 => x"38",
          2433 => x"3d",
          2434 => x"75",
          2435 => x"2e",
          2436 => x"52",
          2437 => x"83",
          2438 => x"fa",
          2439 => x"13",
          2440 => x"81",
          2441 => x"52",
          2442 => x"70",
          2443 => x"26",
          2444 => x"fd",
          2445 => x"06",
          2446 => x"fe",
          2447 => x"fe",
          2448 => x"de",
          2449 => x"89",
          2450 => x"09",
          2451 => x"b5",
          2452 => x"05",
          2453 => x"83",
          2454 => x"fc",
          2455 => x"81",
          2456 => x"fe",
          2457 => x"b5",
          2458 => x"fa",
          2459 => x"e2",
          2460 => x"51",
          2461 => x"3d",
          2462 => x"ba",
          2463 => x"81",
          2464 => x"38",
          2465 => x"8a",
          2466 => x"84",
          2467 => x"38",
          2468 => x"33",
          2469 => x"05",
          2470 => x"33",
          2471 => x"b8",
          2472 => x"fa",
          2473 => x"5a",
          2474 => x"34",
          2475 => x"62",
          2476 => x"7f",
          2477 => x"b8",
          2478 => x"fa",
          2479 => x"72",
          2480 => x"83",
          2481 => x"34",
          2482 => x"58",
          2483 => x"b8",
          2484 => x"ff",
          2485 => x"80",
          2486 => x"0d",
          2487 => x"b7",
          2488 => x"2e",
          2489 => x"89",
          2490 => x"0c",
          2491 => x"33",
          2492 => x"05",
          2493 => x"33",
          2494 => x"b8",
          2495 => x"fa",
          2496 => x"5f",
          2497 => x"34",
          2498 => x"19",
          2499 => x"c7",
          2500 => x"33",
          2501 => x"22",
          2502 => x"11",
          2503 => x"b0",
          2504 => x"81",
          2505 => x"60",
          2506 => x"fa",
          2507 => x"0c",
          2508 => x"82",
          2509 => x"38",
          2510 => x"a8",
          2511 => x"80",
          2512 => x"0d",
          2513 => x"d0",
          2514 => x"38",
          2515 => x"57",
          2516 => x"ba",
          2517 => x"59",
          2518 => x"80",
          2519 => x"0d",
          2520 => x"80",
          2521 => x"f8",
          2522 => x"b5",
          2523 => x"40",
          2524 => x"a0",
          2525 => x"83",
          2526 => x"72",
          2527 => x"78",
          2528 => x"b4",
          2529 => x"83",
          2530 => x"1b",
          2531 => x"ff",
          2532 => x"b5",
          2533 => x"43",
          2534 => x"84",
          2535 => x"fe",
          2536 => x"fa",
          2537 => x"fe",
          2538 => x"fa",
          2539 => x"fa",
          2540 => x"c7",
          2541 => x"40",
          2542 => x"83",
          2543 => x"5a",
          2544 => x"86",
          2545 => x"1a",
          2546 => x"56",
          2547 => x"39",
          2548 => x"0b",
          2549 => x"ba",
          2550 => x"34",
          2551 => x"0b",
          2552 => x"04",
          2553 => x"34",
          2554 => x"34",
          2555 => x"34",
          2556 => x"0b",
          2557 => x"04",
          2558 => x"fa",
          2559 => x"b8",
          2560 => x"fa",
          2561 => x"75",
          2562 => x"83",
          2563 => x"29",
          2564 => x"f9",
          2565 => x"5b",
          2566 => x"78",
          2567 => x"75",
          2568 => x"b5",
          2569 => x"ff",
          2570 => x"29",
          2571 => x"33",
          2572 => x"b8",
          2573 => x"fa",
          2574 => x"5e",
          2575 => x"18",
          2576 => x"29",
          2577 => x"33",
          2578 => x"b8",
          2579 => x"fa",
          2580 => x"72",
          2581 => x"83",
          2582 => x"05",
          2583 => x"5c",
          2584 => x"84",
          2585 => x"38",
          2586 => x"34",
          2587 => x"06",
          2588 => x"78",
          2589 => x"2e",
          2590 => x"a8",
          2591 => x"83",
          2592 => x"b4",
          2593 => x"83",
          2594 => x"80",
          2595 => x"81",
          2596 => x"bb",
          2597 => x"fa",
          2598 => x"81",
          2599 => x"81",
          2600 => x"c7",
          2601 => x"5c",
          2602 => x"ff",
          2603 => x"53",
          2604 => x"2e",
          2605 => x"ff",
          2606 => x"ff",
          2607 => x"40",
          2608 => x"80",
          2609 => x"fa",
          2610 => x"71",
          2611 => x"0b",
          2612 => x"b4",
          2613 => x"83",
          2614 => x"1a",
          2615 => x"ff",
          2616 => x"b5",
          2617 => x"5a",
          2618 => x"99",
          2619 => x"81",
          2620 => x"81",
          2621 => x"77",
          2622 => x"83",
          2623 => x"ff",
          2624 => x"a7",
          2625 => x"f8",
          2626 => x"ff",
          2627 => x"ff",
          2628 => x"43",
          2629 => x"86",
          2630 => x"f8",
          2631 => x"b2",
          2632 => x"5e",
          2633 => x"34",
          2634 => x"1e",
          2635 => x"c7",
          2636 => x"33",
          2637 => x"22",
          2638 => x"11",
          2639 => x"b0",
          2640 => x"81",
          2641 => x"79",
          2642 => x"fa",
          2643 => x"84",
          2644 => x"84",
          2645 => x"b6",
          2646 => x"33",
          2647 => x"81",
          2648 => x"ca",
          2649 => x"80",
          2650 => x"0d",
          2651 => x"84",
          2652 => x"fa",
          2653 => x"fa",
          2654 => x"fc",
          2655 => x"3d",
          2656 => x"88",
          2657 => x"2e",
          2658 => x"81",
          2659 => x"34",
          2660 => x"80",
          2661 => x"05",
          2662 => x"17",
          2663 => x"7b",
          2664 => x"f8",
          2665 => x"5c",
          2666 => x"83",
          2667 => x"72",
          2668 => x"b9",
          2669 => x"80",
          2670 => x"fa",
          2671 => x"71",
          2672 => x"83",
          2673 => x"33",
          2674 => x"fa",
          2675 => x"05",
          2676 => x"ff",
          2677 => x"b5",
          2678 => x"5a",
          2679 => x"99",
          2680 => x"ff",
          2681 => x"a2",
          2682 => x"90",
          2683 => x"fa",
          2684 => x"0c",
          2685 => x"2e",
          2686 => x"56",
          2687 => x"51",
          2688 => x"84",
          2689 => x"ec",
          2690 => x"ed",
          2691 => x"ee",
          2692 => x"ff",
          2693 => x"ba",
          2694 => x"ba",
          2695 => x"ba",
          2696 => x"85",
          2697 => x"38",
          2698 => x"2e",
          2699 => x"fa",
          2700 => x"b4",
          2701 => x"e5",
          2702 => x"fe",
          2703 => x"aa",
          2704 => x"06",
          2705 => x"41",
          2706 => x"52",
          2707 => x"3f",
          2708 => x"85",
          2709 => x"5b",
          2710 => x"10",
          2711 => x"57",
          2712 => x"75",
          2713 => x"7e",
          2714 => x"7d",
          2715 => x"b4",
          2716 => x"31",
          2717 => x"5a",
          2718 => x"b4",
          2719 => x"33",
          2720 => x"84",
          2721 => x"ff",
          2722 => x"5f",
          2723 => x"83",
          2724 => x"0b",
          2725 => x"33",
          2726 => x"80",
          2727 => x"75",
          2728 => x"80",
          2729 => x"b4",
          2730 => x"57",
          2731 => x"81",
          2732 => x"fc",
          2733 => x"7f",
          2734 => x"b5",
          2735 => x"31",
          2736 => x"5a",
          2737 => x"b5",
          2738 => x"33",
          2739 => x"84",
          2740 => x"09",
          2741 => x"f8",
          2742 => x"b4",
          2743 => x"a0",
          2744 => x"51",
          2745 => x"83",
          2746 => x"87",
          2747 => x"5d",
          2748 => x"38",
          2749 => x"f2",
          2750 => x"80",
          2751 => x"22",
          2752 => x"fb",
          2753 => x"34",
          2754 => x"56",
          2755 => x"ba",
          2756 => x"7c",
          2757 => x"59",
          2758 => x"75",
          2759 => x"a2",
          2760 => x"80",
          2761 => x"33",
          2762 => x"84",
          2763 => x"56",
          2764 => x"76",
          2765 => x"83",
          2766 => x"80",
          2767 => x"76",
          2768 => x"84",
          2769 => x"83",
          2770 => x"81",
          2771 => x"85",
          2772 => x"0b",
          2773 => x"80",
          2774 => x"56",
          2775 => x"81",
          2776 => x"f3",
          2777 => x"33",
          2778 => x"84",
          2779 => x"ff",
          2780 => x"70",
          2781 => x"70",
          2782 => x"52",
          2783 => x"83",
          2784 => x"23",
          2785 => x"5f",
          2786 => x"76",
          2787 => x"33",
          2788 => x"f9",
          2789 => x"b5",
          2790 => x"33",
          2791 => x"84",
          2792 => x"40",
          2793 => x"83",
          2794 => x"70",
          2795 => x"71",
          2796 => x"05",
          2797 => x"7e",
          2798 => x"83",
          2799 => x"5f",
          2800 => x"79",
          2801 => x"5d",
          2802 => x"84",
          2803 => x"8e",
          2804 => x"fa",
          2805 => x"7c",
          2806 => x"e5",
          2807 => x"76",
          2808 => x"75",
          2809 => x"06",
          2810 => x"5a",
          2811 => x"31",
          2812 => x"71",
          2813 => x"c7",
          2814 => x"7f",
          2815 => x"71",
          2816 => x"79",
          2817 => x"d6",
          2818 => x"84",
          2819 => x"05",
          2820 => x"33",
          2821 => x"18",
          2822 => x"33",
          2823 => x"58",
          2824 => x"e0",
          2825 => x"33",
          2826 => x"70",
          2827 => x"05",
          2828 => x"33",
          2829 => x"1d",
          2830 => x"ff",
          2831 => x"85",
          2832 => x"38",
          2833 => x"d8",
          2834 => x"84",
          2835 => x"85",
          2836 => x"2e",
          2837 => x"75",
          2838 => x"38",
          2839 => x"ff",
          2840 => x"5c",
          2841 => x"84",
          2842 => x"f6",
          2843 => x"60",
          2844 => x"26",
          2845 => x"f2",
          2846 => x"29",
          2847 => x"70",
          2848 => x"05",
          2849 => x"8b",
          2850 => x"8b",
          2851 => x"98",
          2852 => x"2b",
          2853 => x"5f",
          2854 => x"77",
          2855 => x"70",
          2856 => x"ee",
          2857 => x"f7",
          2858 => x"60",
          2859 => x"7d",
          2860 => x"5a",
          2861 => x"31",
          2862 => x"40",
          2863 => x"26",
          2864 => x"84",
          2865 => x"e0",
          2866 => x"05",
          2867 => x"26",
          2868 => x"19",
          2869 => x"34",
          2870 => x"38",
          2871 => x"ff",
          2872 => x"fa",
          2873 => x"84",
          2874 => x"07",
          2875 => x"09",
          2876 => x"83",
          2877 => x"ff",
          2878 => x"fa",
          2879 => x"1e",
          2880 => x"84",
          2881 => x"84",
          2882 => x"fa",
          2883 => x"07",
          2884 => x"18",
          2885 => x"fb",
          2886 => x"06",
          2887 => x"34",
          2888 => x"fb",
          2889 => x"b0",
          2890 => x"81",
          2891 => x"fa",
          2892 => x"33",
          2893 => x"83",
          2894 => x"f1",
          2895 => x"70",
          2896 => x"39",
          2897 => x"56",
          2898 => x"39",
          2899 => x"90",
          2900 => x"fe",
          2901 => x"ef",
          2902 => x"fa",
          2903 => x"b0",
          2904 => x"56",
          2905 => x"39",
          2906 => x"a0",
          2907 => x"fe",
          2908 => x"fe",
          2909 => x"b0",
          2910 => x"33",
          2911 => x"83",
          2912 => x"fa",
          2913 => x"56",
          2914 => x"39",
          2915 => x"56",
          2916 => x"39",
          2917 => x"56",
          2918 => x"39",
          2919 => x"56",
          2920 => x"39",
          2921 => x"80",
          2922 => x"34",
          2923 => x"81",
          2924 => x"fa",
          2925 => x"83",
          2926 => x"d2",
          2927 => x"ec",
          2928 => x"ed",
          2929 => x"ee",
          2930 => x"80",
          2931 => x"39",
          2932 => x"0b",
          2933 => x"04",
          2934 => x"b5",
          2935 => x"05",
          2936 => x"42",
          2937 => x"51",
          2938 => x"08",
          2939 => x"ba",
          2940 => x"34",
          2941 => x"3d",
          2942 => x"ef",
          2943 => x"11",
          2944 => x"7b",
          2945 => x"ca",
          2946 => x"80",
          2947 => x"80",
          2948 => x"81",
          2949 => x"33",
          2950 => x"56",
          2951 => x"b5",
          2952 => x"3f",
          2953 => x"90",
          2954 => x"33",
          2955 => x"72",
          2956 => x"75",
          2957 => x"f8",
          2958 => x"38",
          2959 => x"39",
          2960 => x"09",
          2961 => x"57",
          2962 => x"81",
          2963 => x"59",
          2964 => x"38",
          2965 => x"f7",
          2966 => x"81",
          2967 => x"b4",
          2968 => x"ff",
          2969 => x"29",
          2970 => x"fa",
          2971 => x"05",
          2972 => x"8a",
          2973 => x"77",
          2974 => x"ff",
          2975 => x"7b",
          2976 => x"33",
          2977 => x"ff",
          2978 => x"7c",
          2979 => x"80",
          2980 => x"f7",
          2981 => x"38",
          2982 => x"34",
          2983 => x"22",
          2984 => x"90",
          2985 => x"81",
          2986 => x"5f",
          2987 => x"86",
          2988 => x"7f",
          2989 => x"41",
          2990 => x"ea",
          2991 => x"e0",
          2992 => x"33",
          2993 => x"70",
          2994 => x"05",
          2995 => x"33",
          2996 => x"1d",
          2997 => x"ec",
          2998 => x"84",
          2999 => x"05",
          3000 => x"33",
          3001 => x"18",
          3002 => x"33",
          3003 => x"58",
          3004 => x"fa",
          3005 => x"84",
          3006 => x"fa",
          3007 => x"fa",
          3008 => x"5c",
          3009 => x"d2",
          3010 => x"ff",
          3011 => x"61",
          3012 => x"fa",
          3013 => x"19",
          3014 => x"80",
          3015 => x"b8",
          3016 => x"12",
          3017 => x"8d",
          3018 => x"34",
          3019 => x"81",
          3020 => x"59",
          3021 => x"38",
          3022 => x"2e",
          3023 => x"fa",
          3024 => x"fa",
          3025 => x"76",
          3026 => x"38",
          3027 => x"83",
          3028 => x"1a",
          3029 => x"e7",
          3030 => x"fa",
          3031 => x"58",
          3032 => x"80",
          3033 => x"fa",
          3034 => x"34",
          3035 => x"76",
          3036 => x"b0",
          3037 => x"79",
          3038 => x"79",
          3039 => x"23",
          3040 => x"b4",
          3041 => x"b2",
          3042 => x"fa",
          3043 => x"83",
          3044 => x"fa",
          3045 => x"1a",
          3046 => x"89",
          3047 => x"02",
          3048 => x"54",
          3049 => x"51",
          3050 => x"84",
          3051 => x"73",
          3052 => x"bb",
          3053 => x"3d",
          3054 => x"0b",
          3055 => x"06",
          3056 => x"55",
          3057 => x"81",
          3058 => x"74",
          3059 => x"3d",
          3060 => x"82",
          3061 => x"73",
          3062 => x"70",
          3063 => x"83",
          3064 => x"7b",
          3065 => x"7b",
          3066 => x"80",
          3067 => x"80",
          3068 => x"33",
          3069 => x"33",
          3070 => x"80",
          3071 => x"5d",
          3072 => x"ff",
          3073 => x"55",
          3074 => x"81",
          3075 => x"34",
          3076 => x"87",
          3077 => x"2e",
          3078 => x"57",
          3079 => x"14",
          3080 => x"f9",
          3081 => x"f8",
          3082 => x"83",
          3083 => x"72",
          3084 => x"ff",
          3085 => x"b8",
          3086 => x"79",
          3087 => x"83",
          3088 => x"14",
          3089 => x"14",
          3090 => x"74",
          3091 => x"33",
          3092 => x"56",
          3093 => x"81",
          3094 => x"70",
          3095 => x"2e",
          3096 => x"dd",
          3097 => x"80",
          3098 => x"f8",
          3099 => x"33",
          3100 => x"33",
          3101 => x"df",
          3102 => x"56",
          3103 => x"81",
          3104 => x"16",
          3105 => x"38",
          3106 => x"81",
          3107 => x"16",
          3108 => x"81",
          3109 => x"8d",
          3110 => x"72",
          3111 => x"ff",
          3112 => x"8c",
          3113 => x"81",
          3114 => x"d8",
          3115 => x"9c",
          3116 => x"ec",
          3117 => x"08",
          3118 => x"70",
          3119 => x"27",
          3120 => x"34",
          3121 => x"19",
          3122 => x"72",
          3123 => x"79",
          3124 => x"73",
          3125 => x"87",
          3126 => x"7d",
          3127 => x"f9",
          3128 => x"83",
          3129 => x"34",
          3130 => x"8c",
          3131 => x"81",
          3132 => x"33",
          3133 => x"34",
          3134 => x"f8",
          3135 => x"9c",
          3136 => x"80",
          3137 => x"8a",
          3138 => x"74",
          3139 => x"9b",
          3140 => x"83",
          3141 => x"38",
          3142 => x"81",
          3143 => x"98",
          3144 => x"38",
          3145 => x"70",
          3146 => x"06",
          3147 => x"53",
          3148 => x"38",
          3149 => x"76",
          3150 => x"94",
          3151 => x"87",
          3152 => x"0c",
          3153 => x"81",
          3154 => x"06",
          3155 => x"9b",
          3156 => x"80",
          3157 => x"72",
          3158 => x"32",
          3159 => x"40",
          3160 => x"2e",
          3161 => x"ff",
          3162 => x"10",
          3163 => x"33",
          3164 => x"38",
          3165 => x"57",
          3166 => x"fb",
          3167 => x"38",
          3168 => x"91",
          3169 => x"51",
          3170 => x"0c",
          3171 => x"81",
          3172 => x"ff",
          3173 => x"33",
          3174 => x"15",
          3175 => x"f8",
          3176 => x"b8",
          3177 => x"15",
          3178 => x"06",
          3179 => x"38",
          3180 => x"75",
          3181 => x"06",
          3182 => x"fb",
          3183 => x"fa",
          3184 => x"55",
          3185 => x"c0",
          3186 => x"76",
          3187 => x"ff",
          3188 => x"ca",
          3189 => x"09",
          3190 => x"72",
          3191 => x"f8",
          3192 => x"f8",
          3193 => x"83",
          3194 => x"5c",
          3195 => x"2e",
          3196 => x"59",
          3197 => x"81",
          3198 => x"fd",
          3199 => x"54",
          3200 => x"fb",
          3201 => x"54",
          3202 => x"f7",
          3203 => x"33",
          3204 => x"73",
          3205 => x"95",
          3206 => x"84",
          3207 => x"f8",
          3208 => x"f7",
          3209 => x"57",
          3210 => x"80",
          3211 => x"81",
          3212 => x"73",
          3213 => x"fa",
          3214 => x"81",
          3215 => x"75",
          3216 => x"fa",
          3217 => x"81",
          3218 => x"ff",
          3219 => x"95",
          3220 => x"e8",
          3221 => x"83",
          3222 => x"59",
          3223 => x"51",
          3224 => x"fa",
          3225 => x"08",
          3226 => x"13",
          3227 => x"e0",
          3228 => x"08",
          3229 => x"80",
          3230 => x"c0",
          3231 => x"55",
          3232 => x"98",
          3233 => x"08",
          3234 => x"14",
          3235 => x"52",
          3236 => x"fe",
          3237 => x"08",
          3238 => x"c8",
          3239 => x"c0",
          3240 => x"ce",
          3241 => x"08",
          3242 => x"74",
          3243 => x"87",
          3244 => x"73",
          3245 => x"db",
          3246 => x"72",
          3247 => x"55",
          3248 => x"53",
          3249 => x"ff",
          3250 => x"ff",
          3251 => x"0c",
          3252 => x"bb",
          3253 => x"3d",
          3254 => x"33",
          3255 => x"08",
          3256 => x"06",
          3257 => x"55",
          3258 => x"2a",
          3259 => x"2a",
          3260 => x"15",
          3261 => x"82",
          3262 => x"80",
          3263 => x"90",
          3264 => x"34",
          3265 => x"87",
          3266 => x"08",
          3267 => x"c0",
          3268 => x"9c",
          3269 => x"81",
          3270 => x"56",
          3271 => x"81",
          3272 => x"a4",
          3273 => x"80",
          3274 => x"80",
          3275 => x"80",
          3276 => x"9c",
          3277 => x"55",
          3278 => x"33",
          3279 => x"70",
          3280 => x"2e",
          3281 => x"55",
          3282 => x"71",
          3283 => x"57",
          3284 => x"74",
          3285 => x"38",
          3286 => x"75",
          3287 => x"80",
          3288 => x"92",
          3289 => x"71",
          3290 => x"26",
          3291 => x"88",
          3292 => x"84",
          3293 => x"c2",
          3294 => x"05",
          3295 => x"83",
          3296 => x"fc",
          3297 => x"07",
          3298 => x"34",
          3299 => x"34",
          3300 => x"34",
          3301 => x"90",
          3302 => x"56",
          3303 => x"38",
          3304 => x"70",
          3305 => x"f0",
          3306 => x"82",
          3307 => x"80",
          3308 => x"90",
          3309 => x"34",
          3310 => x"87",
          3311 => x"08",
          3312 => x"c0",
          3313 => x"9c",
          3314 => x"81",
          3315 => x"56",
          3316 => x"81",
          3317 => x"a4",
          3318 => x"80",
          3319 => x"80",
          3320 => x"80",
          3321 => x"9c",
          3322 => x"55",
          3323 => x"33",
          3324 => x"70",
          3325 => x"2e",
          3326 => x"55",
          3327 => x"71",
          3328 => x"57",
          3329 => x"81",
          3330 => x"74",
          3331 => x"80",
          3332 => x"bb",
          3333 => x"51",
          3334 => x"90",
          3335 => x"0b",
          3336 => x"0b",
          3337 => x"80",
          3338 => x"83",
          3339 => x"05",
          3340 => x"87",
          3341 => x"2e",
          3342 => x"98",
          3343 => x"87",
          3344 => x"87",
          3345 => x"70",
          3346 => x"71",
          3347 => x"98",
          3348 => x"87",
          3349 => x"98",
          3350 => x"38",
          3351 => x"08",
          3352 => x"71",
          3353 => x"98",
          3354 => x"38",
          3355 => x"81",
          3356 => x"8a",
          3357 => x"fe",
          3358 => x"83",
          3359 => x"82",
          3360 => x"ba",
          3361 => x"70",
          3362 => x"73",
          3363 => x"8b",
          3364 => x"70",
          3365 => x"71",
          3366 => x"53",
          3367 => x"80",
          3368 => x"82",
          3369 => x"2b",
          3370 => x"33",
          3371 => x"90",
          3372 => x"56",
          3373 => x"84",
          3374 => x"2b",
          3375 => x"88",
          3376 => x"13",
          3377 => x"87",
          3378 => x"17",
          3379 => x"88",
          3380 => x"59",
          3381 => x"85",
          3382 => x"52",
          3383 => x"87",
          3384 => x"74",
          3385 => x"84",
          3386 => x"12",
          3387 => x"80",
          3388 => x"52",
          3389 => x"89",
          3390 => x"13",
          3391 => x"07",
          3392 => x"33",
          3393 => x"58",
          3394 => x"84",
          3395 => x"ba",
          3396 => x"85",
          3397 => x"2b",
          3398 => x"86",
          3399 => x"2b",
          3400 => x"52",
          3401 => x"34",
          3402 => x"81",
          3403 => x"ff",
          3404 => x"54",
          3405 => x"34",
          3406 => x"33",
          3407 => x"83",
          3408 => x"12",
          3409 => x"2b",
          3410 => x"88",
          3411 => x"57",
          3412 => x"83",
          3413 => x"17",
          3414 => x"2b",
          3415 => x"33",
          3416 => x"81",
          3417 => x"52",
          3418 => x"73",
          3419 => x"f4",
          3420 => x"12",
          3421 => x"07",
          3422 => x"71",
          3423 => x"53",
          3424 => x"80",
          3425 => x"13",
          3426 => x"80",
          3427 => x"76",
          3428 => x"ba",
          3429 => x"12",
          3430 => x"07",
          3431 => x"33",
          3432 => x"57",
          3433 => x"72",
          3434 => x"89",
          3435 => x"84",
          3436 => x"2e",
          3437 => x"77",
          3438 => x"04",
          3439 => x"0c",
          3440 => x"82",
          3441 => x"f4",
          3442 => x"f4",
          3443 => x"81",
          3444 => x"76",
          3445 => x"34",
          3446 => x"17",
          3447 => x"ba",
          3448 => x"05",
          3449 => x"ff",
          3450 => x"56",
          3451 => x"34",
          3452 => x"10",
          3453 => x"55",
          3454 => x"83",
          3455 => x"0d",
          3456 => x"72",
          3457 => x"82",
          3458 => x"51",
          3459 => x"f4",
          3460 => x"71",
          3461 => x"58",
          3462 => x"2e",
          3463 => x"17",
          3464 => x"2b",
          3465 => x"31",
          3466 => x"27",
          3467 => x"74",
          3468 => x"38",
          3469 => x"85",
          3470 => x"5a",
          3471 => x"2e",
          3472 => x"76",
          3473 => x"12",
          3474 => x"ff",
          3475 => x"59",
          3476 => x"80",
          3477 => x"78",
          3478 => x"72",
          3479 => x"70",
          3480 => x"80",
          3481 => x"56",
          3482 => x"34",
          3483 => x"2a",
          3484 => x"83",
          3485 => x"19",
          3486 => x"2b",
          3487 => x"06",
          3488 => x"70",
          3489 => x"52",
          3490 => x"ff",
          3491 => x"ba",
          3492 => x"72",
          3493 => x"70",
          3494 => x"71",
          3495 => x"05",
          3496 => x"15",
          3497 => x"f4",
          3498 => x"11",
          3499 => x"07",
          3500 => x"70",
          3501 => x"84",
          3502 => x"33",
          3503 => x"83",
          3504 => x"5a",
          3505 => x"15",
          3506 => x"55",
          3507 => x"33",
          3508 => x"54",
          3509 => x"79",
          3510 => x"18",
          3511 => x"0c",
          3512 => x"87",
          3513 => x"2b",
          3514 => x"18",
          3515 => x"2a",
          3516 => x"84",
          3517 => x"ba",
          3518 => x"85",
          3519 => x"2b",
          3520 => x"15",
          3521 => x"2a",
          3522 => x"52",
          3523 => x"34",
          3524 => x"81",
          3525 => x"ff",
          3526 => x"54",
          3527 => x"34",
          3528 => x"51",
          3529 => x"84",
          3530 => x"2e",
          3531 => x"73",
          3532 => x"04",
          3533 => x"84",
          3534 => x"0d",
          3535 => x"f4",
          3536 => x"23",
          3537 => x"ff",
          3538 => x"ba",
          3539 => x"0b",
          3540 => x"54",
          3541 => x"15",
          3542 => x"86",
          3543 => x"84",
          3544 => x"ff",
          3545 => x"ff",
          3546 => x"55",
          3547 => x"17",
          3548 => x"10",
          3549 => x"05",
          3550 => x"0b",
          3551 => x"2e",
          3552 => x"3d",
          3553 => x"84",
          3554 => x"61",
          3555 => x"85",
          3556 => x"38",
          3557 => x"7f",
          3558 => x"83",
          3559 => x"ff",
          3560 => x"70",
          3561 => x"7a",
          3562 => x"88",
          3563 => x"ff",
          3564 => x"05",
          3565 => x"81",
          3566 => x"90",
          3567 => x"46",
          3568 => x"59",
          3569 => x"85",
          3570 => x"33",
          3571 => x"10",
          3572 => x"98",
          3573 => x"53",
          3574 => x"c9",
          3575 => x"63",
          3576 => x"38",
          3577 => x"1b",
          3578 => x"63",
          3579 => x"38",
          3580 => x"71",
          3581 => x"11",
          3582 => x"2b",
          3583 => x"52",
          3584 => x"8c",
          3585 => x"83",
          3586 => x"2b",
          3587 => x"12",
          3588 => x"07",
          3589 => x"33",
          3590 => x"59",
          3591 => x"5c",
          3592 => x"85",
          3593 => x"17",
          3594 => x"8b",
          3595 => x"86",
          3596 => x"2b",
          3597 => x"52",
          3598 => x"34",
          3599 => x"08",
          3600 => x"88",
          3601 => x"88",
          3602 => x"34",
          3603 => x"08",
          3604 => x"33",
          3605 => x"74",
          3606 => x"88",
          3607 => x"45",
          3608 => x"34",
          3609 => x"08",
          3610 => x"71",
          3611 => x"05",
          3612 => x"88",
          3613 => x"45",
          3614 => x"1a",
          3615 => x"f4",
          3616 => x"12",
          3617 => x"62",
          3618 => x"5d",
          3619 => x"a4",
          3620 => x"05",
          3621 => x"ff",
          3622 => x"81",
          3623 => x"84",
          3624 => x"f4",
          3625 => x"0b",
          3626 => x"53",
          3627 => x"c6",
          3628 => x"60",
          3629 => x"84",
          3630 => x"34",
          3631 => x"f4",
          3632 => x"0b",
          3633 => x"84",
          3634 => x"80",
          3635 => x"88",
          3636 => x"18",
          3637 => x"f0",
          3638 => x"f4",
          3639 => x"82",
          3640 => x"84",
          3641 => x"38",
          3642 => x"54",
          3643 => x"51",
          3644 => x"84",
          3645 => x"61",
          3646 => x"2b",
          3647 => x"33",
          3648 => x"81",
          3649 => x"44",
          3650 => x"81",
          3651 => x"05",
          3652 => x"19",
          3653 => x"f4",
          3654 => x"33",
          3655 => x"8f",
          3656 => x"ff",
          3657 => x"47",
          3658 => x"05",
          3659 => x"63",
          3660 => x"1e",
          3661 => x"34",
          3662 => x"05",
          3663 => x"bc",
          3664 => x"ff",
          3665 => x"81",
          3666 => x"ff",
          3667 => x"33",
          3668 => x"10",
          3669 => x"98",
          3670 => x"53",
          3671 => x"25",
          3672 => x"78",
          3673 => x"8b",
          3674 => x"5b",
          3675 => x"8f",
          3676 => x"f4",
          3677 => x"23",
          3678 => x"ff",
          3679 => x"ba",
          3680 => x"0b",
          3681 => x"59",
          3682 => x"1a",
          3683 => x"86",
          3684 => x"84",
          3685 => x"ff",
          3686 => x"ff",
          3687 => x"57",
          3688 => x"64",
          3689 => x"70",
          3690 => x"05",
          3691 => x"05",
          3692 => x"ee",
          3693 => x"61",
          3694 => x"27",
          3695 => x"80",
          3696 => x"fb",
          3697 => x"0c",
          3698 => x"11",
          3699 => x"71",
          3700 => x"33",
          3701 => x"83",
          3702 => x"85",
          3703 => x"88",
          3704 => x"58",
          3705 => x"05",
          3706 => x"ba",
          3707 => x"85",
          3708 => x"2b",
          3709 => x"15",
          3710 => x"2a",
          3711 => x"41",
          3712 => x"87",
          3713 => x"70",
          3714 => x"07",
          3715 => x"5f",
          3716 => x"81",
          3717 => x"1f",
          3718 => x"8b",
          3719 => x"73",
          3720 => x"07",
          3721 => x"43",
          3722 => x"81",
          3723 => x"1f",
          3724 => x"2b",
          3725 => x"14",
          3726 => x"07",
          3727 => x"40",
          3728 => x"60",
          3729 => x"70",
          3730 => x"71",
          3731 => x"70",
          3732 => x"05",
          3733 => x"84",
          3734 => x"83",
          3735 => x"39",
          3736 => x"0c",
          3737 => x"82",
          3738 => x"f4",
          3739 => x"f4",
          3740 => x"81",
          3741 => x"7f",
          3742 => x"34",
          3743 => x"15",
          3744 => x"ba",
          3745 => x"05",
          3746 => x"ff",
          3747 => x"5e",
          3748 => x"34",
          3749 => x"10",
          3750 => x"5c",
          3751 => x"83",
          3752 => x"7f",
          3753 => x"87",
          3754 => x"2b",
          3755 => x"1d",
          3756 => x"2a",
          3757 => x"61",
          3758 => x"34",
          3759 => x"11",
          3760 => x"71",
          3761 => x"33",
          3762 => x"70",
          3763 => x"56",
          3764 => x"78",
          3765 => x"08",
          3766 => x"88",
          3767 => x"88",
          3768 => x"34",
          3769 => x"08",
          3770 => x"71",
          3771 => x"05",
          3772 => x"2b",
          3773 => x"06",
          3774 => x"5d",
          3775 => x"82",
          3776 => x"ba",
          3777 => x"12",
          3778 => x"07",
          3779 => x"71",
          3780 => x"70",
          3781 => x"5a",
          3782 => x"81",
          3783 => x"5b",
          3784 => x"16",
          3785 => x"07",
          3786 => x"33",
          3787 => x"5e",
          3788 => x"1e",
          3789 => x"f4",
          3790 => x"12",
          3791 => x"07",
          3792 => x"33",
          3793 => x"44",
          3794 => x"7c",
          3795 => x"05",
          3796 => x"33",
          3797 => x"81",
          3798 => x"5b",
          3799 => x"16",
          3800 => x"70",
          3801 => x"71",
          3802 => x"81",
          3803 => x"83",
          3804 => x"63",
          3805 => x"59",
          3806 => x"7b",
          3807 => x"70",
          3808 => x"8b",
          3809 => x"70",
          3810 => x"07",
          3811 => x"5d",
          3812 => x"75",
          3813 => x"ba",
          3814 => x"83",
          3815 => x"2b",
          3816 => x"12",
          3817 => x"07",
          3818 => x"33",
          3819 => x"59",
          3820 => x"5d",
          3821 => x"79",
          3822 => x"70",
          3823 => x"71",
          3824 => x"05",
          3825 => x"88",
          3826 => x"5e",
          3827 => x"16",
          3828 => x"f4",
          3829 => x"71",
          3830 => x"70",
          3831 => x"79",
          3832 => x"f4",
          3833 => x"12",
          3834 => x"07",
          3835 => x"71",
          3836 => x"5c",
          3837 => x"79",
          3838 => x"f4",
          3839 => x"33",
          3840 => x"74",
          3841 => x"71",
          3842 => x"5c",
          3843 => x"82",
          3844 => x"ba",
          3845 => x"83",
          3846 => x"57",
          3847 => x"5a",
          3848 => x"b4",
          3849 => x"84",
          3850 => x"ff",
          3851 => x"39",
          3852 => x"8b",
          3853 => x"84",
          3854 => x"2b",
          3855 => x"43",
          3856 => x"63",
          3857 => x"08",
          3858 => x"33",
          3859 => x"74",
          3860 => x"71",
          3861 => x"41",
          3862 => x"64",
          3863 => x"34",
          3864 => x"81",
          3865 => x"ff",
          3866 => x"42",
          3867 => x"34",
          3868 => x"33",
          3869 => x"83",
          3870 => x"12",
          3871 => x"2b",
          3872 => x"88",
          3873 => x"45",
          3874 => x"83",
          3875 => x"1f",
          3876 => x"2b",
          3877 => x"33",
          3878 => x"81",
          3879 => x"5f",
          3880 => x"7d",
          3881 => x"ff",
          3882 => x"60",
          3883 => x"84",
          3884 => x"2e",
          3885 => x"bb",
          3886 => x"73",
          3887 => x"7b",
          3888 => x"f9",
          3889 => x"f4",
          3890 => x"38",
          3891 => x"bb",
          3892 => x"51",
          3893 => x"54",
          3894 => x"38",
          3895 => x"08",
          3896 => x"bb",
          3897 => x"ff",
          3898 => x"80",
          3899 => x"80",
          3900 => x"fe",
          3901 => x"55",
          3902 => x"34",
          3903 => x"15",
          3904 => x"ba",
          3905 => x"81",
          3906 => x"08",
          3907 => x"80",
          3908 => x"70",
          3909 => x"88",
          3910 => x"ba",
          3911 => x"ba",
          3912 => x"76",
          3913 => x"34",
          3914 => x"38",
          3915 => x"8f",
          3916 => x"26",
          3917 => x"52",
          3918 => x"0d",
          3919 => x"33",
          3920 => x"38",
          3921 => x"84",
          3922 => x"38",
          3923 => x"bb",
          3924 => x"84",
          3925 => x"0d",
          3926 => x"05",
          3927 => x"76",
          3928 => x"17",
          3929 => x"55",
          3930 => x"87",
          3931 => x"52",
          3932 => x"84",
          3933 => x"2e",
          3934 => x"54",
          3935 => x"38",
          3936 => x"80",
          3937 => x"74",
          3938 => x"04",
          3939 => x"ff",
          3940 => x"ff",
          3941 => x"7c",
          3942 => x"33",
          3943 => x"74",
          3944 => x"33",
          3945 => x"73",
          3946 => x"c0",
          3947 => x"76",
          3948 => x"08",
          3949 => x"a7",
          3950 => x"73",
          3951 => x"74",
          3952 => x"2e",
          3953 => x"84",
          3954 => x"84",
          3955 => x"06",
          3956 => x"ac",
          3957 => x"02",
          3958 => x"05",
          3959 => x"53",
          3960 => x"80",
          3961 => x"83",
          3962 => x"c0",
          3963 => x"2e",
          3964 => x"70",
          3965 => x"84",
          3966 => x"88",
          3967 => x"84",
          3968 => x"75",
          3969 => x"86",
          3970 => x"c0",
          3971 => x"38",
          3972 => x"51",
          3973 => x"c0",
          3974 => x"87",
          3975 => x"38",
          3976 => x"14",
          3977 => x"80",
          3978 => x"06",
          3979 => x"f6",
          3980 => x"19",
          3981 => x"2e",
          3982 => x"56",
          3983 => x"53",
          3984 => x"a3",
          3985 => x"83",
          3986 => x"0c",
          3987 => x"18",
          3988 => x"19",
          3989 => x"59",
          3990 => x"81",
          3991 => x"83",
          3992 => x"1a",
          3993 => x"84",
          3994 => x"27",
          3995 => x"74",
          3996 => x"38",
          3997 => x"81",
          3998 => x"78",
          3999 => x"81",
          4000 => x"57",
          4001 => x"ee",
          4002 => x"56",
          4003 => x"34",
          4004 => x"d5",
          4005 => x"0b",
          4006 => x"34",
          4007 => x"e1",
          4008 => x"bb",
          4009 => x"19",
          4010 => x"34",
          4011 => x"80",
          4012 => x"18",
          4013 => x"74",
          4014 => x"34",
          4015 => x"19",
          4016 => x"a3",
          4017 => x"84",
          4018 => x"74",
          4019 => x"56",
          4020 => x"2a",
          4021 => x"18",
          4022 => x"5b",
          4023 => x"18",
          4024 => x"19",
          4025 => x"33",
          4026 => x"08",
          4027 => x"39",
          4028 => x"59",
          4029 => x"9c",
          4030 => x"58",
          4031 => x"0d",
          4032 => x"82",
          4033 => x"82",
          4034 => x"06",
          4035 => x"89",
          4036 => x"80",
          4037 => x"38",
          4038 => x"09",
          4039 => x"78",
          4040 => x"51",
          4041 => x"80",
          4042 => x"78",
          4043 => x"79",
          4044 => x"81",
          4045 => x"05",
          4046 => x"79",
          4047 => x"33",
          4048 => x"09",
          4049 => x"78",
          4050 => x"51",
          4051 => x"80",
          4052 => x"78",
          4053 => x"7a",
          4054 => x"70",
          4055 => x"71",
          4056 => x"79",
          4057 => x"84",
          4058 => x"75",
          4059 => x"b4",
          4060 => x"0b",
          4061 => x"7b",
          4062 => x"38",
          4063 => x"81",
          4064 => x"bb",
          4065 => x"59",
          4066 => x"fd",
          4067 => x"77",
          4068 => x"33",
          4069 => x"0c",
          4070 => x"83",
          4071 => x"75",
          4072 => x"b4",
          4073 => x"0b",
          4074 => x"7c",
          4075 => x"38",
          4076 => x"81",
          4077 => x"bb",
          4078 => x"59",
          4079 => x"fc",
          4080 => x"06",
          4081 => x"82",
          4082 => x"2b",
          4083 => x"88",
          4084 => x"fe",
          4085 => x"41",
          4086 => x"0d",
          4087 => x"b8",
          4088 => x"5c",
          4089 => x"84",
          4090 => x"be",
          4091 => x"34",
          4092 => x"84",
          4093 => x"18",
          4094 => x"33",
          4095 => x"fd",
          4096 => x"a0",
          4097 => x"17",
          4098 => x"fd",
          4099 => x"53",
          4100 => x"52",
          4101 => x"08",
          4102 => x"38",
          4103 => x"b4",
          4104 => x"7c",
          4105 => x"17",
          4106 => x"38",
          4107 => x"39",
          4108 => x"17",
          4109 => x"f5",
          4110 => x"08",
          4111 => x"38",
          4112 => x"b4",
          4113 => x"bb",
          4114 => x"08",
          4115 => x"55",
          4116 => x"b8",
          4117 => x"18",
          4118 => x"33",
          4119 => x"a0",
          4120 => x"b8",
          4121 => x"5e",
          4122 => x"84",
          4123 => x"cb",
          4124 => x"34",
          4125 => x"84",
          4126 => x"18",
          4127 => x"33",
          4128 => x"fb",
          4129 => x"a0",
          4130 => x"17",
          4131 => x"fa",
          4132 => x"a0",
          4133 => x"17",
          4134 => x"39",
          4135 => x"9f",
          4136 => x"5d",
          4137 => x"9c",
          4138 => x"38",
          4139 => x"38",
          4140 => x"81",
          4141 => x"84",
          4142 => x"2a",
          4143 => x"b4",
          4144 => x"86",
          4145 => x"5d",
          4146 => x"fa",
          4147 => x"52",
          4148 => x"84",
          4149 => x"ff",
          4150 => x"79",
          4151 => x"83",
          4152 => x"ff",
          4153 => x"76",
          4154 => x"81",
          4155 => x"84",
          4156 => x"2e",
          4157 => x"87",
          4158 => x"0b",
          4159 => x"2e",
          4160 => x"5b",
          4161 => x"84",
          4162 => x"19",
          4163 => x"3f",
          4164 => x"38",
          4165 => x"0c",
          4166 => x"82",
          4167 => x"11",
          4168 => x"0a",
          4169 => x"57",
          4170 => x"2a",
          4171 => x"2a",
          4172 => x"2a",
          4173 => x"83",
          4174 => x"2a",
          4175 => x"05",
          4176 => x"78",
          4177 => x"33",
          4178 => x"09",
          4179 => x"77",
          4180 => x"51",
          4181 => x"80",
          4182 => x"77",
          4183 => x"ac",
          4184 => x"05",
          4185 => x"57",
          4186 => x"7a",
          4187 => x"8f",
          4188 => x"34",
          4189 => x"2a",
          4190 => x"b4",
          4191 => x"83",
          4192 => x"19",
          4193 => x"f0",
          4194 => x"08",
          4195 => x"38",
          4196 => x"b4",
          4197 => x"a0",
          4198 => x"5c",
          4199 => x"82",
          4200 => x"e4",
          4201 => x"81",
          4202 => x"bb",
          4203 => x"56",
          4204 => x"fc",
          4205 => x"b8",
          4206 => x"8f",
          4207 => x"f0",
          4208 => x"74",
          4209 => x"fc",
          4210 => x"19",
          4211 => x"ef",
          4212 => x"08",
          4213 => x"38",
          4214 => x"b4",
          4215 => x"a0",
          4216 => x"59",
          4217 => x"38",
          4218 => x"09",
          4219 => x"76",
          4220 => x"51",
          4221 => x"39",
          4222 => x"53",
          4223 => x"3f",
          4224 => x"2e",
          4225 => x"bb",
          4226 => x"08",
          4227 => x"08",
          4228 => x"5f",
          4229 => x"19",
          4230 => x"06",
          4231 => x"53",
          4232 => x"e4",
          4233 => x"54",
          4234 => x"1a",
          4235 => x"5a",
          4236 => x"81",
          4237 => x"08",
          4238 => x"a8",
          4239 => x"bb",
          4240 => x"7d",
          4241 => x"55",
          4242 => x"fa",
          4243 => x"52",
          4244 => x"7b",
          4245 => x"1c",
          4246 => x"ec",
          4247 => x"7b",
          4248 => x"7c",
          4249 => x"76",
          4250 => x"79",
          4251 => x"58",
          4252 => x"83",
          4253 => x"11",
          4254 => x"7f",
          4255 => x"5d",
          4256 => x"56",
          4257 => x"5a",
          4258 => x"5b",
          4259 => x"f6",
          4260 => x"5c",
          4261 => x"08",
          4262 => x"76",
          4263 => x"94",
          4264 => x"2e",
          4265 => x"93",
          4266 => x"19",
          4267 => x"75",
          4268 => x"79",
          4269 => x"08",
          4270 => x"84",
          4271 => x"84",
          4272 => x"72",
          4273 => x"51",
          4274 => x"77",
          4275 => x"73",
          4276 => x"3d",
          4277 => x"84",
          4278 => x"52",
          4279 => x"74",
          4280 => x"84",
          4281 => x"08",
          4282 => x"84",
          4283 => x"57",
          4284 => x"19",
          4285 => x"75",
          4286 => x"58",
          4287 => x"a0",
          4288 => x"30",
          4289 => x"07",
          4290 => x"55",
          4291 => x"84",
          4292 => x"08",
          4293 => x"73",
          4294 => x"73",
          4295 => x"80",
          4296 => x"52",
          4297 => x"84",
          4298 => x"84",
          4299 => x"58",
          4300 => x"e3",
          4301 => x"08",
          4302 => x"74",
          4303 => x"1a",
          4304 => x"79",
          4305 => x"bb",
          4306 => x"0b",
          4307 => x"04",
          4308 => x"39",
          4309 => x"53",
          4310 => x"84",
          4311 => x"84",
          4312 => x"8c",
          4313 => x"2e",
          4314 => x"39",
          4315 => x"59",
          4316 => x"80",
          4317 => x"80",
          4318 => x"18",
          4319 => x"33",
          4320 => x"73",
          4321 => x"22",
          4322 => x"ac",
          4323 => x"19",
          4324 => x"72",
          4325 => x"13",
          4326 => x"17",
          4327 => x"75",
          4328 => x"04",
          4329 => x"3d",
          4330 => x"80",
          4331 => x"70",
          4332 => x"a5",
          4333 => x"fe",
          4334 => x"27",
          4335 => x"29",
          4336 => x"98",
          4337 => x"77",
          4338 => x"08",
          4339 => x"a4",
          4340 => x"27",
          4341 => x"84",
          4342 => x"38",
          4343 => x"cd",
          4344 => x"bb",
          4345 => x"3d",
          4346 => x"a0",
          4347 => x"7a",
          4348 => x"0c",
          4349 => x"80",
          4350 => x"5b",
          4351 => x"08",
          4352 => x"2a",
          4353 => x"27",
          4354 => x"79",
          4355 => x"9c",
          4356 => x"84",
          4357 => x"18",
          4358 => x"89",
          4359 => x"52",
          4360 => x"84",
          4361 => x"bb",
          4362 => x"84",
          4363 => x"9c",
          4364 => x"82",
          4365 => x"38",
          4366 => x"a7",
          4367 => x"56",
          4368 => x"9c",
          4369 => x"81",
          4370 => x"bb",
          4371 => x"84",
          4372 => x"58",
          4373 => x"1a",
          4374 => x"75",
          4375 => x"76",
          4376 => x"5e",
          4377 => x"84",
          4378 => x"81",
          4379 => x"f4",
          4380 => x"75",
          4381 => x"75",
          4382 => x"51",
          4383 => x"80",
          4384 => x"7a",
          4385 => x"84",
          4386 => x"b4",
          4387 => x"81",
          4388 => x"84",
          4389 => x"bb",
          4390 => x"08",
          4391 => x"1a",
          4392 => x"33",
          4393 => x"fe",
          4394 => x"a0",
          4395 => x"19",
          4396 => x"39",
          4397 => x"ff",
          4398 => x"06",
          4399 => x"1d",
          4400 => x"80",
          4401 => x"8a",
          4402 => x"08",
          4403 => x"39",
          4404 => x"3d",
          4405 => x"41",
          4406 => x"ff",
          4407 => x"75",
          4408 => x"5f",
          4409 => x"76",
          4410 => x"78",
          4411 => x"06",
          4412 => x"b8",
          4413 => x"bd",
          4414 => x"85",
          4415 => x"1a",
          4416 => x"9c",
          4417 => x"80",
          4418 => x"bf",
          4419 => x"60",
          4420 => x"70",
          4421 => x"80",
          4422 => x"45",
          4423 => x"df",
          4424 => x"bf",
          4425 => x"81",
          4426 => x"f6",
          4427 => x"bb",
          4428 => x"08",
          4429 => x"bb",
          4430 => x"54",
          4431 => x"19",
          4432 => x"84",
          4433 => x"06",
          4434 => x"83",
          4435 => x"08",
          4436 => x"7a",
          4437 => x"82",
          4438 => x"81",
          4439 => x"19",
          4440 => x"52",
          4441 => x"77",
          4442 => x"09",
          4443 => x"2a",
          4444 => x"38",
          4445 => x"70",
          4446 => x"59",
          4447 => x"81",
          4448 => x"81",
          4449 => x"fe",
          4450 => x"0b",
          4451 => x"0c",
          4452 => x"df",
          4453 => x"2e",
          4454 => x"08",
          4455 => x"88",
          4456 => x"b7",
          4457 => x"8d",
          4458 => x"58",
          4459 => x"05",
          4460 => x"2b",
          4461 => x"80",
          4462 => x"87",
          4463 => x"42",
          4464 => x"17",
          4465 => x"33",
          4466 => x"77",
          4467 => x"26",
          4468 => x"43",
          4469 => x"ff",
          4470 => x"83",
          4471 => x"55",
          4472 => x"55",
          4473 => x"80",
          4474 => x"33",
          4475 => x"ff",
          4476 => x"74",
          4477 => x"ac",
          4478 => x"94",
          4479 => x"70",
          4480 => x"f5",
          4481 => x"84",
          4482 => x"ff",
          4483 => x"0c",
          4484 => x"80",
          4485 => x"cc",
          4486 => x"74",
          4487 => x"38",
          4488 => x"81",
          4489 => x"bb",
          4490 => x"56",
          4491 => x"5a",
          4492 => x"70",
          4493 => x"99",
          4494 => x"81",
          4495 => x"34",
          4496 => x"75",
          4497 => x"2e",
          4498 => x"75",
          4499 => x"38",
          4500 => x"81",
          4501 => x"70",
          4502 => x"70",
          4503 => x"5d",
          4504 => x"cd",
          4505 => x"76",
          4506 => x"57",
          4507 => x"70",
          4508 => x"ff",
          4509 => x"2e",
          4510 => x"38",
          4511 => x"0c",
          4512 => x"84",
          4513 => x"08",
          4514 => x"bb",
          4515 => x"54",
          4516 => x"1b",
          4517 => x"84",
          4518 => x"06",
          4519 => x"83",
          4520 => x"08",
          4521 => x"78",
          4522 => x"82",
          4523 => x"81",
          4524 => x"1b",
          4525 => x"52",
          4526 => x"77",
          4527 => x"e4",
          4528 => x"81",
          4529 => x"76",
          4530 => x"2e",
          4531 => x"bf",
          4532 => x"05",
          4533 => x"af",
          4534 => x"52",
          4535 => x"84",
          4536 => x"2e",
          4537 => x"80",
          4538 => x"ff",
          4539 => x"8d",
          4540 => x"81",
          4541 => x"1a",
          4542 => x"07",
          4543 => x"78",
          4544 => x"05",
          4545 => x"e7",
          4546 => x"33",
          4547 => x"42",
          4548 => x"79",
          4549 => x"51",
          4550 => x"08",
          4551 => x"43",
          4552 => x"3f",
          4553 => x"81",
          4554 => x"18",
          4555 => x"78",
          4556 => x"59",
          4557 => x"2e",
          4558 => x"22",
          4559 => x"1d",
          4560 => x"ae",
          4561 => x"93",
          4562 => x"2e",
          4563 => x"94",
          4564 => x"70",
          4565 => x"5a",
          4566 => x"38",
          4567 => x"57",
          4568 => x"1d",
          4569 => x"5d",
          4570 => x"5b",
          4571 => x"75",
          4572 => x"81",
          4573 => x"ef",
          4574 => x"81",
          4575 => x"aa",
          4576 => x"81",
          4577 => x"08",
          4578 => x"57",
          4579 => x"76",
          4580 => x"55",
          4581 => x"c2",
          4582 => x"80",
          4583 => x"56",
          4584 => x"07",
          4585 => x"06",
          4586 => x"56",
          4587 => x"84",
          4588 => x"77",
          4589 => x"74",
          4590 => x"cf",
          4591 => x"06",
          4592 => x"15",
          4593 => x"19",
          4594 => x"e3",
          4595 => x"34",
          4596 => x"a0",
          4597 => x"98",
          4598 => x"88",
          4599 => x"57",
          4600 => x"38",
          4601 => x"26",
          4602 => x"05",
          4603 => x"74",
          4604 => x"38",
          4605 => x"84",
          4606 => x"e3",
          4607 => x"7a",
          4608 => x"bb",
          4609 => x"84",
          4610 => x"02",
          4611 => x"7d",
          4612 => x"33",
          4613 => x"5f",
          4614 => x"8d",
          4615 => x"3f",
          4616 => x"52",
          4617 => x"84",
          4618 => x"82",
          4619 => x"5e",
          4620 => x"b4",
          4621 => x"83",
          4622 => x"81",
          4623 => x"53",
          4624 => x"d4",
          4625 => x"2e",
          4626 => x"b4",
          4627 => x"9c",
          4628 => x"81",
          4629 => x"70",
          4630 => x"80",
          4631 => x"78",
          4632 => x"7d",
          4633 => x"08",
          4634 => x"ff",
          4635 => x"81",
          4636 => x"38",
          4637 => x"98",
          4638 => x"2e",
          4639 => x"40",
          4640 => x"53",
          4641 => x"d3",
          4642 => x"2e",
          4643 => x"b4",
          4644 => x"38",
          4645 => x"80",
          4646 => x"15",
          4647 => x"1f",
          4648 => x"81",
          4649 => x"59",
          4650 => x"9c",
          4651 => x"5e",
          4652 => x"83",
          4653 => x"84",
          4654 => x"30",
          4655 => x"57",
          4656 => x"52",
          4657 => x"84",
          4658 => x"2e",
          4659 => x"54",
          4660 => x"18",
          4661 => x"84",
          4662 => x"bf",
          4663 => x"34",
          4664 => x"55",
          4665 => x"82",
          4666 => x"ac",
          4667 => x"9c",
          4668 => x"71",
          4669 => x"3f",
          4670 => x"84",
          4671 => x"84",
          4672 => x"2a",
          4673 => x"81",
          4674 => x"81",
          4675 => x"76",
          4676 => x"1d",
          4677 => x"56",
          4678 => x"83",
          4679 => x"81",
          4680 => x"53",
          4681 => x"d0",
          4682 => x"2e",
          4683 => x"b4",
          4684 => x"38",
          4685 => x"81",
          4686 => x"1c",
          4687 => x"8c",
          4688 => x"9b",
          4689 => x"76",
          4690 => x"ff",
          4691 => x"22",
          4692 => x"84",
          4693 => x"70",
          4694 => x"56",
          4695 => x"ff",
          4696 => x"27",
          4697 => x"81",
          4698 => x"58",
          4699 => x"7c",
          4700 => x"80",
          4701 => x"bb",
          4702 => x"fc",
          4703 => x"fe",
          4704 => x"b4",
          4705 => x"81",
          4706 => x"81",
          4707 => x"38",
          4708 => x"b4",
          4709 => x"bb",
          4710 => x"08",
          4711 => x"42",
          4712 => x"bc",
          4713 => x"1d",
          4714 => x"33",
          4715 => x"a4",
          4716 => x"57",
          4717 => x"81",
          4718 => x"81",
          4719 => x"9f",
          4720 => x"07",
          4721 => x"1c",
          4722 => x"51",
          4723 => x"76",
          4724 => x"bb",
          4725 => x"08",
          4726 => x"1d",
          4727 => x"5f",
          4728 => x"84",
          4729 => x"1c",
          4730 => x"38",
          4731 => x"e8",
          4732 => x"2e",
          4733 => x"54",
          4734 => x"53",
          4735 => x"ac",
          4736 => x"18",
          4737 => x"52",
          4738 => x"f8",
          4739 => x"71",
          4740 => x"1e",
          4741 => x"b5",
          4742 => x"d9",
          4743 => x"08",
          4744 => x"72",
          4745 => x"14",
          4746 => x"7a",
          4747 => x"70",
          4748 => x"8f",
          4749 => x"1a",
          4750 => x"5b",
          4751 => x"25",
          4752 => x"7c",
          4753 => x"18",
          4754 => x"58",
          4755 => x"18",
          4756 => x"38",
          4757 => x"89",
          4758 => x"25",
          4759 => x"38",
          4760 => x"70",
          4761 => x"74",
          4762 => x"18",
          4763 => x"7c",
          4764 => x"16",
          4765 => x"38",
          4766 => x"1e",
          4767 => x"56",
          4768 => x"08",
          4769 => x"38",
          4770 => x"53",
          4771 => x"1c",
          4772 => x"12",
          4773 => x"07",
          4774 => x"2b",
          4775 => x"97",
          4776 => x"2b",
          4777 => x"5b",
          4778 => x"33",
          4779 => x"5d",
          4780 => x"0d",
          4781 => x"77",
          4782 => x"58",
          4783 => x"2b",
          4784 => x"84",
          4785 => x"55",
          4786 => x"76",
          4787 => x"54",
          4788 => x"82",
          4789 => x"08",
          4790 => x"22",
          4791 => x"fd",
          4792 => x"78",
          4793 => x"58",
          4794 => x"7a",
          4795 => x"8c",
          4796 => x"73",
          4797 => x"80",
          4798 => x"7e",
          4799 => x"bf",
          4800 => x"38",
          4801 => x"5b",
          4802 => x"2a",
          4803 => x"2e",
          4804 => x"ff",
          4805 => x"05",
          4806 => x"19",
          4807 => x"56",
          4808 => x"39",
          4809 => x"7b",
          4810 => x"06",
          4811 => x"ef",
          4812 => x"57",
          4813 => x"53",
          4814 => x"74",
          4815 => x"80",
          4816 => x"88",
          4817 => x"3d",
          4818 => x"a7",
          4819 => x"80",
          4820 => x"33",
          4821 => x"7f",
          4822 => x"83",
          4823 => x"10",
          4824 => x"57",
          4825 => x"32",
          4826 => x"25",
          4827 => x"90",
          4828 => x"38",
          4829 => x"e6",
          4830 => x"81",
          4831 => x"2e",
          4832 => x"38",
          4833 => x"06",
          4834 => x"81",
          4835 => x"76",
          4836 => x"10",
          4837 => x"62",
          4838 => x"54",
          4839 => x"80",
          4840 => x"70",
          4841 => x"55",
          4842 => x"81",
          4843 => x"54",
          4844 => x"80",
          4845 => x"77",
          4846 => x"72",
          4847 => x"94",
          4848 => x"fe",
          4849 => x"73",
          4850 => x"84",
          4851 => x"fe",
          4852 => x"84",
          4853 => x"a0",
          4854 => x"7a",
          4855 => x"ff",
          4856 => x"7b",
          4857 => x"08",
          4858 => x"04",
          4859 => x"70",
          4860 => x"56",
          4861 => x"42",
          4862 => x"72",
          4863 => x"32",
          4864 => x"40",
          4865 => x"0c",
          4866 => x"81",
          4867 => x"83",
          4868 => x"2e",
          4869 => x"05",
          4870 => x"70",
          4871 => x"59",
          4872 => x"38",
          4873 => x"59",
          4874 => x"80",
          4875 => x"70",
          4876 => x"55",
          4877 => x"73",
          4878 => x"2e",
          4879 => x"38",
          4880 => x"54",
          4881 => x"18",
          4882 => x"80",
          4883 => x"5e",
          4884 => x"eb",
          4885 => x"a0",
          4886 => x"13",
          4887 => x"5e",
          4888 => x"59",
          4889 => x"ed",
          4890 => x"74",
          4891 => x"55",
          4892 => x"38",
          4893 => x"7b",
          4894 => x"32",
          4895 => x"70",
          4896 => x"80",
          4897 => x"86",
          4898 => x"79",
          4899 => x"38",
          4900 => x"2b",
          4901 => x"5d",
          4902 => x"56",
          4903 => x"33",
          4904 => x"38",
          4905 => x"8c",
          4906 => x"38",
          4907 => x"82",
          4908 => x"56",
          4909 => x"7c",
          4910 => x"5a",
          4911 => x"80",
          4912 => x"79",
          4913 => x"3f",
          4914 => x"56",
          4915 => x"81",
          4916 => x"2e",
          4917 => x"85",
          4918 => x"84",
          4919 => x"59",
          4920 => x"55",
          4921 => x"80",
          4922 => x"11",
          4923 => x"56",
          4924 => x"2e",
          4925 => x"fd",
          4926 => x"ae",
          4927 => x"77",
          4928 => x"06",
          4929 => x"80",
          4930 => x"53",
          4931 => x"a0",
          4932 => x"34",
          4933 => x"38",
          4934 => x"34",
          4935 => x"84",
          4936 => x"bb",
          4937 => x"2a",
          4938 => x"86",
          4939 => x"56",
          4940 => x"90",
          4941 => x"80",
          4942 => x"71",
          4943 => x"54",
          4944 => x"74",
          4945 => x"56",
          4946 => x"ae",
          4947 => x"76",
          4948 => x"83",
          4949 => x"39",
          4950 => x"8c",
          4951 => x"81",
          4952 => x"5a",
          4953 => x"34",
          4954 => x"f6",
          4955 => x"1d",
          4956 => x"93",
          4957 => x"9d",
          4958 => x"38",
          4959 => x"f7",
          4960 => x"57",
          4961 => x"07",
          4962 => x"85",
          4963 => x"ff",
          4964 => x"5a",
          4965 => x"80",
          4966 => x"56",
          4967 => x"38",
          4968 => x"e6",
          4969 => x"81",
          4970 => x"2e",
          4971 => x"38",
          4972 => x"06",
          4973 => x"81",
          4974 => x"ff",
          4975 => x"38",
          4976 => x"5f",
          4977 => x"26",
          4978 => x"ff",
          4979 => x"06",
          4980 => x"05",
          4981 => x"75",
          4982 => x"fa",
          4983 => x"81",
          4984 => x"ff",
          4985 => x"7d",
          4986 => x"79",
          4987 => x"cd",
          4988 => x"98",
          4989 => x"88",
          4990 => x"7b",
          4991 => x"54",
          4992 => x"a0",
          4993 => x"1b",
          4994 => x"a0",
          4995 => x"2e",
          4996 => x"a3",
          4997 => x"7b",
          4998 => x"84",
          4999 => x"0d",
          5000 => x"05",
          5001 => x"ff",
          5002 => x"80",
          5003 => x"05",
          5004 => x"75",
          5005 => x"38",
          5006 => x"e2",
          5007 => x"b2",
          5008 => x"05",
          5009 => x"80",
          5010 => x"7f",
          5011 => x"7b",
          5012 => x"51",
          5013 => x"08",
          5014 => x"58",
          5015 => x"77",
          5016 => x"1d",
          5017 => x"17",
          5018 => x"bb",
          5019 => x"06",
          5020 => x"38",
          5021 => x"2a",
          5022 => x"b1",
          5023 => x"ff",
          5024 => x"55",
          5025 => x"53",
          5026 => x"95",
          5027 => x"85",
          5028 => x"18",
          5029 => x"b7",
          5030 => x"88",
          5031 => x"82",
          5032 => x"81",
          5033 => x"33",
          5034 => x"75",
          5035 => x"75",
          5036 => x"17",
          5037 => x"2b",
          5038 => x"09",
          5039 => x"17",
          5040 => x"2b",
          5041 => x"dc",
          5042 => x"71",
          5043 => x"14",
          5044 => x"33",
          5045 => x"5f",
          5046 => x"17",
          5047 => x"33",
          5048 => x"40",
          5049 => x"d9",
          5050 => x"29",
          5051 => x"77",
          5052 => x"2e",
          5053 => x"42",
          5054 => x"33",
          5055 => x"07",
          5056 => x"75",
          5057 => x"82",
          5058 => x"cb",
          5059 => x"5c",
          5060 => x"11",
          5061 => x"71",
          5062 => x"72",
          5063 => x"53",
          5064 => x"c7",
          5065 => x"88",
          5066 => x"80",
          5067 => x"84",
          5068 => x"c1",
          5069 => x"fd",
          5070 => x"56",
          5071 => x"a9",
          5072 => x"ff",
          5073 => x"75",
          5074 => x"5d",
          5075 => x"81",
          5076 => x"7b",
          5077 => x"1a",
          5078 => x"59",
          5079 => x"17",
          5080 => x"80",
          5081 => x"78",
          5082 => x"78",
          5083 => x"06",
          5084 => x"2a",
          5085 => x"26",
          5086 => x"ff",
          5087 => x"84",
          5088 => x"38",
          5089 => x"81",
          5090 => x"7c",
          5091 => x"8c",
          5092 => x"80",
          5093 => x"3d",
          5094 => x"0c",
          5095 => x"11",
          5096 => x"74",
          5097 => x"81",
          5098 => x"7a",
          5099 => x"83",
          5100 => x"7f",
          5101 => x"33",
          5102 => x"9f",
          5103 => x"89",
          5104 => x"57",
          5105 => x"26",
          5106 => x"06",
          5107 => x"59",
          5108 => x"85",
          5109 => x"32",
          5110 => x"7a",
          5111 => x"87",
          5112 => x"5c",
          5113 => x"56",
          5114 => x"cf",
          5115 => x"8a",
          5116 => x"fe",
          5117 => x"75",
          5118 => x"38",
          5119 => x"30",
          5120 => x"5c",
          5121 => x"2e",
          5122 => x"5a",
          5123 => x"59",
          5124 => x"81",
          5125 => x"90",
          5126 => x"19",
          5127 => x"fe",
          5128 => x"40",
          5129 => x"5c",
          5130 => x"78",
          5131 => x"f9",
          5132 => x"72",
          5133 => x"05",
          5134 => x"52",
          5135 => x"56",
          5136 => x"0b",
          5137 => x"0c",
          5138 => x"a5",
          5139 => x"52",
          5140 => x"3f",
          5141 => x"38",
          5142 => x"0c",
          5143 => x"33",
          5144 => x"5e",
          5145 => x"09",
          5146 => x"18",
          5147 => x"82",
          5148 => x"30",
          5149 => x"42",
          5150 => x"b6",
          5151 => x"56",
          5152 => x"5d",
          5153 => x"83",
          5154 => x"bd",
          5155 => x"81",
          5156 => x"27",
          5157 => x"0b",
          5158 => x"5d",
          5159 => x"7e",
          5160 => x"31",
          5161 => x"80",
          5162 => x"e1",
          5163 => x"e6",
          5164 => x"05",
          5165 => x"33",
          5166 => x"42",
          5167 => x"75",
          5168 => x"f3",
          5169 => x"77",
          5170 => x"04",
          5171 => x"38",
          5172 => x"b8",
          5173 => x"0b",
          5174 => x"04",
          5175 => x"b4",
          5176 => x"5a",
          5177 => x"71",
          5178 => x"5f",
          5179 => x"80",
          5180 => x"18",
          5181 => x"70",
          5182 => x"05",
          5183 => x"5b",
          5184 => x"91",
          5185 => x"3d",
          5186 => x"39",
          5187 => x"17",
          5188 => x"2b",
          5189 => x"81",
          5190 => x"80",
          5191 => x"38",
          5192 => x"09",
          5193 => x"77",
          5194 => x"51",
          5195 => x"08",
          5196 => x"5a",
          5197 => x"38",
          5198 => x"33",
          5199 => x"07",
          5200 => x"09",
          5201 => x"83",
          5202 => x"2b",
          5203 => x"70",
          5204 => x"07",
          5205 => x"77",
          5206 => x"81",
          5207 => x"83",
          5208 => x"2b",
          5209 => x"70",
          5210 => x"07",
          5211 => x"60",
          5212 => x"81",
          5213 => x"83",
          5214 => x"2b",
          5215 => x"70",
          5216 => x"07",
          5217 => x"83",
          5218 => x"2b",
          5219 => x"70",
          5220 => x"07",
          5221 => x"46",
          5222 => x"7c",
          5223 => x"05",
          5224 => x"86",
          5225 => x"18",
          5226 => x"cf",
          5227 => x"7b",
          5228 => x"75",
          5229 => x"70",
          5230 => x"af",
          5231 => x"2e",
          5232 => x"bb",
          5233 => x"08",
          5234 => x"18",
          5235 => x"41",
          5236 => x"bb",
          5237 => x"56",
          5238 => x"0b",
          5239 => x"5a",
          5240 => x"33",
          5241 => x"07",
          5242 => x"38",
          5243 => x"38",
          5244 => x"12",
          5245 => x"07",
          5246 => x"2b",
          5247 => x"5a",
          5248 => x"59",
          5249 => x"80",
          5250 => x"e3",
          5251 => x"93",
          5252 => x"f2",
          5253 => x"fc",
          5254 => x"a0",
          5255 => x"17",
          5256 => x"85",
          5257 => x"05",
          5258 => x"57",
          5259 => x"2e",
          5260 => x"5a",
          5261 => x"ba",
          5262 => x"74",
          5263 => x"e0",
          5264 => x"38",
          5265 => x"70",
          5266 => x"38",
          5267 => x"2e",
          5268 => x"73",
          5269 => x"92",
          5270 => x"84",
          5271 => x"84",
          5272 => x"92",
          5273 => x"84",
          5274 => x"d0",
          5275 => x"57",
          5276 => x"77",
          5277 => x"77",
          5278 => x"08",
          5279 => x"08",
          5280 => x"5b",
          5281 => x"ff",
          5282 => x"26",
          5283 => x"06",
          5284 => x"99",
          5285 => x"ff",
          5286 => x"2a",
          5287 => x"06",
          5288 => x"79",
          5289 => x"2a",
          5290 => x"2e",
          5291 => x"5b",
          5292 => x"54",
          5293 => x"38",
          5294 => x"39",
          5295 => x"80",
          5296 => x"79",
          5297 => x"70",
          5298 => x"3d",
          5299 => x"84",
          5300 => x"08",
          5301 => x"76",
          5302 => x"3d",
          5303 => x"3d",
          5304 => x"bb",
          5305 => x"80",
          5306 => x"5d",
          5307 => x"80",
          5308 => x"84",
          5309 => x"ff",
          5310 => x"58",
          5311 => x"9b",
          5312 => x"2b",
          5313 => x"5e",
          5314 => x"80",
          5315 => x"17",
          5316 => x"cc",
          5317 => x"0b",
          5318 => x"80",
          5319 => x"17",
          5320 => x"85",
          5321 => x"19",
          5322 => x"0b",
          5323 => x"34",
          5324 => x"7a",
          5325 => x"11",
          5326 => x"57",
          5327 => x"08",
          5328 => x"80",
          5329 => x"e7",
          5330 => x"7a",
          5331 => x"9c",
          5332 => x"76",
          5333 => x"33",
          5334 => x"7b",
          5335 => x"06",
          5336 => x"81",
          5337 => x"83",
          5338 => x"86",
          5339 => x"b4",
          5340 => x"1c",
          5341 => x"33",
          5342 => x"5b",
          5343 => x"fb",
          5344 => x"83",
          5345 => x"2b",
          5346 => x"70",
          5347 => x"07",
          5348 => x"0c",
          5349 => x"22",
          5350 => x"80",
          5351 => x"1b",
          5352 => x"1a",
          5353 => x"76",
          5354 => x"55",
          5355 => x"06",
          5356 => x"8c",
          5357 => x"bf",
          5358 => x"22",
          5359 => x"59",
          5360 => x"07",
          5361 => x"83",
          5362 => x"5b",
          5363 => x"52",
          5364 => x"bb",
          5365 => x"81",
          5366 => x"84",
          5367 => x"31",
          5368 => x"33",
          5369 => x"82",
          5370 => x"fc",
          5371 => x"fb",
          5372 => x"fb",
          5373 => x"fb",
          5374 => x"57",
          5375 => x"17",
          5376 => x"07",
          5377 => x"83",
          5378 => x"2b",
          5379 => x"70",
          5380 => x"07",
          5381 => x"0c",
          5382 => x"86",
          5383 => x"1b",
          5384 => x"0b",
          5385 => x"0c",
          5386 => x"55",
          5387 => x"3f",
          5388 => x"5a",
          5389 => x"39",
          5390 => x"3f",
          5391 => x"84",
          5392 => x"bb",
          5393 => x"84",
          5394 => x"38",
          5395 => x"b1",
          5396 => x"8f",
          5397 => x"18",
          5398 => x"90",
          5399 => x"16",
          5400 => x"34",
          5401 => x"38",
          5402 => x"5d",
          5403 => x"83",
          5404 => x"81",
          5405 => x"53",
          5406 => x"ff",
          5407 => x"80",
          5408 => x"76",
          5409 => x"1c",
          5410 => x"fb",
          5411 => x"39",
          5412 => x"95",
          5413 => x"33",
          5414 => x"90",
          5415 => x"80",
          5416 => x"17",
          5417 => x"cc",
          5418 => x"0b",
          5419 => x"80",
          5420 => x"17",
          5421 => x"09",
          5422 => x"39",
          5423 => x"38",
          5424 => x"2e",
          5425 => x"12",
          5426 => x"7e",
          5427 => x"78",
          5428 => x"5b",
          5429 => x"89",
          5430 => x"81",
          5431 => x"33",
          5432 => x"84",
          5433 => x"57",
          5434 => x"54",
          5435 => x"53",
          5436 => x"c4",
          5437 => x"09",
          5438 => x"84",
          5439 => x"a8",
          5440 => x"5d",
          5441 => x"dc",
          5442 => x"2e",
          5443 => x"54",
          5444 => x"53",
          5445 => x"a1",
          5446 => x"84",
          5447 => x"f6",
          5448 => x"f2",
          5449 => x"40",
          5450 => x"78",
          5451 => x"75",
          5452 => x"74",
          5453 => x"84",
          5454 => x"83",
          5455 => x"55",
          5456 => x"55",
          5457 => x"81",
          5458 => x"81",
          5459 => x"08",
          5460 => x"81",
          5461 => x"38",
          5462 => x"99",
          5463 => x"77",
          5464 => x"38",
          5465 => x"55",
          5466 => x"ff",
          5467 => x"0c",
          5468 => x"9c",
          5469 => x"7b",
          5470 => x"70",
          5471 => x"56",
          5472 => x"15",
          5473 => x"2e",
          5474 => x"75",
          5475 => x"7a",
          5476 => x"33",
          5477 => x"84",
          5478 => x"70",
          5479 => x"82",
          5480 => x"77",
          5481 => x"1e",
          5482 => x"1c",
          5483 => x"80",
          5484 => x"3d",
          5485 => x"90",
          5486 => x"39",
          5487 => x"80",
          5488 => x"2b",
          5489 => x"25",
          5490 => x"52",
          5491 => x"3f",
          5492 => x"90",
          5493 => x"90",
          5494 => x"53",
          5495 => x"9d",
          5496 => x"c1",
          5497 => x"08",
          5498 => x"71",
          5499 => x"38",
          5500 => x"05",
          5501 => x"d6",
          5502 => x"78",
          5503 => x"56",
          5504 => x"70",
          5505 => x"05",
          5506 => x"38",
          5507 => x"78",
          5508 => x"84",
          5509 => x"33",
          5510 => x"84",
          5511 => x"38",
          5512 => x"39",
          5513 => x"7b",
          5514 => x"71",
          5515 => x"75",
          5516 => x"81",
          5517 => x"80",
          5518 => x"05",
          5519 => x"34",
          5520 => x"ba",
          5521 => x"0b",
          5522 => x"04",
          5523 => x"84",
          5524 => x"f1",
          5525 => x"41",
          5526 => x"78",
          5527 => x"75",
          5528 => x"74",
          5529 => x"84",
          5530 => x"84",
          5531 => x"55",
          5532 => x"55",
          5533 => x"70",
          5534 => x"56",
          5535 => x"19",
          5536 => x"27",
          5537 => x"2e",
          5538 => x"5d",
          5539 => x"22",
          5540 => x"58",
          5541 => x"88",
          5542 => x"8c",
          5543 => x"74",
          5544 => x"1a",
          5545 => x"88",
          5546 => x"70",
          5547 => x"82",
          5548 => x"9c",
          5549 => x"7c",
          5550 => x"70",
          5551 => x"56",
          5552 => x"15",
          5553 => x"2e",
          5554 => x"75",
          5555 => x"79",
          5556 => x"33",
          5557 => x"84",
          5558 => x"7c",
          5559 => x"84",
          5560 => x"60",
          5561 => x"05",
          5562 => x"34",
          5563 => x"19",
          5564 => x"1a",
          5565 => x"31",
          5566 => x"94",
          5567 => x"0c",
          5568 => x"5b",
          5569 => x"74",
          5570 => x"90",
          5571 => x"5b",
          5572 => x"84",
          5573 => x"74",
          5574 => x"04",
          5575 => x"94",
          5576 => x"27",
          5577 => x"19",
          5578 => x"d5",
          5579 => x"38",
          5580 => x"0c",
          5581 => x"31",
          5582 => x"7a",
          5583 => x"59",
          5584 => x"76",
          5585 => x"81",
          5586 => x"ef",
          5587 => x"5a",
          5588 => x"98",
          5589 => x"ef",
          5590 => x"bb",
          5591 => x"33",
          5592 => x"51",
          5593 => x"08",
          5594 => x"38",
          5595 => x"53",
          5596 => x"ff",
          5597 => x"ac",
          5598 => x"56",
          5599 => x"e2",
          5600 => x"d3",
          5601 => x"55",
          5602 => x"56",
          5603 => x"1a",
          5604 => x"91",
          5605 => x"34",
          5606 => x"3d",
          5607 => x"89",
          5608 => x"08",
          5609 => x"33",
          5610 => x"16",
          5611 => x"79",
          5612 => x"5c",
          5613 => x"18",
          5614 => x"57",
          5615 => x"98",
          5616 => x"38",
          5617 => x"16",
          5618 => x"83",
          5619 => x"7a",
          5620 => x"81",
          5621 => x"16",
          5622 => x"bb",
          5623 => x"57",
          5624 => x"56",
          5625 => x"8b",
          5626 => x"8b",
          5627 => x"70",
          5628 => x"7a",
          5629 => x"79",
          5630 => x"96",
          5631 => x"81",
          5632 => x"7b",
          5633 => x"18",
          5634 => x"18",
          5635 => x"18",
          5636 => x"18",
          5637 => x"cc",
          5638 => x"18",
          5639 => x"5b",
          5640 => x"ff",
          5641 => x"90",
          5642 => x"79",
          5643 => x"bb",
          5644 => x"54",
          5645 => x"53",
          5646 => x"b4",
          5647 => x"7a",
          5648 => x"84",
          5649 => x"16",
          5650 => x"84",
          5651 => x"27",
          5652 => x"74",
          5653 => x"38",
          5654 => x"08",
          5655 => x"51",
          5656 => x"df",
          5657 => x"18",
          5658 => x"18",
          5659 => x"34",
          5660 => x"34",
          5661 => x"34",
          5662 => x"34",
          5663 => x"34",
          5664 => x"0b",
          5665 => x"34",
          5666 => x"81",
          5667 => x"96",
          5668 => x"19",
          5669 => x"90",
          5670 => x"33",
          5671 => x"84",
          5672 => x"38",
          5673 => x"39",
          5674 => x"18",
          5675 => x"ff",
          5676 => x"84",
          5677 => x"80",
          5678 => x"7b",
          5679 => x"08",
          5680 => x"38",
          5681 => x"70",
          5682 => x"84",
          5683 => x"38",
          5684 => x"74",
          5685 => x"72",
          5686 => x"86",
          5687 => x"71",
          5688 => x"58",
          5689 => x"0c",
          5690 => x"0d",
          5691 => x"fb",
          5692 => x"53",
          5693 => x"56",
          5694 => x"70",
          5695 => x"38",
          5696 => x"9f",
          5697 => x"38",
          5698 => x"38",
          5699 => x"24",
          5700 => x"80",
          5701 => x"0d",
          5702 => x"8c",
          5703 => x"70",
          5704 => x"89",
          5705 => x"ff",
          5706 => x"2e",
          5707 => x"f4",
          5708 => x"76",
          5709 => x"81",
          5710 => x"54",
          5711 => x"12",
          5712 => x"9f",
          5713 => x"e0",
          5714 => x"71",
          5715 => x"73",
          5716 => x"ff",
          5717 => x"70",
          5718 => x"52",
          5719 => x"18",
          5720 => x"ff",
          5721 => x"77",
          5722 => x"51",
          5723 => x"53",
          5724 => x"51",
          5725 => x"55",
          5726 => x"38",
          5727 => x"0d",
          5728 => x"d0",
          5729 => x"84",
          5730 => x"c6",
          5731 => x"98",
          5732 => x"e2",
          5733 => x"2a",
          5734 => x"b2",
          5735 => x"12",
          5736 => x"5e",
          5737 => x"a4",
          5738 => x"bb",
          5739 => x"bb",
          5740 => x"ff",
          5741 => x"0c",
          5742 => x"94",
          5743 => x"2b",
          5744 => x"54",
          5745 => x"58",
          5746 => x"0d",
          5747 => x"3d",
          5748 => x"80",
          5749 => x"fd",
          5750 => x"d1",
          5751 => x"84",
          5752 => x"80",
          5753 => x"08",
          5754 => x"3d",
          5755 => x"cc",
          5756 => x"5b",
          5757 => x"3f",
          5758 => x"84",
          5759 => x"3d",
          5760 => x"2e",
          5761 => x"17",
          5762 => x"81",
          5763 => x"16",
          5764 => x"bb",
          5765 => x"57",
          5766 => x"82",
          5767 => x"11",
          5768 => x"07",
          5769 => x"56",
          5770 => x"80",
          5771 => x"ff",
          5772 => x"59",
          5773 => x"80",
          5774 => x"84",
          5775 => x"08",
          5776 => x"11",
          5777 => x"07",
          5778 => x"56",
          5779 => x"7a",
          5780 => x"52",
          5781 => x"bb",
          5782 => x"80",
          5783 => x"83",
          5784 => x"e4",
          5785 => x"ff",
          5786 => x"33",
          5787 => x"82",
          5788 => x"33",
          5789 => x"17",
          5790 => x"76",
          5791 => x"05",
          5792 => x"11",
          5793 => x"58",
          5794 => x"ff",
          5795 => x"58",
          5796 => x"5a",
          5797 => x"82",
          5798 => x"33",
          5799 => x"70",
          5800 => x"5a",
          5801 => x"70",
          5802 => x"f5",
          5803 => x"ab",
          5804 => x"38",
          5805 => x"81",
          5806 => x"77",
          5807 => x"05",
          5808 => x"06",
          5809 => x"34",
          5810 => x"3d",
          5811 => x"33",
          5812 => x"79",
          5813 => x"95",
          5814 => x"2b",
          5815 => x"dd",
          5816 => x"51",
          5817 => x"08",
          5818 => x"fd",
          5819 => x"b4",
          5820 => x"81",
          5821 => x"3f",
          5822 => x"be",
          5823 => x"34",
          5824 => x"84",
          5825 => x"17",
          5826 => x"33",
          5827 => x"fb",
          5828 => x"a0",
          5829 => x"16",
          5830 => x"59",
          5831 => x"3d",
          5832 => x"80",
          5833 => x"10",
          5834 => x"33",
          5835 => x"2e",
          5836 => x"f1",
          5837 => x"19",
          5838 => x"05",
          5839 => x"38",
          5840 => x"59",
          5841 => x"5e",
          5842 => x"f5",
          5843 => x"84",
          5844 => x"04",
          5845 => x"89",
          5846 => x"08",
          5847 => x"33",
          5848 => x"16",
          5849 => x"7a",
          5850 => x"5c",
          5851 => x"17",
          5852 => x"17",
          5853 => x"38",
          5854 => x"7a",
          5855 => x"22",
          5856 => x"7a",
          5857 => x"19",
          5858 => x"84",
          5859 => x"57",
          5860 => x"84",
          5861 => x"30",
          5862 => x"71",
          5863 => x"75",
          5864 => x"27",
          5865 => x"18",
          5866 => x"33",
          5867 => x"59",
          5868 => x"52",
          5869 => x"bb",
          5870 => x"80",
          5871 => x"d1",
          5872 => x"7b",
          5873 => x"f8",
          5874 => x"39",
          5875 => x"08",
          5876 => x"06",
          5877 => x"fe",
          5878 => x"57",
          5879 => x"8a",
          5880 => x"08",
          5881 => x"55",
          5882 => x"17",
          5883 => x"76",
          5884 => x"90",
          5885 => x"90",
          5886 => x"7a",
          5887 => x"08",
          5888 => x"90",
          5889 => x"5a",
          5890 => x"81",
          5891 => x"11",
          5892 => x"84",
          5893 => x"33",
          5894 => x"34",
          5895 => x"81",
          5896 => x"3f",
          5897 => x"d3",
          5898 => x"55",
          5899 => x"0d",
          5900 => x"81",
          5901 => x"77",
          5902 => x"78",
          5903 => x"38",
          5904 => x"80",
          5905 => x"56",
          5906 => x"98",
          5907 => x"38",
          5908 => x"80",
          5909 => x"0d",
          5910 => x"a8",
          5911 => x"bb",
          5912 => x"93",
          5913 => x"55",
          5914 => x"56",
          5915 => x"51",
          5916 => x"08",
          5917 => x"98",
          5918 => x"fe",
          5919 => x"18",
          5920 => x"39",
          5921 => x"84",
          5922 => x"f6",
          5923 => x"80",
          5924 => x"fc",
          5925 => x"c6",
          5926 => x"84",
          5927 => x"80",
          5928 => x"84",
          5929 => x"0c",
          5930 => x"3f",
          5931 => x"84",
          5932 => x"70",
          5933 => x"af",
          5934 => x"81",
          5935 => x"c5",
          5936 => x"9a",
          5937 => x"70",
          5938 => x"83",
          5939 => x"7a",
          5940 => x"74",
          5941 => x"84",
          5942 => x"8d",
          5943 => x"80",
          5944 => x"80",
          5945 => x"33",
          5946 => x"90",
          5947 => x"5a",
          5948 => x"78",
          5949 => x"38",
          5950 => x"38",
          5951 => x"38",
          5952 => x"52",
          5953 => x"71",
          5954 => x"73",
          5955 => x"04",
          5956 => x"3f",
          5957 => x"71",
          5958 => x"d7",
          5959 => x"55",
          5960 => x"74",
          5961 => x"73",
          5962 => x"86",
          5963 => x"72",
          5964 => x"72",
          5965 => x"76",
          5966 => x"74",
          5967 => x"84",
          5968 => x"2e",
          5969 => x"38",
          5970 => x"3f",
          5971 => x"3f",
          5972 => x"30",
          5973 => x"84",
          5974 => x"bb",
          5975 => x"77",
          5976 => x"3f",
          5977 => x"3f",
          5978 => x"30",
          5979 => x"84",
          5980 => x"75",
          5981 => x"84",
          5982 => x"8a",
          5983 => x"fe",
          5984 => x"81",
          5985 => x"75",
          5986 => x"3d",
          5987 => x"70",
          5988 => x"3f",
          5989 => x"84",
          5990 => x"bb",
          5991 => x"52",
          5992 => x"bb",
          5993 => x"e5",
          5994 => x"98",
          5995 => x"38",
          5996 => x"75",
          5997 => x"bb",
          5998 => x"0b",
          5999 => x"04",
          6000 => x"80",
          6001 => x"3d",
          6002 => x"08",
          6003 => x"7f",
          6004 => x"fe",
          6005 => x"57",
          6006 => x"0c",
          6007 => x"0d",
          6008 => x"5a",
          6009 => x"77",
          6010 => x"5a",
          6011 => x"81",
          6012 => x"08",
          6013 => x"33",
          6014 => x"81",
          6015 => x"17",
          6016 => x"bb",
          6017 => x"5a",
          6018 => x"7e",
          6019 => x"33",
          6020 => x"77",
          6021 => x"12",
          6022 => x"07",
          6023 => x"2b",
          6024 => x"80",
          6025 => x"63",
          6026 => x"62",
          6027 => x"52",
          6028 => x"f2",
          6029 => x"0c",
          6030 => x"84",
          6031 => x"95",
          6032 => x"08",
          6033 => x"33",
          6034 => x"5e",
          6035 => x"84",
          6036 => x"17",
          6037 => x"84",
          6038 => x"27",
          6039 => x"74",
          6040 => x"38",
          6041 => x"08",
          6042 => x"51",
          6043 => x"97",
          6044 => x"56",
          6045 => x"3f",
          6046 => x"e8",
          6047 => x"80",
          6048 => x"70",
          6049 => x"7c",
          6050 => x"5c",
          6051 => x"7a",
          6052 => x"17",
          6053 => x"34",
          6054 => x"81",
          6055 => x"07",
          6056 => x"1d",
          6057 => x"5f",
          6058 => x"38",
          6059 => x"39",
          6060 => x"7a",
          6061 => x"07",
          6062 => x"39",
          6063 => x"3d",
          6064 => x"2e",
          6065 => x"2e",
          6066 => x"2e",
          6067 => x"22",
          6068 => x"38",
          6069 => x"38",
          6070 => x"38",
          6071 => x"06",
          6072 => x"80",
          6073 => x"8c",
          6074 => x"81",
          6075 => x"58",
          6076 => x"17",
          6077 => x"57",
          6078 => x"08",
          6079 => x"55",
          6080 => x"74",
          6081 => x"38",
          6082 => x"18",
          6083 => x"fe",
          6084 => x"80",
          6085 => x"91",
          6086 => x"84",
          6087 => x"79",
          6088 => x"77",
          6089 => x"84",
          6090 => x"2e",
          6091 => x"81",
          6092 => x"08",
          6093 => x"74",
          6094 => x"84",
          6095 => x"17",
          6096 => x"56",
          6097 => x"81",
          6098 => x"81",
          6099 => x"55",
          6100 => x"39",
          6101 => x"3f",
          6102 => x"74",
          6103 => x"57",
          6104 => x"33",
          6105 => x"19",
          6106 => x"52",
          6107 => x"bb",
          6108 => x"84",
          6109 => x"38",
          6110 => x"bb",
          6111 => x"a1",
          6112 => x"08",
          6113 => x"84",
          6114 => x"84",
          6115 => x"81",
          6116 => x"ff",
          6117 => x"91",
          6118 => x"bb",
          6119 => x"77",
          6120 => x"84",
          6121 => x"2e",
          6122 => x"81",
          6123 => x"08",
          6124 => x"74",
          6125 => x"84",
          6126 => x"17",
          6127 => x"56",
          6128 => x"16",
          6129 => x"07",
          6130 => x"78",
          6131 => x"75",
          6132 => x"39",
          6133 => x"90",
          6134 => x"82",
          6135 => x"ff",
          6136 => x"56",
          6137 => x"33",
          6138 => x"84",
          6139 => x"ea",
          6140 => x"55",
          6141 => x"57",
          6142 => x"39",
          6143 => x"ff",
          6144 => x"b8",
          6145 => x"84",
          6146 => x"75",
          6147 => x"04",
          6148 => x"3d",
          6149 => x"84",
          6150 => x"08",
          6151 => x"70",
          6152 => x"56",
          6153 => x"80",
          6154 => x"05",
          6155 => x"56",
          6156 => x"08",
          6157 => x"88",
          6158 => x"57",
          6159 => x"76",
          6160 => x"2e",
          6161 => x"08",
          6162 => x"7a",
          6163 => x"3d",
          6164 => x"84",
          6165 => x"08",
          6166 => x"52",
          6167 => x"bb",
          6168 => x"a0",
          6169 => x"a7",
          6170 => x"17",
          6171 => x"07",
          6172 => x"39",
          6173 => x"38",
          6174 => x"78",
          6175 => x"57",
          6176 => x"52",
          6177 => x"bb",
          6178 => x"80",
          6179 => x"07",
          6180 => x"9a",
          6181 => x"79",
          6182 => x"38",
          6183 => x"38",
          6184 => x"51",
          6185 => x"08",
          6186 => x"04",
          6187 => x"80",
          6188 => x"b9",
          6189 => x"74",
          6190 => x"38",
          6191 => x"81",
          6192 => x"84",
          6193 => x"ff",
          6194 => x"77",
          6195 => x"58",
          6196 => x"34",
          6197 => x"38",
          6198 => x"3f",
          6199 => x"84",
          6200 => x"84",
          6201 => x"82",
          6202 => x"17",
          6203 => x"51",
          6204 => x"bb",
          6205 => x"ff",
          6206 => x"18",
          6207 => x"31",
          6208 => x"a0",
          6209 => x"17",
          6210 => x"06",
          6211 => x"08",
          6212 => x"81",
          6213 => x"79",
          6214 => x"78",
          6215 => x"51",
          6216 => x"08",
          6217 => x"80",
          6218 => x"2e",
          6219 => x"ff",
          6220 => x"52",
          6221 => x"bb",
          6222 => x"fe",
          6223 => x"75",
          6224 => x"94",
          6225 => x"5c",
          6226 => x"7a",
          6227 => x"a2",
          6228 => x"bb",
          6229 => x"56",
          6230 => x"53",
          6231 => x"3d",
          6232 => x"84",
          6233 => x"2e",
          6234 => x"9f",
          6235 => x"93",
          6236 => x"3f",
          6237 => x"84",
          6238 => x"84",
          6239 => x"84",
          6240 => x"38",
          6241 => x"2a",
          6242 => x"ff",
          6243 => x"3d",
          6244 => x"84",
          6245 => x"bb",
          6246 => x"bb",
          6247 => x"84",
          6248 => x"38",
          6249 => x"84",
          6250 => x"7a",
          6251 => x"08",
          6252 => x"79",
          6253 => x"71",
          6254 => x"7a",
          6255 => x"80",
          6256 => x"05",
          6257 => x"38",
          6258 => x"75",
          6259 => x"1b",
          6260 => x"fe",
          6261 => x"81",
          6262 => x"82",
          6263 => x"17",
          6264 => x"18",
          6265 => x"81",
          6266 => x"84",
          6267 => x"17",
          6268 => x"a0",
          6269 => x"17",
          6270 => x"06",
          6271 => x"08",
          6272 => x"81",
          6273 => x"fe",
          6274 => x"58",
          6275 => x"7b",
          6276 => x"74",
          6277 => x"84",
          6278 => x"08",
          6279 => x"84",
          6280 => x"bb",
          6281 => x"80",
          6282 => x"e9",
          6283 => x"38",
          6284 => x"08",
          6285 => x"38",
          6286 => x"33",
          6287 => x"79",
          6288 => x"75",
          6289 => x"04",
          6290 => x"ff",
          6291 => x"09",
          6292 => x"b8",
          6293 => x"05",
          6294 => x"38",
          6295 => x"7d",
          6296 => x"7d",
          6297 => x"80",
          6298 => x"1a",
          6299 => x"34",
          6300 => x"56",
          6301 => x"2a",
          6302 => x"33",
          6303 => x"7d",
          6304 => x"1b",
          6305 => x"56",
          6306 => x"ff",
          6307 => x"ae",
          6308 => x"71",
          6309 => x"78",
          6310 => x"5b",
          6311 => x"55",
          6312 => x"5b",
          6313 => x"ff",
          6314 => x"56",
          6315 => x"69",
          6316 => x"34",
          6317 => x"a1",
          6318 => x"99",
          6319 => x"9a",
          6320 => x"9b",
          6321 => x"2e",
          6322 => x"8b",
          6323 => x"18",
          6324 => x"84",
          6325 => x"84",
          6326 => x"2a",
          6327 => x"88",
          6328 => x"fe",
          6329 => x"80",
          6330 => x"74",
          6331 => x"0b",
          6332 => x"56",
          6333 => x"77",
          6334 => x"7b",
          6335 => x"8b",
          6336 => x"18",
          6337 => x"84",
          6338 => x"d1",
          6339 => x"70",
          6340 => x"38",
          6341 => x"9f",
          6342 => x"b8",
          6343 => x"81",
          6344 => x"fc",
          6345 => x"ed",
          6346 => x"bb",
          6347 => x"84",
          6348 => x"7f",
          6349 => x"a5",
          6350 => x"3f",
          6351 => x"84",
          6352 => x"33",
          6353 => x"ce",
          6354 => x"08",
          6355 => x"57",
          6356 => x"ff",
          6357 => x"58",
          6358 => x"70",
          6359 => x"05",
          6360 => x"38",
          6361 => x"9f",
          6362 => x"84",
          6363 => x"a8",
          6364 => x"0b",
          6365 => x"04",
          6366 => x"06",
          6367 => x"38",
          6368 => x"05",
          6369 => x"38",
          6370 => x"08",
          6371 => x"70",
          6372 => x"05",
          6373 => x"56",
          6374 => x"70",
          6375 => x"17",
          6376 => x"17",
          6377 => x"30",
          6378 => x"2e",
          6379 => x"be",
          6380 => x"72",
          6381 => x"55",
          6382 => x"84",
          6383 => x"c2",
          6384 => x"96",
          6385 => x"79",
          6386 => x"fc",
          6387 => x"9d",
          6388 => x"bb",
          6389 => x"39",
          6390 => x"06",
          6391 => x"e1",
          6392 => x"bb",
          6393 => x"93",
          6394 => x"cd",
          6395 => x"05",
          6396 => x"34",
          6397 => x"80",
          6398 => x"18",
          6399 => x"56",
          6400 => x"76",
          6401 => x"83",
          6402 => x"2a",
          6403 => x"81",
          6404 => x"81",
          6405 => x"1a",
          6406 => x"41",
          6407 => x"e0",
          6408 => x"05",
          6409 => x"38",
          6410 => x"19",
          6411 => x"82",
          6412 => x"17",
          6413 => x"33",
          6414 => x"75",
          6415 => x"51",
          6416 => x"08",
          6417 => x"5c",
          6418 => x"80",
          6419 => x"38",
          6420 => x"09",
          6421 => x"ff",
          6422 => x"18",
          6423 => x"f3",
          6424 => x"2e",
          6425 => x"2a",
          6426 => x"88",
          6427 => x"7f",
          6428 => x"08",
          6429 => x"5c",
          6430 => x"52",
          6431 => x"bb",
          6432 => x"80",
          6433 => x"08",
          6434 => x"2e",
          6435 => x"5f",
          6436 => x"a8",
          6437 => x"52",
          6438 => x"3f",
          6439 => x"38",
          6440 => x"0c",
          6441 => x"08",
          6442 => x"17",
          6443 => x"38",
          6444 => x"3f",
          6445 => x"84",
          6446 => x"56",
          6447 => x"56",
          6448 => x"e5",
          6449 => x"bb",
          6450 => x"0b",
          6451 => x"04",
          6452 => x"98",
          6453 => x"58",
          6454 => x"84",
          6455 => x"bb",
          6456 => x"75",
          6457 => x"04",
          6458 => x"52",
          6459 => x"3f",
          6460 => x"2e",
          6461 => x"bb",
          6462 => x"08",
          6463 => x"08",
          6464 => x"fe",
          6465 => x"82",
          6466 => x"81",
          6467 => x"05",
          6468 => x"fe",
          6469 => x"39",
          6470 => x"17",
          6471 => x"fe",
          6472 => x"84",
          6473 => x"08",
          6474 => x"18",
          6475 => x"55",
          6476 => x"38",
          6477 => x"09",
          6478 => x"b4",
          6479 => x"7a",
          6480 => x"a4",
          6481 => x"3d",
          6482 => x"84",
          6483 => x"82",
          6484 => x"3d",
          6485 => x"84",
          6486 => x"2e",
          6487 => x"96",
          6488 => x"96",
          6489 => x"3f",
          6490 => x"84",
          6491 => x"33",
          6492 => x"d2",
          6493 => x"8b",
          6494 => x"07",
          6495 => x"34",
          6496 => x"78",
          6497 => x"84",
          6498 => x"0d",
          6499 => x"53",
          6500 => x"51",
          6501 => x"08",
          6502 => x"8a",
          6503 => x"3d",
          6504 => x"3d",
          6505 => x"84",
          6506 => x"08",
          6507 => x"81",
          6508 => x"38",
          6509 => x"71",
          6510 => x"96",
          6511 => x"97",
          6512 => x"98",
          6513 => x"99",
          6514 => x"18",
          6515 => x"84",
          6516 => x"96",
          6517 => x"6d",
          6518 => x"05",
          6519 => x"3f",
          6520 => x"08",
          6521 => x"80",
          6522 => x"8b",
          6523 => x"78",
          6524 => x"07",
          6525 => x"81",
          6526 => x"58",
          6527 => x"a4",
          6528 => x"16",
          6529 => x"16",
          6530 => x"09",
          6531 => x"76",
          6532 => x"51",
          6533 => x"08",
          6534 => x"59",
          6535 => x"bd",
          6536 => x"c3",
          6537 => x"e4",
          6538 => x"56",
          6539 => x"82",
          6540 => x"2b",
          6541 => x"88",
          6542 => x"5f",
          6543 => x"bb",
          6544 => x"5e",
          6545 => x"52",
          6546 => x"84",
          6547 => x"2e",
          6548 => x"81",
          6549 => x"80",
          6550 => x"16",
          6551 => x"17",
          6552 => x"77",
          6553 => x"09",
          6554 => x"84",
          6555 => x"a8",
          6556 => x"5a",
          6557 => x"ad",
          6558 => x"2e",
          6559 => x"54",
          6560 => x"53",
          6561 => x"dc",
          6562 => x"53",
          6563 => x"fe",
          6564 => x"80",
          6565 => x"75",
          6566 => x"84",
          6567 => x"08",
          6568 => x"84",
          6569 => x"79",
          6570 => x"56",
          6571 => x"8a",
          6572 => x"57",
          6573 => x"fc",
          6574 => x"33",
          6575 => x"38",
          6576 => x"39",
          6577 => x"ff",
          6578 => x"9d",
          6579 => x"84",
          6580 => x"3d",
          6581 => x"70",
          6582 => x"74",
          6583 => x"33",
          6584 => x"5a",
          6585 => x"3d",
          6586 => x"06",
          6587 => x"38",
          6588 => x"26",
          6589 => x"3f",
          6590 => x"51",
          6591 => x"83",
          6592 => x"81",
          6593 => x"e8",
          6594 => x"56",
          6595 => x"74",
          6596 => x"18",
          6597 => x"57",
          6598 => x"77",
          6599 => x"81",
          6600 => x"81",
          6601 => x"89",
          6602 => x"27",
          6603 => x"7b",
          6604 => x"5a",
          6605 => x"81",
          6606 => x"81",
          6607 => x"9f",
          6608 => x"57",
          6609 => x"38",
          6610 => x"05",
          6611 => x"7a",
          6612 => x"ff",
          6613 => x"80",
          6614 => x"56",
          6615 => x"08",
          6616 => x"b4",
          6617 => x"0c",
          6618 => x"74",
          6619 => x"08",
          6620 => x"f8",
          6621 => x"0c",
          6622 => x"33",
          6623 => x"51",
          6624 => x"08",
          6625 => x"38",
          6626 => x"6c",
          6627 => x"05",
          6628 => x"34",
          6629 => x"5d",
          6630 => x"fe",
          6631 => x"55",
          6632 => x"27",
          6633 => x"39",
          6634 => x"81",
          6635 => x"75",
          6636 => x"53",
          6637 => x"84",
          6638 => x"08",
          6639 => x"38",
          6640 => x"5a",
          6641 => x"18",
          6642 => x"33",
          6643 => x"81",
          6644 => x"18",
          6645 => x"fd",
          6646 => x"85",
          6647 => x"19",
          6648 => x"9c",
          6649 => x"74",
          6650 => x"30",
          6651 => x"74",
          6652 => x"5a",
          6653 => x"75",
          6654 => x"84",
          6655 => x"2e",
          6656 => x"2e",
          6657 => x"b9",
          6658 => x"70",
          6659 => x"74",
          6660 => x"17",
          6661 => x"76",
          6662 => x"81",
          6663 => x"80",
          6664 => x"05",
          6665 => x"34",
          6666 => x"d6",
          6667 => x"5d",
          6668 => x"fe",
          6669 => x"55",
          6670 => x"39",
          6671 => x"52",
          6672 => x"3f",
          6673 => x"81",
          6674 => x"08",
          6675 => x"19",
          6676 => x"27",
          6677 => x"82",
          6678 => x"59",
          6679 => x"75",
          6680 => x"84",
          6681 => x"2e",
          6682 => x"70",
          6683 => x"38",
          6684 => x"08",
          6685 => x"81",
          6686 => x"fd",
          6687 => x"02",
          6688 => x"5b",
          6689 => x"38",
          6690 => x"38",
          6691 => x"38",
          6692 => x"59",
          6693 => x"54",
          6694 => x"17",
          6695 => x"80",
          6696 => x"81",
          6697 => x"2a",
          6698 => x"81",
          6699 => x"89",
          6700 => x"59",
          6701 => x"06",
          6702 => x"84",
          6703 => x"79",
          6704 => x"27",
          6705 => x"83",
          6706 => x"80",
          6707 => x"c0",
          6708 => x"14",
          6709 => x"84",
          6710 => x"38",
          6711 => x"d8",
          6712 => x"38",
          6713 => x"38",
          6714 => x"38",
          6715 => x"84",
          6716 => x"84",
          6717 => x"81",
          6718 => x"84",
          6719 => x"fe",
          6720 => x"fe",
          6721 => x"38",
          6722 => x"ab",
          6723 => x"80",
          6724 => x"51",
          6725 => x"08",
          6726 => x"38",
          6727 => x"5e",
          6728 => x"0c",
          6729 => x"7a",
          6730 => x"90",
          6731 => x"90",
          6732 => x"94",
          6733 => x"fe",
          6734 => x"0c",
          6735 => x"84",
          6736 => x"ff",
          6737 => x"59",
          6738 => x"39",
          6739 => x"5e",
          6740 => x"e3",
          6741 => x"08",
          6742 => x"44",
          6743 => x"70",
          6744 => x"8a",
          6745 => x"70",
          6746 => x"85",
          6747 => x"2e",
          6748 => x"56",
          6749 => x"10",
          6750 => x"56",
          6751 => x"75",
          6752 => x"33",
          6753 => x"5d",
          6754 => x"3f",
          6755 => x"70",
          6756 => x"84",
          6757 => x"40",
          6758 => x"3d",
          6759 => x"fe",
          6760 => x"84",
          6761 => x"84",
          6762 => x"84",
          6763 => x"74",
          6764 => x"38",
          6765 => x"7e",
          6766 => x"ff",
          6767 => x"38",
          6768 => x"2a",
          6769 => x"5b",
          6770 => x"30",
          6771 => x"91",
          6772 => x"2e",
          6773 => x"60",
          6774 => x"81",
          6775 => x"38",
          6776 => x"fe",
          6777 => x"56",
          6778 => x"09",
          6779 => x"29",
          6780 => x"58",
          6781 => x"b6",
          6782 => x"71",
          6783 => x"14",
          6784 => x"33",
          6785 => x"33",
          6786 => x"88",
          6787 => x"07",
          6788 => x"a2",
          6789 => x"3d",
          6790 => x"41",
          6791 => x"ff",
          6792 => x"7a",
          6793 => x"81",
          6794 => x"80",
          6795 => x"45",
          6796 => x"06",
          6797 => x"70",
          6798 => x"83",
          6799 => x"78",
          6800 => x"a8",
          6801 => x"38",
          6802 => x"a8",
          6803 => x"57",
          6804 => x"76",
          6805 => x"51",
          6806 => x"08",
          6807 => x"08",
          6808 => x"84",
          6809 => x"08",
          6810 => x"57",
          6811 => x"5d",
          6812 => x"11",
          6813 => x"6b",
          6814 => x"62",
          6815 => x"5d",
          6816 => x"56",
          6817 => x"78",
          6818 => x"68",
          6819 => x"84",
          6820 => x"89",
          6821 => x"06",
          6822 => x"84",
          6823 => x"7a",
          6824 => x"80",
          6825 => x"fe",
          6826 => x"84",
          6827 => x"0c",
          6828 => x"0b",
          6829 => x"84",
          6830 => x"11",
          6831 => x"74",
          6832 => x"81",
          6833 => x"7a",
          6834 => x"e6",
          6835 => x"5b",
          6836 => x"70",
          6837 => x"45",
          6838 => x"e0",
          6839 => x"ff",
          6840 => x"38",
          6841 => x"46",
          6842 => x"76",
          6843 => x"78",
          6844 => x"30",
          6845 => x"5d",
          6846 => x"38",
          6847 => x"7c",
          6848 => x"e0",
          6849 => x"52",
          6850 => x"57",
          6851 => x"61",
          6852 => x"08",
          6853 => x"6c",
          6854 => x"9c",
          6855 => x"39",
          6856 => x"24",
          6857 => x"0c",
          6858 => x"48",
          6859 => x"38",
          6860 => x"fc",
          6861 => x"f5",
          6862 => x"18",
          6863 => x"38",
          6864 => x"9f",
          6865 => x"80",
          6866 => x"9f",
          6867 => x"06",
          6868 => x"84",
          6869 => x"81",
          6870 => x"f4",
          6871 => x"57",
          6872 => x"76",
          6873 => x"55",
          6874 => x"74",
          6875 => x"77",
          6876 => x"ff",
          6877 => x"6a",
          6878 => x"34",
          6879 => x"32",
          6880 => x"05",
          6881 => x"68",
          6882 => x"83",
          6883 => x"83",
          6884 => x"05",
          6885 => x"94",
          6886 => x"bf",
          6887 => x"05",
          6888 => x"61",
          6889 => x"34",
          6890 => x"05",
          6891 => x"9e",
          6892 => x"90",
          6893 => x"05",
          6894 => x"80",
          6895 => x"05",
          6896 => x"cc",
          6897 => x"ff",
          6898 => x"74",
          6899 => x"34",
          6900 => x"61",
          6901 => x"83",
          6902 => x"81",
          6903 => x"58",
          6904 => x"60",
          6905 => x"34",
          6906 => x"6b",
          6907 => x"79",
          6908 => x"84",
          6909 => x"17",
          6910 => x"69",
          6911 => x"05",
          6912 => x"38",
          6913 => x"86",
          6914 => x"62",
          6915 => x"61",
          6916 => x"74",
          6917 => x"90",
          6918 => x"46",
          6919 => x"34",
          6920 => x"83",
          6921 => x"60",
          6922 => x"84",
          6923 => x"80",
          6924 => x"05",
          6925 => x"38",
          6926 => x"76",
          6927 => x"80",
          6928 => x"83",
          6929 => x"75",
          6930 => x"54",
          6931 => x"c5",
          6932 => x"9b",
          6933 => x"5b",
          6934 => x"2e",
          6935 => x"ff",
          6936 => x"2e",
          6937 => x"38",
          6938 => x"81",
          6939 => x"80",
          6940 => x"19",
          6941 => x"34",
          6942 => x"05",
          6943 => x"05",
          6944 => x"67",
          6945 => x"34",
          6946 => x"1f",
          6947 => x"85",
          6948 => x"2a",
          6949 => x"34",
          6950 => x"34",
          6951 => x"61",
          6952 => x"c8",
          6953 => x"83",
          6954 => x"05",
          6955 => x"83",
          6956 => x"77",
          6957 => x"2a",
          6958 => x"81",
          6959 => x"fe",
          6960 => x"84",
          6961 => x"52",
          6962 => x"57",
          6963 => x"84",
          6964 => x"9f",
          6965 => x"62",
          6966 => x"16",
          6967 => x"38",
          6968 => x"e8",
          6969 => x"9d",
          6970 => x"e8",
          6971 => x"22",
          6972 => x"38",
          6973 => x"78",
          6974 => x"84",
          6975 => x"89",
          6976 => x"84",
          6977 => x"58",
          6978 => x"f5",
          6979 => x"84",
          6980 => x"f8",
          6981 => x"81",
          6982 => x"57",
          6983 => x"63",
          6984 => x"f4",
          6985 => x"75",
          6986 => x"34",
          6987 => x"05",
          6988 => x"a3",
          6989 => x"80",
          6990 => x"05",
          6991 => x"80",
          6992 => x"61",
          6993 => x"7b",
          6994 => x"59",
          6995 => x"2a",
          6996 => x"61",
          6997 => x"34",
          6998 => x"af",
          6999 => x"80",
          7000 => x"05",
          7001 => x"80",
          7002 => x"80",
          7003 => x"05",
          7004 => x"70",
          7005 => x"05",
          7006 => x"2e",
          7007 => x"58",
          7008 => x"ff",
          7009 => x"39",
          7010 => x"51",
          7011 => x"bb",
          7012 => x"29",
          7013 => x"05",
          7014 => x"53",
          7015 => x"3f",
          7016 => x"84",
          7017 => x"0c",
          7018 => x"6a",
          7019 => x"70",
          7020 => x"ff",
          7021 => x"05",
          7022 => x"61",
          7023 => x"34",
          7024 => x"8a",
          7025 => x"f9",
          7026 => x"60",
          7027 => x"84",
          7028 => x"81",
          7029 => x"f4",
          7030 => x"81",
          7031 => x"75",
          7032 => x"75",
          7033 => x"75",
          7034 => x"34",
          7035 => x"80",
          7036 => x"e1",
          7037 => x"05",
          7038 => x"7a",
          7039 => x"05",
          7040 => x"83",
          7041 => x"7f",
          7042 => x"83",
          7043 => x"05",
          7044 => x"76",
          7045 => x"69",
          7046 => x"87",
          7047 => x"bd",
          7048 => x"60",
          7049 => x"69",
          7050 => x"3d",
          7051 => x"61",
          7052 => x"25",
          7053 => x"f8",
          7054 => x"51",
          7055 => x"09",
          7056 => x"55",
          7057 => x"70",
          7058 => x"74",
          7059 => x"cd",
          7060 => x"83",
          7061 => x"0c",
          7062 => x"7b",
          7063 => x"57",
          7064 => x"17",
          7065 => x"88",
          7066 => x"59",
          7067 => x"bb",
          7068 => x"81",
          7069 => x"04",
          7070 => x"8c",
          7071 => x"a7",
          7072 => x"72",
          7073 => x"0c",
          7074 => x"56",
          7075 => x"94",
          7076 => x"02",
          7077 => x"58",
          7078 => x"70",
          7079 => x"74",
          7080 => x"77",
          7081 => x"80",
          7082 => x"17",
          7083 => x"81",
          7084 => x"74",
          7085 => x"0c",
          7086 => x"9f",
          7087 => x"c0",
          7088 => x"9f",
          7089 => x"7c",
          7090 => x"bb",
          7091 => x"3d",
          7092 => x"05",
          7093 => x"3f",
          7094 => x"07",
          7095 => x"56",
          7096 => x"fd",
          7097 => x"bb",
          7098 => x"3d",
          7099 => x"22",
          7100 => x"26",
          7101 => x"52",
          7102 => x"0d",
          7103 => x"70",
          7104 => x"38",
          7105 => x"c8",
          7106 => x"81",
          7107 => x"54",
          7108 => x"10",
          7109 => x"51",
          7110 => x"ff",
          7111 => x"3d",
          7112 => x"05",
          7113 => x"53",
          7114 => x"8c",
          7115 => x"0c",
          7116 => x"2e",
          7117 => x"ff",
          7118 => x"c8",
          7119 => x"51",
          7120 => x"77",
          7121 => x"e1",
          7122 => x"ea",
          7123 => x"80",
          7124 => x"22",
          7125 => x"7a",
          7126 => x"b7",
          7127 => x"72",
          7128 => x"06",
          7129 => x"b1",
          7130 => x"70",
          7131 => x"30",
          7132 => x"53",
          7133 => x"75",
          7134 => x"3d",
          7135 => x"a2",
          7136 => x"10",
          7137 => x"08",
          7138 => x"ff",
          7139 => x"ff",
          7140 => x"57",
          7141 => x"ff",
          7142 => x"16",
          7143 => x"db",
          7144 => x"06",
          7145 => x"83",
          7146 => x"f0",
          7147 => x"51",
          7148 => x"06",
          7149 => x"06",
          7150 => x"73",
          7151 => x"52",
          7152 => x"ff",
          7153 => x"ff",
          7154 => x"00",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"00",
          7372 => x"00",
          7373 => x"00",
          7374 => x"00",
          7375 => x"00",
          7376 => x"00",
          7377 => x"00",
          7378 => x"00",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"00",
          7383 => x"00",
          7384 => x"00",
          7385 => x"00",
          7386 => x"00",
          7387 => x"00",
          7388 => x"00",
          7389 => x"00",
          7390 => x"00",
          7391 => x"00",
          7392 => x"6c",
          7393 => x"00",
          7394 => x"00",
          7395 => x"00",
          7396 => x"72",
          7397 => x"00",
          7398 => x"00",
          7399 => x"00",
          7400 => x"65",
          7401 => x"69",
          7402 => x"66",
          7403 => x"61",
          7404 => x"6d",
          7405 => x"72",
          7406 => x"00",
          7407 => x"00",
          7408 => x"00",
          7409 => x"38",
          7410 => x"63",
          7411 => x"63",
          7412 => x"00",
          7413 => x"6e",
          7414 => x"72",
          7415 => x"61",
          7416 => x"73",
          7417 => x"65",
          7418 => x"6f",
          7419 => x"6f",
          7420 => x"65",
          7421 => x"6e",
          7422 => x"65",
          7423 => x"72",
          7424 => x"69",
          7425 => x"6f",
          7426 => x"69",
          7427 => x"6f",
          7428 => x"6e",
          7429 => x"6c",
          7430 => x"6f",
          7431 => x"6f",
          7432 => x"6f",
          7433 => x"69",
          7434 => x"65",
          7435 => x"66",
          7436 => x"20",
          7437 => x"69",
          7438 => x"65",
          7439 => x"00",
          7440 => x"20",
          7441 => x"69",
          7442 => x"69",
          7443 => x"44",
          7444 => x"74",
          7445 => x"63",
          7446 => x"69",
          7447 => x"6c",
          7448 => x"69",
          7449 => x"69",
          7450 => x"61",
          7451 => x"74",
          7452 => x"63",
          7453 => x"6e",
          7454 => x"6e",
          7455 => x"69",
          7456 => x"00",
          7457 => x"74",
          7458 => x"2e",
          7459 => x"6c",
          7460 => x"2e",
          7461 => x"6e",
          7462 => x"79",
          7463 => x"6e",
          7464 => x"72",
          7465 => x"45",
          7466 => x"75",
          7467 => x"00",
          7468 => x"62",
          7469 => x"20",
          7470 => x"62",
          7471 => x"63",
          7472 => x"65",
          7473 => x"30",
          7474 => x"20",
          7475 => x"00",
          7476 => x"00",
          7477 => x"30",
          7478 => x"20",
          7479 => x"00",
          7480 => x"2a",
          7481 => x"35",
          7482 => x"31",
          7483 => x"00",
          7484 => x"20",
          7485 => x"78",
          7486 => x"20",
          7487 => x"53",
          7488 => x"61",
          7489 => x"65",
          7490 => x"20",
          7491 => x"3d",
          7492 => x"00",
          7493 => x"70",
          7494 => x"73",
          7495 => x"20",
          7496 => x"3d",
          7497 => x"00",
          7498 => x"6e",
          7499 => x"20",
          7500 => x"00",
          7501 => x"20",
          7502 => x"72",
          7503 => x"41",
          7504 => x"69",
          7505 => x"74",
          7506 => x"20",
          7507 => x"72",
          7508 => x"41",
          7509 => x"69",
          7510 => x"74",
          7511 => x"20",
          7512 => x"72",
          7513 => x"4f",
          7514 => x"69",
          7515 => x"74",
          7516 => x"6e",
          7517 => x"00",
          7518 => x"20",
          7519 => x"70",
          7520 => x"6e",
          7521 => x"6d",
          7522 => x"6e",
          7523 => x"74",
          7524 => x"00",
          7525 => x"78",
          7526 => x"00",
          7527 => x"70",
          7528 => x"61",
          7529 => x"20",
          7530 => x"69",
          7531 => x"61",
          7532 => x"6c",
          7533 => x"69",
          7534 => x"6c",
          7535 => x"20",
          7536 => x"73",
          7537 => x"61",
          7538 => x"6e",
          7539 => x"50",
          7540 => x"64",
          7541 => x"2e",
          7542 => x"6f",
          7543 => x"6f",
          7544 => x"00",
          7545 => x"72",
          7546 => x"70",
          7547 => x"6e",
          7548 => x"61",
          7549 => x"6f",
          7550 => x"38",
          7551 => x"00",
          7552 => x"72",
          7553 => x"20",
          7554 => x"64",
          7555 => x"78",
          7556 => x"20",
          7557 => x"25",
          7558 => x"2e",
          7559 => x"20",
          7560 => x"00",
          7561 => x"20",
          7562 => x"6f",
          7563 => x"2e",
          7564 => x"30",
          7565 => x"78",
          7566 => x"78",
          7567 => x"00",
          7568 => x"6e",
          7569 => x"30",
          7570 => x"58",
          7571 => x"69",
          7572 => x"00",
          7573 => x"4d",
          7574 => x"43",
          7575 => x"2e",
          7576 => x"73",
          7577 => x"65",
          7578 => x"68",
          7579 => x"20",
          7580 => x"70",
          7581 => x"63",
          7582 => x"00",
          7583 => x"64",
          7584 => x"25",
          7585 => x"2e",
          7586 => x"6f",
          7587 => x"67",
          7588 => x"00",
          7589 => x"69",
          7590 => x"6c",
          7591 => x"3a",
          7592 => x"73",
          7593 => x"20",
          7594 => x"65",
          7595 => x"74",
          7596 => x"65",
          7597 => x"38",
          7598 => x"20",
          7599 => x"65",
          7600 => x"61",
          7601 => x"65",
          7602 => x"38",
          7603 => x"20",
          7604 => x"20",
          7605 => x"64",
          7606 => x"20",
          7607 => x"38",
          7608 => x"69",
          7609 => x"20",
          7610 => x"64",
          7611 => x"20",
          7612 => x"20",
          7613 => x"34",
          7614 => x"20",
          7615 => x"6d",
          7616 => x"46",
          7617 => x"20",
          7618 => x"2e",
          7619 => x"0a",
          7620 => x"69",
          7621 => x"53",
          7622 => x"6f",
          7623 => x"3d",
          7624 => x"64",
          7625 => x"20",
          7626 => x"20",
          7627 => x"72",
          7628 => x"20",
          7629 => x"2e",
          7630 => x"0a",
          7631 => x"50",
          7632 => x"53",
          7633 => x"4f",
          7634 => x"20",
          7635 => x"43",
          7636 => x"49",
          7637 => x"42",
          7638 => x"20",
          7639 => x"43",
          7640 => x"61",
          7641 => x"30",
          7642 => x"20",
          7643 => x"31",
          7644 => x"6d",
          7645 => x"30",
          7646 => x"20",
          7647 => x"52",
          7648 => x"76",
          7649 => x"30",
          7650 => x"20",
          7651 => x"20",
          7652 => x"38",
          7653 => x"2e",
          7654 => x"52",
          7655 => x"20",
          7656 => x"30",
          7657 => x"20",
          7658 => x"42",
          7659 => x"38",
          7660 => x"2e",
          7661 => x"44",
          7662 => x"20",
          7663 => x"30",
          7664 => x"20",
          7665 => x"52",
          7666 => x"38",
          7667 => x"2e",
          7668 => x"6d",
          7669 => x"6e",
          7670 => x"6e",
          7671 => x"56",
          7672 => x"6d",
          7673 => x"65",
          7674 => x"6c",
          7675 => x"56",
          7676 => x"00",
          7677 => x"00",
          7678 => x"00",
          7679 => x"00",
          7680 => x"00",
          7681 => x"00",
          7682 => x"00",
          7683 => x"00",
          7684 => x"00",
          7685 => x"00",
          7686 => x"00",
          7687 => x"00",
          7688 => x"00",
          7689 => x"00",
          7690 => x"00",
          7691 => x"00",
          7692 => x"00",
          7693 => x"00",
          7694 => x"00",
          7695 => x"00",
          7696 => x"00",
          7697 => x"00",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"00",
          7703 => x"00",
          7704 => x"00",
          7705 => x"00",
          7706 => x"00",
          7707 => x"00",
          7708 => x"00",
          7709 => x"5b",
          7710 => x"5b",
          7711 => x"5b",
          7712 => x"30",
          7713 => x"5b",
          7714 => x"00",
          7715 => x"00",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"72",
          7721 => x"25",
          7722 => x"61",
          7723 => x"65",
          7724 => x"65",
          7725 => x"79",
          7726 => x"64",
          7727 => x"67",
          7728 => x"72",
          7729 => x"00",
          7730 => x"69",
          7731 => x"75",
          7732 => x"38",
          7733 => x"30",
          7734 => x"0a",
          7735 => x"64",
          7736 => x"65",
          7737 => x"69",
          7738 => x"69",
          7739 => x"4f",
          7740 => x"25",
          7741 => x"5b",
          7742 => x"5b",
          7743 => x"5b",
          7744 => x"5b",
          7745 => x"5b",
          7746 => x"5b",
          7747 => x"5b",
          7748 => x"5b",
          7749 => x"5b",
          7750 => x"5b",
          7751 => x"5b",
          7752 => x"5b",
          7753 => x"5b",
          7754 => x"5b",
          7755 => x"5b",
          7756 => x"5b",
          7757 => x"00",
          7758 => x"00",
          7759 => x"25",
          7760 => x"2c",
          7761 => x"30",
          7762 => x"3a",
          7763 => x"64",
          7764 => x"25",
          7765 => x"64",
          7766 => x"00",
          7767 => x"00",
          7768 => x"3b",
          7769 => x"65",
          7770 => x"72",
          7771 => x"70",
          7772 => x"30",
          7773 => x"77",
          7774 => x"30",
          7775 => x"64",
          7776 => x"00",
          7777 => x"73",
          7778 => x"65",
          7779 => x"44",
          7780 => x"3f",
          7781 => x"2c",
          7782 => x"41",
          7783 => x"00",
          7784 => x"44",
          7785 => x"4f",
          7786 => x"20",
          7787 => x"20",
          7788 => x"4d",
          7789 => x"54",
          7790 => x"00",
          7791 => x"00",
          7792 => x"03",
          7793 => x"16",
          7794 => x"9a",
          7795 => x"45",
          7796 => x"92",
          7797 => x"99",
          7798 => x"49",
          7799 => x"a9",
          7800 => x"b1",
          7801 => x"b9",
          7802 => x"c1",
          7803 => x"c9",
          7804 => x"d1",
          7805 => x"d9",
          7806 => x"e1",
          7807 => x"e9",
          7808 => x"f1",
          7809 => x"f9",
          7810 => x"2e",
          7811 => x"22",
          7812 => x"00",
          7813 => x"10",
          7814 => x"00",
          7815 => x"04",
          7816 => x"00",
          7817 => x"e9",
          7818 => x"e5",
          7819 => x"e8",
          7820 => x"c4",
          7821 => x"c6",
          7822 => x"fb",
          7823 => x"dc",
          7824 => x"a7",
          7825 => x"f3",
          7826 => x"aa",
          7827 => x"ac",
          7828 => x"ab",
          7829 => x"93",
          7830 => x"62",
          7831 => x"51",
          7832 => x"5b",
          7833 => x"2c",
          7834 => x"5e",
          7835 => x"69",
          7836 => x"6c",
          7837 => x"65",
          7838 => x"53",
          7839 => x"0c",
          7840 => x"90",
          7841 => x"93",
          7842 => x"b5",
          7843 => x"a9",
          7844 => x"b5",
          7845 => x"65",
          7846 => x"f7",
          7847 => x"b7",
          7848 => x"a0",
          7849 => x"e0",
          7850 => x"ff",
          7851 => x"30",
          7852 => x"10",
          7853 => x"06",
          7854 => x"81",
          7855 => x"84",
          7856 => x"89",
          7857 => x"8d",
          7858 => x"91",
          7859 => x"f6",
          7860 => x"98",
          7861 => x"9d",
          7862 => x"a0",
          7863 => x"a4",
          7864 => x"a9",
          7865 => x"ac",
          7866 => x"b1",
          7867 => x"b5",
          7868 => x"b8",
          7869 => x"bc",
          7870 => x"c1",
          7871 => x"c5",
          7872 => x"c7",
          7873 => x"cd",
          7874 => x"8e",
          7875 => x"03",
          7876 => x"f8",
          7877 => x"3a",
          7878 => x"3b",
          7879 => x"40",
          7880 => x"0a",
          7881 => x"86",
          7882 => x"58",
          7883 => x"5c",
          7884 => x"93",
          7885 => x"64",
          7886 => x"97",
          7887 => x"6c",
          7888 => x"70",
          7889 => x"74",
          7890 => x"78",
          7891 => x"7c",
          7892 => x"a6",
          7893 => x"84",
          7894 => x"ae",
          7895 => x"45",
          7896 => x"90",
          7897 => x"03",
          7898 => x"ac",
          7899 => x"89",
          7900 => x"c2",
          7901 => x"c4",
          7902 => x"8c",
          7903 => x"18",
          7904 => x"f3",
          7905 => x"f7",
          7906 => x"fa",
          7907 => x"10",
          7908 => x"36",
          7909 => x"01",
          7910 => x"61",
          7911 => x"7d",
          7912 => x"96",
          7913 => x"08",
          7914 => x"08",
          7915 => x"06",
          7916 => x"52",
          7917 => x"56",
          7918 => x"70",
          7919 => x"c8",
          7920 => x"da",
          7921 => x"ea",
          7922 => x"80",
          7923 => x"a0",
          7924 => x"b8",
          7925 => x"cc",
          7926 => x"02",
          7927 => x"01",
          7928 => x"fc",
          7929 => x"70",
          7930 => x"83",
          7931 => x"2f",
          7932 => x"06",
          7933 => x"64",
          7934 => x"1a",
          7935 => x"00",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"00",
          7940 => x"00",
          7941 => x"00",
          7942 => x"00",
          7943 => x"00",
          7944 => x"00",
          7945 => x"00",
          7946 => x"00",
          7947 => x"00",
          7948 => x"00",
          7949 => x"00",
          7950 => x"00",
          7951 => x"00",
          7952 => x"00",
          7953 => x"00",
          7954 => x"00",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"00",
          7959 => x"00",
          7960 => x"00",
          7961 => x"00",
          7962 => x"00",
          7963 => x"00",
          7964 => x"00",
          7965 => x"00",
          7966 => x"00",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"00",
          7983 => x"00",
          7984 => x"00",
          7985 => x"00",
          7986 => x"00",
          7987 => x"00",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"81",
          7996 => x"7f",
          7997 => x"00",
          7998 => x"00",
          7999 => x"f5",
          8000 => x"00",
          8001 => x"01",
          8002 => x"00",
          8003 => x"00",
          8004 => x"00",
          8005 => x"00",
          8006 => x"00",
          8007 => x"00",
          8008 => x"00",
          8009 => x"00",
          8010 => x"00",
          8011 => x"00",
          8012 => x"00",
          8013 => x"00",
          8014 => x"00",
          8015 => x"00",
          8016 => x"00",
          8017 => x"00",
          8018 => x"fc",
          8019 => x"7a",
          8020 => x"72",
          8021 => x"6a",
          8022 => x"62",
          8023 => x"32",
          8024 => x"f3",
          8025 => x"7f",
          8026 => x"f0",
          8027 => x"81",
          8028 => x"fc",
          8029 => x"5a",
          8030 => x"52",
          8031 => x"4a",
          8032 => x"42",
          8033 => x"32",
          8034 => x"f3",
          8035 => x"7f",
          8036 => x"f0",
          8037 => x"81",
          8038 => x"fc",
          8039 => x"5a",
          8040 => x"52",
          8041 => x"4a",
          8042 => x"42",
          8043 => x"22",
          8044 => x"7e",
          8045 => x"e2",
          8046 => x"f0",
          8047 => x"86",
          8048 => x"fe",
          8049 => x"1a",
          8050 => x"12",
          8051 => x"0a",
          8052 => x"02",
          8053 => x"f0",
          8054 => x"1e",
          8055 => x"f0",
          8056 => x"f0",
          8057 => x"81",
          8058 => x"f0",
          8059 => x"77",
          8060 => x"70",
          8061 => x"5d",
          8062 => x"6e",
          8063 => x"36",
          8064 => x"9f",
          8065 => x"c5",
          8066 => x"f0",
          8067 => x"81",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"cf",
          9105 => x"fd",
          9106 => x"c5",
          9107 => x"ee",
          9108 => x"65",
          9109 => x"2a",
          9110 => x"25",
          9111 => x"2b",
          9112 => x"05",
          9113 => x"0d",
          9114 => x"15",
          9115 => x"54",
          9116 => x"85",
          9117 => x"8d",
          9118 => x"95",
          9119 => x"40",
          9120 => x"00",
          9121 => x"00",
          9122 => x"00",
          9123 => x"00",
          9124 => x"00",
          9125 => x"00",
          9126 => x"00",
          9127 => x"00",
          9128 => x"00",
          9129 => x"00",
          9130 => x"00",
          9131 => x"00",
          9132 => x"00",
          9133 => x"00",
          9134 => x"00",
          9135 => x"04",
          9136 => x"04",
        others => X"00"
    );

    shared variable RAM7 : ramArray :=
    (
             0 => x"f8",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"90",
             5 => x"8c",
             6 => x"00",
             7 => x"00",
             8 => x"72",
             9 => x"83",
            10 => x"04",
            11 => x"00",
            12 => x"83",
            13 => x"05",
            14 => x"73",
            15 => x"83",
            16 => x"72",
            17 => x"73",
            18 => x"53",
            19 => x"00",
            20 => x"73",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"0a",
            26 => x"05",
            27 => x"04",
            28 => x"73",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"cd",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"0a",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"09",
            45 => x"05",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"81",
            50 => x"04",
            51 => x"00",
            52 => x"04",
            53 => x"82",
            54 => x"fc",
            55 => x"00",
            56 => x"72",
            57 => x"0a",
            58 => x"00",
            59 => x"00",
            60 => x"72",
            61 => x"0a",
            62 => x"00",
            63 => x"00",
            64 => x"52",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"05",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"73",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"72",
            77 => x"10",
            78 => x"04",
            79 => x"00",
            80 => x"0b",
            81 => x"10",
            82 => x"93",
            83 => x"00",
            84 => x"90",
            85 => x"cc",
            86 => x"0c",
            87 => x"00",
            88 => x"90",
            89 => x"ab",
            90 => x"0c",
            91 => x"00",
            92 => x"05",
            93 => x"70",
            94 => x"05",
            95 => x"04",
            96 => x"05",
            97 => x"05",
            98 => x"74",
            99 => x"51",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"04",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"10",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"05",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"81",
           133 => x"0b",
           134 => x"0b",
           135 => x"b6",
           136 => x"0b",
           137 => x"0b",
           138 => x"f6",
           139 => x"0b",
           140 => x"0b",
           141 => x"b6",
           142 => x"0b",
           143 => x"0b",
           144 => x"f9",
           145 => x"0b",
           146 => x"0b",
           147 => x"bd",
           148 => x"0b",
           149 => x"0b",
           150 => x"81",
           151 => x"0b",
           152 => x"0b",
           153 => x"c5",
           154 => x"0b",
           155 => x"0b",
           156 => x"89",
           157 => x"0b",
           158 => x"0b",
           159 => x"cd",
           160 => x"0b",
           161 => x"0b",
           162 => x"91",
           163 => x"0b",
           164 => x"0b",
           165 => x"d5",
           166 => x"0b",
           167 => x"0b",
           168 => x"99",
           169 => x"0b",
           170 => x"0b",
           171 => x"dc",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"04",
           193 => x"2d",
           194 => x"90",
           195 => x"2d",
           196 => x"90",
           197 => x"2d",
           198 => x"90",
           199 => x"2d",
           200 => x"90",
           201 => x"2d",
           202 => x"90",
           203 => x"2d",
           204 => x"90",
           205 => x"2d",
           206 => x"90",
           207 => x"2d",
           208 => x"90",
           209 => x"2d",
           210 => x"90",
           211 => x"2d",
           212 => x"90",
           213 => x"2d",
           214 => x"90",
           215 => x"2d",
           216 => x"90",
           217 => x"fc",
           218 => x"80",
           219 => x"d5",
           220 => x"c0",
           221 => x"80",
           222 => x"80",
           223 => x"0c",
           224 => x"08",
           225 => x"90",
           226 => x"90",
           227 => x"bb",
           228 => x"bb",
           229 => x"84",
           230 => x"84",
           231 => x"04",
           232 => x"2d",
           233 => x"90",
           234 => x"a6",
           235 => x"80",
           236 => x"fa",
           237 => x"c0",
           238 => x"82",
           239 => x"80",
           240 => x"0c",
           241 => x"08",
           242 => x"90",
           243 => x"90",
           244 => x"bb",
           245 => x"bb",
           246 => x"84",
           247 => x"84",
           248 => x"04",
           249 => x"2d",
           250 => x"90",
           251 => x"95",
           252 => x"80",
           253 => x"f6",
           254 => x"c0",
           255 => x"83",
           256 => x"80",
           257 => x"0c",
           258 => x"08",
           259 => x"90",
           260 => x"90",
           261 => x"bb",
           262 => x"bb",
           263 => x"84",
           264 => x"84",
           265 => x"04",
           266 => x"2d",
           267 => x"90",
           268 => x"a9",
           269 => x"80",
           270 => x"9b",
           271 => x"c0",
           272 => x"83",
           273 => x"80",
           274 => x"0c",
           275 => x"08",
           276 => x"90",
           277 => x"90",
           278 => x"bb",
           279 => x"bb",
           280 => x"84",
           281 => x"84",
           282 => x"04",
           283 => x"2d",
           284 => x"90",
           285 => x"aa",
           286 => x"80",
           287 => x"f7",
           288 => x"c0",
           289 => x"80",
           290 => x"80",
           291 => x"0c",
           292 => x"08",
           293 => x"90",
           294 => x"90",
           295 => x"bb",
           296 => x"90",
           297 => x"bb",
           298 => x"bb",
           299 => x"84",
           300 => x"84",
           301 => x"04",
           302 => x"2d",
           303 => x"90",
           304 => x"d9",
           305 => x"80",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"00",
           311 => x"09",
           312 => x"2b",
           313 => x"04",
           314 => x"05",
           315 => x"72",
           316 => x"51",
           317 => x"70",
           318 => x"71",
           319 => x"0b",
           320 => x"ce",
           321 => x"3d",
           322 => x"53",
           323 => x"81",
           324 => x"3d",
           325 => x"81",
           326 => x"56",
           327 => x"2e",
           328 => x"14",
           329 => x"72",
           330 => x"54",
           331 => x"2e",
           332 => x"84",
           333 => x"08",
           334 => x"08",
           335 => x"14",
           336 => x"07",
           337 => x"80",
           338 => x"52",
           339 => x"0d",
           340 => x"88",
           341 => x"54",
           342 => x"73",
           343 => x"05",
           344 => x"51",
           345 => x"34",
           346 => x"86",
           347 => x"51",
           348 => x"3d",
           349 => x"80",
           350 => x"70",
           351 => x"55",
           352 => x"81",
           353 => x"76",
           354 => x"7b",
           355 => x"81",
           356 => x"26",
           357 => x"30",
           358 => x"ae",
           359 => x"83",
           360 => x"54",
           361 => x"80",
           362 => x"bd",
           363 => x"bb",
           364 => x"83",
           365 => x"10",
           366 => x"19",
           367 => x"05",
           368 => x"5f",
           369 => x"81",
           370 => x"7c",
           371 => x"ff",
           372 => x"06",
           373 => x"5b",
           374 => x"dd",
           375 => x"51",
           376 => x"fe",
           377 => x"2a",
           378 => x"38",
           379 => x"95",
           380 => x"26",
           381 => x"94",
           382 => x"18",
           383 => x"38",
           384 => x"80",
           385 => x"38",
           386 => x"f6",
           387 => x"71",
           388 => x"58",
           389 => x"52",
           390 => x"84",
           391 => x"08",
           392 => x"26",
           393 => x"05",
           394 => x"34",
           395 => x"84",
           396 => x"08",
           397 => x"98",
           398 => x"80",
           399 => x"29",
           400 => x"59",
           401 => x"55",
           402 => x"84",
           403 => x"53",
           404 => x"80",
           405 => x"72",
           406 => x"81",
           407 => x"38",
           408 => x"54",
           409 => x"7a",
           410 => x"71",
           411 => x"06",
           412 => x"77",
           413 => x"7c",
           414 => x"80",
           415 => x"81",
           416 => x"84",
           417 => x"38",
           418 => x"86",
           419 => x"85",
           420 => x"5f",
           421 => x"84",
           422 => x"70",
           423 => x"25",
           424 => x"a9",
           425 => x"fc",
           426 => x"40",
           427 => x"81",
           428 => x"78",
           429 => x"0a",
           430 => x"80",
           431 => x"51",
           432 => x"0a",
           433 => x"2c",
           434 => x"38",
           435 => x"55",
           436 => x"80",
           437 => x"f3",
           438 => x"2e",
           439 => x"2e",
           440 => x"33",
           441 => x"bb",
           442 => x"74",
           443 => x"a7",
           444 => x"fc",
           445 => x"40",
           446 => x"7c",
           447 => x"39",
           448 => x"7c",
           449 => x"fa",
           450 => x"80",
           451 => x"71",
           452 => x"59",
           453 => x"60",
           454 => x"83",
           455 => x"7c",
           456 => x"05",
           457 => x"57",
           458 => x"06",
           459 => x"78",
           460 => x"05",
           461 => x"7f",
           462 => x"51",
           463 => x"70",
           464 => x"83",
           465 => x"52",
           466 => x"85",
           467 => x"83",
           468 => x"ff",
           469 => x"75",
           470 => x"b9",
           471 => x"81",
           472 => x"29",
           473 => x"5a",
           474 => x"70",
           475 => x"c6",
           476 => x"05",
           477 => x"80",
           478 => x"ff",
           479 => x"fa",
           480 => x"58",
           481 => x"39",
           482 => x"58",
           483 => x"39",
           484 => x"81",
           485 => x"8a",
           486 => x"bb",
           487 => x"71",
           488 => x"2c",
           489 => x"07",
           490 => x"38",
           491 => x"71",
           492 => x"54",
           493 => x"bb",
           494 => x"ff",
           495 => x"5a",
           496 => x"33",
           497 => x"c9",
           498 => x"fc",
           499 => x"54",
           500 => x"7c",
           501 => x"39",
           502 => x"79",
           503 => x"38",
           504 => x"7a",
           505 => x"2e",
           506 => x"98",
           507 => x"90",
           508 => x"51",
           509 => x"39",
           510 => x"7e",
           511 => x"a2",
           512 => x"98",
           513 => x"06",
           514 => x"fb",
           515 => x"70",
           516 => x"7c",
           517 => x"39",
           518 => x"ff",
           519 => x"8b",
           520 => x"ff",
           521 => x"5a",
           522 => x"30",
           523 => x"5b",
           524 => x"e6",
           525 => x"f3",
           526 => x"3d",
           527 => x"e8",
           528 => x"81",
           529 => x"55",
           530 => x"81",
           531 => x"05",
           532 => x"38",
           533 => x"90",
           534 => x"84",
           535 => x"74",
           536 => x"80",
           537 => x"54",
           538 => x"84",
           539 => x"14",
           540 => x"08",
           541 => x"56",
           542 => x"0d",
           543 => x"54",
           544 => x"2a",
           545 => x"57",
           546 => x"81",
           547 => x"55",
           548 => x"06",
           549 => x"84",
           550 => x"81",
           551 => x"ea",
           552 => x"08",
           553 => x"80",
           554 => x"05",
           555 => x"ca",
           556 => x"08",
           557 => x"0d",
           558 => x"11",
           559 => x"06",
           560 => x"ae",
           561 => x"73",
           562 => x"53",
           563 => x"74",
           564 => x"81",
           565 => x"81",
           566 => x"84",
           567 => x"74",
           568 => x"15",
           569 => x"bb",
           570 => x"81",
           571 => x"39",
           572 => x"70",
           573 => x"06",
           574 => x"b3",
           575 => x"71",
           576 => x"52",
           577 => x"08",
           578 => x"80",
           579 => x"16",
           580 => x"81",
           581 => x"0c",
           582 => x"06",
           583 => x"08",
           584 => x"33",
           585 => x"04",
           586 => x"2d",
           587 => x"84",
           588 => x"16",
           589 => x"bb",
           590 => x"a0",
           591 => x"54",
           592 => x"0d",
           593 => x"17",
           594 => x"0d",
           595 => x"70",
           596 => x"38",
           597 => x"54",
           598 => x"54",
           599 => x"84",
           600 => x"0d",
           601 => x"54",
           602 => x"27",
           603 => x"71",
           604 => x"81",
           605 => x"ef",
           606 => x"3d",
           607 => x"27",
           608 => x"ff",
           609 => x"73",
           610 => x"d9",
           611 => x"71",
           612 => x"df",
           613 => x"70",
           614 => x"33",
           615 => x"74",
           616 => x"3d",
           617 => x"71",
           618 => x"54",
           619 => x"54",
           620 => x"84",
           621 => x"0d",
           622 => x"54",
           623 => x"81",
           624 => x"55",
           625 => x"73",
           626 => x"04",
           627 => x"56",
           628 => x"33",
           629 => x"52",
           630 => x"38",
           631 => x"38",
           632 => x"51",
           633 => x"0d",
           634 => x"33",
           635 => x"38",
           636 => x"80",
           637 => x"bb",
           638 => x"84",
           639 => x"fb",
           640 => x"56",
           641 => x"84",
           642 => x"81",
           643 => x"54",
           644 => x"38",
           645 => x"74",
           646 => x"84",
           647 => x"84",
           648 => x"87",
           649 => x"77",
           650 => x"80",
           651 => x"54",
           652 => x"ff",
           653 => x"06",
           654 => x"52",
           655 => x"3d",
           656 => x"79",
           657 => x"2e",
           658 => x"54",
           659 => x"73",
           660 => x"04",
           661 => x"a0",
           662 => x"51",
           663 => x"52",
           664 => x"38",
           665 => x"bb",
           666 => x"9f",
           667 => x"9f",
           668 => x"71",
           669 => x"57",
           670 => x"2e",
           671 => x"07",
           672 => x"ff",
           673 => x"72",
           674 => x"56",
           675 => x"da",
           676 => x"84",
           677 => x"fc",
           678 => x"06",
           679 => x"70",
           680 => x"2a",
           681 => x"70",
           682 => x"74",
           683 => x"30",
           684 => x"31",
           685 => x"05",
           686 => x"25",
           687 => x"70",
           688 => x"70",
           689 => x"05",
           690 => x"55",
           691 => x"55",
           692 => x"56",
           693 => x"3d",
           694 => x"54",
           695 => x"08",
           696 => x"84",
           697 => x"3d",
           698 => x"76",
           699 => x"cf",
           700 => x"13",
           701 => x"51",
           702 => x"08",
           703 => x"80",
           704 => x"be",
           705 => x"72",
           706 => x"55",
           707 => x"72",
           708 => x"77",
           709 => x"2c",
           710 => x"71",
           711 => x"55",
           712 => x"84",
           713 => x"fa",
           714 => x"2c",
           715 => x"2c",
           716 => x"31",
           717 => x"59",
           718 => x"84",
           719 => x"84",
           720 => x"0d",
           721 => x"0c",
           722 => x"73",
           723 => x"81",
           724 => x"55",
           725 => x"2e",
           726 => x"83",
           727 => x"89",
           728 => x"56",
           729 => x"e0",
           730 => x"81",
           731 => x"81",
           732 => x"8f",
           733 => x"54",
           734 => x"72",
           735 => x"29",
           736 => x"33",
           737 => x"be",
           738 => x"30",
           739 => x"84",
           740 => x"81",
           741 => x"56",
           742 => x"06",
           743 => x"0c",
           744 => x"2e",
           745 => x"2e",
           746 => x"c6",
           747 => x"58",
           748 => x"84",
           749 => x"82",
           750 => x"33",
           751 => x"80",
           752 => x"0d",
           753 => x"57",
           754 => x"33",
           755 => x"81",
           756 => x"0c",
           757 => x"f3",
           758 => x"73",
           759 => x"58",
           760 => x"38",
           761 => x"80",
           762 => x"38",
           763 => x"53",
           764 => x"53",
           765 => x"70",
           766 => x"27",
           767 => x"83",
           768 => x"70",
           769 => x"73",
           770 => x"2e",
           771 => x"0c",
           772 => x"8b",
           773 => x"79",
           774 => x"b0",
           775 => x"81",
           776 => x"55",
           777 => x"58",
           778 => x"56",
           779 => x"53",
           780 => x"fe",
           781 => x"8b",
           782 => x"70",
           783 => x"56",
           784 => x"84",
           785 => x"aa",
           786 => x"06",
           787 => x"0d",
           788 => x"71",
           789 => x"71",
           790 => x"be",
           791 => x"bc",
           792 => x"04",
           793 => x"83",
           794 => x"ef",
           795 => x"d0",
           796 => x"0d",
           797 => x"3f",
           798 => x"51",
           799 => x"83",
           800 => x"3d",
           801 => x"e6",
           802 => x"80",
           803 => x"04",
           804 => x"83",
           805 => x"ee",
           806 => x"d1",
           807 => x"0d",
           808 => x"3f",
           809 => x"51",
           810 => x"83",
           811 => x"3d",
           812 => x"8e",
           813 => x"a8",
           814 => x"04",
           815 => x"83",
           816 => x"ed",
           817 => x"d2",
           818 => x"0d",
           819 => x"3d",
           820 => x"33",
           821 => x"08",
           822 => x"51",
           823 => x"ff",
           824 => x"07",
           825 => x"57",
           826 => x"52",
           827 => x"99",
           828 => x"bb",
           829 => x"77",
           830 => x"70",
           831 => x"9f",
           832 => x"77",
           833 => x"88",
           834 => x"e3",
           835 => x"51",
           836 => x"54",
           837 => x"d2",
           838 => x"bb",
           839 => x"84",
           840 => x"0c",
           841 => x"3d",
           842 => x"75",
           843 => x"84",
           844 => x"08",
           845 => x"2e",
           846 => x"57",
           847 => x"51",
           848 => x"52",
           849 => x"84",
           850 => x"52",
           851 => x"ff",
           852 => x"84",
           853 => x"58",
           854 => x"e1",
           855 => x"76",
           856 => x"8a",
           857 => x"3d",
           858 => x"56",
           859 => x"53",
           860 => x"bb",
           861 => x"3d",
           862 => x"63",
           863 => x"73",
           864 => x"5f",
           865 => x"38",
           866 => x"f3",
           867 => x"3f",
           868 => x"7c",
           869 => x"2e",
           870 => x"7a",
           871 => x"83",
           872 => x"14",
           873 => x"51",
           874 => x"38",
           875 => x"80",
           876 => x"75",
           877 => x"72",
           878 => x"53",
           879 => x"74",
           880 => x"57",
           881 => x"74",
           882 => x"08",
           883 => x"16",
           884 => x"d3",
           885 => x"79",
           886 => x"3f",
           887 => x"98",
           888 => x"ee",
           889 => x"7b",
           890 => x"38",
           891 => x"3d",
           892 => x"a3",
           893 => x"53",
           894 => x"74",
           895 => x"83",
           896 => x"14",
           897 => x"51",
           898 => x"c0",
           899 => x"df",
           900 => x"51",
           901 => x"e8",
           902 => x"3f",
           903 => x"39",
           904 => x"84",
           905 => x"a0",
           906 => x"fd",
           907 => x"27",
           908 => x"8c",
           909 => x"e6",
           910 => x"f9",
           911 => x"d8",
           912 => x"51",
           913 => x"91",
           914 => x"84",
           915 => x"72",
           916 => x"72",
           917 => x"e0",
           918 => x"51",
           919 => x"98",
           920 => x"70",
           921 => x"72",
           922 => x"58",
           923 => x"fd",
           924 => x"84",
           925 => x"2c",
           926 => x"32",
           927 => x"07",
           928 => x"53",
           929 => x"b9",
           930 => x"8f",
           931 => x"c0",
           932 => x"81",
           933 => x"51",
           934 => x"3f",
           935 => x"52",
           936 => x"70",
           937 => x"38",
           938 => x"52",
           939 => x"70",
           940 => x"38",
           941 => x"52",
           942 => x"70",
           943 => x"38",
           944 => x"52",
           945 => x"06",
           946 => x"84",
           947 => x"3f",
           948 => x"80",
           949 => x"84",
           950 => x"3f",
           951 => x"80",
           952 => x"81",
           953 => x"cb",
           954 => x"d5",
           955 => x"9b",
           956 => x"06",
           957 => x"38",
           958 => x"83",
           959 => x"51",
           960 => x"81",
           961 => x"f0",
           962 => x"a0",
           963 => x"3f",
           964 => x"2a",
           965 => x"2e",
           966 => x"51",
           967 => x"9b",
           968 => x"72",
           969 => x"71",
           970 => x"39",
           971 => x"e0",
           972 => x"d0",
           973 => x"51",
           974 => x"ff",
           975 => x"83",
           976 => x"51",
           977 => x"81",
           978 => x"b8",
           979 => x"80",
           980 => x"90",
           981 => x"b7",
           982 => x"ff",
           983 => x"2e",
           984 => x"e3",
           985 => x"fc",
           986 => x"f8",
           987 => x"3f",
           988 => x"81",
           989 => x"82",
           990 => x"38",
           991 => x"2e",
           992 => x"79",
           993 => x"5c",
           994 => x"38",
           995 => x"a0",
           996 => x"26",
           997 => x"fc",
           998 => x"3f",
           999 => x"08",
          1000 => x"e8",
          1001 => x"38",
          1002 => x"83",
          1003 => x"06",
          1004 => x"9a",
          1005 => x"dd",
          1006 => x"87",
          1007 => x"bb",
          1008 => x"84",
          1009 => x"80",
          1010 => x"84",
          1011 => x"80",
          1012 => x"08",
          1013 => x"08",
          1014 => x"a5",
          1015 => x"8a",
          1016 => x"7a",
          1017 => x"80",
          1018 => x"d5",
          1019 => x"bb",
          1020 => x"54",
          1021 => x"52",
          1022 => x"84",
          1023 => x"30",
          1024 => x"5b",
          1025 => x"38",
          1026 => x"80",
          1027 => x"ff",
          1028 => x"7f",
          1029 => x"7c",
          1030 => x"ec",
          1031 => x"83",
          1032 => x"48",
          1033 => x"e8",
          1034 => x"33",
          1035 => x"fd",
          1036 => x"52",
          1037 => x"3f",
          1038 => x"81",
          1039 => x"84",
          1040 => x"51",
          1041 => x"08",
          1042 => x"08",
          1043 => x"ef",
          1044 => x"59",
          1045 => x"d3",
          1046 => x"82",
          1047 => x"83",
          1048 => x"b8",
          1049 => x"51",
          1050 => x"79",
          1051 => x"63",
          1052 => x"89",
          1053 => x"83",
          1054 => x"83",
          1055 => x"e4",
          1056 => x"c8",
          1057 => x"bb",
          1058 => x"fb",
          1059 => x"41",
          1060 => x"51",
          1061 => x"ac",
          1062 => x"56",
          1063 => x"53",
          1064 => x"e3",
          1065 => x"3f",
          1066 => x"f5",
          1067 => x"dc",
          1068 => x"3f",
          1069 => x"de",
          1070 => x"d7",
          1071 => x"3f",
          1072 => x"11",
          1073 => x"3f",
          1074 => x"b5",
          1075 => x"d0",
          1076 => x"bb",
          1077 => x"84",
          1078 => x"51",
          1079 => x"3d",
          1080 => x"51",
          1081 => x"80",
          1082 => x"d8",
          1083 => x"78",
          1084 => x"ff",
          1085 => x"bb",
          1086 => x"b8",
          1087 => x"05",
          1088 => x"08",
          1089 => x"53",
          1090 => x"f3",
          1091 => x"f8",
          1092 => x"48",
          1093 => x"9d",
          1094 => x"64",
          1095 => x"b8",
          1096 => x"05",
          1097 => x"08",
          1098 => x"fe",
          1099 => x"e8",
          1100 => x"b0",
          1101 => x"52",
          1102 => x"84",
          1103 => x"7e",
          1104 => x"33",
          1105 => x"78",
          1106 => x"05",
          1107 => x"ff",
          1108 => x"e9",
          1109 => x"2e",
          1110 => x"11",
          1111 => x"3f",
          1112 => x"85",
          1113 => x"ff",
          1114 => x"bb",
          1115 => x"83",
          1116 => x"67",
          1117 => x"38",
          1118 => x"5a",
          1119 => x"79",
          1120 => x"d8",
          1121 => x"5b",
          1122 => x"d2",
          1123 => x"ff",
          1124 => x"bb",
          1125 => x"b8",
          1126 => x"05",
          1127 => x"08",
          1128 => x"fe",
          1129 => x"e8",
          1130 => x"2e",
          1131 => x"cd",
          1132 => x"82",
          1133 => x"05",
          1134 => x"46",
          1135 => x"53",
          1136 => x"84",
          1137 => x"38",
          1138 => x"80",
          1139 => x"84",
          1140 => x"52",
          1141 => x"84",
          1142 => x"7e",
          1143 => x"33",
          1144 => x"78",
          1145 => x"05",
          1146 => x"db",
          1147 => x"49",
          1148 => x"80",
          1149 => x"84",
          1150 => x"59",
          1151 => x"68",
          1152 => x"11",
          1153 => x"3f",
          1154 => x"f5",
          1155 => x"53",
          1156 => x"84",
          1157 => x"38",
          1158 => x"80",
          1159 => x"84",
          1160 => x"3d",
          1161 => x"51",
          1162 => x"86",
          1163 => x"d9",
          1164 => x"5b",
          1165 => x"5b",
          1166 => x"79",
          1167 => x"e1",
          1168 => x"80",
          1169 => x"84",
          1170 => x"59",
          1171 => x"84",
          1172 => x"84",
          1173 => x"38",
          1174 => x"3f",
          1175 => x"11",
          1176 => x"3f",
          1177 => x"f4",
          1178 => x"c0",
          1179 => x"3d",
          1180 => x"51",
          1181 => x"91",
          1182 => x"80",
          1183 => x"08",
          1184 => x"ff",
          1185 => x"bb",
          1186 => x"66",
          1187 => x"81",
          1188 => x"72",
          1189 => x"5d",
          1190 => x"2e",
          1191 => x"51",
          1192 => x"65",
          1193 => x"3f",
          1194 => x"f2",
          1195 => x"64",
          1196 => x"11",
          1197 => x"3f",
          1198 => x"d5",
          1199 => x"84",
          1200 => x"53",
          1201 => x"84",
          1202 => x"39",
          1203 => x"7e",
          1204 => x"b8",
          1205 => x"05",
          1206 => x"08",
          1207 => x"02",
          1208 => x"05",
          1209 => x"f0",
          1210 => x"ad",
          1211 => x"38",
          1212 => x"11",
          1213 => x"3f",
          1214 => x"dc",
          1215 => x"33",
          1216 => x"9b",
          1217 => x"ff",
          1218 => x"bb",
          1219 => x"64",
          1220 => x"70",
          1221 => x"2e",
          1222 => x"55",
          1223 => x"d9",
          1224 => x"f3",
          1225 => x"fa",
          1226 => x"51",
          1227 => x"3d",
          1228 => x"51",
          1229 => x"80",
          1230 => x"ce",
          1231 => x"23",
          1232 => x"89",
          1233 => x"38",
          1234 => x"39",
          1235 => x"2e",
          1236 => x"fc",
          1237 => x"c6",
          1238 => x"d9",
          1239 => x"f6",
          1240 => x"78",
          1241 => x"08",
          1242 => x"51",
          1243 => x"f4",
          1244 => x"38",
          1245 => x"39",
          1246 => x"2e",
          1247 => x"fb",
          1248 => x"7d",
          1249 => x"08",
          1250 => x"33",
          1251 => x"f3",
          1252 => x"f4",
          1253 => x"38",
          1254 => x"39",
          1255 => x"49",
          1256 => x"88",
          1257 => x"0d",
          1258 => x"c0",
          1259 => x"84",
          1260 => x"84",
          1261 => x"57",
          1262 => x"da",
          1263 => x"07",
          1264 => x"08",
          1265 => x"51",
          1266 => x"90",
          1267 => x"80",
          1268 => x"84",
          1269 => x"80",
          1270 => x"8c",
          1271 => x"0c",
          1272 => x"5d",
          1273 => x"80",
          1274 => x"70",
          1275 => x"e6",
          1276 => x"9e",
          1277 => x"95",
          1278 => x"d3",
          1279 => x"f4",
          1280 => x"83",
          1281 => x"81",
          1282 => x"c3",
          1283 => x"fc",
          1284 => x"d4",
          1285 => x"0a",
          1286 => x"3f",
          1287 => x"0d",
          1288 => x"52",
          1289 => x"74",
          1290 => x"70",
          1291 => x"81",
          1292 => x"53",
          1293 => x"71",
          1294 => x"81",
          1295 => x"80",
          1296 => x"ff",
          1297 => x"83",
          1298 => x"38",
          1299 => x"52",
          1300 => x"52",
          1301 => x"83",
          1302 => x"30",
          1303 => x"53",
          1304 => x"70",
          1305 => x"74",
          1306 => x"3d",
          1307 => x"73",
          1308 => x"52",
          1309 => x"53",
          1310 => x"81",
          1311 => x"75",
          1312 => x"06",
          1313 => x"0d",
          1314 => x"0b",
          1315 => x"04",
          1316 => x"da",
          1317 => x"2e",
          1318 => x"86",
          1319 => x"82",
          1320 => x"52",
          1321 => x"13",
          1322 => x"9e",
          1323 => x"51",
          1324 => x"38",
          1325 => x"bb",
          1326 => x"55",
          1327 => x"38",
          1328 => x"87",
          1329 => x"22",
          1330 => x"80",
          1331 => x"9c",
          1332 => x"0c",
          1333 => x"0c",
          1334 => x"0c",
          1335 => x"0c",
          1336 => x"0c",
          1337 => x"0c",
          1338 => x"87",
          1339 => x"c0",
          1340 => x"bb",
          1341 => x"3d",
          1342 => x"5d",
          1343 => x"08",
          1344 => x"b8",
          1345 => x"c0",
          1346 => x"34",
          1347 => x"84",
          1348 => x"5a",
          1349 => x"a8",
          1350 => x"c0",
          1351 => x"23",
          1352 => x"8a",
          1353 => x"ff",
          1354 => x"06",
          1355 => x"33",
          1356 => x"33",
          1357 => x"ff",
          1358 => x"ff",
          1359 => x"fe",
          1360 => x"72",
          1361 => x"e9",
          1362 => x"2b",
          1363 => x"2e",
          1364 => x"2e",
          1365 => x"84",
          1366 => x"b7",
          1367 => x"70",
          1368 => x"09",
          1369 => x"e9",
          1370 => x"2b",
          1371 => x"2e",
          1372 => x"80",
          1373 => x"81",
          1374 => x"84",
          1375 => x"52",
          1376 => x"07",
          1377 => x"db",
          1378 => x"3d",
          1379 => x"05",
          1380 => x"ff",
          1381 => x"80",
          1382 => x"70",
          1383 => x"52",
          1384 => x"2a",
          1385 => x"38",
          1386 => x"80",
          1387 => x"06",
          1388 => x"06",
          1389 => x"80",
          1390 => x"52",
          1391 => x"0c",
          1392 => x"70",
          1393 => x"72",
          1394 => x"2e",
          1395 => x"52",
          1396 => x"94",
          1397 => x"06",
          1398 => x"39",
          1399 => x"70",
          1400 => x"70",
          1401 => x"04",
          1402 => x"33",
          1403 => x"80",
          1404 => x"33",
          1405 => x"71",
          1406 => x"94",
          1407 => x"06",
          1408 => x"38",
          1409 => x"51",
          1410 => x"06",
          1411 => x"93",
          1412 => x"75",
          1413 => x"80",
          1414 => x"c0",
          1415 => x"17",
          1416 => x"38",
          1417 => x"0d",
          1418 => x"51",
          1419 => x"81",
          1420 => x"71",
          1421 => x"2e",
          1422 => x"08",
          1423 => x"54",
          1424 => x"3d",
          1425 => x"9c",
          1426 => x"2e",
          1427 => x"08",
          1428 => x"a8",
          1429 => x"9e",
          1430 => x"c0",
          1431 => x"87",
          1432 => x"0c",
          1433 => x"d4",
          1434 => x"f3",
          1435 => x"83",
          1436 => x"08",
          1437 => x"b8",
          1438 => x"9e",
          1439 => x"c0",
          1440 => x"87",
          1441 => x"0c",
          1442 => x"83",
          1443 => x"08",
          1444 => x"88",
          1445 => x"9e",
          1446 => x"0b",
          1447 => x"c0",
          1448 => x"06",
          1449 => x"71",
          1450 => x"c0",
          1451 => x"06",
          1452 => x"38",
          1453 => x"80",
          1454 => x"90",
          1455 => x"80",
          1456 => x"f4",
          1457 => x"90",
          1458 => x"52",
          1459 => x"52",
          1460 => x"87",
          1461 => x"80",
          1462 => x"83",
          1463 => x"34",
          1464 => x"70",
          1465 => x"70",
          1466 => x"83",
          1467 => x"9e",
          1468 => x"51",
          1469 => x"81",
          1470 => x"0b",
          1471 => x"80",
          1472 => x"2e",
          1473 => x"8c",
          1474 => x"08",
          1475 => x"52",
          1476 => x"71",
          1477 => x"c0",
          1478 => x"06",
          1479 => x"38",
          1480 => x"80",
          1481 => x"a0",
          1482 => x"2e",
          1483 => x"8f",
          1484 => x"80",
          1485 => x"83",
          1486 => x"9e",
          1487 => x"52",
          1488 => x"52",
          1489 => x"9e",
          1490 => x"2a",
          1491 => x"80",
          1492 => x"88",
          1493 => x"83",
          1494 => x"34",
          1495 => x"51",
          1496 => x"0d",
          1497 => x"3d",
          1498 => x"b3",
          1499 => x"86",
          1500 => x"8e",
          1501 => x"85",
          1502 => x"73",
          1503 => x"56",
          1504 => x"33",
          1505 => x"8a",
          1506 => x"f4",
          1507 => x"83",
          1508 => x"38",
          1509 => x"e3",
          1510 => x"83",
          1511 => x"73",
          1512 => x"55",
          1513 => x"33",
          1514 => x"8e",
          1515 => x"da",
          1516 => x"e8",
          1517 => x"b5",
          1518 => x"83",
          1519 => x"83",
          1520 => x"51",
          1521 => x"51",
          1522 => x"52",
          1523 => x"3f",
          1524 => x"c0",
          1525 => x"bb",
          1526 => x"71",
          1527 => x"52",
          1528 => x"3f",
          1529 => x"38",
          1530 => x"38",
          1531 => x"08",
          1532 => x"c9",
          1533 => x"84",
          1534 => x"84",
          1535 => x"51",
          1536 => x"04",
          1537 => x"c0",
          1538 => x"bb",
          1539 => x"71",
          1540 => x"52",
          1541 => x"3f",
          1542 => x"2e",
          1543 => x"dc",
          1544 => x"c0",
          1545 => x"08",
          1546 => x"b3",
          1547 => x"da",
          1548 => x"f3",
          1549 => x"ff",
          1550 => x"ff",
          1551 => x"52",
          1552 => x"3f",
          1553 => x"c0",
          1554 => x"bb",
          1555 => x"71",
          1556 => x"52",
          1557 => x"3f",
          1558 => x"2e",
          1559 => x"dd",
          1560 => x"f4",
          1561 => x"8e",
          1562 => x"51",
          1563 => x"33",
          1564 => x"d6",
          1565 => x"86",
          1566 => x"80",
          1567 => x"dd",
          1568 => x"f4",
          1569 => x"b3",
          1570 => x"52",
          1571 => x"3f",
          1572 => x"2e",
          1573 => x"94",
          1574 => x"b1",
          1575 => x"74",
          1576 => x"83",
          1577 => x"51",
          1578 => x"33",
          1579 => x"cd",
          1580 => x"d4",
          1581 => x"51",
          1582 => x"33",
          1583 => x"c7",
          1584 => x"cc",
          1585 => x"51",
          1586 => x"33",
          1587 => x"c1",
          1588 => x"c4",
          1589 => x"51",
          1590 => x"33",
          1591 => x"c1",
          1592 => x"dc",
          1593 => x"51",
          1594 => x"33",
          1595 => x"c1",
          1596 => x"e4",
          1597 => x"51",
          1598 => x"33",
          1599 => x"c1",
          1600 => x"83",
          1601 => x"e6",
          1602 => x"80",
          1603 => x"3d",
          1604 => x"85",
          1605 => x"c4",
          1606 => x"df",
          1607 => x"3d",
          1608 => x"af",
          1609 => x"df",
          1610 => x"3d",
          1611 => x"af",
          1612 => x"df",
          1613 => x"3d",
          1614 => x"af",
          1615 => x"88",
          1616 => x"96",
          1617 => x"87",
          1618 => x"0d",
          1619 => x"5a",
          1620 => x"f4",
          1621 => x"84",
          1622 => x"3d",
          1623 => x"54",
          1624 => x"d3",
          1625 => x"2e",
          1626 => x"84",
          1627 => x"80",
          1628 => x"38",
          1629 => x"18",
          1630 => x"70",
          1631 => x"55",
          1632 => x"ff",
          1633 => x"11",
          1634 => x"84",
          1635 => x"2e",
          1636 => x"a9",
          1637 => x"ff",
          1638 => x"81",
          1639 => x"c0",
          1640 => x"3f",
          1641 => x"08",
          1642 => x"51",
          1643 => x"bb",
          1644 => x"3d",
          1645 => x"71",
          1646 => x"57",
          1647 => x"0b",
          1648 => x"10",
          1649 => x"54",
          1650 => x"08",
          1651 => x"bf",
          1652 => x"38",
          1653 => x"81",
          1654 => x"81",
          1655 => x"82",
          1656 => x"84",
          1657 => x"81",
          1658 => x"53",
          1659 => x"84",
          1660 => x"ff",
          1661 => x"a5",
          1662 => x"06",
          1663 => x"16",
          1664 => x"76",
          1665 => x"78",
          1666 => x"fe",
          1667 => x"33",
          1668 => x"06",
          1669 => x"38",
          1670 => x"cc",
          1671 => x"83",
          1672 => x"e1",
          1673 => x"38",
          1674 => x"52",
          1675 => x"bb",
          1676 => x"51",
          1677 => x"08",
          1678 => x"25",
          1679 => x"05",
          1680 => x"77",
          1681 => x"ac",
          1682 => x"ff",
          1683 => x"81",
          1684 => x"0d",
          1685 => x"b8",
          1686 => x"08",
          1687 => x"5c",
          1688 => x"f4",
          1689 => x"83",
          1690 => x"74",
          1691 => x"80",
          1692 => x"91",
          1693 => x"56",
          1694 => x"90",
          1695 => x"40",
          1696 => x"84",
          1697 => x"57",
          1698 => x"81",
          1699 => x"98",
          1700 => x"33",
          1701 => x"98",
          1702 => x"e0",
          1703 => x"53",
          1704 => x"59",
          1705 => x"38",
          1706 => x"81",
          1707 => x"70",
          1708 => x"81",
          1709 => x"2b",
          1710 => x"16",
          1711 => x"38",
          1712 => x"33",
          1713 => x"38",
          1714 => x"e2",
          1715 => x"81",
          1716 => x"70",
          1717 => x"98",
          1718 => x"05",
          1719 => x"33",
          1720 => x"57",
          1721 => x"84",
          1722 => x"3f",
          1723 => x"98",
          1724 => x"81",
          1725 => x"fe",
          1726 => x"81",
          1727 => x"80",
          1728 => x"98",
          1729 => x"42",
          1730 => x"10",
          1731 => x"0b",
          1732 => x"77",
          1733 => x"15",
          1734 => x"62",
          1735 => x"ff",
          1736 => x"76",
          1737 => x"39",
          1738 => x"76",
          1739 => x"34",
          1740 => x"34",
          1741 => x"26",
          1742 => x"c4",
          1743 => x"df",
          1744 => x"84",
          1745 => x"bc",
          1746 => x"56",
          1747 => x"e6",
          1748 => x"c9",
          1749 => x"5b",
          1750 => x"39",
          1751 => x"06",
          1752 => x"75",
          1753 => x"e8",
          1754 => x"e2",
          1755 => x"55",
          1756 => x"7c",
          1757 => x"26",
          1758 => x"a0",
          1759 => x"a5",
          1760 => x"80",
          1761 => x"e2",
          1762 => x"b6",
          1763 => x"51",
          1764 => x"08",
          1765 => x"84",
          1766 => x"b4",
          1767 => x"05",
          1768 => x"81",
          1769 => x"51",
          1770 => x"c8",
          1771 => x"83",
          1772 => x"38",
          1773 => x"58",
          1774 => x"10",
          1775 => x"55",
          1776 => x"fa",
          1777 => x"9c",
          1778 => x"2e",
          1779 => x"8b",
          1780 => x"c4",
          1781 => x"06",
          1782 => x"ff",
          1783 => x"84",
          1784 => x"2e",
          1785 => x"52",
          1786 => x"e6",
          1787 => x"91",
          1788 => x"51",
          1789 => x"33",
          1790 => x"34",
          1791 => x"84",
          1792 => x"84",
          1793 => x"7a",
          1794 => x"08",
          1795 => x"c8",
          1796 => x"ff",
          1797 => x"70",
          1798 => x"5a",
          1799 => x"38",
          1800 => x"57",
          1801 => x"70",
          1802 => x"84",
          1803 => x"84",
          1804 => x"76",
          1805 => x"84",
          1806 => x"56",
          1807 => x"ff",
          1808 => x"75",
          1809 => x"ff",
          1810 => x"80",
          1811 => x"a0",
          1812 => x"c8",
          1813 => x"84",
          1814 => x"74",
          1815 => x"e8",
          1816 => x"3f",
          1817 => x"0a",
          1818 => x"33",
          1819 => x"a0",
          1820 => x"51",
          1821 => x"0a",
          1822 => x"2c",
          1823 => x"7a",
          1824 => x"39",
          1825 => x"34",
          1826 => x"51",
          1827 => x"0a",
          1828 => x"2c",
          1829 => x"75",
          1830 => x"58",
          1831 => x"e8",
          1832 => x"a9",
          1833 => x"80",
          1834 => x"c4",
          1835 => x"ff",
          1836 => x"c8",
          1837 => x"38",
          1838 => x"ff",
          1839 => x"ff",
          1840 => x"76",
          1841 => x"e2",
          1842 => x"34",
          1843 => x"ff",
          1844 => x"7b",
          1845 => x"08",
          1846 => x"38",
          1847 => x"2e",
          1848 => x"70",
          1849 => x"08",
          1850 => x"75",
          1851 => x"9c",
          1852 => x"80",
          1853 => x"79",
          1854 => x"10",
          1855 => x"43",
          1856 => x"83",
          1857 => x"10",
          1858 => x"5e",
          1859 => x"ec",
          1860 => x"83",
          1861 => x"8b",
          1862 => x"34",
          1863 => x"84",
          1864 => x"84",
          1865 => x"b6",
          1866 => x"51",
          1867 => x"08",
          1868 => x"84",
          1869 => x"ae",
          1870 => x"05",
          1871 => x"81",
          1872 => x"d3",
          1873 => x"0b",
          1874 => x"e2",
          1875 => x"c8",
          1876 => x"7a",
          1877 => x"c4",
          1878 => x"c4",
          1879 => x"c8",
          1880 => x"51",
          1881 => x"33",
          1882 => x"e2",
          1883 => x"76",
          1884 => x"08",
          1885 => x"84",
          1886 => x"98",
          1887 => x"59",
          1888 => x"84",
          1889 => x"ac",
          1890 => x"81",
          1891 => x"e2",
          1892 => x"24",
          1893 => x"52",
          1894 => x"81",
          1895 => x"70",
          1896 => x"51",
          1897 => x"f3",
          1898 => x"33",
          1899 => x"76",
          1900 => x"81",
          1901 => x"70",
          1902 => x"57",
          1903 => x"7b",
          1904 => x"84",
          1905 => x"ff",
          1906 => x"29",
          1907 => x"84",
          1908 => x"76",
          1909 => x"83",
          1910 => x"84",
          1911 => x"b6",
          1912 => x"51",
          1913 => x"08",
          1914 => x"84",
          1915 => x"ab",
          1916 => x"05",
          1917 => x"81",
          1918 => x"d3",
          1919 => x"0b",
          1920 => x"e2",
          1921 => x"b5",
          1922 => x"70",
          1923 => x"2e",
          1924 => x"55",
          1925 => x"2b",
          1926 => x"24",
          1927 => x"81",
          1928 => x"81",
          1929 => x"e2",
          1930 => x"25",
          1931 => x"e2",
          1932 => x"05",
          1933 => x"e2",
          1934 => x"38",
          1935 => x"34",
          1936 => x"81",
          1937 => x"70",
          1938 => x"58",
          1939 => x"38",
          1940 => x"81",
          1941 => x"25",
          1942 => x"52",
          1943 => x"81",
          1944 => x"70",
          1945 => x"57",
          1946 => x"84",
          1947 => x"a9",
          1948 => x"81",
          1949 => x"e2",
          1950 => x"24",
          1951 => x"a8",
          1952 => x"84",
          1953 => x"84",
          1954 => x"99",
          1955 => x"74",
          1956 => x"34",
          1957 => x"84",
          1958 => x"33",
          1959 => x"81",
          1960 => x"70",
          1961 => x"57",
          1962 => x"e2",
          1963 => x"2c",
          1964 => x"58",
          1965 => x"c3",
          1966 => x"ef",
          1967 => x"56",
          1968 => x"16",
          1969 => x"f0",
          1970 => x"83",
          1971 => x"ee",
          1972 => x"3f",
          1973 => x"ac",
          1974 => x"94",
          1975 => x"39",
          1976 => x"77",
          1977 => x"75",
          1978 => x"39",
          1979 => x"bb",
          1980 => x"bb",
          1981 => x"53",
          1982 => x"3f",
          1983 => x"e2",
          1984 => x"2e",
          1985 => x"52",
          1986 => x"e6",
          1987 => x"d1",
          1988 => x"51",
          1989 => x"33",
          1990 => x"34",
          1991 => x"75",
          1992 => x"84",
          1993 => x"84",
          1994 => x"75",
          1995 => x"76",
          1996 => x"33",
          1997 => x"de",
          1998 => x"51",
          1999 => x"08",
          2000 => x"84",
          2001 => x"a5",
          2002 => x"05",
          2003 => x"81",
          2004 => x"ff",
          2005 => x"84",
          2006 => x"81",
          2007 => x"7b",
          2008 => x"70",
          2009 => x"84",
          2010 => x"74",
          2011 => x"e8",
          2012 => x"3f",
          2013 => x"ff",
          2014 => x"52",
          2015 => x"e2",
          2016 => x"e2",
          2017 => x"c7",
          2018 => x"e2",
          2019 => x"34",
          2020 => x"0d",
          2021 => x"80",
          2022 => x"a7",
          2023 => x"e2",
          2024 => x"ff",
          2025 => x"51",
          2026 => x"33",
          2027 => x"80",
          2028 => x"08",
          2029 => x"84",
          2030 => x"a3",
          2031 => x"88",
          2032 => x"c8",
          2033 => x"c8",
          2034 => x"39",
          2035 => x"f4",
          2036 => x"06",
          2037 => x"54",
          2038 => x"84",
          2039 => x"f4",
          2040 => x"05",
          2041 => x"52",
          2042 => x"f4",
          2043 => x"05",
          2044 => x"2e",
          2045 => x"74",
          2046 => x"f4",
          2047 => x"56",
          2048 => x"77",
          2049 => x"b5",
          2050 => x"7b",
          2051 => x"83",
          2052 => x"b9",
          2053 => x"81",
          2054 => x"c8",
          2055 => x"7b",
          2056 => x"04",
          2057 => x"ca",
          2058 => x"d5",
          2059 => x"5c",
          2060 => x"f8",
          2061 => x"84",
          2062 => x"08",
          2063 => x"38",
          2064 => x"a3",
          2065 => x"0b",
          2066 => x"38",
          2067 => x"1b",
          2068 => x"ff",
          2069 => x"10",
          2070 => x"41",
          2071 => x"82",
          2072 => x"05",
          2073 => x"da",
          2074 => x"0c",
          2075 => x"83",
          2076 => x"83",
          2077 => x"3f",
          2078 => x"83",
          2079 => x"42",
          2080 => x"ff",
          2081 => x"38",
          2082 => x"06",
          2083 => x"f8",
          2084 => x"51",
          2085 => x"33",
          2086 => x"56",
          2087 => x"0b",
          2088 => x"74",
          2089 => x"f4",
          2090 => x"83",
          2091 => x"52",
          2092 => x"bb",
          2093 => x"33",
          2094 => x"70",
          2095 => x"59",
          2096 => x"33",
          2097 => x"70",
          2098 => x"fe",
          2099 => x"f4",
          2100 => x"f4",
          2101 => x"d4",
          2102 => x"c2",
          2103 => x"02",
          2104 => x"80",
          2105 => x"26",
          2106 => x"8b",
          2107 => x"72",
          2108 => x"a0",
          2109 => x"5e",
          2110 => x"76",
          2111 => x"34",
          2112 => x"fa",
          2113 => x"98",
          2114 => x"2b",
          2115 => x"56",
          2116 => x"74",
          2117 => x"70",
          2118 => x"ee",
          2119 => x"fa",
          2120 => x"78",
          2121 => x"e0",
          2122 => x"56",
          2123 => x"90",
          2124 => x"0b",
          2125 => x"11",
          2126 => x"11",
          2127 => x"86",
          2128 => x"33",
          2129 => x"33",
          2130 => x"22",
          2131 => x"29",
          2132 => x"5d",
          2133 => x"31",
          2134 => x"7e",
          2135 => x"7a",
          2136 => x"06",
          2137 => x"57",
          2138 => x"83",
          2139 => x"70",
          2140 => x"06",
          2141 => x"78",
          2142 => x"c1",
          2143 => x"34",
          2144 => x"05",
          2145 => x"80",
          2146 => x"b8",
          2147 => x"b8",
          2148 => x"fa",
          2149 => x"5d",
          2150 => x"27",
          2151 => x"73",
          2152 => x"5a",
          2153 => x"38",
          2154 => x"0b",
          2155 => x"33",
          2156 => x"71",
          2157 => x"56",
          2158 => x"ae",
          2159 => x"38",
          2160 => x"06",
          2161 => x"33",
          2162 => x"80",
          2163 => x"86",
          2164 => x"f8",
          2165 => x"f7",
          2166 => x"b2",
          2167 => x"75",
          2168 => x"58",
          2169 => x"8b",
          2170 => x"29",
          2171 => x"74",
          2172 => x"83",
          2173 => x"70",
          2174 => x"55",
          2175 => x"29",
          2176 => x"06",
          2177 => x"83",
          2178 => x"f2",
          2179 => x"fe",
          2180 => x"80",
          2181 => x"73",
          2182 => x"87",
          2183 => x"34",
          2184 => x"98",
          2185 => x"87",
          2186 => x"80",
          2187 => x"52",
          2188 => x"87",
          2189 => x"56",
          2190 => x"84",
          2191 => x"08",
          2192 => x"51",
          2193 => x"cc",
          2194 => x"53",
          2195 => x"08",
          2196 => x"75",
          2197 => x"34",
          2198 => x"3d",
          2199 => x"bb",
          2200 => x"af",
          2201 => x"33",
          2202 => x"81",
          2203 => x"84",
          2204 => x"83",
          2205 => x"86",
          2206 => x"22",
          2207 => x"05",
          2208 => x"8a",
          2209 => x"2e",
          2210 => x"76",
          2211 => x"83",
          2212 => x"ff",
          2213 => x"55",
          2214 => x"19",
          2215 => x"fa",
          2216 => x"84",
          2217 => x"74",
          2218 => x"33",
          2219 => x"72",
          2220 => x"d6",
          2221 => x"33",
          2222 => x"05",
          2223 => x"34",
          2224 => x"27",
          2225 => x"38",
          2226 => x"15",
          2227 => x"34",
          2228 => x"81",
          2229 => x"38",
          2230 => x"75",
          2231 => x"81",
          2232 => x"54",
          2233 => x"72",
          2234 => x"33",
          2235 => x"55",
          2236 => x"b0",
          2237 => x"ff",
          2238 => x"54",
          2239 => x"99",
          2240 => x"53",
          2241 => x"81",
          2242 => x"55",
          2243 => x"81",
          2244 => x"f7",
          2245 => x"5a",
          2246 => x"53",
          2247 => x"0d",
          2248 => x"fa",
          2249 => x"84",
          2250 => x"7a",
          2251 => x"fe",
          2252 => x"05",
          2253 => x"75",
          2254 => x"73",
          2255 => x"33",
          2256 => x"56",
          2257 => x"ae",
          2258 => x"d6",
          2259 => x"a0",
          2260 => x"70",
          2261 => x"72",
          2262 => x"e0",
          2263 => x"05",
          2264 => x"38",
          2265 => x"f8",
          2266 => x"fa",
          2267 => x"19",
          2268 => x"59",
          2269 => x"02",
          2270 => x"70",
          2271 => x"83",
          2272 => x"84",
          2273 => x"86",
          2274 => x"0b",
          2275 => x"04",
          2276 => x"fa",
          2277 => x"52",
          2278 => x"51",
          2279 => x"84",
          2280 => x"83",
          2281 => x"09",
          2282 => x"53",
          2283 => x"39",
          2284 => x"b8",
          2285 => x"70",
          2286 => x"83",
          2287 => x"84",
          2288 => x"b5",
          2289 => x"9f",
          2290 => x"70",
          2291 => x"bb",
          2292 => x"fa",
          2293 => x"33",
          2294 => x"25",
          2295 => x"b5",
          2296 => x"86",
          2297 => x"b5",
          2298 => x"f7",
          2299 => x"25",
          2300 => x"83",
          2301 => x"3d",
          2302 => x"b1",
          2303 => x"c5",
          2304 => x"fa",
          2305 => x"84",
          2306 => x"2a",
          2307 => x"f0",
          2308 => x"f2",
          2309 => x"84",
          2310 => x"83",
          2311 => x"07",
          2312 => x"0b",
          2313 => x"04",
          2314 => x"51",
          2315 => x"83",
          2316 => x"07",
          2317 => x"39",
          2318 => x"80",
          2319 => x"0d",
          2320 => x"06",
          2321 => x"34",
          2322 => x"87",
          2323 => x"ff",
          2324 => x"fd",
          2325 => x"b0",
          2326 => x"33",
          2327 => x"83",
          2328 => x"fa",
          2329 => x"51",
          2330 => x"39",
          2331 => x"51",
          2332 => x"39",
          2333 => x"80",
          2334 => x"34",
          2335 => x"81",
          2336 => x"fa",
          2337 => x"b0",
          2338 => x"51",
          2339 => x"39",
          2340 => x"80",
          2341 => x"34",
          2342 => x"81",
          2343 => x"fa",
          2344 => x"b0",
          2345 => x"fa",
          2346 => x"b0",
          2347 => x"70",
          2348 => x"f3",
          2349 => x"84",
          2350 => x"b4",
          2351 => x"b5",
          2352 => x"5f",
          2353 => x"a1",
          2354 => x"81",
          2355 => x"fa",
          2356 => x"7a",
          2357 => x"b2",
          2358 => x"3d",
          2359 => x"06",
          2360 => x"34",
          2361 => x"0b",
          2362 => x"fa",
          2363 => x"23",
          2364 => x"84",
          2365 => x"33",
          2366 => x"83",
          2367 => x"7d",
          2368 => x"b8",
          2369 => x"7b",
          2370 => x"b5",
          2371 => x"84",
          2372 => x"fc",
          2373 => x"a8",
          2374 => x"83",
          2375 => x"58",
          2376 => x"85",
          2377 => x"53",
          2378 => x"ff",
          2379 => x"33",
          2380 => x"79",
          2381 => x"53",
          2382 => x"93",
          2383 => x"84",
          2384 => x"7a",
          2385 => x"fe",
          2386 => x"34",
          2387 => x"83",
          2388 => x"23",
          2389 => x"0d",
          2390 => x"81",
          2391 => x"83",
          2392 => x"b5",
          2393 => x"83",
          2394 => x"84",
          2395 => x"51",
          2396 => x"f8",
          2397 => x"84",
          2398 => x"83",
          2399 => x"b8",
          2400 => x"70",
          2401 => x"f9",
          2402 => x"05",
          2403 => x"b5",
          2404 => x"29",
          2405 => x"fa",
          2406 => x"7c",
          2407 => x"83",
          2408 => x"57",
          2409 => x"75",
          2410 => x"24",
          2411 => x"85",
          2412 => x"84",
          2413 => x"83",
          2414 => x"55",
          2415 => x"86",
          2416 => x"f8",
          2417 => x"b2",
          2418 => x"56",
          2419 => x"83",
          2420 => x"58",
          2421 => x"b0",
          2422 => x"70",
          2423 => x"83",
          2424 => x"57",
          2425 => x"33",
          2426 => x"70",
          2427 => x"26",
          2428 => x"58",
          2429 => x"72",
          2430 => x"33",
          2431 => x"b8",
          2432 => x"fb",
          2433 => x"89",
          2434 => x"38",
          2435 => x"8a",
          2436 => x"81",
          2437 => x"0b",
          2438 => x"83",
          2439 => x"80",
          2440 => x"09",
          2441 => x"76",
          2442 => x"13",
          2443 => x"83",
          2444 => x"51",
          2445 => x"ff",
          2446 => x"38",
          2447 => x"34",
          2448 => x"f9",
          2449 => x"0c",
          2450 => x"2e",
          2451 => x"fa",
          2452 => x"ff",
          2453 => x"72",
          2454 => x"51",
          2455 => x"70",
          2456 => x"73",
          2457 => x"fa",
          2458 => x"83",
          2459 => x"ef",
          2460 => x"75",
          2461 => x"e6",
          2462 => x"84",
          2463 => x"2e",
          2464 => x"82",
          2465 => x"78",
          2466 => x"2e",
          2467 => x"8f",
          2468 => x"b4",
          2469 => x"29",
          2470 => x"19",
          2471 => x"84",
          2472 => x"83",
          2473 => x"5a",
          2474 => x"18",
          2475 => x"29",
          2476 => x"33",
          2477 => x"84",
          2478 => x"83",
          2479 => x"72",
          2480 => x"59",
          2481 => x"1f",
          2482 => x"42",
          2483 => x"84",
          2484 => x"38",
          2485 => x"34",
          2486 => x"3d",
          2487 => x"38",
          2488 => x"b8",
          2489 => x"2e",
          2490 => x"80",
          2491 => x"b4",
          2492 => x"29",
          2493 => x"19",
          2494 => x"84",
          2495 => x"83",
          2496 => x"41",
          2497 => x"1f",
          2498 => x"29",
          2499 => x"86",
          2500 => x"f8",
          2501 => x"b2",
          2502 => x"29",
          2503 => x"fa",
          2504 => x"34",
          2505 => x"41",
          2506 => x"83",
          2507 => x"84",
          2508 => x"2e",
          2509 => x"81",
          2510 => x"fd",
          2511 => x"34",
          2512 => x"3d",
          2513 => x"38",
          2514 => x"d0",
          2515 => x"59",
          2516 => x"84",
          2517 => x"06",
          2518 => x"34",
          2519 => x"3d",
          2520 => x"38",
          2521 => x"b8",
          2522 => x"fa",
          2523 => x"40",
          2524 => x"c7",
          2525 => x"33",
          2526 => x"22",
          2527 => x"56",
          2528 => x"fa",
          2529 => x"57",
          2530 => x"80",
          2531 => x"81",
          2532 => x"fa",
          2533 => x"42",
          2534 => x"60",
          2535 => x"58",
          2536 => x"ea",
          2537 => x"34",
          2538 => x"83",
          2539 => x"83",
          2540 => x"86",
          2541 => x"22",
          2542 => x"70",
          2543 => x"33",
          2544 => x"2e",
          2545 => x"ff",
          2546 => x"76",
          2547 => x"90",
          2548 => x"80",
          2549 => x"84",
          2550 => x"87",
          2551 => x"80",
          2552 => x"0d",
          2553 => x"ec",
          2554 => x"ed",
          2555 => x"ee",
          2556 => x"80",
          2557 => x"0d",
          2558 => x"06",
          2559 => x"84",
          2560 => x"83",
          2561 => x"72",
          2562 => x"05",
          2563 => x"7b",
          2564 => x"83",
          2565 => x"42",
          2566 => x"38",
          2567 => x"56",
          2568 => x"fa",
          2569 => x"81",
          2570 => x"72",
          2571 => x"a0",
          2572 => x"84",
          2573 => x"83",
          2574 => x"5a",
          2575 => x"b6",
          2576 => x"71",
          2577 => x"b0",
          2578 => x"84",
          2579 => x"83",
          2580 => x"72",
          2581 => x"59",
          2582 => x"d6",
          2583 => x"06",
          2584 => x"38",
          2585 => x"d0",
          2586 => x"b5",
          2587 => x"ff",
          2588 => x"39",
          2589 => x"bd",
          2590 => x"95",
          2591 => x"7e",
          2592 => x"75",
          2593 => x"10",
          2594 => x"04",
          2595 => x"52",
          2596 => x"84",
          2597 => x"83",
          2598 => x"70",
          2599 => x"70",
          2600 => x"86",
          2601 => x"22",
          2602 => x"83",
          2603 => x"46",
          2604 => x"81",
          2605 => x"81",
          2606 => x"81",
          2607 => x"58",
          2608 => x"a0",
          2609 => x"83",
          2610 => x"72",
          2611 => x"a0",
          2612 => x"fa",
          2613 => x"5e",
          2614 => x"80",
          2615 => x"81",
          2616 => x"fa",
          2617 => x"44",
          2618 => x"84",
          2619 => x"70",
          2620 => x"26",
          2621 => x"58",
          2622 => x"75",
          2623 => x"81",
          2624 => x"f7",
          2625 => x"b8",
          2626 => x"81",
          2627 => x"81",
          2628 => x"5b",
          2629 => x"33",
          2630 => x"b8",
          2631 => x"fa",
          2632 => x"41",
          2633 => x"1c",
          2634 => x"29",
          2635 => x"86",
          2636 => x"f8",
          2637 => x"b2",
          2638 => x"29",
          2639 => x"fa",
          2640 => x"60",
          2641 => x"58",
          2642 => x"83",
          2643 => x"0b",
          2644 => x"bb",
          2645 => x"fa",
          2646 => x"19",
          2647 => x"70",
          2648 => x"f9",
          2649 => x"34",
          2650 => x"3d",
          2651 => x"5b",
          2652 => x"83",
          2653 => x"83",
          2654 => x"5c",
          2655 => x"9c",
          2656 => x"ff",
          2657 => x"80",
          2658 => x"33",
          2659 => x"85",
          2660 => x"02",
          2661 => x"d8",
          2662 => x"b6",
          2663 => x"33",
          2664 => x"b8",
          2665 => x"5b",
          2666 => x"33",
          2667 => x"33",
          2668 => x"84",
          2669 => x"a0",
          2670 => x"83",
          2671 => x"72",
          2672 => x"78",
          2673 => x"b4",
          2674 => x"83",
          2675 => x"80",
          2676 => x"81",
          2677 => x"fa",
          2678 => x"5f",
          2679 => x"84",
          2680 => x"81",
          2681 => x"90",
          2682 => x"77",
          2683 => x"83",
          2684 => x"80",
          2685 => x"80",
          2686 => x"33",
          2687 => x"81",
          2688 => x"bb",
          2689 => x"ba",
          2690 => x"ba",
          2691 => x"ba",
          2692 => x"23",
          2693 => x"84",
          2694 => x"84",
          2695 => x"84",
          2696 => x"ba",
          2697 => x"93",
          2698 => x"86",
          2699 => x"83",
          2700 => x"fa",
          2701 => x"83",
          2702 => x"57",
          2703 => x"fd",
          2704 => x"ff",
          2705 => x"05",
          2706 => x"76",
          2707 => x"f5",
          2708 => x"ba",
          2709 => x"06",
          2710 => x"77",
          2711 => x"33",
          2712 => x"38",
          2713 => x"5f",
          2714 => x"5e",
          2715 => x"fa",
          2716 => x"71",
          2717 => x"06",
          2718 => x"fa",
          2719 => x"85",
          2720 => x"38",
          2721 => x"81",
          2722 => x"57",
          2723 => x"75",
          2724 => x"80",
          2725 => x"b4",
          2726 => x"7b",
          2727 => x"56",
          2728 => x"39",
          2729 => x"fa",
          2730 => x"05",
          2731 => x"38",
          2732 => x"34",
          2733 => x"40",
          2734 => x"fa",
          2735 => x"71",
          2736 => x"06",
          2737 => x"fa",
          2738 => x"85",
          2739 => x"38",
          2740 => x"2e",
          2741 => x"b8",
          2742 => x"fa",
          2743 => x"c7",
          2744 => x"43",
          2745 => x"70",
          2746 => x"08",
          2747 => x"5d",
          2748 => x"bf",
          2749 => x"fb",
          2750 => x"79",
          2751 => x"d8",
          2752 => x"06",
          2753 => x"89",
          2754 => x"33",
          2755 => x"84",
          2756 => x"5d",
          2757 => x"11",
          2758 => x"38",
          2759 => x"fb",
          2760 => x"76",
          2761 => x"d9",
          2762 => x"05",
          2763 => x"41",
          2764 => x"57",
          2765 => x"39",
          2766 => x"3f",
          2767 => x"57",
          2768 => x"10",
          2769 => x"5a",
          2770 => x"3f",
          2771 => x"ba",
          2772 => x"82",
          2773 => x"7d",
          2774 => x"22",
          2775 => x"57",
          2776 => x"d5",
          2777 => x"85",
          2778 => x"38",
          2779 => x"81",
          2780 => x"05",
          2781 => x"33",
          2782 => x"43",
          2783 => x"27",
          2784 => x"b2",
          2785 => x"58",
          2786 => x"57",
          2787 => x"f8",
          2788 => x"27",
          2789 => x"fa",
          2790 => x"85",
          2791 => x"38",
          2792 => x"33",
          2793 => x"38",
          2794 => x"33",
          2795 => x"33",
          2796 => x"80",
          2797 => x"71",
          2798 => x"06",
          2799 => x"59",
          2800 => x"38",
          2801 => x"31",
          2802 => x"38",
          2803 => x"27",
          2804 => x"83",
          2805 => x"70",
          2806 => x"8e",
          2807 => x"76",
          2808 => x"56",
          2809 => x"ff",
          2810 => x"80",
          2811 => x"77",
          2812 => x"71",
          2813 => x"86",
          2814 => x"80",
          2815 => x"06",
          2816 => x"5c",
          2817 => x"99",
          2818 => x"5f",
          2819 => x"81",
          2820 => x"58",
          2821 => x"81",
          2822 => x"f7",
          2823 => x"5e",
          2824 => x"e0",
          2825 => x"1f",
          2826 => x"76",
          2827 => x"81",
          2828 => x"f8",
          2829 => x"29",
          2830 => x"26",
          2831 => x"ba",
          2832 => x"e0",
          2833 => x"51",
          2834 => x"0b",
          2835 => x"ba",
          2836 => x"78",
          2837 => x"56",
          2838 => x"be",
          2839 => x"81",
          2840 => x"43",
          2841 => x"38",
          2842 => x"26",
          2843 => x"56",
          2844 => x"76",
          2845 => x"f5",
          2846 => x"90",
          2847 => x"11",
          2848 => x"80",
          2849 => x"75",
          2850 => x"76",
          2851 => x"70",
          2852 => x"88",
          2853 => x"52",
          2854 => x"80",
          2855 => x"76",
          2856 => x"26",
          2857 => x"b8",
          2858 => x"06",
          2859 => x"22",
          2860 => x"59",
          2861 => x"78",
          2862 => x"57",
          2863 => x"76",
          2864 => x"33",
          2865 => x"0b",
          2866 => x"81",
          2867 => x"76",
          2868 => x"e0",
          2869 => x"5a",
          2870 => x"d6",
          2871 => x"81",
          2872 => x"83",
          2873 => x"71",
          2874 => x"2a",
          2875 => x"2e",
          2876 => x"0b",
          2877 => x"81",
          2878 => x"83",
          2879 => x"80",
          2880 => x"33",
          2881 => x"22",
          2882 => x"5d",
          2883 => x"87",
          2884 => x"81",
          2885 => x"f4",
          2886 => x"fd",
          2887 => x"b0",
          2888 => x"81",
          2889 => x"fa",
          2890 => x"33",
          2891 => x"83",
          2892 => x"b0",
          2893 => x"75",
          2894 => x"80",
          2895 => x"18",
          2896 => x"a4",
          2897 => x"06",
          2898 => x"8f",
          2899 => x"06",
          2900 => x"34",
          2901 => x"81",
          2902 => x"83",
          2903 => x"fa",
          2904 => x"07",
          2905 => x"d7",
          2906 => x"06",
          2907 => x"34",
          2908 => x"81",
          2909 => x"fa",
          2910 => x"b0",
          2911 => x"75",
          2912 => x"83",
          2913 => x"07",
          2914 => x"8f",
          2915 => x"06",
          2916 => x"ff",
          2917 => x"07",
          2918 => x"ef",
          2919 => x"07",
          2920 => x"df",
          2921 => x"06",
          2922 => x"b0",
          2923 => x"33",
          2924 => x"83",
          2925 => x"0b",
          2926 => x"51",
          2927 => x"ba",
          2928 => x"ba",
          2929 => x"ba",
          2930 => x"23",
          2931 => x"c7",
          2932 => x"80",
          2933 => x"0d",
          2934 => x"fa",
          2935 => x"ff",
          2936 => x"88",
          2937 => x"05",
          2938 => x"84",
          2939 => x"84",
          2940 => x"84",
          2941 => x"9c",
          2942 => x"34",
          2943 => x"81",
          2944 => x"34",
          2945 => x"80",
          2946 => x"23",
          2947 => x"39",
          2948 => x"52",
          2949 => x"b5",
          2950 => x"05",
          2951 => x"fa",
          2952 => x"fb",
          2953 => x"ea",
          2954 => x"b5",
          2955 => x"2c",
          2956 => x"39",
          2957 => x"b8",
          2958 => x"eb",
          2959 => x"e3",
          2960 => x"70",
          2961 => x"40",
          2962 => x"33",
          2963 => x"11",
          2964 => x"c0",
          2965 => x"b8",
          2966 => x"5c",
          2967 => x"fa",
          2968 => x"81",
          2969 => x"74",
          2970 => x"83",
          2971 => x"29",
          2972 => x"f9",
          2973 => x"5d",
          2974 => x"83",
          2975 => x"80",
          2976 => x"f7",
          2977 => x"38",
          2978 => x"23",
          2979 => x"57",
          2980 => x"b8",
          2981 => x"ec",
          2982 => x"b4",
          2983 => x"b2",
          2984 => x"26",
          2985 => x"7e",
          2986 => x"5e",
          2987 => x"5b",
          2988 => x"06",
          2989 => x"1d",
          2990 => x"ec",
          2991 => x"e0",
          2992 => x"1e",
          2993 => x"76",
          2994 => x"81",
          2995 => x"f8",
          2996 => x"29",
          2997 => x"27",
          2998 => x"5e",
          2999 => x"81",
          3000 => x"58",
          3001 => x"81",
          3002 => x"f7",
          3003 => x"5d",
          3004 => x"eb",
          3005 => x"5c",
          3006 => x"83",
          3007 => x"83",
          3008 => x"5f",
          3009 => x"eb",
          3010 => x"81",
          3011 => x"76",
          3012 => x"83",
          3013 => x"ff",
          3014 => x"38",
          3015 => x"84",
          3016 => x"ff",
          3017 => x"eb",
          3018 => x"b5",
          3019 => x"33",
          3020 => x"11",
          3021 => x"ca",
          3022 => x"81",
          3023 => x"83",
          3024 => x"83",
          3025 => x"57",
          3026 => x"b8",
          3027 => x"75",
          3028 => x"ff",
          3029 => x"fc",
          3030 => x"83",
          3031 => x"7d",
          3032 => x"38",
          3033 => x"83",
          3034 => x"59",
          3035 => x"80",
          3036 => x"fa",
          3037 => x"34",
          3038 => x"39",
          3039 => x"b2",
          3040 => x"fa",
          3041 => x"fa",
          3042 => x"83",
          3043 => x"0b",
          3044 => x"83",
          3045 => x"80",
          3046 => x"f9",
          3047 => x"0d",
          3048 => x"33",
          3049 => x"73",
          3050 => x"bb",
          3051 => x"52",
          3052 => x"84",
          3053 => x"f3",
          3054 => x"ff",
          3055 => x"ff",
          3056 => x"55",
          3057 => x"38",
          3058 => x"34",
          3059 => x"8f",
          3060 => x"54",
          3061 => x"73",
          3062 => x"09",
          3063 => x"72",
          3064 => x"54",
          3065 => x"38",
          3066 => x"70",
          3067 => x"79",
          3068 => x"f8",
          3069 => x"b4",
          3070 => x"a0",
          3071 => x"59",
          3072 => x"ff",
          3073 => x"59",
          3074 => x"38",
          3075 => x"80",
          3076 => x"0c",
          3077 => x"80",
          3078 => x"08",
          3079 => x"81",
          3080 => x"81",
          3081 => x"83",
          3082 => x"06",
          3083 => x"55",
          3084 => x"81",
          3085 => x"f8",
          3086 => x"5a",
          3087 => x"75",
          3088 => x"a4",
          3089 => x"81",
          3090 => x"89",
          3091 => x"ac",
          3092 => x"58",
          3093 => x"73",
          3094 => x"32",
          3095 => x"80",
          3096 => x"f8",
          3097 => x"72",
          3098 => x"83",
          3099 => x"dd",
          3100 => x"de",
          3101 => x"f8",
          3102 => x"5e",
          3103 => x"74",
          3104 => x"cc",
          3105 => x"82",
          3106 => x"72",
          3107 => x"cc",
          3108 => x"74",
          3109 => x"2e",
          3110 => x"53",
          3111 => x"81",
          3112 => x"84",
          3113 => x"54",
          3114 => x"f8",
          3115 => x"98",
          3116 => x"83",
          3117 => x"9c",
          3118 => x"16",
          3119 => x"76",
          3120 => x"df",
          3121 => x"9e",
          3122 => x"38",
          3123 => x"5a",
          3124 => x"54",
          3125 => x"14",
          3126 => x"7d",
          3127 => x"83",
          3128 => x"2e",
          3129 => x"8a",
          3130 => x"f9",
          3131 => x"77",
          3132 => x"17",
          3133 => x"76",
          3134 => x"83",
          3135 => x"82",
          3136 => x"38",
          3137 => x"fc",
          3138 => x"80",
          3139 => x"2e",
          3140 => x"06",
          3141 => x"ed",
          3142 => x"79",
          3143 => x"75",
          3144 => x"a1",
          3145 => x"17",
          3146 => x"fe",
          3147 => x"57",
          3148 => x"e1",
          3149 => x"05",
          3150 => x"f5",
          3151 => x"78",
          3152 => x"d8",
          3153 => x"7d",
          3154 => x"ff",
          3155 => x"ff",
          3156 => x"38",
          3157 => x"54",
          3158 => x"82",
          3159 => x"07",
          3160 => x"83",
          3161 => x"78",
          3162 => x"72",
          3163 => x"70",
          3164 => x"ba",
          3165 => x"54",
          3166 => x"b8",
          3167 => x"9a",
          3168 => x"f9",
          3169 => x"82",
          3170 => x"84",
          3171 => x"34",
          3172 => x"81",
          3173 => x"14",
          3174 => x"cc",
          3175 => x"83",
          3176 => x"f8",
          3177 => x"c2",
          3178 => x"ff",
          3179 => x"96",
          3180 => x"81",
          3181 => x"ff",
          3182 => x"06",
          3183 => x"81",
          3184 => x"54",
          3185 => x"87",
          3186 => x"0c",
          3187 => x"39",
          3188 => x"f9",
          3189 => x"73",
          3190 => x"38",
          3191 => x"83",
          3192 => x"83",
          3193 => x"33",
          3194 => x"5e",
          3195 => x"82",
          3196 => x"7a",
          3197 => x"79",
          3198 => x"38",
          3199 => x"f0",
          3200 => x"b8",
          3201 => x"81",
          3202 => x"59",
          3203 => x"fa",
          3204 => x"54",
          3205 => x"f7",
          3206 => x"08",
          3207 => x"83",
          3208 => x"b8",
          3209 => x"11",
          3210 => x"38",
          3211 => x"73",
          3212 => x"80",
          3213 => x"83",
          3214 => x"70",
          3215 => x"80",
          3216 => x"83",
          3217 => x"39",
          3218 => x"3f",
          3219 => x"fc",
          3220 => x"f8",
          3221 => x"0b",
          3222 => x"33",
          3223 => x"81",
          3224 => x"04",
          3225 => x"90",
          3226 => x"82",
          3227 => x"80",
          3228 => x"90",
          3229 => x"34",
          3230 => x"87",
          3231 => x"08",
          3232 => x"c0",
          3233 => x"9c",
          3234 => x"81",
          3235 => x"56",
          3236 => x"81",
          3237 => x"a4",
          3238 => x"80",
          3239 => x"80",
          3240 => x"80",
          3241 => x"9c",
          3242 => x"55",
          3243 => x"33",
          3244 => x"70",
          3245 => x"2e",
          3246 => x"55",
          3247 => x"71",
          3248 => x"57",
          3249 => x"81",
          3250 => x"74",
          3251 => x"84",
          3252 => x"84",
          3253 => x"fa",
          3254 => x"05",
          3255 => x"90",
          3256 => x"80",
          3257 => x"55",
          3258 => x"90",
          3259 => x"90",
          3260 => x"86",
          3261 => x"74",
          3262 => x"51",
          3263 => x"f5",
          3264 => x"15",
          3265 => x"34",
          3266 => x"90",
          3267 => x"87",
          3268 => x"98",
          3269 => x"38",
          3270 => x"08",
          3271 => x"71",
          3272 => x"98",
          3273 => x"27",
          3274 => x"2e",
          3275 => x"08",
          3276 => x"98",
          3277 => x"08",
          3278 => x"14",
          3279 => x"52",
          3280 => x"ff",
          3281 => x"08",
          3282 => x"52",
          3283 => x"06",
          3284 => x"38",
          3285 => x"d4",
          3286 => x"56",
          3287 => x"84",
          3288 => x"27",
          3289 => x"33",
          3290 => x"71",
          3291 => x"0c",
          3292 => x"bb",
          3293 => x"51",
          3294 => x"84",
          3295 => x"0b",
          3296 => x"87",
          3297 => x"2a",
          3298 => x"15",
          3299 => x"15",
          3300 => x"15",
          3301 => x"f5",
          3302 => x"13",
          3303 => x"97",
          3304 => x"72",
          3305 => x"26",
          3306 => x"74",
          3307 => x"55",
          3308 => x"f5",
          3309 => x"15",
          3310 => x"34",
          3311 => x"90",
          3312 => x"87",
          3313 => x"98",
          3314 => x"38",
          3315 => x"08",
          3316 => x"71",
          3317 => x"98",
          3318 => x"27",
          3319 => x"2e",
          3320 => x"08",
          3321 => x"98",
          3322 => x"08",
          3323 => x"14",
          3324 => x"52",
          3325 => x"ff",
          3326 => x"08",
          3327 => x"52",
          3328 => x"06",
          3329 => x"74",
          3330 => x"38",
          3331 => x"73",
          3332 => x"84",
          3333 => x"ff",
          3334 => x"f5",
          3335 => x"85",
          3336 => x"fe",
          3337 => x"90",
          3338 => x"08",
          3339 => x"90",
          3340 => x"52",
          3341 => x"72",
          3342 => x"c0",
          3343 => x"27",
          3344 => x"38",
          3345 => x"53",
          3346 => x"53",
          3347 => x"c0",
          3348 => x"53",
          3349 => x"c0",
          3350 => x"f6",
          3351 => x"9c",
          3352 => x"38",
          3353 => x"c0",
          3354 => x"83",
          3355 => x"70",
          3356 => x"2e",
          3357 => x"73",
          3358 => x"0d",
          3359 => x"3f",
          3360 => x"84",
          3361 => x"2a",
          3362 => x"2b",
          3363 => x"71",
          3364 => x"11",
          3365 => x"2b",
          3366 => x"53",
          3367 => x"53",
          3368 => x"16",
          3369 => x"8b",
          3370 => x"70",
          3371 => x"71",
          3372 => x"59",
          3373 => x"38",
          3374 => x"8b",
          3375 => x"76",
          3376 => x"86",
          3377 => x"73",
          3378 => x"70",
          3379 => x"71",
          3380 => x"55",
          3381 => x"71",
          3382 => x"16",
          3383 => x"0b",
          3384 => x"53",
          3385 => x"34",
          3386 => x"81",
          3387 => x"80",
          3388 => x"52",
          3389 => x"34",
          3390 => x"87",
          3391 => x"2b",
          3392 => x"17",
          3393 => x"2a",
          3394 => x"71",
          3395 => x"84",
          3396 => x"33",
          3397 => x"83",
          3398 => x"05",
          3399 => x"88",
          3400 => x"59",
          3401 => x"13",
          3402 => x"33",
          3403 => x"81",
          3404 => x"5a",
          3405 => x"13",
          3406 => x"70",
          3407 => x"71",
          3408 => x"81",
          3409 => x"83",
          3410 => x"7b",
          3411 => x"5a",
          3412 => x"73",
          3413 => x"70",
          3414 => x"8b",
          3415 => x"70",
          3416 => x"07",
          3417 => x"5f",
          3418 => x"77",
          3419 => x"ba",
          3420 => x"83",
          3421 => x"2b",
          3422 => x"33",
          3423 => x"58",
          3424 => x"70",
          3425 => x"81",
          3426 => x"80",
          3427 => x"54",
          3428 => x"84",
          3429 => x"81",
          3430 => x"2b",
          3431 => x"15",
          3432 => x"2a",
          3433 => x"53",
          3434 => x"34",
          3435 => x"79",
          3436 => x"80",
          3437 => x"38",
          3438 => x"0d",
          3439 => x"f4",
          3440 => x"23",
          3441 => x"ff",
          3442 => x"ba",
          3443 => x"0b",
          3444 => x"54",
          3445 => x"15",
          3446 => x"86",
          3447 => x"84",
          3448 => x"ff",
          3449 => x"ff",
          3450 => x"55",
          3451 => x"17",
          3452 => x"10",
          3453 => x"05",
          3454 => x"0b",
          3455 => x"3d",
          3456 => x"84",
          3457 => x"2a",
          3458 => x"51",
          3459 => x"ba",
          3460 => x"33",
          3461 => x"5a",
          3462 => x"80",
          3463 => x"10",
          3464 => x"88",
          3465 => x"79",
          3466 => x"7a",
          3467 => x"72",
          3468 => x"85",
          3469 => x"33",
          3470 => x"57",
          3471 => x"ff",
          3472 => x"80",
          3473 => x"81",
          3474 => x"81",
          3475 => x"59",
          3476 => x"59",
          3477 => x"38",
          3478 => x"38",
          3479 => x"16",
          3480 => x"80",
          3481 => x"56",
          3482 => x"15",
          3483 => x"88",
          3484 => x"75",
          3485 => x"70",
          3486 => x"88",
          3487 => x"f8",
          3488 => x"06",
          3489 => x"59",
          3490 => x"81",
          3491 => x"84",
          3492 => x"34",
          3493 => x"08",
          3494 => x"33",
          3495 => x"74",
          3496 => x"84",
          3497 => x"ba",
          3498 => x"86",
          3499 => x"2b",
          3500 => x"59",
          3501 => x"34",
          3502 => x"11",
          3503 => x"71",
          3504 => x"5c",
          3505 => x"87",
          3506 => x"16",
          3507 => x"12",
          3508 => x"2a",
          3509 => x"34",
          3510 => x"08",
          3511 => x"84",
          3512 => x"33",
          3513 => x"83",
          3514 => x"85",
          3515 => x"88",
          3516 => x"74",
          3517 => x"84",
          3518 => x"33",
          3519 => x"83",
          3520 => x"87",
          3521 => x"88",
          3522 => x"57",
          3523 => x"1a",
          3524 => x"33",
          3525 => x"81",
          3526 => x"57",
          3527 => x"18",
          3528 => x"05",
          3529 => x"79",
          3530 => x"80",
          3531 => x"38",
          3532 => x"0d",
          3533 => x"bb",
          3534 => x"3d",
          3535 => x"ba",
          3536 => x"f0",
          3537 => x"84",
          3538 => x"84",
          3539 => x"81",
          3540 => x"08",
          3541 => x"85",
          3542 => x"76",
          3543 => x"34",
          3544 => x"22",
          3545 => x"83",
          3546 => x"51",
          3547 => x"89",
          3548 => x"10",
          3549 => x"f8",
          3550 => x"81",
          3551 => x"80",
          3552 => x"ed",
          3553 => x"70",
          3554 => x"76",
          3555 => x"2e",
          3556 => x"d7",
          3557 => x"38",
          3558 => x"70",
          3559 => x"83",
          3560 => x"2a",
          3561 => x"2b",
          3562 => x"71",
          3563 => x"83",
          3564 => x"fc",
          3565 => x"33",
          3566 => x"70",
          3567 => x"45",
          3568 => x"48",
          3569 => x"24",
          3570 => x"16",
          3571 => x"10",
          3572 => x"71",
          3573 => x"5c",
          3574 => x"85",
          3575 => x"38",
          3576 => x"a2",
          3577 => x"60",
          3578 => x"38",
          3579 => x"f7",
          3580 => x"33",
          3581 => x"7a",
          3582 => x"98",
          3583 => x"59",
          3584 => x"24",
          3585 => x"33",
          3586 => x"83",
          3587 => x"87",
          3588 => x"2b",
          3589 => x"15",
          3590 => x"2a",
          3591 => x"53",
          3592 => x"79",
          3593 => x"70",
          3594 => x"71",
          3595 => x"05",
          3596 => x"88",
          3597 => x"5e",
          3598 => x"16",
          3599 => x"f4",
          3600 => x"71",
          3601 => x"70",
          3602 => x"79",
          3603 => x"f4",
          3604 => x"12",
          3605 => x"07",
          3606 => x"71",
          3607 => x"5c",
          3608 => x"79",
          3609 => x"f4",
          3610 => x"33",
          3611 => x"74",
          3612 => x"71",
          3613 => x"5c",
          3614 => x"82",
          3615 => x"ba",
          3616 => x"83",
          3617 => x"57",
          3618 => x"5a",
          3619 => x"c3",
          3620 => x"84",
          3621 => x"ff",
          3622 => x"26",
          3623 => x"bb",
          3624 => x"ff",
          3625 => x"80",
          3626 => x"80",
          3627 => x"fe",
          3628 => x"5e",
          3629 => x"34",
          3630 => x"1e",
          3631 => x"ba",
          3632 => x"81",
          3633 => x"08",
          3634 => x"80",
          3635 => x"70",
          3636 => x"88",
          3637 => x"ba",
          3638 => x"ba",
          3639 => x"60",
          3640 => x"34",
          3641 => x"d3",
          3642 => x"7e",
          3643 => x"7f",
          3644 => x"08",
          3645 => x"04",
          3646 => x"83",
          3647 => x"70",
          3648 => x"07",
          3649 => x"48",
          3650 => x"60",
          3651 => x"08",
          3652 => x"82",
          3653 => x"ba",
          3654 => x"12",
          3655 => x"2b",
          3656 => x"83",
          3657 => x"5c",
          3658 => x"82",
          3659 => x"60",
          3660 => x"08",
          3661 => x"1c",
          3662 => x"84",
          3663 => x"fd",
          3664 => x"ff",
          3665 => x"77",
          3666 => x"83",
          3667 => x"18",
          3668 => x"10",
          3669 => x"71",
          3670 => x"5e",
          3671 => x"80",
          3672 => x"61",
          3673 => x"24",
          3674 => x"06",
          3675 => x"fe",
          3676 => x"ba",
          3677 => x"f0",
          3678 => x"84",
          3679 => x"84",
          3680 => x"81",
          3681 => x"08",
          3682 => x"85",
          3683 => x"7e",
          3684 => x"34",
          3685 => x"22",
          3686 => x"83",
          3687 => x"56",
          3688 => x"73",
          3689 => x"22",
          3690 => x"08",
          3691 => x"82",
          3692 => x"fc",
          3693 => x"38",
          3694 => x"7b",
          3695 => x"76",
          3696 => x"ea",
          3697 => x"84",
          3698 => x"82",
          3699 => x"2b",
          3700 => x"11",
          3701 => x"71",
          3702 => x"33",
          3703 => x"70",
          3704 => x"46",
          3705 => x"84",
          3706 => x"84",
          3707 => x"33",
          3708 => x"83",
          3709 => x"87",
          3710 => x"88",
          3711 => x"5d",
          3712 => x"64",
          3713 => x"16",
          3714 => x"2b",
          3715 => x"2a",
          3716 => x"79",
          3717 => x"70",
          3718 => x"71",
          3719 => x"05",
          3720 => x"2b",
          3721 => x"40",
          3722 => x"75",
          3723 => x"70",
          3724 => x"8b",
          3725 => x"82",
          3726 => x"2b",
          3727 => x"5b",
          3728 => x"34",
          3729 => x"08",
          3730 => x"33",
          3731 => x"56",
          3732 => x"7e",
          3733 => x"3f",
          3734 => x"78",
          3735 => x"99",
          3736 => x"f4",
          3737 => x"23",
          3738 => x"ff",
          3739 => x"ba",
          3740 => x"0b",
          3741 => x"55",
          3742 => x"16",
          3743 => x"86",
          3744 => x"84",
          3745 => x"ff",
          3746 => x"ff",
          3747 => x"44",
          3748 => x"1f",
          3749 => x"10",
          3750 => x"05",
          3751 => x"0b",
          3752 => x"3f",
          3753 => x"33",
          3754 => x"83",
          3755 => x"85",
          3756 => x"88",
          3757 => x"76",
          3758 => x"05",
          3759 => x"84",
          3760 => x"2b",
          3761 => x"14",
          3762 => x"07",
          3763 => x"59",
          3764 => x"34",
          3765 => x"f4",
          3766 => x"71",
          3767 => x"70",
          3768 => x"78",
          3769 => x"f4",
          3770 => x"33",
          3771 => x"74",
          3772 => x"88",
          3773 => x"f8",
          3774 => x"5d",
          3775 => x"7f",
          3776 => x"84",
          3777 => x"81",
          3778 => x"2b",
          3779 => x"33",
          3780 => x"06",
          3781 => x"46",
          3782 => x"60",
          3783 => x"06",
          3784 => x"87",
          3785 => x"2b",
          3786 => x"19",
          3787 => x"2a",
          3788 => x"84",
          3789 => x"ba",
          3790 => x"85",
          3791 => x"2b",
          3792 => x"15",
          3793 => x"2a",
          3794 => x"56",
          3795 => x"87",
          3796 => x"70",
          3797 => x"07",
          3798 => x"5b",
          3799 => x"81",
          3800 => x"1f",
          3801 => x"2b",
          3802 => x"33",
          3803 => x"70",
          3804 => x"05",
          3805 => x"58",
          3806 => x"34",
          3807 => x"08",
          3808 => x"71",
          3809 => x"05",
          3810 => x"2b",
          3811 => x"2a",
          3812 => x"55",
          3813 => x"84",
          3814 => x"33",
          3815 => x"83",
          3816 => x"87",
          3817 => x"2b",
          3818 => x"15",
          3819 => x"2a",
          3820 => x"53",
          3821 => x"34",
          3822 => x"08",
          3823 => x"33",
          3824 => x"74",
          3825 => x"71",
          3826 => x"42",
          3827 => x"86",
          3828 => x"ba",
          3829 => x"33",
          3830 => x"06",
          3831 => x"76",
          3832 => x"ba",
          3833 => x"83",
          3834 => x"2b",
          3835 => x"33",
          3836 => x"41",
          3837 => x"79",
          3838 => x"ba",
          3839 => x"12",
          3840 => x"07",
          3841 => x"33",
          3842 => x"41",
          3843 => x"79",
          3844 => x"84",
          3845 => x"33",
          3846 => x"66",
          3847 => x"52",
          3848 => x"fe",
          3849 => x"1e",
          3850 => x"83",
          3851 => x"d5",
          3852 => x"71",
          3853 => x"05",
          3854 => x"88",
          3855 => x"5d",
          3856 => x"34",
          3857 => x"f4",
          3858 => x"12",
          3859 => x"07",
          3860 => x"33",
          3861 => x"5b",
          3862 => x"73",
          3863 => x"05",
          3864 => x"33",
          3865 => x"81",
          3866 => x"5f",
          3867 => x"16",
          3868 => x"70",
          3869 => x"71",
          3870 => x"81",
          3871 => x"83",
          3872 => x"63",
          3873 => x"5e",
          3874 => x"7b",
          3875 => x"70",
          3876 => x"8b",
          3877 => x"70",
          3878 => x"07",
          3879 => x"47",
          3880 => x"7f",
          3881 => x"83",
          3882 => x"7e",
          3883 => x"bb",
          3884 => x"80",
          3885 => x"84",
          3886 => x"3f",
          3887 => x"61",
          3888 => x"39",
          3889 => x"ba",
          3890 => x"b7",
          3891 => x"84",
          3892 => x"77",
          3893 => x"08",
          3894 => x"e6",
          3895 => x"84",
          3896 => x"84",
          3897 => x"84",
          3898 => x"a0",
          3899 => x"80",
          3900 => x"51",
          3901 => x"08",
          3902 => x"16",
          3903 => x"84",
          3904 => x"84",
          3905 => x"34",
          3906 => x"f4",
          3907 => x"fe",
          3908 => x"06",
          3909 => x"74",
          3910 => x"84",
          3911 => x"84",
          3912 => x"55",
          3913 => x"15",
          3914 => x"c6",
          3915 => x"02",
          3916 => x"72",
          3917 => x"33",
          3918 => x"3d",
          3919 => x"05",
          3920 => x"9d",
          3921 => x"bb",
          3922 => x"87",
          3923 => x"84",
          3924 => x"bb",
          3925 => x"3d",
          3926 => x"af",
          3927 => x"54",
          3928 => x"80",
          3929 => x"83",
          3930 => x"0b",
          3931 => x"75",
          3932 => x"bb",
          3933 => x"80",
          3934 => x"08",
          3935 => x"d6",
          3936 => x"73",
          3937 => x"55",
          3938 => x"0d",
          3939 => x"81",
          3940 => x"26",
          3941 => x"0d",
          3942 => x"05",
          3943 => x"76",
          3944 => x"17",
          3945 => x"55",
          3946 => x"87",
          3947 => x"52",
          3948 => x"84",
          3949 => x"2e",
          3950 => x"54",
          3951 => x"38",
          3952 => x"80",
          3953 => x"74",
          3954 => x"04",
          3955 => x"ff",
          3956 => x"ff",
          3957 => x"78",
          3958 => x"88",
          3959 => x"81",
          3960 => x"bb",
          3961 => x"54",
          3962 => x"87",
          3963 => x"73",
          3964 => x"38",
          3965 => x"72",
          3966 => x"04",
          3967 => x"bb",
          3968 => x"80",
          3969 => x"0c",
          3970 => x"87",
          3971 => x"cd",
          3972 => x"06",
          3973 => x"87",
          3974 => x"38",
          3975 => x"ca",
          3976 => x"8c",
          3977 => x"73",
          3978 => x"82",
          3979 => x"39",
          3980 => x"83",
          3981 => x"77",
          3982 => x"33",
          3983 => x"80",
          3984 => x"fe",
          3985 => x"2e",
          3986 => x"84",
          3987 => x"b4",
          3988 => x"81",
          3989 => x"81",
          3990 => x"09",
          3991 => x"08",
          3992 => x"a8",
          3993 => x"bb",
          3994 => x"76",
          3995 => x"55",
          3996 => x"8e",
          3997 => x"52",
          3998 => x"76",
          3999 => x"09",
          4000 => x"33",
          4001 => x"fe",
          4002 => x"7a",
          4003 => x"57",
          4004 => x"80",
          4005 => x"aa",
          4006 => x"7a",
          4007 => x"80",
          4008 => x"0b",
          4009 => x"9c",
          4010 => x"19",
          4011 => x"34",
          4012 => x"94",
          4013 => x"34",
          4014 => x"19",
          4015 => x"a2",
          4016 => x"84",
          4017 => x"7a",
          4018 => x"55",
          4019 => x"2a",
          4020 => x"98",
          4021 => x"a4",
          4022 => x"0c",
          4023 => x"81",
          4024 => x"84",
          4025 => x"18",
          4026 => x"84",
          4027 => x"b2",
          4028 => x"08",
          4029 => x"38",
          4030 => x"81",
          4031 => x"3d",
          4032 => x"74",
          4033 => x"24",
          4034 => x"81",
          4035 => x"70",
          4036 => x"5a",
          4037 => x"b0",
          4038 => x"2e",
          4039 => x"54",
          4040 => x"33",
          4041 => x"08",
          4042 => x"5b",
          4043 => x"38",
          4044 => x"33",
          4045 => x"08",
          4046 => x"08",
          4047 => x"18",
          4048 => x"2e",
          4049 => x"54",
          4050 => x"33",
          4051 => x"08",
          4052 => x"5a",
          4053 => x"38",
          4054 => x"33",
          4055 => x"06",
          4056 => x"5d",
          4057 => x"06",
          4058 => x"04",
          4059 => x"59",
          4060 => x"80",
          4061 => x"5b",
          4062 => x"c2",
          4063 => x"52",
          4064 => x"84",
          4065 => x"ff",
          4066 => x"79",
          4067 => x"06",
          4068 => x"71",
          4069 => x"84",
          4070 => x"74",
          4071 => x"38",
          4072 => x"59",
          4073 => x"80",
          4074 => x"5b",
          4075 => x"81",
          4076 => x"52",
          4077 => x"84",
          4078 => x"ff",
          4079 => x"79",
          4080 => x"fc",
          4081 => x"33",
          4082 => x"88",
          4083 => x"07",
          4084 => x"ff",
          4085 => x"0c",
          4086 => x"3d",
          4087 => x"53",
          4088 => x"52",
          4089 => x"bb",
          4090 => x"fe",
          4091 => x"18",
          4092 => x"31",
          4093 => x"a0",
          4094 => x"17",
          4095 => x"06",
          4096 => x"08",
          4097 => x"81",
          4098 => x"5a",
          4099 => x"08",
          4100 => x"33",
          4101 => x"84",
          4102 => x"81",
          4103 => x"34",
          4104 => x"5d",
          4105 => x"82",
          4106 => x"cb",
          4107 => x"de",
          4108 => x"b8",
          4109 => x"5c",
          4110 => x"84",
          4111 => x"ff",
          4112 => x"34",
          4113 => x"84",
          4114 => x"18",
          4115 => x"33",
          4116 => x"fd",
          4117 => x"a0",
          4118 => x"17",
          4119 => x"fd",
          4120 => x"53",
          4121 => x"52",
          4122 => x"bb",
          4123 => x"fb",
          4124 => x"18",
          4125 => x"31",
          4126 => x"a0",
          4127 => x"17",
          4128 => x"06",
          4129 => x"08",
          4130 => x"81",
          4131 => x"5a",
          4132 => x"08",
          4133 => x"81",
          4134 => x"86",
          4135 => x"fa",
          4136 => x"64",
          4137 => x"27",
          4138 => x"95",
          4139 => x"96",
          4140 => x"74",
          4141 => x"bb",
          4142 => x"88",
          4143 => x"0b",
          4144 => x"2e",
          4145 => x"5b",
          4146 => x"83",
          4147 => x"19",
          4148 => x"3f",
          4149 => x"38",
          4150 => x"0c",
          4151 => x"10",
          4152 => x"ff",
          4153 => x"34",
          4154 => x"34",
          4155 => x"bb",
          4156 => x"83",
          4157 => x"75",
          4158 => x"80",
          4159 => x"78",
          4160 => x"7c",
          4161 => x"06",
          4162 => x"b8",
          4163 => x"8e",
          4164 => x"85",
          4165 => x"1a",
          4166 => x"75",
          4167 => x"b8",
          4168 => x"8f",
          4169 => x"41",
          4170 => x"88",
          4171 => x"90",
          4172 => x"98",
          4173 => x"0b",
          4174 => x"81",
          4175 => x"08",
          4176 => x"76",
          4177 => x"1a",
          4178 => x"2e",
          4179 => x"54",
          4180 => x"33",
          4181 => x"08",
          4182 => x"5c",
          4183 => x"fd",
          4184 => x"b8",
          4185 => x"5f",
          4186 => x"38",
          4187 => x"33",
          4188 => x"77",
          4189 => x"89",
          4190 => x"0b",
          4191 => x"2e",
          4192 => x"b8",
          4193 => x"57",
          4194 => x"84",
          4195 => x"c7",
          4196 => x"34",
          4197 => x"31",
          4198 => x"5b",
          4199 => x"38",
          4200 => x"82",
          4201 => x"52",
          4202 => x"84",
          4203 => x"ff",
          4204 => x"77",
          4205 => x"19",
          4206 => x"7c",
          4207 => x"81",
          4208 => x"5c",
          4209 => x"34",
          4210 => x"b8",
          4211 => x"5d",
          4212 => x"84",
          4213 => x"88",
          4214 => x"34",
          4215 => x"31",
          4216 => x"5d",
          4217 => x"ca",
          4218 => x"2e",
          4219 => x"54",
          4220 => x"33",
          4221 => x"aa",
          4222 => x"70",
          4223 => x"ad",
          4224 => x"7d",
          4225 => x"84",
          4226 => x"19",
          4227 => x"1b",
          4228 => x"56",
          4229 => x"82",
          4230 => x"81",
          4231 => x"1f",
          4232 => x"ed",
          4233 => x"81",
          4234 => x"81",
          4235 => x"81",
          4236 => x"09",
          4237 => x"84",
          4238 => x"70",
          4239 => x"84",
          4240 => x"7e",
          4241 => x"33",
          4242 => x"fa",
          4243 => x"76",
          4244 => x"3f",
          4245 => x"79",
          4246 => x"51",
          4247 => x"39",
          4248 => x"05",
          4249 => x"58",
          4250 => x"5a",
          4251 => x"7e",
          4252 => x"2b",
          4253 => x"83",
          4254 => x"06",
          4255 => x"5f",
          4256 => x"2a",
          4257 => x"2a",
          4258 => x"2a",
          4259 => x"39",
          4260 => x"5b",
          4261 => x"19",
          4262 => x"38",
          4263 => x"38",
          4264 => x"80",
          4265 => x"81",
          4266 => x"9c",
          4267 => x"56",
          4268 => x"52",
          4269 => x"84",
          4270 => x"58",
          4271 => x"38",
          4272 => x"70",
          4273 => x"51",
          4274 => x"75",
          4275 => x"38",
          4276 => x"8c",
          4277 => x"39",
          4278 => x"7a",
          4279 => x"55",
          4280 => x"38",
          4281 => x"84",
          4282 => x"08",
          4283 => x"7a",
          4284 => x"9c",
          4285 => x"56",
          4286 => x"80",
          4287 => x"81",
          4288 => x"70",
          4289 => x"7b",
          4290 => x"51",
          4291 => x"bb",
          4292 => x"19",
          4293 => x"38",
          4294 => x"38",
          4295 => x"75",
          4296 => x"75",
          4297 => x"bb",
          4298 => x"70",
          4299 => x"56",
          4300 => x"80",
          4301 => x"19",
          4302 => x"58",
          4303 => x"94",
          4304 => x"5a",
          4305 => x"84",
          4306 => x"80",
          4307 => x"0d",
          4308 => x"da",
          4309 => x"75",
          4310 => x"3f",
          4311 => x"39",
          4312 => x"0c",
          4313 => x"81",
          4314 => x"b6",
          4315 => x"08",
          4316 => x"26",
          4317 => x"72",
          4318 => x"88",
          4319 => x"76",
          4320 => x"38",
          4321 => x"18",
          4322 => x"38",
          4323 => x"94",
          4324 => x"56",
          4325 => x"2a",
          4326 => x"06",
          4327 => x"56",
          4328 => x"0d",
          4329 => x"8a",
          4330 => x"74",
          4331 => x"22",
          4332 => x"27",
          4333 => x"15",
          4334 => x"73",
          4335 => x"71",
          4336 => x"78",
          4337 => x"52",
          4338 => x"84",
          4339 => x"2e",
          4340 => x"08",
          4341 => x"53",
          4342 => x"91",
          4343 => x"27",
          4344 => x"84",
          4345 => x"f3",
          4346 => x"08",
          4347 => x"0a",
          4348 => x"18",
          4349 => x"74",
          4350 => x"06",
          4351 => x"18",
          4352 => x"85",
          4353 => x"76",
          4354 => x"0c",
          4355 => x"05",
          4356 => x"bb",
          4357 => x"98",
          4358 => x"7a",
          4359 => x"75",
          4360 => x"bb",
          4361 => x"84",
          4362 => x"56",
          4363 => x"38",
          4364 => x"26",
          4365 => x"98",
          4366 => x"f9",
          4367 => x"87",
          4368 => x"ff",
          4369 => x"08",
          4370 => x"84",
          4371 => x"38",
          4372 => x"5f",
          4373 => x"9c",
          4374 => x"5c",
          4375 => x"22",
          4376 => x"5d",
          4377 => x"58",
          4378 => x"70",
          4379 => x"74",
          4380 => x"55",
          4381 => x"54",
          4382 => x"33",
          4383 => x"08",
          4384 => x"39",
          4385 => x"bb",
          4386 => x"54",
          4387 => x"53",
          4388 => x"3f",
          4389 => x"84",
          4390 => x"19",
          4391 => x"a0",
          4392 => x"19",
          4393 => x"06",
          4394 => x"08",
          4395 => x"81",
          4396 => x"c5",
          4397 => x"ff",
          4398 => x"81",
          4399 => x"fe",
          4400 => x"56",
          4401 => x"38",
          4402 => x"1b",
          4403 => x"f8",
          4404 => x"8f",
          4405 => x"66",
          4406 => x"81",
          4407 => x"5e",
          4408 => x"19",
          4409 => x"08",
          4410 => x"33",
          4411 => x"81",
          4412 => x"53",
          4413 => x"e1",
          4414 => x"2e",
          4415 => x"b4",
          4416 => x"38",
          4417 => x"76",
          4418 => x"33",
          4419 => x"41",
          4420 => x"32",
          4421 => x"72",
          4422 => x"45",
          4423 => x"7a",
          4424 => x"81",
          4425 => x"38",
          4426 => x"fa",
          4427 => x"84",
          4428 => x"1c",
          4429 => x"84",
          4430 => x"81",
          4431 => x"81",
          4432 => x"57",
          4433 => x"81",
          4434 => x"08",
          4435 => x"1a",
          4436 => x"5b",
          4437 => x"38",
          4438 => x"09",
          4439 => x"b4",
          4440 => x"7e",
          4441 => x"3f",
          4442 => x"2e",
          4443 => x"86",
          4444 => x"93",
          4445 => x"06",
          4446 => x"0c",
          4447 => x"38",
          4448 => x"39",
          4449 => x"06",
          4450 => x"80",
          4451 => x"84",
          4452 => x"fd",
          4453 => x"77",
          4454 => x"19",
          4455 => x"71",
          4456 => x"ff",
          4457 => x"06",
          4458 => x"76",
          4459 => x"78",
          4460 => x"88",
          4461 => x"2e",
          4462 => x"ff",
          4463 => x"5c",
          4464 => x"81",
          4465 => x"77",
          4466 => x"57",
          4467 => x"fe",
          4468 => x"05",
          4469 => x"81",
          4470 => x"75",
          4471 => x"ff",
          4472 => x"7c",
          4473 => x"81",
          4474 => x"5a",
          4475 => x"06",
          4476 => x"38",
          4477 => x"0b",
          4478 => x"0c",
          4479 => x"63",
          4480 => x"51",
          4481 => x"5a",
          4482 => x"81",
          4483 => x"1d",
          4484 => x"56",
          4485 => x"82",
          4486 => x"55",
          4487 => x"df",
          4488 => x"52",
          4489 => x"84",
          4490 => x"ff",
          4491 => x"76",
          4492 => x"08",
          4493 => x"84",
          4494 => x"70",
          4495 => x"1d",
          4496 => x"38",
          4497 => x"8f",
          4498 => x"38",
          4499 => x"aa",
          4500 => x"74",
          4501 => x"78",
          4502 => x"05",
          4503 => x"56",
          4504 => x"80",
          4505 => x"57",
          4506 => x"59",
          4507 => x"78",
          4508 => x"31",
          4509 => x"80",
          4510 => x"e1",
          4511 => x"1d",
          4512 => x"3f",
          4513 => x"84",
          4514 => x"84",
          4515 => x"81",
          4516 => x"81",
          4517 => x"57",
          4518 => x"81",
          4519 => x"08",
          4520 => x"1c",
          4521 => x"59",
          4522 => x"38",
          4523 => x"09",
          4524 => x"b4",
          4525 => x"7d",
          4526 => x"3f",
          4527 => x"fd",
          4528 => x"2a",
          4529 => x"38",
          4530 => x"80",
          4531 => x"81",
          4532 => x"ac",
          4533 => x"2e",
          4534 => x"80",
          4535 => x"bb",
          4536 => x"80",
          4537 => x"75",
          4538 => x"5d",
          4539 => x"39",
          4540 => x"09",
          4541 => x"9b",
          4542 => x"2b",
          4543 => x"38",
          4544 => x"f3",
          4545 => x"83",
          4546 => x"11",
          4547 => x"52",
          4548 => x"38",
          4549 => x"76",
          4550 => x"84",
          4551 => x"53",
          4552 => x"bd",
          4553 => x"09",
          4554 => x"81",
          4555 => x"38",
          4556 => x"56",
          4557 => x"80",
          4558 => x"70",
          4559 => x"ff",
          4560 => x"fe",
          4561 => x"0c",
          4562 => x"ff",
          4563 => x"fe",
          4564 => x"08",
          4565 => x"58",
          4566 => x"b5",
          4567 => x"57",
          4568 => x"81",
          4569 => x"56",
          4570 => x"1f",
          4571 => x"55",
          4572 => x"70",
          4573 => x"74",
          4574 => x"70",
          4575 => x"82",
          4576 => x"34",
          4577 => x"1c",
          4578 => x"5a",
          4579 => x"33",
          4580 => x"15",
          4581 => x"80",
          4582 => x"74",
          4583 => x"5a",
          4584 => x"10",
          4585 => x"ff",
          4586 => x"58",
          4587 => x"76",
          4588 => x"58",
          4589 => x"55",
          4590 => x"80",
          4591 => x"bf",
          4592 => x"87",
          4593 => x"ff",
          4594 => x"76",
          4595 => x"79",
          4596 => x"27",
          4597 => x"2e",
          4598 => x"27",
          4599 => x"56",
          4600 => x"ea",
          4601 => x"87",
          4602 => x"ec",
          4603 => x"41",
          4604 => x"f4",
          4605 => x"bb",
          4606 => x"80",
          4607 => x"56",
          4608 => x"84",
          4609 => x"08",
          4610 => x"38",
          4611 => x"34",
          4612 => x"05",
          4613 => x"06",
          4614 => x"38",
          4615 => x"e8",
          4616 => x"80",
          4617 => x"bb",
          4618 => x"81",
          4619 => x"19",
          4620 => x"57",
          4621 => x"38",
          4622 => x"09",
          4623 => x"75",
          4624 => x"51",
          4625 => x"80",
          4626 => x"75",
          4627 => x"38",
          4628 => x"74",
          4629 => x"30",
          4630 => x"74",
          4631 => x"59",
          4632 => x"52",
          4633 => x"84",
          4634 => x"2e",
          4635 => x"2e",
          4636 => x"83",
          4637 => x"38",
          4638 => x"77",
          4639 => x"57",
          4640 => x"76",
          4641 => x"51",
          4642 => x"80",
          4643 => x"76",
          4644 => x"c3",
          4645 => x"55",
          4646 => x"ff",
          4647 => x"9c",
          4648 => x"70",
          4649 => x"05",
          4650 => x"38",
          4651 => x"06",
          4652 => x"0b",
          4653 => x"bb",
          4654 => x"75",
          4655 => x"40",
          4656 => x"81",
          4657 => x"bb",
          4658 => x"80",
          4659 => x"81",
          4660 => x"81",
          4661 => x"bb",
          4662 => x"83",
          4663 => x"19",
          4664 => x"31",
          4665 => x"38",
          4666 => x"84",
          4667 => x"fd",
          4668 => x"08",
          4669 => x"e9",
          4670 => x"bb",
          4671 => x"bb",
          4672 => x"81",
          4673 => x"70",
          4674 => x"70",
          4675 => x"5d",
          4676 => x"b8",
          4677 => x"80",
          4678 => x"38",
          4679 => x"09",
          4680 => x"76",
          4681 => x"51",
          4682 => x"80",
          4683 => x"76",
          4684 => x"83",
          4685 => x"61",
          4686 => x"8d",
          4687 => x"75",
          4688 => x"75",
          4689 => x"05",
          4690 => x"ff",
          4691 => x"70",
          4692 => x"e7",
          4693 => x"75",
          4694 => x"2a",
          4695 => x"83",
          4696 => x"78",
          4697 => x"2e",
          4698 => x"22",
          4699 => x"38",
          4700 => x"34",
          4701 => x"84",
          4702 => x"08",
          4703 => x"7f",
          4704 => x"54",
          4705 => x"53",
          4706 => x"3f",
          4707 => x"83",
          4708 => x"34",
          4709 => x"84",
          4710 => x"1d",
          4711 => x"33",
          4712 => x"fb",
          4713 => x"a0",
          4714 => x"1c",
          4715 => x"fb",
          4716 => x"33",
          4717 => x"09",
          4718 => x"39",
          4719 => x"fa",
          4720 => x"c0",
          4721 => x"b4",
          4722 => x"33",
          4723 => x"08",
          4724 => x"84",
          4725 => x"1c",
          4726 => x"a0",
          4727 => x"33",
          4728 => x"bb",
          4729 => x"ff",
          4730 => x"98",
          4731 => x"f7",
          4732 => x"80",
          4733 => x"81",
          4734 => x"05",
          4735 => x"ce",
          4736 => x"b4",
          4737 => x"7c",
          4738 => x"3f",
          4739 => x"61",
          4740 => x"96",
          4741 => x"82",
          4742 => x"80",
          4743 => x"05",
          4744 => x"58",
          4745 => x"74",
          4746 => x"56",
          4747 => x"14",
          4748 => x"76",
          4749 => x"79",
          4750 => x"55",
          4751 => x"80",
          4752 => x"5e",
          4753 => x"82",
          4754 => x"57",
          4755 => x"81",
          4756 => x"b2",
          4757 => x"75",
          4758 => x"80",
          4759 => x"90",
          4760 => x"77",
          4761 => x"58",
          4762 => x"81",
          4763 => x"38",
          4764 => x"81",
          4765 => x"a5",
          4766 => x"96",
          4767 => x"05",
          4768 => x"1c",
          4769 => x"89",
          4770 => x"08",
          4771 => x"9c",
          4772 => x"82",
          4773 => x"2b",
          4774 => x"88",
          4775 => x"59",
          4776 => x"88",
          4777 => x"56",
          4778 => x"15",
          4779 => x"07",
          4780 => x"3d",
          4781 => x"39",
          4782 => x"31",
          4783 => x"90",
          4784 => x"3f",
          4785 => x"06",
          4786 => x"81",
          4787 => x"2a",
          4788 => x"34",
          4789 => x"1f",
          4790 => x"70",
          4791 => x"38",
          4792 => x"70",
          4793 => x"07",
          4794 => x"74",
          4795 => x"0b",
          4796 => x"72",
          4797 => x"77",
          4798 => x"1e",
          4799 => x"ff",
          4800 => x"a4",
          4801 => x"54",
          4802 => x"84",
          4803 => x"80",
          4804 => x"ff",
          4805 => x"81",
          4806 => x"81",
          4807 => x"59",
          4808 => x"b4",
          4809 => x"80",
          4810 => x"73",
          4811 => x"39",
          4812 => x"42",
          4813 => x"55",
          4814 => x"53",
          4815 => x"72",
          4816 => x"08",
          4817 => x"94",
          4818 => x"82",
          4819 => x"58",
          4820 => x"52",
          4821 => x"72",
          4822 => x"38",
          4823 => x"76",
          4824 => x"17",
          4825 => x"af",
          4826 => x"80",
          4827 => x"82",
          4828 => x"89",
          4829 => x"83",
          4830 => x"70",
          4831 => x"80",
          4832 => x"8f",
          4833 => x"ff",
          4834 => x"72",
          4835 => x"38",
          4836 => x"76",
          4837 => x"17",
          4838 => x"56",
          4839 => x"38",
          4840 => x"32",
          4841 => x"51",
          4842 => x"38",
          4843 => x"33",
          4844 => x"72",
          4845 => x"25",
          4846 => x"38",
          4847 => x"3d",
          4848 => x"26",
          4849 => x"52",
          4850 => x"bb",
          4851 => x"73",
          4852 => x"bb",
          4853 => x"e6",
          4854 => x"53",
          4855 => x"39",
          4856 => x"52",
          4857 => x"84",
          4858 => x"0d",
          4859 => x"30",
          4860 => x"5a",
          4861 => x"14",
          4862 => x"56",
          4863 => x"dc",
          4864 => x"07",
          4865 => x"61",
          4866 => x"76",
          4867 => x"2e",
          4868 => x"80",
          4869 => x"fe",
          4870 => x"30",
          4871 => x"56",
          4872 => x"89",
          4873 => x"76",
          4874 => x"76",
          4875 => x"22",
          4876 => x"5d",
          4877 => x"38",
          4878 => x"ae",
          4879 => x"aa",
          4880 => x"5a",
          4881 => x"10",
          4882 => x"76",
          4883 => x"22",
          4884 => x"06",
          4885 => x"53",
          4886 => x"ff",
          4887 => x"5c",
          4888 => x"19",
          4889 => x"80",
          4890 => x"38",
          4891 => x"25",
          4892 => x"ce",
          4893 => x"7c",
          4894 => x"77",
          4895 => x"25",
          4896 => x"72",
          4897 => x"2e",
          4898 => x"38",
          4899 => x"9e",
          4900 => x"82",
          4901 => x"5f",
          4902 => x"58",
          4903 => x"1c",
          4904 => x"84",
          4905 => x"7d",
          4906 => x"ed",
          4907 => x"2e",
          4908 => x"06",
          4909 => x"5d",
          4910 => x"07",
          4911 => x"7d",
          4912 => x"5a",
          4913 => x"ec",
          4914 => x"33",
          4915 => x"2e",
          4916 => x"84",
          4917 => x"74",
          4918 => x"2e",
          4919 => x"06",
          4920 => x"65",
          4921 => x"58",
          4922 => x"70",
          4923 => x"56",
          4924 => x"80",
          4925 => x"5a",
          4926 => x"75",
          4927 => x"38",
          4928 => x"81",
          4929 => x"5b",
          4930 => x"56",
          4931 => x"38",
          4932 => x"57",
          4933 => x"e9",
          4934 => x"1d",
          4935 => x"bb",
          4936 => x"84",
          4937 => x"82",
          4938 => x"38",
          4939 => x"06",
          4940 => x"38",
          4941 => x"05",
          4942 => x"33",
          4943 => x"57",
          4944 => x"38",
          4945 => x"55",
          4946 => x"74",
          4947 => x"59",
          4948 => x"79",
          4949 => x"81",
          4950 => x"70",
          4951 => x"09",
          4952 => x"07",
          4953 => x"1d",
          4954 => x"fc",
          4955 => x"ab",
          4956 => x"0c",
          4957 => x"26",
          4958 => x"c9",
          4959 => x"81",
          4960 => x"18",
          4961 => x"82",
          4962 => x"81",
          4963 => x"83",
          4964 => x"06",
          4965 => x"74",
          4966 => x"33",
          4967 => x"b9",
          4968 => x"83",
          4969 => x"70",
          4970 => x"80",
          4971 => x"8f",
          4972 => x"ff",
          4973 => x"72",
          4974 => x"38",
          4975 => x"8a",
          4976 => x"06",
          4977 => x"99",
          4978 => x"81",
          4979 => x"ff",
          4980 => x"a0",
          4981 => x"5b",
          4982 => x"53",
          4983 => x"70",
          4984 => x"2e",
          4985 => x"07",
          4986 => x"74",
          4987 => x"80",
          4988 => x"71",
          4989 => x"07",
          4990 => x"39",
          4991 => x"54",
          4992 => x"11",
          4993 => x"81",
          4994 => x"07",
          4995 => x"e5",
          4996 => x"fd",
          4997 => x"5c",
          4998 => x"bb",
          4999 => x"3d",
          5000 => x"e7",
          5001 => x"0c",
          5002 => x"79",
          5003 => x"81",
          5004 => x"56",
          5005 => x"ed",
          5006 => x"84",
          5007 => x"85",
          5008 => x"cc",
          5009 => x"76",
          5010 => x"0c",
          5011 => x"59",
          5012 => x"33",
          5013 => x"84",
          5014 => x"5e",
          5015 => x"80",
          5016 => x"f8",
          5017 => x"81",
          5018 => x"84",
          5019 => x"81",
          5020 => x"c2",
          5021 => x"82",
          5022 => x"84",
          5023 => x"34",
          5024 => x"5a",
          5025 => x"70",
          5026 => x"bb",
          5027 => x"2e",
          5028 => x"b4",
          5029 => x"84",
          5030 => x"71",
          5031 => x"74",
          5032 => x"75",
          5033 => x"1d",
          5034 => x"58",
          5035 => x"58",
          5036 => x"c4",
          5037 => x"88",
          5038 => x"2e",
          5039 => x"cf",
          5040 => x"88",
          5041 => x"80",
          5042 => x"33",
          5043 => x"81",
          5044 => x"75",
          5045 => x"5e",
          5046 => x"c8",
          5047 => x"17",
          5048 => x"5f",
          5049 => x"82",
          5050 => x"71",
          5051 => x"5a",
          5052 => x"80",
          5053 => x"06",
          5054 => x"17",
          5055 => x"2b",
          5056 => x"74",
          5057 => x"7c",
          5058 => x"80",
          5059 => x"56",
          5060 => x"83",
          5061 => x"2b",
          5062 => x"70",
          5063 => x"07",
          5064 => x"80",
          5065 => x"71",
          5066 => x"7b",
          5067 => x"7a",
          5068 => x"81",
          5069 => x"51",
          5070 => x"08",
          5071 => x"81",
          5072 => x"ff",
          5073 => x"5d",
          5074 => x"82",
          5075 => x"38",
          5076 => x"0c",
          5077 => x"a8",
          5078 => x"57",
          5079 => x"88",
          5080 => x"2e",
          5081 => x"0c",
          5082 => x"38",
          5083 => x"81",
          5084 => x"89",
          5085 => x"08",
          5086 => x"0c",
          5087 => x"0b",
          5088 => x"96",
          5089 => x"22",
          5090 => x"23",
          5091 => x"0b",
          5092 => x"0c",
          5093 => x"97",
          5094 => x"84",
          5095 => x"d0",
          5096 => x"58",
          5097 => x"78",
          5098 => x"78",
          5099 => x"08",
          5100 => x"08",
          5101 => x"5c",
          5102 => x"ff",
          5103 => x"26",
          5104 => x"06",
          5105 => x"99",
          5106 => x"ff",
          5107 => x"2a",
          5108 => x"06",
          5109 => x"7a",
          5110 => x"2a",
          5111 => x"2e",
          5112 => x"5e",
          5113 => x"61",
          5114 => x"fe",
          5115 => x"5e",
          5116 => x"58",
          5117 => x"59",
          5118 => x"83",
          5119 => x"70",
          5120 => x"5b",
          5121 => x"e8",
          5122 => x"57",
          5123 => x"70",
          5124 => x"84",
          5125 => x"71",
          5126 => x"ff",
          5127 => x"83",
          5128 => x"5b",
          5129 => x"05",
          5130 => x"59",
          5131 => x"ba",
          5132 => x"2a",
          5133 => x"10",
          5134 => x"5d",
          5135 => x"83",
          5136 => x"80",
          5137 => x"18",
          5138 => x"2e",
          5139 => x"17",
          5140 => x"86",
          5141 => x"85",
          5142 => x"18",
          5143 => x"1f",
          5144 => x"5d",
          5145 => x"2e",
          5146 => x"b8",
          5147 => x"2e",
          5148 => x"70",
          5149 => x"42",
          5150 => x"2e",
          5151 => x"06",
          5152 => x"33",
          5153 => x"06",
          5154 => x"f8",
          5155 => x"38",
          5156 => x"7a",
          5157 => x"83",
          5158 => x"40",
          5159 => x"33",
          5160 => x"71",
          5161 => x"77",
          5162 => x"2e",
          5163 => x"83",
          5164 => x"81",
          5165 => x"40",
          5166 => x"58",
          5167 => x"38",
          5168 => x"fe",
          5169 => x"38",
          5170 => x"0d",
          5171 => x"dc",
          5172 => x"e6",
          5173 => x"8d",
          5174 => x"0d",
          5175 => x"e6",
          5176 => x"05",
          5177 => x"33",
          5178 => x"5f",
          5179 => x"74",
          5180 => x"8a",
          5181 => x"78",
          5182 => x"81",
          5183 => x"1b",
          5184 => x"84",
          5185 => x"93",
          5186 => x"83",
          5187 => x"e9",
          5188 => x"88",
          5189 => x"09",
          5190 => x"58",
          5191 => x"b1",
          5192 => x"2e",
          5193 => x"54",
          5194 => x"33",
          5195 => x"84",
          5196 => x"81",
          5197 => x"99",
          5198 => x"17",
          5199 => x"2b",
          5200 => x"2e",
          5201 => x"17",
          5202 => x"90",
          5203 => x"33",
          5204 => x"71",
          5205 => x"59",
          5206 => x"09",
          5207 => x"17",
          5208 => x"90",
          5209 => x"33",
          5210 => x"71",
          5211 => x"5e",
          5212 => x"09",
          5213 => x"17",
          5214 => x"90",
          5215 => x"33",
          5216 => x"71",
          5217 => x"1c",
          5218 => x"90",
          5219 => x"33",
          5220 => x"71",
          5221 => x"49",
          5222 => x"5a",
          5223 => x"81",
          5224 => x"7c",
          5225 => x"8c",
          5226 => x"f7",
          5227 => x"38",
          5228 => x"39",
          5229 => x"17",
          5230 => x"ff",
          5231 => x"7a",
          5232 => x"84",
          5233 => x"17",
          5234 => x"a0",
          5235 => x"33",
          5236 => x"84",
          5237 => x"74",
          5238 => x"85",
          5239 => x"5c",
          5240 => x"17",
          5241 => x"2b",
          5242 => x"d2",
          5243 => x"ca",
          5244 => x"82",
          5245 => x"2b",
          5246 => x"88",
          5247 => x"0c",
          5248 => x"40",
          5249 => x"75",
          5250 => x"f9",
          5251 => x"38",
          5252 => x"f7",
          5253 => x"38",
          5254 => x"08",
          5255 => x"81",
          5256 => x"fc",
          5257 => x"d3",
          5258 => x"41",
          5259 => x"80",
          5260 => x"05",
          5261 => x"74",
          5262 => x"38",
          5263 => x"e2",
          5264 => x"c4",
          5265 => x"05",
          5266 => x"84",
          5267 => x"80",
          5268 => x"54",
          5269 => x"2e",
          5270 => x"53",
          5271 => x"bb",
          5272 => x"0c",
          5273 => x"bb",
          5274 => x"33",
          5275 => x"56",
          5276 => x"16",
          5277 => x"58",
          5278 => x"7f",
          5279 => x"7b",
          5280 => x"05",
          5281 => x"33",
          5282 => x"99",
          5283 => x"ff",
          5284 => x"76",
          5285 => x"81",
          5286 => x"9f",
          5287 => x"81",
          5288 => x"77",
          5289 => x"9f",
          5290 => x"80",
          5291 => x"5d",
          5292 => x"7f",
          5293 => x"f7",
          5294 => x"8b",
          5295 => x"05",
          5296 => x"56",
          5297 => x"06",
          5298 => x"9e",
          5299 => x"3f",
          5300 => x"84",
          5301 => x"0c",
          5302 => x"9c",
          5303 => x"90",
          5304 => x"84",
          5305 => x"08",
          5306 => x"06",
          5307 => x"76",
          5308 => x"2e",
          5309 => x"76",
          5310 => x"06",
          5311 => x"66",
          5312 => x"88",
          5313 => x"5d",
          5314 => x"38",
          5315 => x"8f",
          5316 => x"80",
          5317 => x"a0",
          5318 => x"5e",
          5319 => x"9b",
          5320 => x"2e",
          5321 => x"9c",
          5322 => x"80",
          5323 => x"19",
          5324 => x"34",
          5325 => x"b4",
          5326 => x"5f",
          5327 => x"16",
          5328 => x"57",
          5329 => x"80",
          5330 => x"58",
          5331 => x"79",
          5332 => x"38",
          5333 => x"05",
          5334 => x"56",
          5335 => x"81",
          5336 => x"75",
          5337 => x"78",
          5338 => x"2e",
          5339 => x"7e",
          5340 => x"a4",
          5341 => x"12",
          5342 => x"40",
          5343 => x"81",
          5344 => x"16",
          5345 => x"90",
          5346 => x"33",
          5347 => x"71",
          5348 => x"7f",
          5349 => x"1b",
          5350 => x"34",
          5351 => x"9c",
          5352 => x"a8",
          5353 => x"80",
          5354 => x"15",
          5355 => x"81",
          5356 => x"38",
          5357 => x"fc",
          5358 => x"1b",
          5359 => x"77",
          5360 => x"78",
          5361 => x"27",
          5362 => x"5e",
          5363 => x"77",
          5364 => x"84",
          5365 => x"08",
          5366 => x"bb",
          5367 => x"79",
          5368 => x"05",
          5369 => x"78",
          5370 => x"2e",
          5371 => x"0c",
          5372 => x"0c",
          5373 => x"0c",
          5374 => x"57",
          5375 => x"94",
          5376 => x"2b",
          5377 => x"18",
          5378 => x"90",
          5379 => x"33",
          5380 => x"71",
          5381 => x"61",
          5382 => x"5c",
          5383 => x"90",
          5384 => x"80",
          5385 => x"1b",
          5386 => x"57",
          5387 => x"c2",
          5388 => x"07",
          5389 => x"83",
          5390 => x"e9",
          5391 => x"bb",
          5392 => x"84",
          5393 => x"38",
          5394 => x"b7",
          5395 => x"ff",
          5396 => x"83",
          5397 => x"94",
          5398 => x"27",
          5399 => x"84",
          5400 => x"17",
          5401 => x"a1",
          5402 => x"57",
          5403 => x"38",
          5404 => x"09",
          5405 => x"7d",
          5406 => x"51",
          5407 => x"08",
          5408 => x"5c",
          5409 => x"ff",
          5410 => x"2e",
          5411 => x"90",
          5412 => x"0b",
          5413 => x"16",
          5414 => x"71",
          5415 => x"58",
          5416 => x"8f",
          5417 => x"80",
          5418 => x"a0",
          5419 => x"5e",
          5420 => x"9b",
          5421 => x"2e",
          5422 => x"a9",
          5423 => x"ad",
          5424 => x"80",
          5425 => x"9c",
          5426 => x"77",
          5427 => x"22",
          5428 => x"56",
          5429 => x"75",
          5430 => x"58",
          5431 => x"19",
          5432 => x"bb",
          5433 => x"81",
          5434 => x"81",
          5435 => x"70",
          5436 => x"a2",
          5437 => x"2e",
          5438 => x"bb",
          5439 => x"08",
          5440 => x"08",
          5441 => x"fd",
          5442 => x"82",
          5443 => x"81",
          5444 => x"05",
          5445 => x"ff",
          5446 => x"39",
          5447 => x"0c",
          5448 => x"39",
          5449 => x"40",
          5450 => x"57",
          5451 => x"56",
          5452 => x"55",
          5453 => x"22",
          5454 => x"2e",
          5455 => x"76",
          5456 => x"33",
          5457 => x"33",
          5458 => x"2e",
          5459 => x"1a",
          5460 => x"26",
          5461 => x"b0",
          5462 => x"82",
          5463 => x"05",
          5464 => x"9b",
          5465 => x"08",
          5466 => x"74",
          5467 => x"1a",
          5468 => x"05",
          5469 => x"76",
          5470 => x"22",
          5471 => x"56",
          5472 => x"7b",
          5473 => x"80",
          5474 => x"75",
          5475 => x"5b",
          5476 => x"18",
          5477 => x"bb",
          5478 => x"33",
          5479 => x"24",
          5480 => x"79",
          5481 => x"77",
          5482 => x"94",
          5483 => x"38",
          5484 => x"90",
          5485 => x"0c",
          5486 => x"b3",
          5487 => x"2e",
          5488 => x"98",
          5489 => x"80",
          5490 => x"7a",
          5491 => x"8d",
          5492 => x"38",
          5493 => x"74",
          5494 => x"76",
          5495 => x"ff",
          5496 => x"81",
          5497 => x"19",
          5498 => x"80",
          5499 => x"83",
          5500 => x"a8",
          5501 => x"fe",
          5502 => x"33",
          5503 => x"16",
          5504 => x"74",
          5505 => x"81",
          5506 => x"da",
          5507 => x"52",
          5508 => x"bb",
          5509 => x"16",
          5510 => x"bb",
          5511 => x"bb",
          5512 => x"b5",
          5513 => x"75",
          5514 => x"76",
          5515 => x"55",
          5516 => x"70",
          5517 => x"74",
          5518 => x"81",
          5519 => x"59",
          5520 => x"fd",
          5521 => x"81",
          5522 => x"0d",
          5523 => x"0b",
          5524 => x"04",
          5525 => x"41",
          5526 => x"57",
          5527 => x"56",
          5528 => x"55",
          5529 => x"22",
          5530 => x"2e",
          5531 => x"76",
          5532 => x"33",
          5533 => x"33",
          5534 => x"87",
          5535 => x"94",
          5536 => x"77",
          5537 => x"80",
          5538 => x"06",
          5539 => x"11",
          5540 => x"5e",
          5541 => x"38",
          5542 => x"83",
          5543 => x"38",
          5544 => x"98",
          5545 => x"74",
          5546 => x"33",
          5547 => x"24",
          5548 => x"05",
          5549 => x"76",
          5550 => x"22",
          5551 => x"56",
          5552 => x"7c",
          5553 => x"80",
          5554 => x"75",
          5555 => x"5a",
          5556 => x"18",
          5557 => x"bb",
          5558 => x"08",
          5559 => x"38",
          5560 => x"29",
          5561 => x"81",
          5562 => x"59",
          5563 => x"90",
          5564 => x"90",
          5565 => x"78",
          5566 => x"1f",
          5567 => x"1e",
          5568 => x"5f",
          5569 => x"55",
          5570 => x"38",
          5571 => x"07",
          5572 => x"75",
          5573 => x"04",
          5574 => x"0d",
          5575 => x"38",
          5576 => x"08",
          5577 => x"a8",
          5578 => x"98",
          5579 => x"bd",
          5580 => x"1a",
          5581 => x"71",
          5582 => x"38",
          5583 => x"7f",
          5584 => x"38",
          5585 => x"70",
          5586 => x"75",
          5587 => x"07",
          5588 => x"39",
          5589 => x"ac",
          5590 => x"84",
          5591 => x"19",
          5592 => x"78",
          5593 => x"84",
          5594 => x"e2",
          5595 => x"08",
          5596 => x"51",
          5597 => x"08",
          5598 => x"06",
          5599 => x"fc",
          5600 => x"96",
          5601 => x"06",
          5602 => x"08",
          5603 => x"91",
          5604 => x"0c",
          5605 => x"1a",
          5606 => x"91",
          5607 => x"58",
          5608 => x"77",
          5609 => x"75",
          5610 => x"86",
          5611 => x"79",
          5612 => x"74",
          5613 => x"90",
          5614 => x"5c",
          5615 => x"76",
          5616 => x"c9",
          5617 => x"b4",
          5618 => x"0b",
          5619 => x"7a",
          5620 => x"38",
          5621 => x"81",
          5622 => x"84",
          5623 => x"ff",
          5624 => x"78",
          5625 => x"08",
          5626 => x"74",
          5627 => x"08",
          5628 => x"56",
          5629 => x"5a",
          5630 => x"33",
          5631 => x"2e",
          5632 => x"74",
          5633 => x"9d",
          5634 => x"9e",
          5635 => x"9f",
          5636 => x"97",
          5637 => x"80",
          5638 => x"92",
          5639 => x"7b",
          5640 => x"51",
          5641 => x"08",
          5642 => x"56",
          5643 => x"84",
          5644 => x"81",
          5645 => x"70",
          5646 => x"95",
          5647 => x"08",
          5648 => x"38",
          5649 => x"b4",
          5650 => x"bb",
          5651 => x"08",
          5652 => x"55",
          5653 => x"f8",
          5654 => x"17",
          5655 => x"33",
          5656 => x"fd",
          5657 => x"94",
          5658 => x"95",
          5659 => x"7b",
          5660 => x"18",
          5661 => x"18",
          5662 => x"18",
          5663 => x"18",
          5664 => x"cc",
          5665 => x"18",
          5666 => x"5b",
          5667 => x"ff",
          5668 => x"90",
          5669 => x"79",
          5670 => x"16",
          5671 => x"bb",
          5672 => x"9d",
          5673 => x"97",
          5674 => x"a8",
          5675 => x"57",
          5676 => x"bb",
          5677 => x"33",
          5678 => x"34",
          5679 => x"16",
          5680 => x"8e",
          5681 => x"79",
          5682 => x"bb",
          5683 => x"b1",
          5684 => x"38",
          5685 => x"38",
          5686 => x"38",
          5687 => x"52",
          5688 => x"71",
          5689 => x"75",
          5690 => x"3d",
          5691 => x"90",
          5692 => x"06",
          5693 => x"53",
          5694 => x"7d",
          5695 => x"b2",
          5696 => x"70",
          5697 => x"ac",
          5698 => x"a4",
          5699 => x"71",
          5700 => x"34",
          5701 => x"3d",
          5702 => x"0c",
          5703 => x"11",
          5704 => x"70",
          5705 => x"81",
          5706 => x"76",
          5707 => x"e6",
          5708 => x"57",
          5709 => x"70",
          5710 => x"53",
          5711 => x"e0",
          5712 => x"ff",
          5713 => x"38",
          5714 => x"54",
          5715 => x"71",
          5716 => x"73",
          5717 => x"30",
          5718 => x"59",
          5719 => x"81",
          5720 => x"25",
          5721 => x"39",
          5722 => x"5e",
          5723 => x"80",
          5724 => x"3d",
          5725 => x"08",
          5726 => x"8a",
          5727 => x"3d",
          5728 => x"3d",
          5729 => x"bb",
          5730 => x"80",
          5731 => x"70",
          5732 => x"80",
          5733 => x"84",
          5734 => x"2e",
          5735 => x"9a",
          5736 => x"33",
          5737 => x"2e",
          5738 => x"84",
          5739 => x"84",
          5740 => x"06",
          5741 => x"84",
          5742 => x"33",
          5743 => x"90",
          5744 => x"5b",
          5745 => x"0c",
          5746 => x"3d",
          5747 => x"e6",
          5748 => x"40",
          5749 => x"3d",
          5750 => x"51",
          5751 => x"59",
          5752 => x"60",
          5753 => x"11",
          5754 => x"db",
          5755 => x"82",
          5756 => x"40",
          5757 => x"e9",
          5758 => x"bb",
          5759 => x"df",
          5760 => x"77",
          5761 => x"83",
          5762 => x"38",
          5763 => x"81",
          5764 => x"84",
          5765 => x"ff",
          5766 => x"78",
          5767 => x"9b",
          5768 => x"2b",
          5769 => x"56",
          5770 => x"76",
          5771 => x"51",
          5772 => x"08",
          5773 => x"38",
          5774 => x"3f",
          5775 => x"84",
          5776 => x"9b",
          5777 => x"2b",
          5778 => x"5e",
          5779 => x"76",
          5780 => x"08",
          5781 => x"84",
          5782 => x"08",
          5783 => x"2e",
          5784 => x"80",
          5785 => x"51",
          5786 => x"05",
          5787 => x"38",
          5788 => x"70",
          5789 => x"81",
          5790 => x"38",
          5791 => x"82",
          5792 => x"08",
          5793 => x"56",
          5794 => x"38",
          5795 => x"5f",
          5796 => x"08",
          5797 => x"2e",
          5798 => x"e0",
          5799 => x"05",
          5800 => x"5e",
          5801 => x"1a",
          5802 => x"74",
          5803 => x"26",
          5804 => x"94",
          5805 => x"70",
          5806 => x"79",
          5807 => x"81",
          5808 => x"81",
          5809 => x"7c",
          5810 => x"e4",
          5811 => x"17",
          5812 => x"07",
          5813 => x"39",
          5814 => x"98",
          5815 => x"80",
          5816 => x"7a",
          5817 => x"84",
          5818 => x"2e",
          5819 => x"54",
          5820 => x"53",
          5821 => x"bd",
          5822 => x"fc",
          5823 => x"17",
          5824 => x"31",
          5825 => x"a0",
          5826 => x"16",
          5827 => x"06",
          5828 => x"08",
          5829 => x"81",
          5830 => x"7c",
          5831 => x"e6",
          5832 => x"34",
          5833 => x"10",
          5834 => x"70",
          5835 => x"7a",
          5836 => x"fd",
          5837 => x"81",
          5838 => x"81",
          5839 => x"8e",
          5840 => x"19",
          5841 => x"05",
          5842 => x"fd",
          5843 => x"78",
          5844 => x"0d",
          5845 => x"57",
          5846 => x"76",
          5847 => x"75",
          5848 => x"86",
          5849 => x"7a",
          5850 => x"74",
          5851 => x"91",
          5852 => x"8c",
          5853 => x"f2",
          5854 => x"78",
          5855 => x"11",
          5856 => x"75",
          5857 => x"ff",
          5858 => x"bb",
          5859 => x"53",
          5860 => x"bb",
          5861 => x"77",
          5862 => x"79",
          5863 => x"5b",
          5864 => x"79",
          5865 => x"94",
          5866 => x"18",
          5867 => x"5c",
          5868 => x"75",
          5869 => x"84",
          5870 => x"08",
          5871 => x"81",
          5872 => x"38",
          5873 => x"82",
          5874 => x"ae",
          5875 => x"17",
          5876 => x"ff",
          5877 => x"7b",
          5878 => x"5c",
          5879 => x"38",
          5880 => x"1a",
          5881 => x"5c",
          5882 => x"8c",
          5883 => x"77",
          5884 => x"0c",
          5885 => x"78",
          5886 => x"5b",
          5887 => x"17",
          5888 => x"38",
          5889 => x"19",
          5890 => x"38",
          5891 => x"81",
          5892 => x"3f",
          5893 => x"17",
          5894 => x"18",
          5895 => x"7b",
          5896 => x"e6",
          5897 => x"80",
          5898 => x"81",
          5899 => x"3d",
          5900 => x"2a",
          5901 => x"38",
          5902 => x"5a",
          5903 => x"fd",
          5904 => x"39",
          5905 => x"08",
          5906 => x"75",
          5907 => x"b7",
          5908 => x"0c",
          5909 => x"3d",
          5910 => x"8a",
          5911 => x"fd",
          5912 => x"83",
          5913 => x"06",
          5914 => x"08",
          5915 => x"76",
          5916 => x"84",
          5917 => x"2e",
          5918 => x"2e",
          5919 => x"88",
          5920 => x"93",
          5921 => x"0b",
          5922 => x"04",
          5923 => x"75",
          5924 => x"3d",
          5925 => x"51",
          5926 => x"55",
          5927 => x"38",
          5928 => x"bb",
          5929 => x"76",
          5930 => x"88",
          5931 => x"bb",
          5932 => x"33",
          5933 => x"24",
          5934 => x"2a",
          5935 => x"80",
          5936 => x"33",
          5937 => x"7d",
          5938 => x"78",
          5939 => x"0c",
          5940 => x"23",
          5941 => x"3f",
          5942 => x"2e",
          5943 => x"38",
          5944 => x"55",
          5945 => x"17",
          5946 => x"71",
          5947 => x"0c",
          5948 => x"0d",
          5949 => x"9e",
          5950 => x"96",
          5951 => x"8e",
          5952 => x"57",
          5953 => x"52",
          5954 => x"0c",
          5955 => x"0d",
          5956 => x"b4",
          5957 => x"52",
          5958 => x"54",
          5959 => x"58",
          5960 => x"38",
          5961 => x"38",
          5962 => x"38",
          5963 => x"53",
          5964 => x"53",
          5965 => x"38",
          5966 => x"52",
          5967 => x"bb",
          5968 => x"84",
          5969 => x"a6",
          5970 => x"83",
          5971 => x"af",
          5972 => x"70",
          5973 => x"bb",
          5974 => x"84",
          5975 => x"75",
          5976 => x"d3",
          5977 => x"ff",
          5978 => x"70",
          5979 => x"bb",
          5980 => x"39",
          5981 => x"3f",
          5982 => x"0c",
          5983 => x"51",
          5984 => x"08",
          5985 => x"72",
          5986 => x"ed",
          5987 => x"3d",
          5988 => x"96",
          5989 => x"bb",
          5990 => x"84",
          5991 => x"65",
          5992 => x"84",
          5993 => x"08",
          5994 => x"70",
          5995 => x"97",
          5996 => x"52",
          5997 => x"84",
          5998 => x"86",
          5999 => x"0d",
          6000 => x"5f",
          6001 => x"96",
          6002 => x"84",
          6003 => x"38",
          6004 => x"08",
          6005 => x"59",
          6006 => x"7f",
          6007 => x"3d",
          6008 => x"33",
          6009 => x"38",
          6010 => x"08",
          6011 => x"7b",
          6012 => x"17",
          6013 => x"17",
          6014 => x"38",
          6015 => x"81",
          6016 => x"84",
          6017 => x"ff",
          6018 => x"7f",
          6019 => x"76",
          6020 => x"38",
          6021 => x"82",
          6022 => x"2b",
          6023 => x"88",
          6024 => x"fe",
          6025 => x"25",
          6026 => x"06",
          6027 => x"54",
          6028 => x"fe",
          6029 => x"18",
          6030 => x"77",
          6031 => x"0c",
          6032 => x"17",
          6033 => x"18",
          6034 => x"81",
          6035 => x"38",
          6036 => x"b4",
          6037 => x"bb",
          6038 => x"08",
          6039 => x"55",
          6040 => x"b0",
          6041 => x"18",
          6042 => x"33",
          6043 => x"fe",
          6044 => x"59",
          6045 => x"f1",
          6046 => x"80",
          6047 => x"2e",
          6048 => x"30",
          6049 => x"25",
          6050 => x"5c",
          6051 => x"38",
          6052 => x"84",
          6053 => x"18",
          6054 => x"05",
          6055 => x"2b",
          6056 => x"82",
          6057 => x"5d",
          6058 => x"83",
          6059 => x"bf",
          6060 => x"0c",
          6061 => x"81",
          6062 => x"83",
          6063 => x"f6",
          6064 => x"80",
          6065 => x"80",
          6066 => x"80",
          6067 => x"19",
          6068 => x"81",
          6069 => x"83",
          6070 => x"fb",
          6071 => x"81",
          6072 => x"2e",
          6073 => x"74",
          6074 => x"74",
          6075 => x"08",
          6076 => x"9c",
          6077 => x"82",
          6078 => x"18",
          6079 => x"07",
          6080 => x"38",
          6081 => x"a3",
          6082 => x"a8",
          6083 => x"59",
          6084 => x"08",
          6085 => x"76",
          6086 => x"bb",
          6087 => x"55",
          6088 => x"52",
          6089 => x"bb",
          6090 => x"80",
          6091 => x"08",
          6092 => x"84",
          6093 => x"53",
          6094 => x"3f",
          6095 => x"9c",
          6096 => x"58",
          6097 => x"38",
          6098 => x"33",
          6099 => x"79",
          6100 => x"9c",
          6101 => x"ac",
          6102 => x"55",
          6103 => x"56",
          6104 => x"19",
          6105 => x"88",
          6106 => x"08",
          6107 => x"84",
          6108 => x"38",
          6109 => x"be",
          6110 => x"84",
          6111 => x"81",
          6112 => x"19",
          6113 => x"0b",
          6114 => x"38",
          6115 => x"27",
          6116 => x"38",
          6117 => x"84",
          6118 => x"84",
          6119 => x"52",
          6120 => x"bb",
          6121 => x"80",
          6122 => x"08",
          6123 => x"84",
          6124 => x"53",
          6125 => x"3f",
          6126 => x"9c",
          6127 => x"58",
          6128 => x"81",
          6129 => x"81",
          6130 => x"55",
          6131 => x"56",
          6132 => x"ce",
          6133 => x"0b",
          6134 => x"39",
          6135 => x"80",
          6136 => x"76",
          6137 => x"19",
          6138 => x"bb",
          6139 => x"fd",
          6140 => x"5a",
          6141 => x"08",
          6142 => x"aa",
          6143 => x"3d",
          6144 => x"ff",
          6145 => x"56",
          6146 => x"38",
          6147 => x"0d",
          6148 => x"9b",
          6149 => x"3f",
          6150 => x"84",
          6151 => x"33",
          6152 => x"86",
          6153 => x"5b",
          6154 => x"ee",
          6155 => x"87",
          6156 => x"3d",
          6157 => x"71",
          6158 => x"5c",
          6159 => x"38",
          6160 => x"80",
          6161 => x"18",
          6162 => x"5f",
          6163 => x"8f",
          6164 => x"3f",
          6165 => x"84",
          6166 => x"08",
          6167 => x"84",
          6168 => x"08",
          6169 => x"0c",
          6170 => x"94",
          6171 => x"2b",
          6172 => x"98",
          6173 => x"88",
          6174 => x"38",
          6175 => x"5d",
          6176 => x"74",
          6177 => x"84",
          6178 => x"08",
          6179 => x"77",
          6180 => x"2e",
          6181 => x"7a",
          6182 => x"89",
          6183 => x"fd",
          6184 => x"7d",
          6185 => x"84",
          6186 => x"0d",
          6187 => x"56",
          6188 => x"82",
          6189 => x"55",
          6190 => x"dd",
          6191 => x"52",
          6192 => x"3f",
          6193 => x"38",
          6194 => x"0c",
          6195 => x"08",
          6196 => x"18",
          6197 => x"ec",
          6198 => x"97",
          6199 => x"bb",
          6200 => x"75",
          6201 => x"38",
          6202 => x"b4",
          6203 => x"33",
          6204 => x"84",
          6205 => x"06",
          6206 => x"83",
          6207 => x"08",
          6208 => x"74",
          6209 => x"82",
          6210 => x"81",
          6211 => x"17",
          6212 => x"52",
          6213 => x"3f",
          6214 => x"79",
          6215 => x"78",
          6216 => x"84",
          6217 => x"2e",
          6218 => x"81",
          6219 => x"08",
          6220 => x"74",
          6221 => x"84",
          6222 => x"08",
          6223 => x"58",
          6224 => x"16",
          6225 => x"07",
          6226 => x"77",
          6227 => x"fd",
          6228 => x"84",
          6229 => x"81",
          6230 => x"82",
          6231 => x"a0",
          6232 => x"bb",
          6233 => x"80",
          6234 => x"0c",
          6235 => x"52",
          6236 => x"f8",
          6237 => x"bb",
          6238 => x"bb",
          6239 => x"bb",
          6240 => x"cb",
          6241 => x"85",
          6242 => x"74",
          6243 => x"8f",
          6244 => x"3f",
          6245 => x"84",
          6246 => x"84",
          6247 => x"38",
          6248 => x"cb",
          6249 => x"bb",
          6250 => x"57",
          6251 => x"18",
          6252 => x"75",
          6253 => x"76",
          6254 => x"58",
          6255 => x"84",
          6256 => x"81",
          6257 => x"f4",
          6258 => x"77",
          6259 => x"77",
          6260 => x"51",
          6261 => x"08",
          6262 => x"39",
          6263 => x"b4",
          6264 => x"81",
          6265 => x"3f",
          6266 => x"38",
          6267 => x"b4",
          6268 => x"74",
          6269 => x"82",
          6270 => x"81",
          6271 => x"17",
          6272 => x"52",
          6273 => x"3f",
          6274 => x"08",
          6275 => x"38",
          6276 => x"38",
          6277 => x"3f",
          6278 => x"84",
          6279 => x"bb",
          6280 => x"84",
          6281 => x"38",
          6282 => x"f9",
          6283 => x"f3",
          6284 => x"19",
          6285 => x"90",
          6286 => x"17",
          6287 => x"34",
          6288 => x"38",
          6289 => x"0d",
          6290 => x"ff",
          6291 => x"2e",
          6292 => x"0b",
          6293 => x"81",
          6294 => x"f4",
          6295 => x"34",
          6296 => x"34",
          6297 => x"75",
          6298 => x"d0",
          6299 => x"1a",
          6300 => x"59",
          6301 => x"88",
          6302 => x"75",
          6303 => x"38",
          6304 => x"b8",
          6305 => x"05",
          6306 => x"34",
          6307 => x"56",
          6308 => x"7e",
          6309 => x"57",
          6310 => x"2a",
          6311 => x"33",
          6312 => x"7d",
          6313 => x"51",
          6314 => x"08",
          6315 => x"38",
          6316 => x"17",
          6317 => x"34",
          6318 => x"0b",
          6319 => x"77",
          6320 => x"78",
          6321 => x"83",
          6322 => x"0b",
          6323 => x"83",
          6324 => x"3f",
          6325 => x"bb",
          6326 => x"90",
          6327 => x"74",
          6328 => x"34",
          6329 => x"7a",
          6330 => x"55",
          6331 => x"a0",
          6332 => x"58",
          6333 => x"58",
          6334 => x"5c",
          6335 => x"0b",
          6336 => x"83",
          6337 => x"3f",
          6338 => x"39",
          6339 => x"08",
          6340 => x"9b",
          6341 => x"70",
          6342 => x"81",
          6343 => x"2e",
          6344 => x"fe",
          6345 => x"ab",
          6346 => x"84",
          6347 => x"75",
          6348 => x"04",
          6349 => x"52",
          6350 => x"e8",
          6351 => x"bb",
          6352 => x"05",
          6353 => x"7c",
          6354 => x"3d",
          6355 => x"05",
          6356 => x"34",
          6357 => x"3d",
          6358 => x"75",
          6359 => x"81",
          6360 => x"ef",
          6361 => x"ff",
          6362 => x"56",
          6363 => x"6a",
          6364 => x"88",
          6365 => x"0d",
          6366 => x"ff",
          6367 => x"91",
          6368 => x"d0",
          6369 => x"fa",
          6370 => x"70",
          6371 => x"7a",
          6372 => x"81",
          6373 => x"58",
          6374 => x"16",
          6375 => x"9f",
          6376 => x"e0",
          6377 => x"75",
          6378 => x"77",
          6379 => x"ff",
          6380 => x"70",
          6381 => x"58",
          6382 => x"1c",
          6383 => x"fd",
          6384 => x"ff",
          6385 => x"38",
          6386 => x"fe",
          6387 => x"a9",
          6388 => x"84",
          6389 => x"b8",
          6390 => x"81",
          6391 => x"8d",
          6392 => x"84",
          6393 => x"58",
          6394 => x"80",
          6395 => x"81",
          6396 => x"57",
          6397 => x"02",
          6398 => x"8b",
          6399 => x"40",
          6400 => x"57",
          6401 => x"0b",
          6402 => x"84",
          6403 => x"2e",
          6404 => x"2e",
          6405 => x"9a",
          6406 => x"33",
          6407 => x"82",
          6408 => x"fe",
          6409 => x"c7",
          6410 => x"b0",
          6411 => x"2e",
          6412 => x"b4",
          6413 => x"17",
          6414 => x"54",
          6415 => x"33",
          6416 => x"84",
          6417 => x"81",
          6418 => x"7b",
          6419 => x"bf",
          6420 => x"2e",
          6421 => x"83",
          6422 => x"f2",
          6423 => x"80",
          6424 => x"83",
          6425 => x"90",
          6426 => x"7d",
          6427 => x"34",
          6428 => x"78",
          6429 => x"57",
          6430 => x"74",
          6431 => x"84",
          6432 => x"08",
          6433 => x"19",
          6434 => x"77",
          6435 => x"59",
          6436 => x"81",
          6437 => x"16",
          6438 => x"f6",
          6439 => x"85",
          6440 => x"17",
          6441 => x"19",
          6442 => x"83",
          6443 => x"a5",
          6444 => x"e7",
          6445 => x"bb",
          6446 => x"82",
          6447 => x"74",
          6448 => x"fe",
          6449 => x"84",
          6450 => x"82",
          6451 => x"0d",
          6452 => x"71",
          6453 => x"07",
          6454 => x"bb",
          6455 => x"84",
          6456 => x"38",
          6457 => x"0d",
          6458 => x"7b",
          6459 => x"cd",
          6460 => x"7a",
          6461 => x"84",
          6462 => x"16",
          6463 => x"84",
          6464 => x"27",
          6465 => x"7c",
          6466 => x"38",
          6467 => x"08",
          6468 => x"51",
          6469 => x"fa",
          6470 => x"b8",
          6471 => x"5b",
          6472 => x"bb",
          6473 => x"84",
          6474 => x"a8",
          6475 => x"5d",
          6476 => x"8e",
          6477 => x"2e",
          6478 => x"54",
          6479 => x"53",
          6480 => x"e1",
          6481 => x"ec",
          6482 => x"02",
          6483 => x"57",
          6484 => x"97",
          6485 => x"bb",
          6486 => x"80",
          6487 => x"0c",
          6488 => x"52",
          6489 => x"90",
          6490 => x"bb",
          6491 => x"05",
          6492 => x"73",
          6493 => x"09",
          6494 => x"06",
          6495 => x"17",
          6496 => x"34",
          6497 => x"bb",
          6498 => x"3d",
          6499 => x"82",
          6500 => x"3d",
          6501 => x"84",
          6502 => x"2e",
          6503 => x"96",
          6504 => x"96",
          6505 => x"3f",
          6506 => x"84",
          6507 => x"33",
          6508 => x"d2",
          6509 => x"22",
          6510 => x"76",
          6511 => x"74",
          6512 => x"77",
          6513 => x"73",
          6514 => x"83",
          6515 => x"3f",
          6516 => x"0c",
          6517 => x"6b",
          6518 => x"cc",
          6519 => x"fe",
          6520 => x"84",
          6521 => x"07",
          6522 => x"2e",
          6523 => x"56",
          6524 => x"78",
          6525 => x"2e",
          6526 => x"5a",
          6527 => x"7c",
          6528 => x"b4",
          6529 => x"83",
          6530 => x"2e",
          6531 => x"54",
          6532 => x"33",
          6533 => x"84",
          6534 => x"81",
          6535 => x"78",
          6536 => x"80",
          6537 => x"80",
          6538 => x"a7",
          6539 => x"33",
          6540 => x"88",
          6541 => x"07",
          6542 => x"0c",
          6543 => x"84",
          6544 => x"7c",
          6545 => x"70",
          6546 => x"bb",
          6547 => x"80",
          6548 => x"09",
          6549 => x"34",
          6550 => x"b4",
          6551 => x"81",
          6552 => x"3f",
          6553 => x"2e",
          6554 => x"bb",
          6555 => x"08",
          6556 => x"08",
          6557 => x"fe",
          6558 => x"82",
          6559 => x"77",
          6560 => x"05",
          6561 => x"fe",
          6562 => x"76",
          6563 => x"51",
          6564 => x"08",
          6565 => x"39",
          6566 => x"3f",
          6567 => x"84",
          6568 => x"08",
          6569 => x"59",
          6570 => x"59",
          6571 => x"59",
          6572 => x"1c",
          6573 => x"2e",
          6574 => x"70",
          6575 => x"ea",
          6576 => x"ba",
          6577 => x"3d",
          6578 => x"ff",
          6579 => x"56",
          6580 => x"8f",
          6581 => x"76",
          6582 => x"55",
          6583 => x"70",
          6584 => x"58",
          6585 => x"a2",
          6586 => x"ff",
          6587 => x"f5",
          6588 => x"ff",
          6589 => x"95",
          6590 => x"08",
          6591 => x"08",
          6592 => x"2e",
          6593 => x"83",
          6594 => x"5b",
          6595 => x"38",
          6596 => x"81",
          6597 => x"57",
          6598 => x"74",
          6599 => x"75",
          6600 => x"38",
          6601 => x"79",
          6602 => x"77",
          6603 => x"74",
          6604 => x"1a",
          6605 => x"34",
          6606 => x"70",
          6607 => x"77",
          6608 => x"33",
          6609 => x"bc",
          6610 => x"b7",
          6611 => x"5c",
          6612 => x"38",
          6613 => x"45",
          6614 => x"52",
          6615 => x"84",
          6616 => x"2e",
          6617 => x"84",
          6618 => x"52",
          6619 => x"84",
          6620 => x"fd",
          6621 => x"84",
          6622 => x"94",
          6623 => x"75",
          6624 => x"84",
          6625 => x"c1",
          6626 => x"8b",
          6627 => x"81",
          6628 => x"58",
          6629 => x"7d",
          6630 => x"51",
          6631 => x"08",
          6632 => x"7a",
          6633 => x"9c",
          6634 => x"09",
          6635 => x"79",
          6636 => x"75",
          6637 => x"3f",
          6638 => x"84",
          6639 => x"84",
          6640 => x"5c",
          6641 => x"b4",
          6642 => x"18",
          6643 => x"06",
          6644 => x"b8",
          6645 => x"d5",
          6646 => x"2e",
          6647 => x"b4",
          6648 => x"78",
          6649 => x"57",
          6650 => x"74",
          6651 => x"5c",
          6652 => x"1a",
          6653 => x"52",
          6654 => x"bb",
          6655 => x"80",
          6656 => x"84",
          6657 => x"fd",
          6658 => x"76",
          6659 => x"55",
          6660 => x"8b",
          6661 => x"55",
          6662 => x"70",
          6663 => x"74",
          6664 => x"81",
          6665 => x"58",
          6666 => x"fd",
          6667 => x"7d",
          6668 => x"51",
          6669 => x"08",
          6670 => x"df",
          6671 => x"7a",
          6672 => x"a5",
          6673 => x"09",
          6674 => x"84",
          6675 => x"a8",
          6676 => x"08",
          6677 => x"74",
          6678 => x"08",
          6679 => x"52",
          6680 => x"bb",
          6681 => x"80",
          6682 => x"81",
          6683 => x"e7",
          6684 => x"18",
          6685 => x"52",
          6686 => x"3f",
          6687 => x"62",
          6688 => x"5e",
          6689 => x"9f",
          6690 => x"97",
          6691 => x"8f",
          6692 => x"59",
          6693 => x"80",
          6694 => x"91",
          6695 => x"79",
          6696 => x"08",
          6697 => x"81",
          6698 => x"2e",
          6699 => x"70",
          6700 => x"5c",
          6701 => x"7a",
          6702 => x"2a",
          6703 => x"08",
          6704 => x"78",
          6705 => x"26",
          6706 => x"5b",
          6707 => x"d8",
          6708 => x"9c",
          6709 => x"55",
          6710 => x"dc",
          6711 => x"81",
          6712 => x"c5",
          6713 => x"bb",
          6714 => x"c2",
          6715 => x"bb",
          6716 => x"0b",
          6717 => x"04",
          6718 => x"3f",
          6719 => x"73",
          6720 => x"56",
          6721 => x"8e",
          6722 => x"2e",
          6723 => x"2e",
          6724 => x"7e",
          6725 => x"84",
          6726 => x"a3",
          6727 => x"59",
          6728 => x"12",
          6729 => x"38",
          6730 => x"0c",
          6731 => x"7b",
          6732 => x"05",
          6733 => x"26",
          6734 => x"16",
          6735 => x"7c",
          6736 => x"39",
          6737 => x"80",
          6738 => x"c5",
          6739 => x"1b",
          6740 => x"08",
          6741 => x"3d",
          6742 => x"33",
          6743 => x"08",
          6744 => x"85",
          6745 => x"33",
          6746 => x"2e",
          6747 => x"ba",
          6748 => x"33",
          6749 => x"75",
          6750 => x"08",
          6751 => x"80",
          6752 => x"11",
          6753 => x"5b",
          6754 => x"e2",
          6755 => x"06",
          6756 => x"7b",
          6757 => x"06",
          6758 => x"9f",
          6759 => x"51",
          6760 => x"08",
          6761 => x"2e",
          6762 => x"26",
          6763 => x"55",
          6764 => x"88",
          6765 => x"38",
          6766 => x"38",
          6767 => x"e7",
          6768 => x"89",
          6769 => x"47",
          6770 => x"65",
          6771 => x"5f",
          6772 => x"80",
          6773 => x"53",
          6774 => x"3f",
          6775 => x"95",
          6776 => x"83",
          6777 => x"59",
          6778 => x"2e",
          6779 => x"90",
          6780 => x"44",
          6781 => x"83",
          6782 => x"33",
          6783 => x"81",
          6784 => x"75",
          6785 => x"11",
          6786 => x"71",
          6787 => x"72",
          6788 => x"5c",
          6789 => x"a3",
          6790 => x"4f",
          6791 => x"80",
          6792 => x"57",
          6793 => x"61",
          6794 => x"63",
          6795 => x"06",
          6796 => x"81",
          6797 => x"6e",
          6798 => x"62",
          6799 => x"38",
          6800 => x"e8",
          6801 => x"9d",
          6802 => x"e8",
          6803 => x"22",
          6804 => x"38",
          6805 => x"78",
          6806 => x"84",
          6807 => x"84",
          6808 => x"0b",
          6809 => x"84",
          6810 => x"05",
          6811 => x"2a",
          6812 => x"7d",
          6813 => x"70",
          6814 => x"44",
          6815 => x"1d",
          6816 => x"31",
          6817 => x"38",
          6818 => x"70",
          6819 => x"3f",
          6820 => x"2e",
          6821 => x"81",
          6822 => x"0b",
          6823 => x"38",
          6824 => x"74",
          6825 => x"5b",
          6826 => x"bb",
          6827 => x"90",
          6828 => x"93",
          6829 => x"0d",
          6830 => x"d0",
          6831 => x"57",
          6832 => x"77",
          6833 => x"77",
          6834 => x"83",
          6835 => x"57",
          6836 => x"76",
          6837 => x"12",
          6838 => x"38",
          6839 => x"44",
          6840 => x"89",
          6841 => x"59",
          6842 => x"47",
          6843 => x"38",
          6844 => x"70",
          6845 => x"07",
          6846 => x"ce",
          6847 => x"83",
          6848 => x"f9",
          6849 => x"81",
          6850 => x"81",
          6851 => x"38",
          6852 => x"84",
          6853 => x"5f",
          6854 => x"fe",
          6855 => x"fb",
          6856 => x"83",
          6857 => x"3d",
          6858 => x"06",
          6859 => x"f5",
          6860 => x"43",
          6861 => x"9f",
          6862 => x"77",
          6863 => x"f5",
          6864 => x"0c",
          6865 => x"04",
          6866 => x"38",
          6867 => x"81",
          6868 => x"38",
          6869 => x"70",
          6870 => x"74",
          6871 => x"59",
          6872 => x"33",
          6873 => x"15",
          6874 => x"45",
          6875 => x"34",
          6876 => x"ff",
          6877 => x"34",
          6878 => x"05",
          6879 => x"83",
          6880 => x"91",
          6881 => x"49",
          6882 => x"75",
          6883 => x"75",
          6884 => x"93",
          6885 => x"61",
          6886 => x"34",
          6887 => x"99",
          6888 => x"80",
          6889 => x"05",
          6890 => x"9d",
          6891 => x"61",
          6892 => x"bb",
          6893 => x"9f",
          6894 => x"38",
          6895 => x"a8",
          6896 => x"80",
          6897 => x"ff",
          6898 => x"34",
          6899 => x"05",
          6900 => x"a9",
          6901 => x"05",
          6902 => x"70",
          6903 => x"05",
          6904 => x"38",
          6905 => x"69",
          6906 => x"aa",
          6907 => x"52",
          6908 => x"57",
          6909 => x"60",
          6910 => x"38",
          6911 => x"81",
          6912 => x"f4",
          6913 => x"2e",
          6914 => x"57",
          6915 => x"76",
          6916 => x"55",
          6917 => x"76",
          6918 => x"05",
          6919 => x"64",
          6920 => x"26",
          6921 => x"53",
          6922 => x"3f",
          6923 => x"84",
          6924 => x"81",
          6925 => x"f4",
          6926 => x"5b",
          6927 => x"7f",
          6928 => x"62",
          6929 => x"55",
          6930 => x"74",
          6931 => x"fe",
          6932 => x"85",
          6933 => x"57",
          6934 => x"83",
          6935 => x"ff",
          6936 => x"82",
          6937 => x"c1",
          6938 => x"7d",
          6939 => x"59",
          6940 => x"ff",
          6941 => x"69",
          6942 => x"be",
          6943 => x"81",
          6944 => x"78",
          6945 => x"05",
          6946 => x"62",
          6947 => x"67",
          6948 => x"82",
          6949 => x"05",
          6950 => x"05",
          6951 => x"67",
          6952 => x"83",
          6953 => x"61",
          6954 => x"ca",
          6955 => x"61",
          6956 => x"58",
          6957 => x"98",
          6958 => x"34",
          6959 => x"51",
          6960 => x"bb",
          6961 => x"80",
          6962 => x"81",
          6963 => x"38",
          6964 => x"0c",
          6965 => x"04",
          6966 => x"64",
          6967 => x"ae",
          6968 => x"83",
          6969 => x"2e",
          6970 => x"83",
          6971 => x"70",
          6972 => x"86",
          6973 => x"52",
          6974 => x"bb",
          6975 => x"70",
          6976 => x"0b",
          6977 => x"05",
          6978 => x"27",
          6979 => x"39",
          6980 => x"26",
          6981 => x"77",
          6982 => x"8e",
          6983 => x"44",
          6984 => x"43",
          6985 => x"34",
          6986 => x"05",
          6987 => x"a2",
          6988 => x"61",
          6989 => x"61",
          6990 => x"c4",
          6991 => x"34",
          6992 => x"7c",
          6993 => x"5c",
          6994 => x"2a",
          6995 => x"98",
          6996 => x"82",
          6997 => x"05",
          6998 => x"61",
          6999 => x"34",
          7000 => x"b2",
          7001 => x"ff",
          7002 => x"61",
          7003 => x"c7",
          7004 => x"76",
          7005 => x"81",
          7006 => x"80",
          7007 => x"05",
          7008 => x"34",
          7009 => x"b8",
          7010 => x"79",
          7011 => x"84",
          7012 => x"90",
          7013 => x"b2",
          7014 => x"08",
          7015 => x"ed",
          7016 => x"bb",
          7017 => x"90",
          7018 => x"ff",
          7019 => x"6a",
          7020 => x"34",
          7021 => x"85",
          7022 => x"ff",
          7023 => x"05",
          7024 => x"61",
          7025 => x"57",
          7026 => x"53",
          7027 => x"3f",
          7028 => x"70",
          7029 => x"76",
          7030 => x"70",
          7031 => x"d2",
          7032 => x"e1",
          7033 => x"c1",
          7034 => x"05",
          7035 => x"34",
          7036 => x"80",
          7037 => x"ff",
          7038 => x"34",
          7039 => x"e9",
          7040 => x"61",
          7041 => x"40",
          7042 => x"61",
          7043 => x"ed",
          7044 => x"34",
          7045 => x"d5",
          7046 => x"54",
          7047 => x"fe",
          7048 => x"53",
          7049 => x"3f",
          7050 => x"f4",
          7051 => x"7b",
          7052 => x"78",
          7053 => x"3d",
          7054 => x"79",
          7055 => x"2e",
          7056 => x"33",
          7057 => x"76",
          7058 => x"57",
          7059 => x"24",
          7060 => x"76",
          7061 => x"84",
          7062 => x"0d",
          7063 => x"59",
          7064 => x"84",
          7065 => x"38",
          7066 => x"56",
          7067 => x"74",
          7068 => x"0c",
          7069 => x"0d",
          7070 => x"53",
          7071 => x"9f",
          7072 => x"70",
          7073 => x"1b",
          7074 => x"56",
          7075 => x"ff",
          7076 => x"0d",
          7077 => x"58",
          7078 => x"76",
          7079 => x"55",
          7080 => x"0c",
          7081 => x"56",
          7082 => x"77",
          7083 => x"34",
          7084 => x"38",
          7085 => x"18",
          7086 => x"38",
          7087 => x"54",
          7088 => x"9e",
          7089 => x"38",
          7090 => x"84",
          7091 => x"9f",
          7092 => x"c0",
          7093 => x"f8",
          7094 => x"72",
          7095 => x"56",
          7096 => x"51",
          7097 => x"84",
          7098 => x"fd",
          7099 => x"05",
          7100 => x"ff",
          7101 => x"06",
          7102 => x"3d",
          7103 => x"54",
          7104 => x"e9",
          7105 => x"e8",
          7106 => x"38",
          7107 => x"53",
          7108 => x"71",
          7109 => x"51",
          7110 => x"81",
          7111 => x"85",
          7112 => x"92",
          7113 => x"22",
          7114 => x"26",
          7115 => x"84",
          7116 => x"b5",
          7117 => x"81",
          7118 => x"e6",
          7119 => x"0c",
          7120 => x"0d",
          7121 => x"80",
          7122 => x"83",
          7123 => x"26",
          7124 => x"56",
          7125 => x"73",
          7126 => x"70",
          7127 => x"22",
          7128 => x"ff",
          7129 => x"24",
          7130 => x"15",
          7131 => x"73",
          7132 => x"07",
          7133 => x"38",
          7134 => x"87",
          7135 => x"ff",
          7136 => x"71",
          7137 => x"73",
          7138 => x"ff",
          7139 => x"39",
          7140 => x"06",
          7141 => x"83",
          7142 => x"e6",
          7143 => x"51",
          7144 => x"ff",
          7145 => x"70",
          7146 => x"39",
          7147 => x"57",
          7148 => x"81",
          7149 => x"ff",
          7150 => x"75",
          7151 => x"52",
          7152 => x"00",
          7153 => x"ff",
          7154 => x"00",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"00",
          7372 => x"00",
          7373 => x"00",
          7374 => x"00",
          7375 => x"00",
          7376 => x"00",
          7377 => x"00",
          7378 => x"00",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"00",
          7383 => x"00",
          7384 => x"00",
          7385 => x"00",
          7386 => x"00",
          7387 => x"00",
          7388 => x"00",
          7389 => x"00",
          7390 => x"00",
          7391 => x"74",
          7392 => x"74",
          7393 => x"74",
          7394 => x"64",
          7395 => x"63",
          7396 => x"61",
          7397 => x"79",
          7398 => x"66",
          7399 => x"70",
          7400 => x"6d",
          7401 => x"68",
          7402 => x"68",
          7403 => x"63",
          7404 => x"6a",
          7405 => x"61",
          7406 => x"74",
          7407 => x"00",
          7408 => x"00",
          7409 => x"7a",
          7410 => x"69",
          7411 => x"69",
          7412 => x"00",
          7413 => x"55",
          7414 => x"65",
          7415 => x"50",
          7416 => x"72",
          7417 => x"72",
          7418 => x"54",
          7419 => x"20",
          7420 => x"6c",
          7421 => x"49",
          7422 => x"69",
          7423 => x"6f",
          7424 => x"46",
          7425 => x"6c",
          7426 => x"54",
          7427 => x"20",
          7428 => x"6f",
          7429 => x"6c",
          7430 => x"46",
          7431 => x"62",
          7432 => x"4e",
          7433 => x"74",
          7434 => x"6c",
          7435 => x"20",
          7436 => x"6e",
          7437 => x"44",
          7438 => x"20",
          7439 => x"2e",
          7440 => x"65",
          7441 => x"20",
          7442 => x"6c",
          7443 => x"53",
          7444 => x"69",
          7445 => x"65",
          7446 => x"46",
          7447 => x"64",
          7448 => x"6c",
          7449 => x"46",
          7450 => x"65",
          7451 => x"73",
          7452 => x"41",
          7453 => x"65",
          7454 => x"49",
          7455 => x"66",
          7456 => x"2e",
          7457 => x"61",
          7458 => x"64",
          7459 => x"69",
          7460 => x"64",
          7461 => x"20",
          7462 => x"64",
          7463 => x"72",
          7464 => x"6f",
          7465 => x"20",
          7466 => x"53",
          7467 => x"00",
          7468 => x"20",
          7469 => x"73",
          7470 => x"20",
          7471 => x"65",
          7472 => x"72",
          7473 => x"25",
          7474 => x"3a",
          7475 => x"00",
          7476 => x"7c",
          7477 => x"25",
          7478 => x"20",
          7479 => x"00",
          7480 => x"2a",
          7481 => x"32",
          7482 => x"32",
          7483 => x"32",
          7484 => x"2c",
          7485 => x"32",
          7486 => x"73",
          7487 => x"4f",
          7488 => x"42",
          7489 => x"72",
          7490 => x"20",
          7491 => x"20",
          7492 => x"0a",
          7493 => x"41",
          7494 => x"65",
          7495 => x"20",
          7496 => x"20",
          7497 => x"0a",
          7498 => x"49",
          7499 => x"74",
          7500 => x"72",
          7501 => x"31",
          7502 => x"65",
          7503 => x"55",
          7504 => x"20",
          7505 => x"70",
          7506 => x"30",
          7507 => x"65",
          7508 => x"55",
          7509 => x"20",
          7510 => x"70",
          7511 => x"4c",
          7512 => x"65",
          7513 => x"49",
          7514 => x"20",
          7515 => x"70",
          7516 => x"69",
          7517 => x"74",
          7518 => x"72",
          7519 => x"75",
          7520 => x"69",
          7521 => x"69",
          7522 => x"45",
          7523 => x"20",
          7524 => x"2e",
          7525 => x"65",
          7526 => x"00",
          7527 => x"7a",
          7528 => x"46",
          7529 => x"6f",
          7530 => x"6c",
          7531 => x"63",
          7532 => x"70",
          7533 => x"6e",
          7534 => x"61",
          7535 => x"2a",
          7536 => x"25",
          7537 => x"42",
          7538 => x"61",
          7539 => x"5a",
          7540 => x"25",
          7541 => x"73",
          7542 => x"43",
          7543 => x"6f",
          7544 => x"2e",
          7545 => x"61",
          7546 => x"70",
          7547 => x"6f",
          7548 => x"43",
          7549 => x"63",
          7550 => x"30",
          7551 => x"0a",
          7552 => x"20",
          7553 => x"64",
          7554 => x"25",
          7555 => x"45",
          7556 => x"67",
          7557 => x"20",
          7558 => x"2e",
          7559 => x"58",
          7560 => x"00",
          7561 => x"58",
          7562 => x"43",
          7563 => x"67",
          7564 => x"25",
          7565 => x"38",
          7566 => x"6c",
          7567 => x"0a",
          7568 => x"69",
          7569 => x"25",
          7570 => x"32",
          7571 => x"72",
          7572 => x"00",
          7573 => x"20",
          7574 => x"0a",
          7575 => x"65",
          7576 => x"25",
          7577 => x"4d",
          7578 => x"78",
          7579 => x"2c",
          7580 => x"20",
          7581 => x"20",
          7582 => x"2e",
          7583 => x"25",
          7584 => x"20",
          7585 => x"64",
          7586 => x"53",
          7587 => x"69",
          7588 => x"6e",
          7589 => x"76",
          7590 => x"70",
          7591 => x"64",
          7592 => x"65",
          7593 => x"20",
          7594 => x"52",
          7595 => x"63",
          7596 => x"72",
          7597 => x"30",
          7598 => x"20",
          7599 => x"4d",
          7600 => x"74",
          7601 => x"72",
          7602 => x"30",
          7603 => x"20",
          7604 => x"6b",
          7605 => x"41",
          7606 => x"20",
          7607 => x"30",
          7608 => x"4d",
          7609 => x"20",
          7610 => x"49",
          7611 => x"20",
          7612 => x"20",
          7613 => x"30",
          7614 => x"20",
          7615 => x"65",
          7616 => x"20",
          7617 => x"20",
          7618 => x"64",
          7619 => x"7a",
          7620 => x"57",
          7621 => x"20",
          7622 => x"6c",
          7623 => x"71",
          7624 => x"34",
          7625 => x"20",
          7626 => x"4d",
          7627 => x"46",
          7628 => x"20",
          7629 => x"64",
          7630 => x"7a",
          7631 => x"53",
          7632 => x"50",
          7633 => x"49",
          7634 => x"20",
          7635 => x"32",
          7636 => x"57",
          7637 => x"20",
          7638 => x"20",
          7639 => x"20",
          7640 => x"68",
          7641 => x"25",
          7642 => x"20",
          7643 => x"52",
          7644 => x"69",
          7645 => x"25",
          7646 => x"20",
          7647 => x"41",
          7648 => x"65",
          7649 => x"25",
          7650 => x"20",
          7651 => x"20",
          7652 => x"30",
          7653 => x"29",
          7654 => x"42",
          7655 => x"20",
          7656 => x"25",
          7657 => x"20",
          7658 => x"20",
          7659 => x"30",
          7660 => x"29",
          7661 => x"53",
          7662 => x"20",
          7663 => x"25",
          7664 => x"20",
          7665 => x"44",
          7666 => x"30",
          7667 => x"29",
          7668 => x"6f",
          7669 => x"6f",
          7670 => x"55",
          7671 => x"45",
          7672 => x"53",
          7673 => x"4d",
          7674 => x"46",
          7675 => x"45",
          7676 => x"01",
          7677 => x"00",
          7678 => x"00",
          7679 => x"01",
          7680 => x"00",
          7681 => x"00",
          7682 => x"01",
          7683 => x"00",
          7684 => x"00",
          7685 => x"01",
          7686 => x"00",
          7687 => x"00",
          7688 => x"01",
          7689 => x"00",
          7690 => x"00",
          7691 => x"01",
          7692 => x"00",
          7693 => x"00",
          7694 => x"04",
          7695 => x"00",
          7696 => x"00",
          7697 => x"03",
          7698 => x"00",
          7699 => x"00",
          7700 => x"04",
          7701 => x"00",
          7702 => x"00",
          7703 => x"03",
          7704 => x"00",
          7705 => x"00",
          7706 => x"03",
          7707 => x"00",
          7708 => x"00",
          7709 => x"1b",
          7710 => x"1b",
          7711 => x"1b",
          7712 => x"1b",
          7713 => x"1b",
          7714 => x"10",
          7715 => x"0d",
          7716 => x"08",
          7717 => x"05",
          7718 => x"03",
          7719 => x"01",
          7720 => x"6f",
          7721 => x"3a",
          7722 => x"43",
          7723 => x"70",
          7724 => x"74",
          7725 => x"72",
          7726 => x"20",
          7727 => x"6e",
          7728 => x"6f",
          7729 => x"00",
          7730 => x"48",
          7731 => x"62",
          7732 => x"30",
          7733 => x"25",
          7734 => x"73",
          7735 => x"65",
          7736 => x"73",
          7737 => x"68",
          7738 => x"66",
          7739 => x"45",
          7740 => x"3e",
          7741 => x"1b",
          7742 => x"1b",
          7743 => x"1b",
          7744 => x"1b",
          7745 => x"1b",
          7746 => x"1b",
          7747 => x"1b",
          7748 => x"1b",
          7749 => x"1b",
          7750 => x"1b",
          7751 => x"1b",
          7752 => x"1b",
          7753 => x"1b",
          7754 => x"1b",
          7755 => x"1b",
          7756 => x"1b",
          7757 => x"00",
          7758 => x"00",
          7759 => x"2c",
          7760 => x"64",
          7761 => x"25",
          7762 => x"44",
          7763 => x"25",
          7764 => x"2c",
          7765 => x"25",
          7766 => x"3a",
          7767 => x"2c",
          7768 => x"64",
          7769 => x"52",
          7770 => x"75",
          7771 => x"55",
          7772 => x"25",
          7773 => x"44",
          7774 => x"25",
          7775 => x"48",
          7776 => x"00",
          7777 => x"65",
          7778 => x"6e",
          7779 => x"53",
          7780 => x"3e",
          7781 => x"2b",
          7782 => x"46",
          7783 => x"32",
          7784 => x"53",
          7785 => x"4e",
          7786 => x"20",
          7787 => x"20",
          7788 => x"41",
          7789 => x"41",
          7790 => x"00",
          7791 => x"00",
          7792 => x"01",
          7793 => x"14",
          7794 => x"80",
          7795 => x"45",
          7796 => x"90",
          7797 => x"59",
          7798 => x"41",
          7799 => x"a8",
          7800 => x"b0",
          7801 => x"b8",
          7802 => x"c0",
          7803 => x"c8",
          7804 => x"d0",
          7805 => x"d8",
          7806 => x"e0",
          7807 => x"e8",
          7808 => x"f0",
          7809 => x"f8",
          7810 => x"2b",
          7811 => x"5c",
          7812 => x"7f",
          7813 => x"00",
          7814 => x"00",
          7815 => x"00",
          7816 => x"00",
          7817 => x"00",
          7818 => x"00",
          7819 => x"00",
          7820 => x"00",
          7821 => x"00",
          7822 => x"00",
          7823 => x"00",
          7824 => x"20",
          7825 => x"00",
          7826 => x"00",
          7827 => x"00",
          7828 => x"00",
          7829 => x"25",
          7830 => x"25",
          7831 => x"25",
          7832 => x"25",
          7833 => x"25",
          7834 => x"25",
          7835 => x"25",
          7836 => x"25",
          7837 => x"25",
          7838 => x"25",
          7839 => x"25",
          7840 => x"25",
          7841 => x"03",
          7842 => x"00",
          7843 => x"03",
          7844 => x"03",
          7845 => x"22",
          7846 => x"00",
          7847 => x"00",
          7848 => x"25",
          7849 => x"00",
          7850 => x"00",
          7851 => x"01",
          7852 => x"01",
          7853 => x"01",
          7854 => x"01",
          7855 => x"01",
          7856 => x"01",
          7857 => x"01",
          7858 => x"01",
          7859 => x"01",
          7860 => x"01",
          7861 => x"01",
          7862 => x"01",
          7863 => x"01",
          7864 => x"01",
          7865 => x"01",
          7866 => x"01",
          7867 => x"01",
          7868 => x"01",
          7869 => x"01",
          7870 => x"01",
          7871 => x"01",
          7872 => x"01",
          7873 => x"01",
          7874 => x"01",
          7875 => x"00",
          7876 => x"01",
          7877 => x"02",
          7878 => x"02",
          7879 => x"02",
          7880 => x"01",
          7881 => x"01",
          7882 => x"02",
          7883 => x"02",
          7884 => x"01",
          7885 => x"02",
          7886 => x"01",
          7887 => x"02",
          7888 => x"02",
          7889 => x"02",
          7890 => x"02",
          7891 => x"02",
          7892 => x"01",
          7893 => x"02",
          7894 => x"01",
          7895 => x"02",
          7896 => x"02",
          7897 => x"00",
          7898 => x"03",
          7899 => x"03",
          7900 => x"03",
          7901 => x"03",
          7902 => x"03",
          7903 => x"01",
          7904 => x"03",
          7905 => x"03",
          7906 => x"03",
          7907 => x"07",
          7908 => x"01",
          7909 => x"00",
          7910 => x"05",
          7911 => x"1d",
          7912 => x"01",
          7913 => x"06",
          7914 => x"06",
          7915 => x"06",
          7916 => x"1f",
          7917 => x"1f",
          7918 => x"1f",
          7919 => x"1f",
          7920 => x"1f",
          7921 => x"1f",
          7922 => x"1f",
          7923 => x"1f",
          7924 => x"1f",
          7925 => x"1f",
          7926 => x"06",
          7927 => x"00",
          7928 => x"1f",
          7929 => x"21",
          7930 => x"21",
          7931 => x"04",
          7932 => x"01",
          7933 => x"01",
          7934 => x"03",
          7935 => x"00",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"00",
          7940 => x"00",
          7941 => x"00",
          7942 => x"00",
          7943 => x"00",
          7944 => x"00",
          7945 => x"00",
          7946 => x"00",
          7947 => x"00",
          7948 => x"00",
          7949 => x"00",
          7950 => x"00",
          7951 => x"00",
          7952 => x"00",
          7953 => x"00",
          7954 => x"00",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"00",
          7959 => x"00",
          7960 => x"00",
          7961 => x"00",
          7962 => x"00",
          7963 => x"00",
          7964 => x"00",
          7965 => x"00",
          7966 => x"00",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"00",
          7983 => x"00",
          7984 => x"00",
          7985 => x"00",
          7986 => x"00",
          7987 => x"00",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"00",
          7996 => x"01",
          7997 => x"00",
          7998 => x"00",
          7999 => x"05",
          8000 => x"00",
          8001 => x"01",
          8002 => x"01",
          8003 => x"00",
          8004 => x"00",
          8005 => x"00",
          8006 => x"00",
          8007 => x"00",
          8008 => x"00",
          8009 => x"00",
          8010 => x"00",
          8011 => x"00",
          8012 => x"00",
          8013 => x"00",
          8014 => x"00",
          8015 => x"01",
          8016 => x"01",
          8017 => x"02",
          8018 => x"1b",
          8019 => x"79",
          8020 => x"71",
          8021 => x"69",
          8022 => x"61",
          8023 => x"31",
          8024 => x"5c",
          8025 => x"f6",
          8026 => x"08",
          8027 => x"80",
          8028 => x"1b",
          8029 => x"59",
          8030 => x"51",
          8031 => x"49",
          8032 => x"41",
          8033 => x"31",
          8034 => x"5c",
          8035 => x"f6",
          8036 => x"08",
          8037 => x"80",
          8038 => x"1b",
          8039 => x"59",
          8040 => x"51",
          8041 => x"49",
          8042 => x"41",
          8043 => x"21",
          8044 => x"7c",
          8045 => x"f7",
          8046 => x"fb",
          8047 => x"85",
          8048 => x"1b",
          8049 => x"19",
          8050 => x"11",
          8051 => x"09",
          8052 => x"01",
          8053 => x"f0",
          8054 => x"f0",
          8055 => x"f0",
          8056 => x"f0",
          8057 => x"80",
          8058 => x"bf",
          8059 => x"35",
          8060 => x"7c",
          8061 => x"3d",
          8062 => x"46",
          8063 => x"3f",
          8064 => x"d3",
          8065 => x"c6",
          8066 => x"f0",
          8067 => x"80",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
          9101 => x"00",
          9102 => x"00",
          9103 => x"00",
          9104 => x"ce",
          9105 => x"fc",
          9106 => x"c4",
          9107 => x"eb",
          9108 => x"64",
          9109 => x"2f",
          9110 => x"24",
          9111 => x"51",
          9112 => x"04",
          9113 => x"0c",
          9114 => x"14",
          9115 => x"59",
          9116 => x"84",
          9117 => x"8c",
          9118 => x"94",
          9119 => x"80",
          9120 => x"00",
          9121 => x"00",
          9122 => x"00",
          9123 => x"00",
          9124 => x"00",
          9125 => x"00",
          9126 => x"00",
          9127 => x"00",
          9128 => x"00",
          9129 => x"00",
          9130 => x"00",
          9131 => x"00",
          9132 => x"00",
          9133 => x"00",
          9134 => x"00",
          9135 => x"00",
          9136 => x"00",
        others => X"00"
    );

    signal RAM0_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM1_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM2_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM3_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM4_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM5_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM6_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM7_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM0_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM1_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM2_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM3_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM4_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM5_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM6_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM7_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal lowDataA          :     std_logic_vector(WORD_32BIT_RANGE);   -- Low word in 64 bit output from RAM matrix.
    signal highDataA         :     std_logic_vector(WORD_32BIT_RANGE);   -- High word in 64 bit output from RAM matrix.
    signal lowDataB          :     std_logic_vector(WORD_32BIT_RANGE);   -- Low word in 64 bit output from RAM matrix.
    signal highDataB         :     std_logic_vector(WORD_32BIT_RANGE);   -- High word in 64 bit output from RAM matrix.

begin

    -- Correctly assign the Little Endian value to the correct array, byte writes the data is in '7 downto 0', h-word writes
    -- the data is in '15 downto 0', word writes the data is in '31 downto 0'. Long words (64bits) are treated as two words for Endianness,
    -- and not as one continuous long word, this is because the ZPU is 32bit even when accessing a 64bit chunk.
    --
    RAM0_DATA <= memAWrite(7 downto 0)   when memAAddr(2) = '0'
                 else (others => '0');
    RAM1_DATA <= memAWrite(15 downto 8)  when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(15 downto 8)  when memAAddr(2) = '0' and (memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM4_DATA <= memAWrite(7 downto 0)   when memAAddr(2) = '1'
                 else (others => '0');
    RAM5_DATA <= memAWrite(15 downto 8)  when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM6_DATA <= memAWrite(23 downto 16) when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(7 downto 0);
    RAM7_DATA <= memAWrite(31 downto 24) when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(15 downto 8)  when memAAddr(2) = '1' and (memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "011") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "01"))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "010") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "01"))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "001") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "00"))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "000") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "00"))
                 else '0';
    RAM4_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "111") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "11"))
                 else '0';
    RAM5_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "110") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "11"))
                 else '0';
    RAM6_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "101") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "10"))
                 else '0';
    RAM7_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "100") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "10"))
                 else '0';

    memARead  <= lowDataA  when memAAddr(2) = '0'
                 else
                 highDataA;
    memBRead  <= lowDataB & highDataB;

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM0_DATA;
            else
                lowDataA(7 downto 0)    <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM1_DATA;
            else
                lowDataA(15 downto 8)   <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM2_DATA;
            else
                lowDataA(23 downto 16)  <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM3_DATA;
            else
                lowDataA(31 downto 24)  <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 4 - Port A - bits 39 to 32 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM4_WREN = '1' then
                RAM4(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM4_DATA;
            else
                highDataA(7 downto 0)   <= RAM4(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 5 - Port A - bits 47 to 40 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM5_WREN = '1' then
                RAM5(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM5_DATA;
            else
                highDataA(15 downto 8)  <= RAM5(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 6 - Port A - bits 56 to 48
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM6_WREN = '1' then
                RAM6(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM6_DATA;
            else
                highDataA(23 downto 16) <= RAM6(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 7 - Port A - bits 63 to 57 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM7_WREN = '1' then
                RAM7(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM7_DATA;
            else
                highDataA(31 downto 24) <= RAM7(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;


    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(7 downto 0);
                lowDataB(7 downto 0)    <= memBWrite(7 downto 0);
            else
                lowDataB(7 downto 0)    <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(15 downto 8);
                lowDataB(15 downto 8)    <= memBWrite(15 downto 8);
            else
                lowDataB(15 downto 8)    <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(23 downto 16);
                lowDataB(23 downto 16)  <= memBWrite(23 downto 16);
            else
                lowDataB(23 downto 16)  <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(31 downto 24);
                lowDataB(31 downto 24)  <= memBWrite(31 downto 24);
            else
                lowDataB(31 downto 24)  <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 4 - Port B - bits 39 downto 32
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM4(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(39 downto 32);
                highDataB(7 downto 0)   <= memBWrite(39 downto 32);
            else
                highDataB(7 downto 0)   <= RAM4(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 5 - Port B - bits 47 downto 40
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM5(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(47 downto 40);
                highDataB(15 downto 8)  <= memBWrite(47 downto 40);
            else
                highDataB(15 downto 8)  <= RAM5(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 6 - Port B - bits 55 downto 48
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM6(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(55 downto 48);
                highDataB(23 downto 16)  <= memBWrite(55 downto 48);
            else
                highDataB(23 downto 16)  <= RAM6(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 7 - Port B - bits 63 downto 56 
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM7(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(63 downto 56);
                highDataB(31 downto 24)  <= memBWrite(63 downto 56);
            else
                highDataB(31 downto 24)  <= RAM7(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

end arch;
