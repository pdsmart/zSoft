-- Byte Addressed 32bit/64bit BRAM module for the ZPU Evo implementation.
--
-- This template provides a 32bit wide bus on port A and a 64bit bus
-- on port B. This is typically used for the ZPU Boot BRAM where port B
-- is used exclusively for instruction storage.
--
-- Copyright 2018-2021 - Philip Smart for the ZPU Evo implementation.
-- History:
--   20190618  - Initial 32 bit dual port BRAM described by inference rather than
--               using an IP Megacore. This was to make it more portable but also
--               to allow 8/16/32 bit writes to the memory.
--   20210108  - Updated to 64bit on Port B to allow for the 64bit decoder on the ZPU.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.softZPU_pkg.all;

entity DualPort3264BootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 3);
        memBWrite            : in  std_logic_vector(WORD_64BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_64BIT_RANGE)
    );
end DualPort3264BootBRAM;

architecture arch of DualPort3264BootBRAM is

    -- Declare 8 byte wide arrays for byte level addressing.
    type ramArray is array(natural range 0 to (2**(addrbits-3))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"fa",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"05",
            10 => x"52",
            11 => x"00",
            12 => x"08",
            13 => x"81",
            14 => x"06",
            15 => x"0b",
            16 => x"05",
            17 => x"06",
            18 => x"06",
            19 => x"00",
            20 => x"73",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"09",
            25 => x"72",
            26 => x"31",
            27 => x"51",
            28 => x"73",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"93",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"2b",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"06",
            45 => x"b0",
            46 => x"00",
            47 => x"00",
            48 => x"ff",
            49 => x"0a",
            50 => x"51",
            51 => x"00",
            52 => x"51",
            53 => x"05",
            54 => x"72",
            55 => x"00",
            56 => x"05",
            57 => x"06",
            58 => x"00",
            59 => x"00",
            60 => x"05",
            61 => x"06",
            62 => x"00",
            63 => x"00",
            64 => x"05",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"81",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"06",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"08",
            77 => x"05",
            78 => x"52",
            79 => x"00",
            80 => x"08",
            81 => x"06",
            82 => x"0b",
            83 => x"00",
            84 => x"08",
            85 => x"ac",
            86 => x"90",
            87 => x"00",
            88 => x"08",
            89 => x"ab",
            90 => x"90",
            91 => x"00",
            92 => x"81",
            93 => x"05",
            94 => x"74",
            95 => x"51",
            96 => x"81",
            97 => x"ff",
            98 => x"72",
            99 => x"51",
           100 => x"04",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"52",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"72",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"ff",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"8c",
           133 => x"04",
           134 => x"0b",
           135 => x"8c",
           136 => x"04",
           137 => x"0b",
           138 => x"8c",
           139 => x"04",
           140 => x"0b",
           141 => x"8d",
           142 => x"04",
           143 => x"0b",
           144 => x"8d",
           145 => x"04",
           146 => x"0b",
           147 => x"8e",
           148 => x"04",
           149 => x"0b",
           150 => x"8f",
           151 => x"04",
           152 => x"0b",
           153 => x"8f",
           154 => x"04",
           155 => x"0b",
           156 => x"90",
           157 => x"04",
           158 => x"0b",
           159 => x"90",
           160 => x"04",
           161 => x"0b",
           162 => x"91",
           163 => x"04",
           164 => x"0b",
           165 => x"91",
           166 => x"04",
           167 => x"0b",
           168 => x"92",
           169 => x"04",
           170 => x"0b",
           171 => x"92",
           172 => x"04",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"81",
           193 => x"f6",
           194 => x"80",
           195 => x"ee",
           196 => x"80",
           197 => x"f3",
           198 => x"80",
           199 => x"e0",
           200 => x"80",
           201 => x"a3",
           202 => x"80",
           203 => x"f6",
           204 => x"80",
           205 => x"86",
           206 => x"80",
           207 => x"82",
           208 => x"80",
           209 => x"88",
           210 => x"80",
           211 => x"a8",
           212 => x"80",
           213 => x"d1",
           214 => x"80",
           215 => x"8a",
           216 => x"80",
           217 => x"d4",
           218 => x"c0",
           219 => x"80",
           220 => x"80",
           221 => x"0c",
           222 => x"08",
           223 => x"98",
           224 => x"98",
           225 => x"ba",
           226 => x"ba",
           227 => x"84",
           228 => x"84",
           229 => x"04",
           230 => x"2d",
           231 => x"90",
           232 => x"89",
           233 => x"80",
           234 => x"ed",
           235 => x"c0",
           236 => x"82",
           237 => x"80",
           238 => x"0c",
           239 => x"08",
           240 => x"98",
           241 => x"98",
           242 => x"ba",
           243 => x"ba",
           244 => x"84",
           245 => x"84",
           246 => x"04",
           247 => x"2d",
           248 => x"90",
           249 => x"b0",
           250 => x"80",
           251 => x"8b",
           252 => x"c0",
           253 => x"82",
           254 => x"80",
           255 => x"0c",
           256 => x"08",
           257 => x"98",
           258 => x"98",
           259 => x"ba",
           260 => x"ba",
           261 => x"84",
           262 => x"84",
           263 => x"04",
           264 => x"2d",
           265 => x"90",
           266 => x"f0",
           267 => x"80",
           268 => x"96",
           269 => x"c0",
           270 => x"83",
           271 => x"80",
           272 => x"0c",
           273 => x"08",
           274 => x"98",
           275 => x"98",
           276 => x"ba",
           277 => x"ba",
           278 => x"84",
           279 => x"84",
           280 => x"04",
           281 => x"2d",
           282 => x"90",
           283 => x"ac",
           284 => x"80",
           285 => x"f5",
           286 => x"c0",
           287 => x"81",
           288 => x"80",
           289 => x"0c",
           290 => x"08",
           291 => x"98",
           292 => x"98",
           293 => x"ba",
           294 => x"ba",
           295 => x"84",
           296 => x"ba",
           297 => x"84",
           298 => x"84",
           299 => x"04",
           300 => x"2d",
           301 => x"90",
           302 => x"86",
           303 => x"80",
           304 => x"d5",
           305 => x"c0",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"00",
           311 => x"06",
           312 => x"10",
           313 => x"51",
           314 => x"ff",
           315 => x"52",
           316 => x"38",
           317 => x"8c",
           318 => x"80",
           319 => x"0b",
           320 => x"80",
           321 => x"87",
           322 => x"56",
           323 => x"51",
           324 => x"fa",
           325 => x"33",
           326 => x"07",
           327 => x"72",
           328 => x"ff",
           329 => x"70",
           330 => x"56",
           331 => x"80",
           332 => x"3f",
           333 => x"8c",
           334 => x"8c",
           335 => x"ff",
           336 => x"72",
           337 => x"73",
           338 => x"76",
           339 => x"3d",
           340 => x"0c",
           341 => x"7d",
           342 => x"34",
           343 => x"88",
           344 => x"05",
           345 => x"74",
           346 => x"0d",
           347 => x"75",
           348 => x"f1",
           349 => x"5d",
           350 => x"33",
           351 => x"55",
           352 => x"09",
           353 => x"57",
           354 => x"1c",
           355 => x"2e",
           356 => x"89",
           357 => x"70",
           358 => x"78",
           359 => x"7a",
           360 => x"40",
           361 => x"82",
           362 => x"ff",
           363 => x"84",
           364 => x"7a",
           365 => x"79",
           366 => x"2c",
           367 => x"0a",
           368 => x"56",
           369 => x"73",
           370 => x"78",
           371 => x"38",
           372 => x"81",
           373 => x"5a",
           374 => x"fe",
           375 => x"76",
           376 => x"76",
           377 => x"83",
           378 => x"8a",
           379 => x"7e",
           380 => x"d8",
           381 => x"ca",
           382 => x"e0",
           383 => x"eb",
           384 => x"3f",
           385 => x"86",
           386 => x"fe",
           387 => x"05",
           388 => x"5e",
           389 => x"79",
           390 => x"ba",
           391 => x"8c",
           392 => x"89",
           393 => x"b0",
           394 => x"40",
           395 => x"3f",
           396 => x"8c",
           397 => x"31",
           398 => x"7e",
           399 => x"80",
           400 => x"2c",
           401 => x"06",
           402 => x"77",
           403 => x"05",
           404 => x"84",
           405 => x"53",
           406 => x"70",
           407 => x"9e",
           408 => x"06",
           409 => x"38",
           410 => x"2a",
           411 => x"81",
           412 => x"38",
           413 => x"2c",
           414 => x"73",
           415 => x"2a",
           416 => x"7a",
           417 => x"98",
           418 => x"73",
           419 => x"73",
           420 => x"06",
           421 => x"78",
           422 => x"05",
           423 => x"74",
           424 => x"88",
           425 => x"29",
           426 => x"5a",
           427 => x"74",
           428 => x"38",
           429 => x"ff",
           430 => x"55",
           431 => x"b0",
           432 => x"80",
           433 => x"98",
           434 => x"e5",
           435 => x"5c",
           436 => x"76",
           437 => x"80",
           438 => x"d3",
           439 => x"9c",
           440 => x"70",
           441 => x"84",
           442 => x"38",
           443 => x"fc",
           444 => x"29",
           445 => x"5a",
           446 => x"38",
           447 => x"e2",
           448 => x"07",
           449 => x"38",
           450 => x"5b",
           451 => x"05",
           452 => x"5f",
           453 => x"7f",
           454 => x"06",
           455 => x"07",
           456 => x"80",
           457 => x"56",
           458 => x"81",
           459 => x"77",
           460 => x"80",
           461 => x"80",
           462 => x"a0",
           463 => x"1a",
           464 => x"79",
           465 => x"7c",
           466 => x"51",
           467 => x"70",
           468 => x"83",
           469 => x"52",
           470 => x"85",
           471 => x"06",
           472 => x"80",
           473 => x"2c",
           474 => x"2a",
           475 => x"fd",
           476 => x"84",
           477 => x"56",
           478 => x"83",
           479 => x"5e",
           480 => x"33",
           481 => x"ca",
           482 => x"33",
           483 => x"ba",
           484 => x"77",
           485 => x"82",
           486 => x"84",
           487 => x"78",
           488 => x"90",
           489 => x"c0",
           490 => x"be",
           491 => x"05",
           492 => x"41",
           493 => x"87",
           494 => x"ff",
           495 => x"54",
           496 => x"7c",
           497 => x"f7",
           498 => x"29",
           499 => x"5a",
           500 => x"38",
           501 => x"e2",
           502 => x"3f",
           503 => x"e3",
           504 => x"3f",
           505 => x"80",
           506 => x"75",
           507 => x"70",
           508 => x"5a",
           509 => x"a2",
           510 => x"3f",
           511 => x"fa",
           512 => x"75",
           513 => x"81",
           514 => x"38",
           515 => x"2b",
           516 => x"39",
           517 => x"c8",
           518 => x"3f",
           519 => x"88",
           520 => x"ff",
           521 => x"54",
           522 => x"7e",
           523 => x"57",
           524 => x"84",
           525 => x"51",
           526 => x"fa",
           527 => x"d5",
           528 => x"2a",
           529 => x"58",
           530 => x"09",
           531 => x"81",
           532 => x"b0",
           533 => x"51",
           534 => x"ba",
           535 => x"57",
           536 => x"72",
           537 => x"08",
           538 => x"54",
           539 => x"90",
           540 => x"8c",
           541 => x"76",
           542 => x"3d",
           543 => x"56",
           544 => x"81",
           545 => x"55",
           546 => x"09",
           547 => x"05",
           548 => x"81",
           549 => x"ba",
           550 => x"70",
           551 => x"2e",
           552 => x"15",
           553 => x"08",
           554 => x"81",
           555 => x"38",
           556 => x"f0",
           557 => x"3d",
           558 => x"85",
           559 => x"81",
           560 => x"72",
           561 => x"54",
           562 => x"08",
           563 => x"38",
           564 => x"08",
           565 => x"53",
           566 => x"75",
           567 => x"04",
           568 => x"90",
           569 => x"84",
           570 => x"08",
           571 => x"d7",
           572 => x"33",
           573 => x"81",
           574 => x"71",
           575 => x"52",
           576 => x"06",
           577 => x"75",
           578 => x"2e",
           579 => x"8c",
           580 => x"71",
           581 => x"8c",
           582 => x"bf",
           583 => x"16",
           584 => x"16",
           585 => x"0d",
           586 => x"74",
           587 => x"ba",
           588 => x"85",
           589 => x"84",
           590 => x"71",
           591 => x"ff",
           592 => x"3d",
           593 => x"85",
           594 => x"3d",
           595 => x"71",
           596 => x"f7",
           597 => x"05",
           598 => x"05",
           599 => x"ba",
           600 => x"3d",
           601 => x"52",
           602 => x"72",
           603 => x"38",
           604 => x"70",
           605 => x"70",
           606 => x"86",
           607 => x"75",
           608 => x"53",
           609 => x"33",
           610 => x"2e",
           611 => x"53",
           612 => x"70",
           613 => x"74",
           614 => x"53",
           615 => x"70",
           616 => x"84",
           617 => x"77",
           618 => x"05",
           619 => x"05",
           620 => x"ba",
           621 => x"3d",
           622 => x"52",
           623 => x"70",
           624 => x"05",
           625 => x"38",
           626 => x"0d",
           627 => x"55",
           628 => x"73",
           629 => x"52",
           630 => x"9a",
           631 => x"b7",
           632 => x"80",
           633 => x"3d",
           634 => x"73",
           635 => x"e9",
           636 => x"71",
           637 => x"84",
           638 => x"71",
           639 => x"04",
           640 => x"52",
           641 => x"08",
           642 => x"55",
           643 => x"08",
           644 => x"9b",
           645 => x"80",
           646 => x"ba",
           647 => x"ba",
           648 => x"0c",
           649 => x"75",
           650 => x"71",
           651 => x"05",
           652 => x"38",
           653 => x"81",
           654 => x"31",
           655 => x"85",
           656 => x"77",
           657 => x"80",
           658 => x"05",
           659 => x"38",
           660 => x"0d",
           661 => x"54",
           662 => x"76",
           663 => x"08",
           664 => x"8d",
           665 => x"84",
           666 => x"72",
           667 => x"72",
           668 => x"74",
           669 => x"2b",
           670 => x"76",
           671 => x"2a",
           672 => x"31",
           673 => x"7b",
           674 => x"5c",
           675 => x"74",
           676 => x"71",
           677 => x"04",
           678 => x"80",
           679 => x"25",
           680 => x"71",
           681 => x"30",
           682 => x"31",
           683 => x"70",
           684 => x"71",
           685 => x"1b",
           686 => x"80",
           687 => x"2a",
           688 => x"06",
           689 => x"19",
           690 => x"54",
           691 => x"55",
           692 => x"58",
           693 => x"fd",
           694 => x"53",
           695 => x"8c",
           696 => x"ba",
           697 => x"fa",
           698 => x"53",
           699 => x"fe",
           700 => x"e0",
           701 => x"73",
           702 => x"8c",
           703 => x"26",
           704 => x"2e",
           705 => x"a0",
           706 => x"54",
           707 => x"38",
           708 => x"10",
           709 => x"9f",
           710 => x"75",
           711 => x"52",
           712 => x"72",
           713 => x"04",
           714 => x"9f",
           715 => x"9f",
           716 => x"74",
           717 => x"56",
           718 => x"ba",
           719 => x"ba",
           720 => x"3d",
           721 => x"7b",
           722 => x"59",
           723 => x"38",
           724 => x"55",
           725 => x"ad",
           726 => x"81",
           727 => x"77",
           728 => x"80",
           729 => x"80",
           730 => x"70",
           731 => x"70",
           732 => x"27",
           733 => x"06",
           734 => x"38",
           735 => x"76",
           736 => x"70",
           737 => x"ff",
           738 => x"75",
           739 => x"75",
           740 => x"04",
           741 => x"33",
           742 => x"81",
           743 => x"78",
           744 => x"e2",
           745 => x"f8",
           746 => x"27",
           747 => x"88",
           748 => x"75",
           749 => x"04",
           750 => x"70",
           751 => x"39",
           752 => x"3d",
           753 => x"5b",
           754 => x"70",
           755 => x"09",
           756 => x"78",
           757 => x"2e",
           758 => x"38",
           759 => x"14",
           760 => x"db",
           761 => x"27",
           762 => x"89",
           763 => x"55",
           764 => x"51",
           765 => x"13",
           766 => x"73",
           767 => x"81",
           768 => x"16",
           769 => x"56",
           770 => x"80",
           771 => x"7a",
           772 => x"0c",
           773 => x"70",
           774 => x"73",
           775 => x"38",
           776 => x"55",
           777 => x"90",
           778 => x"81",
           779 => x"14",
           780 => x"27",
           781 => x"0c",
           782 => x"15",
           783 => x"80",
           784 => x"ba",
           785 => x"d6",
           786 => x"ff",
           787 => x"3d",
           788 => x"38",
           789 => x"52",
           790 => x"ef",
           791 => x"ce",
           792 => x"0d",
           793 => x"3f",
           794 => x"51",
           795 => x"83",
           796 => x"3d",
           797 => x"87",
           798 => x"ec",
           799 => x"04",
           800 => x"83",
           801 => x"ee",
           802 => x"d0",
           803 => x"0d",
           804 => x"3f",
           805 => x"51",
           806 => x"83",
           807 => x"3d",
           808 => x"af",
           809 => x"ac",
           810 => x"04",
           811 => x"83",
           812 => x"ee",
           813 => x"d1",
           814 => x"0d",
           815 => x"3f",
           816 => x"51",
           817 => x"83",
           818 => x"3d",
           819 => x"84",
           820 => x"80",
           821 => x"25",
           822 => x"87",
           823 => x"77",
           824 => x"93",
           825 => x"77",
           826 => x"96",
           827 => x"84",
           828 => x"38",
           829 => x"30",
           830 => x"70",
           831 => x"58",
           832 => x"98",
           833 => x"80",
           834 => x"29",
           835 => x"08",
           836 => x"83",
           837 => x"84",
           838 => x"84",
           839 => x"0c",
           840 => x"d4",
           841 => x"77",
           842 => x"8c",
           843 => x"88",
           844 => x"80",
           845 => x"d5",
           846 => x"b1",
           847 => x"51",
           848 => x"54",
           849 => x"d2",
           850 => x"39",
           851 => x"b7",
           852 => x"53",
           853 => x"84",
           854 => x"2e",
           855 => x"77",
           856 => x"04",
           857 => x"55",
           858 => x"52",
           859 => x"08",
           860 => x"04",
           861 => x"8c",
           862 => x"15",
           863 => x"5e",
           864 => x"52",
           865 => x"83",
           866 => x"54",
           867 => x"2e",
           868 => x"a8",
           869 => x"81",
           870 => x"d0",
           871 => x"d5",
           872 => x"aa",
           873 => x"d2",
           874 => x"75",
           875 => x"70",
           876 => x"27",
           877 => x"74",
           878 => x"06",
           879 => x"80",
           880 => x"81",
           881 => x"a0",
           882 => x"78",
           883 => x"51",
           884 => x"5c",
           885 => x"ba",
           886 => x"58",
           887 => x"76",
           888 => x"57",
           889 => x"0b",
           890 => x"04",
           891 => x"81",
           892 => x"a0",
           893 => x"fe",
           894 => x"f0",
           895 => x"d5",
           896 => x"ea",
           897 => x"73",
           898 => x"72",
           899 => x"ec",
           900 => x"53",
           901 => x"74",
           902 => x"d2",
           903 => x"84",
           904 => x"ea",
           905 => x"38",
           906 => x"38",
           907 => x"db",
           908 => x"08",
           909 => x"78",
           910 => x"84",
           911 => x"f2",
           912 => x"80",
           913 => x"81",
           914 => x"2e",
           915 => x"d0",
           916 => x"90",
           917 => x"af",
           918 => x"70",
           919 => x"72",
           920 => x"73",
           921 => x"57",
           922 => x"38",
           923 => x"8c",
           924 => x"a0",
           925 => x"30",
           926 => x"51",
           927 => x"73",
           928 => x"80",
           929 => x"0d",
           930 => x"80",
           931 => x"9c",
           932 => x"88",
           933 => x"81",
           934 => x"82",
           935 => x"06",
           936 => x"83",
           937 => x"81",
           938 => x"06",
           939 => x"85",
           940 => x"80",
           941 => x"06",
           942 => x"87",
           943 => x"a9",
           944 => x"72",
           945 => x"0d",
           946 => x"d3",
           947 => x"9b",
           948 => x"0d",
           949 => x"d3",
           950 => x"9b",
           951 => x"53",
           952 => x"81",
           953 => x"51",
           954 => x"3f",
           955 => x"52",
           956 => x"39",
           957 => x"88",
           958 => x"a0",
           959 => x"51",
           960 => x"ff",
           961 => x"83",
           962 => x"51",
           963 => x"81",
           964 => x"c2",
           965 => x"e8",
           966 => x"3f",
           967 => x"2a",
           968 => x"2e",
           969 => x"51",
           970 => x"9a",
           971 => x"72",
           972 => x"71",
           973 => x"39",
           974 => x"d4",
           975 => x"98",
           976 => x"51",
           977 => x"ff",
           978 => x"41",
           979 => x"42",
           980 => x"3f",
           981 => x"9b",
           982 => x"b1",
           983 => x"3f",
           984 => x"d6",
           985 => x"80",
           986 => x"0b",
           987 => x"06",
           988 => x"38",
           989 => x"81",
           990 => x"c1",
           991 => x"2e",
           992 => x"a0",
           993 => x"1a",
           994 => x"f6",
           995 => x"38",
           996 => x"70",
           997 => x"ba",
           998 => x"7a",
           999 => x"3f",
          1000 => x"1b",
          1001 => x"38",
          1002 => x"5b",
          1003 => x"33",
          1004 => x"80",
          1005 => x"84",
          1006 => x"08",
          1007 => x"8c",
          1008 => x"51",
          1009 => x"60",
          1010 => x"81",
          1011 => x"e7",
          1012 => x"26",
          1013 => x"5e",
          1014 => x"7a",
          1015 => x"2e",
          1016 => x"83",
          1017 => x"3f",
          1018 => x"57",
          1019 => x"80",
          1020 => x"51",
          1021 => x"84",
          1022 => x"72",
          1023 => x"80",
          1024 => x"5a",
          1025 => x"8d",
          1026 => x"5c",
          1027 => x"32",
          1028 => x"f8",
          1029 => x"7d",
          1030 => x"e0",
          1031 => x"f8",
          1032 => x"3f",
          1033 => x"81",
          1034 => x"38",
          1035 => x"d1",
          1036 => x"ba",
          1037 => x"0b",
          1038 => x"9c",
          1039 => x"f7",
          1040 => x"2e",
          1041 => x"df",
          1042 => x"33",
          1043 => x"82",
          1044 => x"91",
          1045 => x"9d",
          1046 => x"80",
          1047 => x"52",
          1048 => x"5a",
          1049 => x"7c",
          1050 => x"78",
          1051 => x"10",
          1052 => x"08",
          1053 => x"3f",
          1054 => x"80",
          1055 => x"53",
          1056 => x"85",
          1057 => x"2e",
          1058 => x"70",
          1059 => x"39",
          1060 => x"7d",
          1061 => x"39",
          1062 => x"d6",
          1063 => x"52",
          1064 => x"39",
          1065 => x"9a",
          1066 => x"83",
          1067 => x"81",
          1068 => x"d6",
          1069 => x"78",
          1070 => x"3f",
          1071 => x"3d",
          1072 => x"51",
          1073 => x"80",
          1074 => x"d6",
          1075 => x"79",
          1076 => x"fa",
          1077 => x"83",
          1078 => x"8b",
          1079 => x"ff",
          1080 => x"ba",
          1081 => x"68",
          1082 => x"3f",
          1083 => x"f4",
          1084 => x"9e",
          1085 => x"f9",
          1086 => x"53",
          1087 => x"84",
          1088 => x"59",
          1089 => x"b0",
          1090 => x"08",
          1091 => x"87",
          1092 => x"ae",
          1093 => x"87",
          1094 => x"59",
          1095 => x"53",
          1096 => x"84",
          1097 => x"38",
          1098 => x"80",
          1099 => x"8c",
          1100 => x"22",
          1101 => x"cf",
          1102 => x"80",
          1103 => x"7e",
          1104 => x"f8",
          1105 => x"38",
          1106 => x"39",
          1107 => x"80",
          1108 => x"8c",
          1109 => x"3d",
          1110 => x"51",
          1111 => x"80",
          1112 => x"f8",
          1113 => x"ba",
          1114 => x"f7",
          1115 => x"ac",
          1116 => x"27",
          1117 => x"33",
          1118 => x"38",
          1119 => x"78",
          1120 => x"3f",
          1121 => x"1b",
          1122 => x"84",
          1123 => x"ea",
          1124 => x"f7",
          1125 => x"53",
          1126 => x"84",
          1127 => x"38",
          1128 => x"80",
          1129 => x"8c",
          1130 => x"d7",
          1131 => x"79",
          1132 => x"79",
          1133 => x"65",
          1134 => x"ff",
          1135 => x"e8",
          1136 => x"2e",
          1137 => x"11",
          1138 => x"3f",
          1139 => x"70",
          1140 => x"cc",
          1141 => x"80",
          1142 => x"7e",
          1143 => x"f6",
          1144 => x"38",
          1145 => x"59",
          1146 => x"68",
          1147 => x"11",
          1148 => x"3f",
          1149 => x"d3",
          1150 => x"33",
          1151 => x"3d",
          1152 => x"51",
          1153 => x"ff",
          1154 => x"ff",
          1155 => x"e6",
          1156 => x"2e",
          1157 => x"11",
          1158 => x"3f",
          1159 => x"83",
          1160 => x"ff",
          1161 => x"ba",
          1162 => x"08",
          1163 => x"3f",
          1164 => x"8f",
          1165 => x"05",
          1166 => x"8a",
          1167 => x"b8",
          1168 => x"3f",
          1169 => x"80",
          1170 => x"53",
          1171 => x"e9",
          1172 => x"2e",
          1173 => x"51",
          1174 => x"3d",
          1175 => x"51",
          1176 => x"91",
          1177 => x"80",
          1178 => x"08",
          1179 => x"ff",
          1180 => x"ba",
          1181 => x"33",
          1182 => x"83",
          1183 => x"f8",
          1184 => x"82",
          1185 => x"a5",
          1186 => x"2e",
          1187 => x"70",
          1188 => x"06",
          1189 => x"38",
          1190 => x"83",
          1191 => x"55",
          1192 => x"51",
          1193 => x"d6",
          1194 => x"71",
          1195 => x"3d",
          1196 => x"51",
          1197 => x"80",
          1198 => x"0c",
          1199 => x"fe",
          1200 => x"e1",
          1201 => x"38",
          1202 => x"ce",
          1203 => x"23",
          1204 => x"53",
          1205 => x"84",
          1206 => x"38",
          1207 => x"7e",
          1208 => x"b8",
          1209 => x"05",
          1210 => x"08",
          1211 => x"3d",
          1212 => x"51",
          1213 => x"80",
          1214 => x"80",
          1215 => x"05",
          1216 => x"f0",
          1217 => x"f6",
          1218 => x"81",
          1219 => x"64",
          1220 => x"39",
          1221 => x"93",
          1222 => x"80",
          1223 => x"c8",
          1224 => x"7c",
          1225 => x"83",
          1226 => x"eb",
          1227 => x"ff",
          1228 => x"ba",
          1229 => x"59",
          1230 => x"82",
          1231 => x"39",
          1232 => x"2e",
          1233 => x"47",
          1234 => x"5c",
          1235 => x"d0",
          1236 => x"f0",
          1237 => x"b6",
          1238 => x"3f",
          1239 => x"92",
          1240 => x"83",
          1241 => x"83",
          1242 => x"c6",
          1243 => x"80",
          1244 => x"47",
          1245 => x"5e",
          1246 => x"e0",
          1247 => x"93",
          1248 => x"83",
          1249 => x"83",
          1250 => x"9b",
          1251 => x"b9",
          1252 => x"80",
          1253 => x"47",
          1254 => x"fc",
          1255 => x"f2",
          1256 => x"39",
          1257 => x"bc",
          1258 => x"56",
          1259 => x"da",
          1260 => x"2b",
          1261 => x"52",
          1262 => x"ba",
          1263 => x"94",
          1264 => x"80",
          1265 => x"ba",
          1266 => x"55",
          1267 => x"89",
          1268 => x"77",
          1269 => x"94",
          1270 => x"c0",
          1271 => x"81",
          1272 => x"a1",
          1273 => x"0b",
          1274 => x"72",
          1275 => x"f5",
          1276 => x"ba",
          1277 => x"f8",
          1278 => x"3f",
          1279 => x"94",
          1280 => x"d3",
          1281 => x"d3",
          1282 => x"3f",
          1283 => x"0d",
          1284 => x"52",
          1285 => x"74",
          1286 => x"70",
          1287 => x"81",
          1288 => x"53",
          1289 => x"71",
          1290 => x"81",
          1291 => x"80",
          1292 => x"ff",
          1293 => x"83",
          1294 => x"38",
          1295 => x"52",
          1296 => x"52",
          1297 => x"83",
          1298 => x"30",
          1299 => x"53",
          1300 => x"70",
          1301 => x"74",
          1302 => x"3d",
          1303 => x"73",
          1304 => x"52",
          1305 => x"53",
          1306 => x"81",
          1307 => x"75",
          1308 => x"06",
          1309 => x"0d",
          1310 => x"0b",
          1311 => x"04",
          1312 => x"da",
          1313 => x"2e",
          1314 => x"86",
          1315 => x"82",
          1316 => x"52",
          1317 => x"13",
          1318 => x"9e",
          1319 => x"51",
          1320 => x"38",
          1321 => x"bb",
          1322 => x"55",
          1323 => x"38",
          1324 => x"87",
          1325 => x"22",
          1326 => x"80",
          1327 => x"9c",
          1328 => x"0c",
          1329 => x"0c",
          1330 => x"0c",
          1331 => x"0c",
          1332 => x"0c",
          1333 => x"0c",
          1334 => x"87",
          1335 => x"c0",
          1336 => x"ba",
          1337 => x"3d",
          1338 => x"5d",
          1339 => x"08",
          1340 => x"b8",
          1341 => x"c0",
          1342 => x"34",
          1343 => x"84",
          1344 => x"5a",
          1345 => x"a8",
          1346 => x"c0",
          1347 => x"23",
          1348 => x"8a",
          1349 => x"ff",
          1350 => x"06",
          1351 => x"33",
          1352 => x"33",
          1353 => x"ff",
          1354 => x"ff",
          1355 => x"fe",
          1356 => x"72",
          1357 => x"e8",
          1358 => x"2b",
          1359 => x"2e",
          1360 => x"2e",
          1361 => x"84",
          1362 => x"8a",
          1363 => x"70",
          1364 => x"09",
          1365 => x"e7",
          1366 => x"2b",
          1367 => x"2e",
          1368 => x"80",
          1369 => x"81",
          1370 => x"8c",
          1371 => x"52",
          1372 => x"07",
          1373 => x"db",
          1374 => x"3d",
          1375 => x"05",
          1376 => x"ff",
          1377 => x"80",
          1378 => x"70",
          1379 => x"52",
          1380 => x"2a",
          1381 => x"38",
          1382 => x"80",
          1383 => x"06",
          1384 => x"06",
          1385 => x"80",
          1386 => x"52",
          1387 => x"0c",
          1388 => x"70",
          1389 => x"72",
          1390 => x"2e",
          1391 => x"52",
          1392 => x"94",
          1393 => x"06",
          1394 => x"39",
          1395 => x"70",
          1396 => x"70",
          1397 => x"04",
          1398 => x"33",
          1399 => x"80",
          1400 => x"33",
          1401 => x"71",
          1402 => x"94",
          1403 => x"06",
          1404 => x"38",
          1405 => x"51",
          1406 => x"06",
          1407 => x"93",
          1408 => x"75",
          1409 => x"80",
          1410 => x"c0",
          1411 => x"17",
          1412 => x"38",
          1413 => x"0d",
          1414 => x"51",
          1415 => x"81",
          1416 => x"71",
          1417 => x"2e",
          1418 => x"08",
          1419 => x"54",
          1420 => x"3d",
          1421 => x"9c",
          1422 => x"2e",
          1423 => x"08",
          1424 => x"a8",
          1425 => x"9e",
          1426 => x"c0",
          1427 => x"87",
          1428 => x"0c",
          1429 => x"dc",
          1430 => x"f2",
          1431 => x"83",
          1432 => x"08",
          1433 => x"b8",
          1434 => x"9e",
          1435 => x"c0",
          1436 => x"87",
          1437 => x"0c",
          1438 => x"83",
          1439 => x"08",
          1440 => x"88",
          1441 => x"9e",
          1442 => x"0b",
          1443 => x"c0",
          1444 => x"06",
          1445 => x"71",
          1446 => x"c0",
          1447 => x"06",
          1448 => x"38",
          1449 => x"80",
          1450 => x"90",
          1451 => x"80",
          1452 => x"f3",
          1453 => x"90",
          1454 => x"52",
          1455 => x"52",
          1456 => x"87",
          1457 => x"80",
          1458 => x"83",
          1459 => x"34",
          1460 => x"70",
          1461 => x"70",
          1462 => x"83",
          1463 => x"9e",
          1464 => x"51",
          1465 => x"81",
          1466 => x"0b",
          1467 => x"80",
          1468 => x"2e",
          1469 => x"94",
          1470 => x"08",
          1471 => x"52",
          1472 => x"71",
          1473 => x"c0",
          1474 => x"06",
          1475 => x"38",
          1476 => x"80",
          1477 => x"a0",
          1478 => x"2e",
          1479 => x"97",
          1480 => x"80",
          1481 => x"83",
          1482 => x"9e",
          1483 => x"52",
          1484 => x"52",
          1485 => x"9e",
          1486 => x"2a",
          1487 => x"80",
          1488 => x"88",
          1489 => x"83",
          1490 => x"34",
          1491 => x"51",
          1492 => x"0d",
          1493 => x"3d",
          1494 => x"d4",
          1495 => x"86",
          1496 => x"af",
          1497 => x"85",
          1498 => x"73",
          1499 => x"56",
          1500 => x"33",
          1501 => x"92",
          1502 => x"f3",
          1503 => x"83",
          1504 => x"38",
          1505 => x"ed",
          1506 => x"83",
          1507 => x"73",
          1508 => x"55",
          1509 => x"33",
          1510 => x"96",
          1511 => x"d9",
          1512 => x"f0",
          1513 => x"b5",
          1514 => x"83",
          1515 => x"83",
          1516 => x"51",
          1517 => x"51",
          1518 => x"52",
          1519 => x"3f",
          1520 => x"c0",
          1521 => x"ba",
          1522 => x"71",
          1523 => x"52",
          1524 => x"3f",
          1525 => x"c3",
          1526 => x"8a",
          1527 => x"3d",
          1528 => x"bd",
          1529 => x"3f",
          1530 => x"29",
          1531 => x"8c",
          1532 => x"b4",
          1533 => x"87",
          1534 => x"56",
          1535 => x"a9",
          1536 => x"c0",
          1537 => x"ba",
          1538 => x"ff",
          1539 => x"55",
          1540 => x"9a",
          1541 => x"3f",
          1542 => x"83",
          1543 => x"51",
          1544 => x"08",
          1545 => x"bc",
          1546 => x"da",
          1547 => x"da",
          1548 => x"fc",
          1549 => x"b3",
          1550 => x"bd",
          1551 => x"3f",
          1552 => x"29",
          1553 => x"8c",
          1554 => x"b2",
          1555 => x"74",
          1556 => x"39",
          1557 => x"3f",
          1558 => x"2e",
          1559 => x"dc",
          1560 => x"f3",
          1561 => x"e5",
          1562 => x"ff",
          1563 => x"55",
          1564 => x"39",
          1565 => x"3f",
          1566 => x"2e",
          1567 => x"9a",
          1568 => x"b2",
          1569 => x"75",
          1570 => x"83",
          1571 => x"51",
          1572 => x"33",
          1573 => x"cd",
          1574 => x"dc",
          1575 => x"f3",
          1576 => x"c0",
          1577 => x"83",
          1578 => x"dd",
          1579 => x"f3",
          1580 => x"97",
          1581 => x"83",
          1582 => x"dd",
          1583 => x"f3",
          1584 => x"ee",
          1585 => x"83",
          1586 => x"dd",
          1587 => x"f3",
          1588 => x"c5",
          1589 => x"83",
          1590 => x"dd",
          1591 => x"f3",
          1592 => x"9c",
          1593 => x"83",
          1594 => x"dd",
          1595 => x"f3",
          1596 => x"f3",
          1597 => x"ff",
          1598 => x"ff",
          1599 => x"55",
          1600 => x"39",
          1601 => x"52",
          1602 => x"10",
          1603 => x"04",
          1604 => x"3f",
          1605 => x"51",
          1606 => x"04",
          1607 => x"3f",
          1608 => x"51",
          1609 => x"04",
          1610 => x"3f",
          1611 => x"51",
          1612 => x"04",
          1613 => x"87",
          1614 => x"a0",
          1615 => x"d9",
          1616 => x"08",
          1617 => x"52",
          1618 => x"d2",
          1619 => x"38",
          1620 => x"f8",
          1621 => x"51",
          1622 => x"08",
          1623 => x"ec",
          1624 => x"57",
          1625 => x"25",
          1626 => x"05",
          1627 => x"74",
          1628 => x"2a",
          1629 => x"38",
          1630 => x"08",
          1631 => x"ea",
          1632 => x"78",
          1633 => x"8c",
          1634 => x"84",
          1635 => x"2e",
          1636 => x"79",
          1637 => x"bf",
          1638 => x"ba",
          1639 => x"e2",
          1640 => x"0b",
          1641 => x"04",
          1642 => x"3d",
          1643 => x"57",
          1644 => x"38",
          1645 => x"10",
          1646 => x"08",
          1647 => x"ba",
          1648 => x"51",
          1649 => x"90",
          1650 => x"2e",
          1651 => x"38",
          1652 => x"54",
          1653 => x"73",
          1654 => x"04",
          1655 => x"11",
          1656 => x"3f",
          1657 => x"38",
          1658 => x"fd",
          1659 => x"ff",
          1660 => x"81",
          1661 => x"82",
          1662 => x"39",
          1663 => x"27",
          1664 => x"70",
          1665 => x"81",
          1666 => x"eb",
          1667 => x"fe",
          1668 => x"53",
          1669 => x"85",
          1670 => x"d0",
          1671 => x"f8",
          1672 => x"84",
          1673 => x"77",
          1674 => x"8c",
          1675 => x"08",
          1676 => x"ff",
          1677 => x"34",
          1678 => x"e1",
          1679 => x"74",
          1680 => x"38",
          1681 => x"3d",
          1682 => x"08",
          1683 => x"41",
          1684 => x"f3",
          1685 => x"5d",
          1686 => x"33",
          1687 => x"38",
          1688 => x"70",
          1689 => x"38",
          1690 => x"3d",
          1691 => x"ff",
          1692 => x"70",
          1693 => x"ec",
          1694 => x"c8",
          1695 => x"84",
          1696 => x"97",
          1697 => x"10",
          1698 => x"70",
          1699 => x"5b",
          1700 => x"2e",
          1701 => x"87",
          1702 => x"ff",
          1703 => x"80",
          1704 => x"16",
          1705 => x"83",
          1706 => x"61",
          1707 => x"08",
          1708 => x"2e",
          1709 => x"38",
          1710 => x"76",
          1711 => x"70",
          1712 => x"c4",
          1713 => x"71",
          1714 => x"de",
          1715 => x"58",
          1716 => x"90",
          1717 => x"ac",
          1718 => x"75",
          1719 => x"05",
          1720 => x"59",
          1721 => x"38",
          1722 => x"55",
          1723 => x"42",
          1724 => x"de",
          1725 => x"55",
          1726 => x"80",
          1727 => x"81",
          1728 => x"fe",
          1729 => x"80",
          1730 => x"d1",
          1731 => x"79",
          1732 => x"74",
          1733 => x"10",
          1734 => x"04",
          1735 => x"80",
          1736 => x"84",
          1737 => x"d0",
          1738 => x"38",
          1739 => x"ff",
          1740 => x"ff",
          1741 => x"fc",
          1742 => x"81",
          1743 => x"57",
          1744 => x"84",
          1745 => x"77",
          1746 => x"33",
          1747 => x"bc",
          1748 => x"7c",
          1749 => x"08",
          1750 => x"84",
          1751 => x"d1",
          1752 => x"56",
          1753 => x"f0",
          1754 => x"3f",
          1755 => x"ff",
          1756 => x"52",
          1757 => x"d1",
          1758 => x"d1",
          1759 => x"74",
          1760 => x"3f",
          1761 => x"39",
          1762 => x"56",
          1763 => x"83",
          1764 => x"55",
          1765 => x"75",
          1766 => x"ff",
          1767 => x"84",
          1768 => x"81",
          1769 => x"7b",
          1770 => x"cc",
          1771 => x"74",
          1772 => x"f0",
          1773 => x"3f",
          1774 => x"ff",
          1775 => x"52",
          1776 => x"d1",
          1777 => x"d1",
          1778 => x"c7",
          1779 => x"ff",
          1780 => x"55",
          1781 => x"d5",
          1782 => x"84",
          1783 => x"52",
          1784 => x"d0",
          1785 => x"cc",
          1786 => x"fa",
          1787 => x"81",
          1788 => x"7b",
          1789 => x"82",
          1790 => x"ff",
          1791 => x"55",
          1792 => x"d4",
          1793 => x"cc",
          1794 => x"c4",
          1795 => x"cc",
          1796 => x"7c",
          1797 => x"76",
          1798 => x"08",
          1799 => x"84",
          1800 => x"98",
          1801 => x"57",
          1802 => x"84",
          1803 => x"b2",
          1804 => x"81",
          1805 => x"d1",
          1806 => x"24",
          1807 => x"52",
          1808 => x"81",
          1809 => x"70",
          1810 => x"56",
          1811 => x"f8",
          1812 => x"33",
          1813 => x"77",
          1814 => x"81",
          1815 => x"70",
          1816 => x"57",
          1817 => x"7b",
          1818 => x"84",
          1819 => x"ff",
          1820 => x"29",
          1821 => x"84",
          1822 => x"76",
          1823 => x"84",
          1824 => x"f7",
          1825 => x"88",
          1826 => x"d0",
          1827 => x"d0",
          1828 => x"39",
          1829 => x"80",
          1830 => x"8a",
          1831 => x"cc",
          1832 => x"ba",
          1833 => x"89",
          1834 => x"76",
          1835 => x"fc",
          1836 => x"05",
          1837 => x"a0",
          1838 => x"83",
          1839 => x"57",
          1840 => x"8c",
          1841 => x"70",
          1842 => x"08",
          1843 => x"83",
          1844 => x"8c",
          1845 => x"80",
          1846 => x"d1",
          1847 => x"34",
          1848 => x"0d",
          1849 => x"80",
          1850 => x"52",
          1851 => x"d5",
          1852 => x"8a",
          1853 => x"51",
          1854 => x"33",
          1855 => x"34",
          1856 => x"38",
          1857 => x"3f",
          1858 => x"0b",
          1859 => x"83",
          1860 => x"84",
          1861 => x"b6",
          1862 => x"51",
          1863 => x"08",
          1864 => x"84",
          1865 => x"ae",
          1866 => x"05",
          1867 => x"81",
          1868 => x"d2",
          1869 => x"0b",
          1870 => x"d1",
          1871 => x"b4",
          1872 => x"70",
          1873 => x"2e",
          1874 => x"ff",
          1875 => x"ff",
          1876 => x"84",
          1877 => x"ad",
          1878 => x"98",
          1879 => x"33",
          1880 => x"80",
          1881 => x"a0",
          1882 => x"d0",
          1883 => x"84",
          1884 => x"74",
          1885 => x"f0",
          1886 => x"3f",
          1887 => x"0a",
          1888 => x"33",
          1889 => x"cc",
          1890 => x"51",
          1891 => x"0a",
          1892 => x"2c",
          1893 => x"78",
          1894 => x"39",
          1895 => x"34",
          1896 => x"51",
          1897 => x"0a",
          1898 => x"2c",
          1899 => x"75",
          1900 => x"57",
          1901 => x"f0",
          1902 => x"fa",
          1903 => x"80",
          1904 => x"cc",
          1905 => x"ff",
          1906 => x"d0",
          1907 => x"76",
          1908 => x"cc",
          1909 => x"74",
          1910 => x"76",
          1911 => x"7a",
          1912 => x"0a",
          1913 => x"2c",
          1914 => x"75",
          1915 => x"74",
          1916 => x"06",
          1917 => x"34",
          1918 => x"25",
          1919 => x"d1",
          1920 => x"33",
          1921 => x"0a",
          1922 => x"06",
          1923 => x"81",
          1924 => x"2c",
          1925 => x"75",
          1926 => x"f0",
          1927 => x"3f",
          1928 => x"0a",
          1929 => x"33",
          1930 => x"84",
          1931 => x"51",
          1932 => x"0a",
          1933 => x"2c",
          1934 => x"74",
          1935 => x"39",
          1936 => x"2e",
          1937 => x"9c",
          1938 => x"cc",
          1939 => x"06",
          1940 => x"ff",
          1941 => x"84",
          1942 => x"2e",
          1943 => x"52",
          1944 => x"d5",
          1945 => x"a2",
          1946 => x"51",
          1947 => x"33",
          1948 => x"34",
          1949 => x"a8",
          1950 => x"8c",
          1951 => x"8c",
          1952 => x"f4",
          1953 => x"39",
          1954 => x"70",
          1955 => x"75",
          1956 => x"05",
          1957 => x"52",
          1958 => x"84",
          1959 => x"98",
          1960 => x"5a",
          1961 => x"fd",
          1962 => x"2e",
          1963 => x"93",
          1964 => x"ff",
          1965 => x"25",
          1966 => x"34",
          1967 => x"2e",
          1968 => x"c5",
          1969 => x"da",
          1970 => x"0c",
          1971 => x"bc",
          1972 => x"80",
          1973 => x"56",
          1974 => x"ba",
          1975 => x"84",
          1976 => x"84",
          1977 => x"05",
          1978 => x"96",
          1979 => x"84",
          1980 => x"80",
          1981 => x"08",
          1982 => x"84",
          1983 => x"a6",
          1984 => x"88",
          1985 => x"d0",
          1986 => x"d0",
          1987 => x"39",
          1988 => x"d0",
          1989 => x"7b",
          1990 => x"04",
          1991 => x"ba",
          1992 => x"ba",
          1993 => x"53",
          1994 => x"3f",
          1995 => x"d1",
          1996 => x"52",
          1997 => x"38",
          1998 => x"ff",
          1999 => x"52",
          2000 => x"d5",
          2001 => x"e2",
          2002 => x"57",
          2003 => x"ff",
          2004 => x"a9",
          2005 => x"d1",
          2006 => x"ff",
          2007 => x"51",
          2008 => x"81",
          2009 => x"d1",
          2010 => x"80",
          2011 => x"08",
          2012 => x"84",
          2013 => x"a5",
          2014 => x"88",
          2015 => x"d0",
          2016 => x"d0",
          2017 => x"39",
          2018 => x"f3",
          2019 => x"06",
          2020 => x"54",
          2021 => x"84",
          2022 => x"fc",
          2023 => x"05",
          2024 => x"2e",
          2025 => x"74",
          2026 => x"fc",
          2027 => x"5a",
          2028 => x"77",
          2029 => x"b4",
          2030 => x"7b",
          2031 => x"83",
          2032 => x"ba",
          2033 => x"81",
          2034 => x"d0",
          2035 => x"7b",
          2036 => x"04",
          2037 => x"08",
          2038 => x"8c",
          2039 => x"08",
          2040 => x"08",
          2041 => x"b8",
          2042 => x"84",
          2043 => x"06",
          2044 => x"51",
          2045 => x"08",
          2046 => x"25",
          2047 => x"ff",
          2048 => x"34",
          2049 => x"33",
          2050 => x"70",
          2051 => x"f2",
          2052 => x"83",
          2053 => x"58",
          2054 => x"8c",
          2055 => x"70",
          2056 => x"08",
          2057 => x"1d",
          2058 => x"7d",
          2059 => x"2e",
          2060 => x"e8",
          2061 => x"79",
          2062 => x"83",
          2063 => x"ff",
          2064 => x"c8",
          2065 => x"ff",
          2066 => x"3f",
          2067 => x"87",
          2068 => x"1b",
          2069 => x"9e",
          2070 => x"83",
          2071 => x"f3",
          2072 => x"74",
          2073 => x"39",
          2074 => x"39",
          2075 => x"39",
          2076 => x"3f",
          2077 => x"f2",
          2078 => x"02",
          2079 => x"53",
          2080 => x"81",
          2081 => x"83",
          2082 => x"38",
          2083 => x"b0",
          2084 => x"a0",
          2085 => x"83",
          2086 => x"34",
          2087 => x"b8",
          2088 => x"07",
          2089 => x"7f",
          2090 => x"94",
          2091 => x"0c",
          2092 => x"76",
          2093 => x"a2",
          2094 => x"de",
          2095 => x"a0",
          2096 => x"70",
          2097 => x"72",
          2098 => x"a3",
          2099 => x"70",
          2100 => x"71",
          2101 => x"58",
          2102 => x"84",
          2103 => x"84",
          2104 => x"83",
          2105 => x"06",
          2106 => x"5e",
          2107 => x"38",
          2108 => x"81",
          2109 => x"81",
          2110 => x"62",
          2111 => x"5d",
          2112 => x"26",
          2113 => x"76",
          2114 => x"5f",
          2115 => x"fe",
          2116 => x"77",
          2117 => x"81",
          2118 => x"74",
          2119 => x"87",
          2120 => x"80",
          2121 => x"ff",
          2122 => x"ff",
          2123 => x"29",
          2124 => x"57",
          2125 => x"81",
          2126 => x"71",
          2127 => x"2e",
          2128 => x"bc",
          2129 => x"83",
          2130 => x"90",
          2131 => x"07",
          2132 => x"79",
          2133 => x"72",
          2134 => x"70",
          2135 => x"83",
          2136 => x"87",
          2137 => x"56",
          2138 => x"14",
          2139 => x"06",
          2140 => x"06",
          2141 => x"ff",
          2142 => x"5a",
          2143 => x"79",
          2144 => x"15",
          2145 => x"81",
          2146 => x"71",
          2147 => x"81",
          2148 => x"5b",
          2149 => x"38",
          2150 => x"16",
          2151 => x"e2",
          2152 => x"da",
          2153 => x"7b",
          2154 => x"0d",
          2155 => x"74",
          2156 => x"80",
          2157 => x"34",
          2158 => x"34",
          2159 => x"86",
          2160 => x"34",
          2161 => x"75",
          2162 => x"3f",
          2163 => x"54",
          2164 => x"73",
          2165 => x"75",
          2166 => x"80",
          2167 => x"87",
          2168 => x"81",
          2169 => x"f3",
          2170 => x"07",
          2171 => x"84",
          2172 => x"8c",
          2173 => x"80",
          2174 => x"3d",
          2175 => x"05",
          2176 => x"5b",
          2177 => x"82",
          2178 => x"f9",
          2179 => x"71",
          2180 => x"83",
          2181 => x"71",
          2182 => x"06",
          2183 => x"53",
          2184 => x"f9",
          2185 => x"f9",
          2186 => x"05",
          2187 => x"06",
          2188 => x"8c",
          2189 => x"bc",
          2190 => x"ff",
          2191 => x"55",
          2192 => x"84",
          2193 => x"58",
          2194 => x"38",
          2195 => x"e0",
          2196 => x"72",
          2197 => x"81",
          2198 => x"b7",
          2199 => x"9f",
          2200 => x"84",
          2201 => x"e0",
          2202 => x"05",
          2203 => x"74",
          2204 => x"ff",
          2205 => x"75",
          2206 => x"ff",
          2207 => x"81",
          2208 => x"84",
          2209 => x"55",
          2210 => x"58",
          2211 => x"06",
          2212 => x"19",
          2213 => x"b9",
          2214 => x"e0",
          2215 => x"33",
          2216 => x"70",
          2217 => x"05",
          2218 => x"33",
          2219 => x"19",
          2220 => x"ce",
          2221 => x"0c",
          2222 => x"bc",
          2223 => x"ff",
          2224 => x"55",
          2225 => x"77",
          2226 => x"ff",
          2227 => x"56",
          2228 => x"fe",
          2229 => x"84",
          2230 => x"72",
          2231 => x"73",
          2232 => x"33",
          2233 => x"55",
          2234 => x"34",
          2235 => x"ff",
          2236 => x"38",
          2237 => x"75",
          2238 => x"53",
          2239 => x"0b",
          2240 => x"89",
          2241 => x"84",
          2242 => x"b7",
          2243 => x"3d",
          2244 => x"33",
          2245 => x"70",
          2246 => x"70",
          2247 => x"71",
          2248 => x"bd",
          2249 => x"86",
          2250 => x"bd",
          2251 => x"ff",
          2252 => x"38",
          2253 => x"34",
          2254 => x"3d",
          2255 => x"73",
          2256 => x"06",
          2257 => x"bc",
          2258 => x"72",
          2259 => x"55",
          2260 => x"70",
          2261 => x"0b",
          2262 => x"04",
          2263 => x"70",
          2264 => x"56",
          2265 => x"80",
          2266 => x"0d",
          2267 => x"84",
          2268 => x"51",
          2269 => x"72",
          2270 => x"ba",
          2271 => x"0b",
          2272 => x"33",
          2273 => x"52",
          2274 => x"12",
          2275 => x"d0",
          2276 => x"33",
          2277 => x"10",
          2278 => x"08",
          2279 => x"f0",
          2280 => x"70",
          2281 => x"51",
          2282 => x"9c",
          2283 => x"34",
          2284 => x"3d",
          2285 => x"9f",
          2286 => x"b8",
          2287 => x"83",
          2288 => x"80",
          2289 => x"34",
          2290 => x"fe",
          2291 => x"b8",
          2292 => x"f9",
          2293 => x"0c",
          2294 => x"33",
          2295 => x"83",
          2296 => x"f9",
          2297 => x"f9",
          2298 => x"b8",
          2299 => x"70",
          2300 => x"83",
          2301 => x"07",
          2302 => x"81",
          2303 => x"06",
          2304 => x"34",
          2305 => x"81",
          2306 => x"34",
          2307 => x"81",
          2308 => x"83",
          2309 => x"f9",
          2310 => x"51",
          2311 => x"39",
          2312 => x"80",
          2313 => x"34",
          2314 => x"81",
          2315 => x"83",
          2316 => x"f9",
          2317 => x"51",
          2318 => x"39",
          2319 => x"51",
          2320 => x"39",
          2321 => x"82",
          2322 => x"fd",
          2323 => x"05",
          2324 => x"33",
          2325 => x"33",
          2326 => x"33",
          2327 => x"82",
          2328 => x"a5",
          2329 => x"7d",
          2330 => x"b8",
          2331 => x"7b",
          2332 => x"bd",
          2333 => x"2e",
          2334 => x"84",
          2335 => x"84",
          2336 => x"a8",
          2337 => x"83",
          2338 => x"80",
          2339 => x"84",
          2340 => x"53",
          2341 => x"81",
          2342 => x"80",
          2343 => x"f9",
          2344 => x"7c",
          2345 => x"04",
          2346 => x"0b",
          2347 => x"f9",
          2348 => x"34",
          2349 => x"b9",
          2350 => x"57",
          2351 => x"7b",
          2352 => x"e0",
          2353 => x"84",
          2354 => x"27",
          2355 => x"05",
          2356 => x"51",
          2357 => x"81",
          2358 => x"5b",
          2359 => x"d2",
          2360 => x"84",
          2361 => x"84",
          2362 => x"83",
          2363 => x"34",
          2364 => x"b8",
          2365 => x"34",
          2366 => x"0b",
          2367 => x"f9",
          2368 => x"92",
          2369 => x"83",
          2370 => x"80",
          2371 => x"8c",
          2372 => x"fd",
          2373 => x"52",
          2374 => x"3f",
          2375 => x"5a",
          2376 => x"84",
          2377 => x"33",
          2378 => x"33",
          2379 => x"80",
          2380 => x"59",
          2381 => x"ff",
          2382 => x"59",
          2383 => x"81",
          2384 => x"38",
          2385 => x"81",
          2386 => x"82",
          2387 => x"f9",
          2388 => x"72",
          2389 => x"88",
          2390 => x"34",
          2391 => x"33",
          2392 => x"12",
          2393 => x"be",
          2394 => x"71",
          2395 => x"33",
          2396 => x"b8",
          2397 => x"f9",
          2398 => x"72",
          2399 => x"83",
          2400 => x"34",
          2401 => x"55",
          2402 => x"b8",
          2403 => x"ff",
          2404 => x"84",
          2405 => x"8c",
          2406 => x"80",
          2407 => x"ba",
          2408 => x"8d",
          2409 => x"f7",
          2410 => x"fe",
          2411 => x"96",
          2412 => x"ff",
          2413 => x"53",
          2414 => x"75",
          2415 => x"38",
          2416 => x"ba",
          2417 => x"54",
          2418 => x"76",
          2419 => x"13",
          2420 => x"73",
          2421 => x"83",
          2422 => x"52",
          2423 => x"84",
          2424 => x"75",
          2425 => x"ca",
          2426 => x"ff",
          2427 => x"38",
          2428 => x"76",
          2429 => x"f9",
          2430 => x"ff",
          2431 => x"53",
          2432 => x"39",
          2433 => x"52",
          2434 => x"39",
          2435 => x"fe",
          2436 => x"f3",
          2437 => x"59",
          2438 => x"82",
          2439 => x"84",
          2440 => x"38",
          2441 => x"89",
          2442 => x"33",
          2443 => x"33",
          2444 => x"84",
          2445 => x"80",
          2446 => x"f9",
          2447 => x"71",
          2448 => x"83",
          2449 => x"33",
          2450 => x"83",
          2451 => x"80",
          2452 => x"81",
          2453 => x"f9",
          2454 => x"40",
          2455 => x"84",
          2456 => x"81",
          2457 => x"81",
          2458 => x"79",
          2459 => x"83",
          2460 => x"8c",
          2461 => x"2e",
          2462 => x"fd",
          2463 => x"78",
          2464 => x"0b",
          2465 => x"33",
          2466 => x"33",
          2467 => x"84",
          2468 => x"80",
          2469 => x"f9",
          2470 => x"71",
          2471 => x"83",
          2472 => x"33",
          2473 => x"f9",
          2474 => x"34",
          2475 => x"06",
          2476 => x"33",
          2477 => x"58",
          2478 => x"98",
          2479 => x"81",
          2480 => x"ca",
          2481 => x"0b",
          2482 => x"04",
          2483 => x"9b",
          2484 => x"09",
          2485 => x"83",
          2486 => x"8c",
          2487 => x"2e",
          2488 => x"89",
          2489 => x"33",
          2490 => x"8c",
          2491 => x"77",
          2492 => x"b9",
          2493 => x"8c",
          2494 => x"2e",
          2495 => x"88",
          2496 => x"bc",
          2497 => x"29",
          2498 => x"19",
          2499 => x"84",
          2500 => x"83",
          2501 => x"41",
          2502 => x"1f",
          2503 => x"29",
          2504 => x"87",
          2505 => x"80",
          2506 => x"ba",
          2507 => x"29",
          2508 => x"f9",
          2509 => x"34",
          2510 => x"52",
          2511 => x"83",
          2512 => x"b8",
          2513 => x"81",
          2514 => x"71",
          2515 => x"83",
          2516 => x"7e",
          2517 => x"83",
          2518 => x"5c",
          2519 => x"81",
          2520 => x"fc",
          2521 => x"bd",
          2522 => x"b9",
          2523 => x"34",
          2524 => x"0b",
          2525 => x"b9",
          2526 => x"0c",
          2527 => x"33",
          2528 => x"33",
          2529 => x"33",
          2530 => x"b9",
          2531 => x"0c",
          2532 => x"2e",
          2533 => x"f9",
          2534 => x"81",
          2535 => x"81",
          2536 => x"a3",
          2537 => x"5c",
          2538 => x"ff",
          2539 => x"5c",
          2540 => x"2e",
          2541 => x"ff",
          2542 => x"57",
          2543 => x"ff",
          2544 => x"ff",
          2545 => x"5b",
          2546 => x"80",
          2547 => x"f9",
          2548 => x"71",
          2549 => x"0b",
          2550 => x"bc",
          2551 => x"56",
          2552 => x"80",
          2553 => x"81",
          2554 => x"f9",
          2555 => x"5d",
          2556 => x"7f",
          2557 => x"70",
          2558 => x"26",
          2559 => x"5a",
          2560 => x"77",
          2561 => x"33",
          2562 => x"56",
          2563 => x"d8",
          2564 => x"78",
          2565 => x"8c",
          2566 => x"bf",
          2567 => x"38",
          2568 => x"58",
          2569 => x"bd",
          2570 => x"3f",
          2571 => x"3d",
          2572 => x"b8",
          2573 => x"f9",
          2574 => x"75",
          2575 => x"83",
          2576 => x"29",
          2577 => x"f8",
          2578 => x"5b",
          2579 => x"80",
          2580 => x"ff",
          2581 => x"29",
          2582 => x"33",
          2583 => x"b8",
          2584 => x"f9",
          2585 => x"41",
          2586 => x"1c",
          2587 => x"29",
          2588 => x"87",
          2589 => x"80",
          2590 => x"ba",
          2591 => x"29",
          2592 => x"f9",
          2593 => x"60",
          2594 => x"58",
          2595 => x"b8",
          2596 => x"ff",
          2597 => x"81",
          2598 => x"7b",
          2599 => x"bc",
          2600 => x"bd",
          2601 => x"ff",
          2602 => x"29",
          2603 => x"84",
          2604 => x"1b",
          2605 => x"bd",
          2606 => x"29",
          2607 => x"83",
          2608 => x"33",
          2609 => x"f9",
          2610 => x"34",
          2611 => x"06",
          2612 => x"33",
          2613 => x"40",
          2614 => x"de",
          2615 => x"ff",
          2616 => x"d6",
          2617 => x"df",
          2618 => x"80",
          2619 => x"0d",
          2620 => x"84",
          2621 => x"f9",
          2622 => x"ff",
          2623 => x"84",
          2624 => x"8c",
          2625 => x"be",
          2626 => x"33",
          2627 => x"b8",
          2628 => x"5b",
          2629 => x"b9",
          2630 => x"d8",
          2631 => x"ba",
          2632 => x"84",
          2633 => x"75",
          2634 => x"fe",
          2635 => x"61",
          2636 => x"39",
          2637 => x"b8",
          2638 => x"bc",
          2639 => x"bd",
          2640 => x"84",
          2641 => x"83",
          2642 => x"41",
          2643 => x"7f",
          2644 => x"b8",
          2645 => x"f9",
          2646 => x"43",
          2647 => x"34",
          2648 => x"1b",
          2649 => x"87",
          2650 => x"80",
          2651 => x"ba",
          2652 => x"29",
          2653 => x"f9",
          2654 => x"81",
          2655 => x"60",
          2656 => x"81",
          2657 => x"1a",
          2658 => x"0b",
          2659 => x"33",
          2660 => x"84",
          2661 => x"38",
          2662 => x"80",
          2663 => x"0d",
          2664 => x"bc",
          2665 => x"bd",
          2666 => x"83",
          2667 => x"f9",
          2668 => x"f9",
          2669 => x"f9",
          2670 => x"9e",
          2671 => x"80",
          2672 => x"22",
          2673 => x"ff",
          2674 => x"05",
          2675 => x"54",
          2676 => x"3d",
          2677 => x"76",
          2678 => x"8c",
          2679 => x"33",
          2680 => x"fe",
          2681 => x"51",
          2682 => x"80",
          2683 => x"79",
          2684 => x"fe",
          2685 => x"05",
          2686 => x"26",
          2687 => x"c7",
          2688 => x"b9",
          2689 => x"a4",
          2690 => x"e1",
          2691 => x"9f",
          2692 => x"5c",
          2693 => x"39",
          2694 => x"2e",
          2695 => x"ff",
          2696 => x"80",
          2697 => x"fd",
          2698 => x"fd",
          2699 => x"34",
          2700 => x"06",
          2701 => x"38",
          2702 => x"34",
          2703 => x"bd",
          2704 => x"ff",
          2705 => x"25",
          2706 => x"83",
          2707 => x"b9",
          2708 => x"e0",
          2709 => x"e1",
          2710 => x"9f",
          2711 => x"5a",
          2712 => x"39",
          2713 => x"2e",
          2714 => x"41",
          2715 => x"b6",
          2716 => x"bd",
          2717 => x"29",
          2718 => x"f9",
          2719 => x"60",
          2720 => x"83",
          2721 => x"06",
          2722 => x"80",
          2723 => x"f8",
          2724 => x"8d",
          2725 => x"38",
          2726 => x"2e",
          2727 => x"0b",
          2728 => x"84",
          2729 => x"90",
          2730 => x"f9",
          2731 => x"80",
          2732 => x"7d",
          2733 => x"f9",
          2734 => x"8d",
          2735 => x"38",
          2736 => x"33",
          2737 => x"ff",
          2738 => x"83",
          2739 => x"34",
          2740 => x"fe",
          2741 => x"8d",
          2742 => x"c7",
          2743 => x"70",
          2744 => x"fe",
          2745 => x"ff",
          2746 => x"58",
          2747 => x"33",
          2748 => x"84",
          2749 => x"83",
          2750 => x"ff",
          2751 => x"39",
          2752 => x"27",
          2753 => x"ff",
          2754 => x"e1",
          2755 => x"84",
          2756 => x"ff",
          2757 => x"5c",
          2758 => x"79",
          2759 => x"06",
          2760 => x"83",
          2761 => x"34",
          2762 => x"40",
          2763 => x"56",
          2764 => x"39",
          2765 => x"2e",
          2766 => x"84",
          2767 => x"26",
          2768 => x"84",
          2769 => x"83",
          2770 => x"87",
          2771 => x"22",
          2772 => x"83",
          2773 => x"46",
          2774 => x"2e",
          2775 => x"06",
          2776 => x"24",
          2777 => x"56",
          2778 => x"16",
          2779 => x"81",
          2780 => x"80",
          2781 => x"ff",
          2782 => x"38",
          2783 => x"34",
          2784 => x"22",
          2785 => x"90",
          2786 => x"81",
          2787 => x"5b",
          2788 => x"87",
          2789 => x"7f",
          2790 => x"42",
          2791 => x"d6",
          2792 => x"e0",
          2793 => x"33",
          2794 => x"70",
          2795 => x"05",
          2796 => x"33",
          2797 => x"1d",
          2798 => x"f7",
          2799 => x"84",
          2800 => x"05",
          2801 => x"33",
          2802 => x"18",
          2803 => x"33",
          2804 => x"58",
          2805 => x"e6",
          2806 => x"80",
          2807 => x"b9",
          2808 => x"ce",
          2809 => x"ff",
          2810 => x"40",
          2811 => x"b9",
          2812 => x"81",
          2813 => x"33",
          2814 => x"bc",
          2815 => x"2e",
          2816 => x"40",
          2817 => x"81",
          2818 => x"fe",
          2819 => x"07",
          2820 => x"10",
          2821 => x"a3",
          2822 => x"87",
          2823 => x"58",
          2824 => x"83",
          2825 => x"f9",
          2826 => x"2b",
          2827 => x"79",
          2828 => x"27",
          2829 => x"59",
          2830 => x"0c",
          2831 => x"80",
          2832 => x"7e",
          2833 => x"83",
          2834 => x"05",
          2835 => x"8c",
          2836 => x"29",
          2837 => x"57",
          2838 => x"83",
          2839 => x"59",
          2840 => x"79",
          2841 => x"17",
          2842 => x"a0",
          2843 => x"70",
          2844 => x"75",
          2845 => x"ff",
          2846 => x"fe",
          2847 => x"80",
          2848 => x"06",
          2849 => x"7b",
          2850 => x"38",
          2851 => x"81",
          2852 => x"f5",
          2853 => x"5e",
          2854 => x"83",
          2855 => x"83",
          2856 => x"42",
          2857 => x"f9",
          2858 => x"f9",
          2859 => x"06",
          2860 => x"b8",
          2861 => x"75",
          2862 => x"f9",
          2863 => x"56",
          2864 => x"83",
          2865 => x"07",
          2866 => x"39",
          2867 => x"90",
          2868 => x"ff",
          2869 => x"b8",
          2870 => x"59",
          2871 => x"33",
          2872 => x"b8",
          2873 => x"33",
          2874 => x"83",
          2875 => x"f9",
          2876 => x"07",
          2877 => x"ea",
          2878 => x"06",
          2879 => x"b8",
          2880 => x"33",
          2881 => x"83",
          2882 => x"f9",
          2883 => x"56",
          2884 => x"39",
          2885 => x"84",
          2886 => x"fe",
          2887 => x"fa",
          2888 => x"b8",
          2889 => x"33",
          2890 => x"b8",
          2891 => x"33",
          2892 => x"b8",
          2893 => x"33",
          2894 => x"b8",
          2895 => x"33",
          2896 => x"75",
          2897 => x"83",
          2898 => x"07",
          2899 => x"ba",
          2900 => x"80",
          2901 => x"ff",
          2902 => x"bc",
          2903 => x"bd",
          2904 => x"83",
          2905 => x"88",
          2906 => x"b9",
          2907 => x"0c",
          2908 => x"bd",
          2909 => x"ff",
          2910 => x"39",
          2911 => x"11",
          2912 => x"3f",
          2913 => x"ba",
          2914 => x"0b",
          2915 => x"ba",
          2916 => x"83",
          2917 => x"b9",
          2918 => x"84",
          2919 => x"06",
          2920 => x"b9",
          2921 => x"8c",
          2922 => x"bd",
          2923 => x"3f",
          2924 => x"06",
          2925 => x"80",
          2926 => x"81",
          2927 => x"8a",
          2928 => x"39",
          2929 => x"09",
          2930 => x"57",
          2931 => x"d9",
          2932 => x"60",
          2933 => x"bd",
          2934 => x"33",
          2935 => x"72",
          2936 => x"83",
          2937 => x"ff",
          2938 => x"78",
          2939 => x"bb",
          2940 => x"ff",
          2941 => x"a6",
          2942 => x"80",
          2943 => x"bd",
          2944 => x"a0",
          2945 => x"5f",
          2946 => x"ff",
          2947 => x"44",
          2948 => x"f5",
          2949 => x"11",
          2950 => x"38",
          2951 => x"27",
          2952 => x"83",
          2953 => x"ff",
          2954 => x"df",
          2955 => x"76",
          2956 => x"75",
          2957 => x"06",
          2958 => x"5a",
          2959 => x"31",
          2960 => x"71",
          2961 => x"a3",
          2962 => x"7c",
          2963 => x"71",
          2964 => x"79",
          2965 => x"de",
          2966 => x"84",
          2967 => x"05",
          2968 => x"33",
          2969 => x"18",
          2970 => x"33",
          2971 => x"58",
          2972 => x"e0",
          2973 => x"33",
          2974 => x"70",
          2975 => x"05",
          2976 => x"33",
          2977 => x"1d",
          2978 => x"ff",
          2979 => x"be",
          2980 => x"33",
          2981 => x"b8",
          2982 => x"b7",
          2983 => x"e9",
          2984 => x"ff",
          2985 => x"5c",
          2986 => x"76",
          2987 => x"81",
          2988 => x"7a",
          2989 => x"f9",
          2990 => x"81",
          2991 => x"80",
          2992 => x"75",
          2993 => x"83",
          2994 => x"80",
          2995 => x"7f",
          2996 => x"c5",
          2997 => x"f4",
          2998 => x"81",
          2999 => x"44",
          3000 => x"81",
          3001 => x"ff",
          3002 => x"fd",
          3003 => x"f9",
          3004 => x"31",
          3005 => x"90",
          3006 => x"26",
          3007 => x"05",
          3008 => x"70",
          3009 => x"f4",
          3010 => x"58",
          3011 => x"81",
          3012 => x"38",
          3013 => x"75",
          3014 => x"80",
          3015 => x"39",
          3016 => x"39",
          3017 => x"8e",
          3018 => x"f1",
          3019 => x"5a",
          3020 => x"80",
          3021 => x"39",
          3022 => x"84",
          3023 => x"2e",
          3024 => x"80",
          3025 => x"0d",
          3026 => x"3f",
          3027 => x"3d",
          3028 => x"05",
          3029 => x"33",
          3030 => x"11",
          3031 => x"2e",
          3032 => x"83",
          3033 => x"ba",
          3034 => x"f7",
          3035 => x"2e",
          3036 => x"71",
          3037 => x"5d",
          3038 => x"ff",
          3039 => x"81",
          3040 => x"32",
          3041 => x"5c",
          3042 => x"38",
          3043 => x"33",
          3044 => x"12",
          3045 => x"ba",
          3046 => x"05",
          3047 => x"91",
          3048 => x"2e",
          3049 => x"86",
          3050 => x"c0",
          3051 => x"08",
          3052 => x"ee",
          3053 => x"bc",
          3054 => x"06",
          3055 => x"38",
          3056 => x"70",
          3057 => x"33",
          3058 => x"c1",
          3059 => x"38",
          3060 => x"81",
          3061 => x"85",
          3062 => x"34",
          3063 => x"b6",
          3064 => x"06",
          3065 => x"38",
          3066 => x"70",
          3067 => x"f7",
          3068 => x"86",
          3069 => x"54",
          3070 => x"81",
          3071 => x"81",
          3072 => x"38",
          3073 => x"0b",
          3074 => x"08",
          3075 => x"e8",
          3076 => x"42",
          3077 => x"16",
          3078 => x"38",
          3079 => x"80",
          3080 => x"16",
          3081 => x"38",
          3082 => x"81",
          3083 => x"73",
          3084 => x"d4",
          3085 => x"da",
          3086 => x"81",
          3087 => x"d4",
          3088 => x"80",
          3089 => x"05",
          3090 => x"73",
          3091 => x"87",
          3092 => x"0c",
          3093 => x"57",
          3094 => x"76",
          3095 => x"e8",
          3096 => x"26",
          3097 => x"c9",
          3098 => x"f8",
          3099 => x"38",
          3100 => x"08",
          3101 => x"38",
          3102 => x"54",
          3103 => x"73",
          3104 => x"9c",
          3105 => x"ff",
          3106 => x"83",
          3107 => x"88",
          3108 => x"fc",
          3109 => x"72",
          3110 => x"2e",
          3111 => x"81",
          3112 => x"fe",
          3113 => x"59",
          3114 => x"2e",
          3115 => x"81",
          3116 => x"80",
          3117 => x"87",
          3118 => x"72",
          3119 => x"9c",
          3120 => x"76",
          3121 => x"71",
          3122 => x"80",
          3123 => x"10",
          3124 => x"78",
          3125 => x"5b",
          3126 => x"08",
          3127 => x"39",
          3128 => x"38",
          3129 => x"39",
          3130 => x"2e",
          3131 => x"82",
          3132 => x"e8",
          3133 => x"80",
          3134 => x"8a",
          3135 => x"f9",
          3136 => x"38",
          3137 => x"f8",
          3138 => x"7c",
          3139 => x"81",
          3140 => x"e2",
          3141 => x"80",
          3142 => x"33",
          3143 => x"ff",
          3144 => x"78",
          3145 => x"04",
          3146 => x"f6",
          3147 => x"83",
          3148 => x"7a",
          3149 => x"39",
          3150 => x"ff",
          3151 => x"0b",
          3152 => x"39",
          3153 => x"ff",
          3154 => x"16",
          3155 => x"38",
          3156 => x"2e",
          3157 => x"f7",
          3158 => x"98",
          3159 => x"fb",
          3160 => x"83",
          3161 => x"59",
          3162 => x"c0",
          3163 => x"f7",
          3164 => x"72",
          3165 => x"34",
          3166 => x"f7",
          3167 => x"83",
          3168 => x"5d",
          3169 => x"9c",
          3170 => x"fc",
          3171 => x"fc",
          3172 => x"06",
          3173 => x"76",
          3174 => x"80",
          3175 => x"75",
          3176 => x"83",
          3177 => x"0b",
          3178 => x"83",
          3179 => x"34",
          3180 => x"83",
          3181 => x"38",
          3182 => x"ff",
          3183 => x"ff",
          3184 => x"79",
          3185 => x"f9",
          3186 => x"15",
          3187 => x"80",
          3188 => x"b8",
          3189 => x"ff",
          3190 => x"80",
          3191 => x"59",
          3192 => x"ff",
          3193 => x"39",
          3194 => x"08",
          3195 => x"eb",
          3196 => x"83",
          3197 => x"80",
          3198 => x"82",
          3199 => x"0b",
          3200 => x"a7",
          3201 => x"98",
          3202 => x"0b",
          3203 => x"0b",
          3204 => x"80",
          3205 => x"83",
          3206 => x"05",
          3207 => x"87",
          3208 => x"2e",
          3209 => x"98",
          3210 => x"87",
          3211 => x"87",
          3212 => x"71",
          3213 => x"72",
          3214 => x"98",
          3215 => x"87",
          3216 => x"98",
          3217 => x"38",
          3218 => x"08",
          3219 => x"72",
          3220 => x"98",
          3221 => x"27",
          3222 => x"9d",
          3223 => x"81",
          3224 => x"75",
          3225 => x"8c",
          3226 => x"70",
          3227 => x"38",
          3228 => x"fe",
          3229 => x"0c",
          3230 => x"7a",
          3231 => x"53",
          3232 => x"88",
          3233 => x"76",
          3234 => x"72",
          3235 => x"71",
          3236 => x"76",
          3237 => x"83",
          3238 => x"34",
          3239 => x"72",
          3240 => x"56",
          3241 => x"0b",
          3242 => x"98",
          3243 => x"80",
          3244 => x"9c",
          3245 => x"52",
          3246 => x"33",
          3247 => x"75",
          3248 => x"2e",
          3249 => x"52",
          3250 => x"38",
          3251 => x"38",
          3252 => x"90",
          3253 => x"53",
          3254 => x"73",
          3255 => x"c0",
          3256 => x"27",
          3257 => x"38",
          3258 => x"56",
          3259 => x"56",
          3260 => x"80",
          3261 => x"06",
          3262 => x"71",
          3263 => x"80",
          3264 => x"53",
          3265 => x"70",
          3266 => x"05",
          3267 => x"77",
          3268 => x"04",
          3269 => x"fe",
          3270 => x"0c",
          3271 => x"81",
          3272 => x"38",
          3273 => x"0d",
          3274 => x"57",
          3275 => x"78",
          3276 => x"70",
          3277 => x"58",
          3278 => x"52",
          3279 => x"53",
          3280 => x"34",
          3281 => x"11",
          3282 => x"71",
          3283 => x"05",
          3284 => x"34",
          3285 => x"98",
          3286 => x"f4",
          3287 => x"85",
          3288 => x"fe",
          3289 => x"f0",
          3290 => x"08",
          3291 => x"90",
          3292 => x"53",
          3293 => x"73",
          3294 => x"c0",
          3295 => x"27",
          3296 => x"38",
          3297 => x"56",
          3298 => x"56",
          3299 => x"c0",
          3300 => x"54",
          3301 => x"c0",
          3302 => x"f6",
          3303 => x"9c",
          3304 => x"38",
          3305 => x"c0",
          3306 => x"74",
          3307 => x"2e",
          3308 => x"75",
          3309 => x"38",
          3310 => x"74",
          3311 => x"89",
          3312 => x"ff",
          3313 => x"70",
          3314 => x"2e",
          3315 => x"52",
          3316 => x"ba",
          3317 => x"3d",
          3318 => x"d0",
          3319 => x"08",
          3320 => x"80",
          3321 => x"c0",
          3322 => x"56",
          3323 => x"98",
          3324 => x"08",
          3325 => x"15",
          3326 => x"52",
          3327 => x"fe",
          3328 => x"08",
          3329 => x"cd",
          3330 => x"c5",
          3331 => x"ce",
          3332 => x"08",
          3333 => x"72",
          3334 => x"87",
          3335 => x"74",
          3336 => x"db",
          3337 => x"ff",
          3338 => x"53",
          3339 => x"2e",
          3340 => x"71",
          3341 => x"70",
          3342 => x"80",
          3343 => x"cf",
          3344 => x"3d",
          3345 => x"31",
          3346 => x"70",
          3347 => x"12",
          3348 => x"07",
          3349 => x"71",
          3350 => x"54",
          3351 => x"56",
          3352 => x"38",
          3353 => x"33",
          3354 => x"76",
          3355 => x"98",
          3356 => x"5c",
          3357 => x"83",
          3358 => x"33",
          3359 => x"75",
          3360 => x"57",
          3361 => x"06",
          3362 => x"fc",
          3363 => x"13",
          3364 => x"2a",
          3365 => x"14",
          3366 => x"fc",
          3367 => x"34",
          3368 => x"fc",
          3369 => x"85",
          3370 => x"70",
          3371 => x"07",
          3372 => x"58",
          3373 => x"81",
          3374 => x"12",
          3375 => x"71",
          3376 => x"33",
          3377 => x"70",
          3378 => x"58",
          3379 => x"12",
          3380 => x"84",
          3381 => x"2b",
          3382 => x"52",
          3383 => x"33",
          3384 => x"52",
          3385 => x"72",
          3386 => x"15",
          3387 => x"2b",
          3388 => x"2a",
          3389 => x"77",
          3390 => x"70",
          3391 => x"8b",
          3392 => x"70",
          3393 => x"07",
          3394 => x"77",
          3395 => x"54",
          3396 => x"14",
          3397 => x"fc",
          3398 => x"33",
          3399 => x"74",
          3400 => x"88",
          3401 => x"88",
          3402 => x"54",
          3403 => x"34",
          3404 => x"11",
          3405 => x"71",
          3406 => x"81",
          3407 => x"2b",
          3408 => x"53",
          3409 => x"71",
          3410 => x"07",
          3411 => x"59",
          3412 => x"16",
          3413 => x"70",
          3414 => x"71",
          3415 => x"33",
          3416 => x"70",
          3417 => x"56",
          3418 => x"83",
          3419 => x"3d",
          3420 => x"58",
          3421 => x"2e",
          3422 => x"89",
          3423 => x"84",
          3424 => x"b9",
          3425 => x"52",
          3426 => x"3f",
          3427 => x"34",
          3428 => x"fc",
          3429 => x"0b",
          3430 => x"56",
          3431 => x"17",
          3432 => x"f8",
          3433 => x"70",
          3434 => x"58",
          3435 => x"73",
          3436 => x"70",
          3437 => x"05",
          3438 => x"34",
          3439 => x"39",
          3440 => x"81",
          3441 => x"12",
          3442 => x"ff",
          3443 => x"06",
          3444 => x"85",
          3445 => x"52",
          3446 => x"54",
          3447 => x"10",
          3448 => x"33",
          3449 => x"ff",
          3450 => x"06",
          3451 => x"54",
          3452 => x"80",
          3453 => x"84",
          3454 => x"2b",
          3455 => x"81",
          3456 => x"54",
          3457 => x"70",
          3458 => x"07",
          3459 => x"5d",
          3460 => x"38",
          3461 => x"82",
          3462 => x"82",
          3463 => x"38",
          3464 => x"74",
          3465 => x"5b",
          3466 => x"78",
          3467 => x"15",
          3468 => x"14",
          3469 => x"fc",
          3470 => x"33",
          3471 => x"8f",
          3472 => x"ff",
          3473 => x"53",
          3474 => x"34",
          3475 => x"12",
          3476 => x"75",
          3477 => x"b9",
          3478 => x"87",
          3479 => x"2b",
          3480 => x"57",
          3481 => x"34",
          3482 => x"78",
          3483 => x"71",
          3484 => x"54",
          3485 => x"87",
          3486 => x"19",
          3487 => x"8b",
          3488 => x"58",
          3489 => x"34",
          3490 => x"08",
          3491 => x"33",
          3492 => x"70",
          3493 => x"84",
          3494 => x"b9",
          3495 => x"84",
          3496 => x"86",
          3497 => x"2b",
          3498 => x"17",
          3499 => x"07",
          3500 => x"54",
          3501 => x"12",
          3502 => x"84",
          3503 => x"2b",
          3504 => x"14",
          3505 => x"07",
          3506 => x"56",
          3507 => x"76",
          3508 => x"18",
          3509 => x"2b",
          3510 => x"2a",
          3511 => x"74",
          3512 => x"18",
          3513 => x"3d",
          3514 => x"58",
          3515 => x"77",
          3516 => x"89",
          3517 => x"3f",
          3518 => x"0c",
          3519 => x"0b",
          3520 => x"84",
          3521 => x"76",
          3522 => x"eb",
          3523 => x"75",
          3524 => x"b9",
          3525 => x"81",
          3526 => x"08",
          3527 => x"87",
          3528 => x"b9",
          3529 => x"07",
          3530 => x"2a",
          3531 => x"34",
          3532 => x"22",
          3533 => x"08",
          3534 => x"15",
          3535 => x"54",
          3536 => x"e3",
          3537 => x"5f",
          3538 => x"45",
          3539 => x"7e",
          3540 => x"2e",
          3541 => x"27",
          3542 => x"82",
          3543 => x"58",
          3544 => x"31",
          3545 => x"70",
          3546 => x"12",
          3547 => x"31",
          3548 => x"10",
          3549 => x"11",
          3550 => x"2b",
          3551 => x"53",
          3552 => x"44",
          3553 => x"80",
          3554 => x"33",
          3555 => x"70",
          3556 => x"12",
          3557 => x"07",
          3558 => x"74",
          3559 => x"82",
          3560 => x"2e",
          3561 => x"f9",
          3562 => x"87",
          3563 => x"24",
          3564 => x"81",
          3565 => x"2b",
          3566 => x"33",
          3567 => x"47",
          3568 => x"80",
          3569 => x"82",
          3570 => x"2b",
          3571 => x"11",
          3572 => x"71",
          3573 => x"33",
          3574 => x"70",
          3575 => x"41",
          3576 => x"1d",
          3577 => x"fc",
          3578 => x"12",
          3579 => x"07",
          3580 => x"33",
          3581 => x"5f",
          3582 => x"77",
          3583 => x"84",
          3584 => x"12",
          3585 => x"ff",
          3586 => x"59",
          3587 => x"84",
          3588 => x"33",
          3589 => x"83",
          3590 => x"15",
          3591 => x"2a",
          3592 => x"55",
          3593 => x"84",
          3594 => x"81",
          3595 => x"2b",
          3596 => x"15",
          3597 => x"2a",
          3598 => x"55",
          3599 => x"34",
          3600 => x"11",
          3601 => x"07",
          3602 => x"42",
          3603 => x"51",
          3604 => x"08",
          3605 => x"70",
          3606 => x"7a",
          3607 => x"73",
          3608 => x"04",
          3609 => x"0c",
          3610 => x"82",
          3611 => x"f4",
          3612 => x"fc",
          3613 => x"81",
          3614 => x"60",
          3615 => x"34",
          3616 => x"1d",
          3617 => x"b9",
          3618 => x"05",
          3619 => x"ff",
          3620 => x"57",
          3621 => x"34",
          3622 => x"10",
          3623 => x"55",
          3624 => x"83",
          3625 => x"7e",
          3626 => x"8c",
          3627 => x"df",
          3628 => x"ba",
          3629 => x"3d",
          3630 => x"08",
          3631 => x"7f",
          3632 => x"88",
          3633 => x"88",
          3634 => x"7b",
          3635 => x"b9",
          3636 => x"58",
          3637 => x"34",
          3638 => x"33",
          3639 => x"70",
          3640 => x"05",
          3641 => x"2a",
          3642 => x"63",
          3643 => x"06",
          3644 => x"b9",
          3645 => x"60",
          3646 => x"08",
          3647 => x"7e",
          3648 => x"70",
          3649 => x"ac",
          3650 => x"31",
          3651 => x"33",
          3652 => x"70",
          3653 => x"12",
          3654 => x"07",
          3655 => x"54",
          3656 => x"bc",
          3657 => x"80",
          3658 => x"ff",
          3659 => x"dd",
          3660 => x"0b",
          3661 => x"84",
          3662 => x"7e",
          3663 => x"83",
          3664 => x"7a",
          3665 => x"b9",
          3666 => x"81",
          3667 => x"08",
          3668 => x"87",
          3669 => x"b9",
          3670 => x"07",
          3671 => x"2a",
          3672 => x"05",
          3673 => x"b9",
          3674 => x"b9",
          3675 => x"7e",
          3676 => x"05",
          3677 => x"83",
          3678 => x"5b",
          3679 => x"f2",
          3680 => x"7e",
          3681 => x"84",
          3682 => x"76",
          3683 => x"71",
          3684 => x"11",
          3685 => x"8b",
          3686 => x"84",
          3687 => x"2b",
          3688 => x"56",
          3689 => x"78",
          3690 => x"05",
          3691 => x"84",
          3692 => x"2b",
          3693 => x"14",
          3694 => x"07",
          3695 => x"5d",
          3696 => x"34",
          3697 => x"fc",
          3698 => x"71",
          3699 => x"70",
          3700 => x"7d",
          3701 => x"fc",
          3702 => x"12",
          3703 => x"07",
          3704 => x"71",
          3705 => x"5c",
          3706 => x"7c",
          3707 => x"fc",
          3708 => x"33",
          3709 => x"74",
          3710 => x"71",
          3711 => x"47",
          3712 => x"82",
          3713 => x"b9",
          3714 => x"83",
          3715 => x"57",
          3716 => x"58",
          3717 => x"bd",
          3718 => x"84",
          3719 => x"5f",
          3720 => x"84",
          3721 => x"b9",
          3722 => x"52",
          3723 => x"3f",
          3724 => x"34",
          3725 => x"fc",
          3726 => x"0b",
          3727 => x"54",
          3728 => x"15",
          3729 => x"f8",
          3730 => x"70",
          3731 => x"45",
          3732 => x"60",
          3733 => x"70",
          3734 => x"05",
          3735 => x"34",
          3736 => x"e7",
          3737 => x"86",
          3738 => x"2b",
          3739 => x"1c",
          3740 => x"07",
          3741 => x"59",
          3742 => x"61",
          3743 => x"70",
          3744 => x"71",
          3745 => x"05",
          3746 => x"88",
          3747 => x"48",
          3748 => x"86",
          3749 => x"84",
          3750 => x"12",
          3751 => x"ff",
          3752 => x"58",
          3753 => x"84",
          3754 => x"81",
          3755 => x"2b",
          3756 => x"33",
          3757 => x"8f",
          3758 => x"2a",
          3759 => x"44",
          3760 => x"17",
          3761 => x"70",
          3762 => x"71",
          3763 => x"81",
          3764 => x"ff",
          3765 => x"5e",
          3766 => x"34",
          3767 => x"ff",
          3768 => x"15",
          3769 => x"71",
          3770 => x"33",
          3771 => x"70",
          3772 => x"5d",
          3773 => x"34",
          3774 => x"11",
          3775 => x"71",
          3776 => x"33",
          3777 => x"70",
          3778 => x"42",
          3779 => x"75",
          3780 => x"08",
          3781 => x"88",
          3782 => x"88",
          3783 => x"34",
          3784 => x"08",
          3785 => x"71",
          3786 => x"05",
          3787 => x"2b",
          3788 => x"06",
          3789 => x"5f",
          3790 => x"82",
          3791 => x"b9",
          3792 => x"12",
          3793 => x"07",
          3794 => x"71",
          3795 => x"70",
          3796 => x"59",
          3797 => x"1d",
          3798 => x"82",
          3799 => x"2b",
          3800 => x"11",
          3801 => x"71",
          3802 => x"33",
          3803 => x"70",
          3804 => x"42",
          3805 => x"84",
          3806 => x"b9",
          3807 => x"85",
          3808 => x"2b",
          3809 => x"15",
          3810 => x"2a",
          3811 => x"57",
          3812 => x"34",
          3813 => x"81",
          3814 => x"ff",
          3815 => x"5e",
          3816 => x"34",
          3817 => x"11",
          3818 => x"71",
          3819 => x"81",
          3820 => x"88",
          3821 => x"55",
          3822 => x"34",
          3823 => x"33",
          3824 => x"83",
          3825 => x"83",
          3826 => x"88",
          3827 => x"55",
          3828 => x"1a",
          3829 => x"82",
          3830 => x"2b",
          3831 => x"2b",
          3832 => x"05",
          3833 => x"fc",
          3834 => x"1c",
          3835 => x"5f",
          3836 => x"1a",
          3837 => x"07",
          3838 => x"33",
          3839 => x"40",
          3840 => x"84",
          3841 => x"84",
          3842 => x"33",
          3843 => x"83",
          3844 => x"87",
          3845 => x"88",
          3846 => x"41",
          3847 => x"64",
          3848 => x"1d",
          3849 => x"2b",
          3850 => x"2a",
          3851 => x"7c",
          3852 => x"70",
          3853 => x"8b",
          3854 => x"70",
          3855 => x"07",
          3856 => x"77",
          3857 => x"49",
          3858 => x"1e",
          3859 => x"fc",
          3860 => x"33",
          3861 => x"74",
          3862 => x"88",
          3863 => x"88",
          3864 => x"5e",
          3865 => x"34",
          3866 => x"83",
          3867 => x"3f",
          3868 => x"8c",
          3869 => x"73",
          3870 => x"b4",
          3871 => x"61",
          3872 => x"f0",
          3873 => x"29",
          3874 => x"80",
          3875 => x"38",
          3876 => x"0d",
          3877 => x"ba",
          3878 => x"80",
          3879 => x"84",
          3880 => x"3f",
          3881 => x"0d",
          3882 => x"fc",
          3883 => x"23",
          3884 => x"ff",
          3885 => x"b9",
          3886 => x"0b",
          3887 => x"54",
          3888 => x"15",
          3889 => x"86",
          3890 => x"84",
          3891 => x"ff",
          3892 => x"ff",
          3893 => x"55",
          3894 => x"17",
          3895 => x"10",
          3896 => x"05",
          3897 => x"0b",
          3898 => x"2e",
          3899 => x"3d",
          3900 => x"52",
          3901 => x"88",
          3902 => x"0c",
          3903 => x"02",
          3904 => x"81",
          3905 => x"3f",
          3906 => x"53",
          3907 => x"13",
          3908 => x"72",
          3909 => x"04",
          3910 => x"8c",
          3911 => x"59",
          3912 => x"84",
          3913 => x"06",
          3914 => x"58",
          3915 => x"78",
          3916 => x"3f",
          3917 => x"55",
          3918 => x"98",
          3919 => x"78",
          3920 => x"06",
          3921 => x"54",
          3922 => x"8b",
          3923 => x"19",
          3924 => x"79",
          3925 => x"f7",
          3926 => x"05",
          3927 => x"81",
          3928 => x"ba",
          3929 => x"54",
          3930 => x"85",
          3931 => x"53",
          3932 => x"84",
          3933 => x"74",
          3934 => x"8c",
          3935 => x"26",
          3936 => x"54",
          3937 => x"73",
          3938 => x"3d",
          3939 => x"70",
          3940 => x"78",
          3941 => x"3d",
          3942 => x"33",
          3943 => x"53",
          3944 => x"38",
          3945 => x"81",
          3946 => x"85",
          3947 => x"53",
          3948 => x"25",
          3949 => x"84",
          3950 => x"3d",
          3951 => x"73",
          3952 => x"04",
          3953 => x"ba",
          3954 => x"84",
          3955 => x"54",
          3956 => x"2a",
          3957 => x"8a",
          3958 => x"74",
          3959 => x"51",
          3960 => x"c0",
          3961 => x"06",
          3962 => x"71",
          3963 => x"ff",
          3964 => x"80",
          3965 => x"57",
          3966 => x"38",
          3967 => x"87",
          3968 => x"33",
          3969 => x"08",
          3970 => x"84",
          3971 => x"81",
          3972 => x"70",
          3973 => x"ff",
          3974 => x"77",
          3975 => x"ba",
          3976 => x"08",
          3977 => x"08",
          3978 => x"5b",
          3979 => x"18",
          3980 => x"06",
          3981 => x"53",
          3982 => x"b7",
          3983 => x"83",
          3984 => x"84",
          3985 => x"81",
          3986 => x"84",
          3987 => x"81",
          3988 => x"f4",
          3989 => x"34",
          3990 => x"80",
          3991 => x"19",
          3992 => x"80",
          3993 => x"0b",
          3994 => x"84",
          3995 => x"9e",
          3996 => x"19",
          3997 => x"a0",
          3998 => x"84",
          3999 => x"75",
          4000 => x"5b",
          4001 => x"08",
          4002 => x"88",
          4003 => x"7a",
          4004 => x"34",
          4005 => x"19",
          4006 => x"b4",
          4007 => x"79",
          4008 => x"3f",
          4009 => x"52",
          4010 => x"84",
          4011 => x"38",
          4012 => x"60",
          4013 => x"27",
          4014 => x"8c",
          4015 => x"0c",
          4016 => x"56",
          4017 => x"74",
          4018 => x"2e",
          4019 => x"2a",
          4020 => x"05",
          4021 => x"79",
          4022 => x"7b",
          4023 => x"38",
          4024 => x"81",
          4025 => x"ba",
          4026 => x"59",
          4027 => x"ff",
          4028 => x"b8",
          4029 => x"a8",
          4030 => x"b4",
          4031 => x"0b",
          4032 => x"74",
          4033 => x"38",
          4034 => x"81",
          4035 => x"ba",
          4036 => x"59",
          4037 => x"fe",
          4038 => x"b8",
          4039 => x"78",
          4040 => x"59",
          4041 => x"9f",
          4042 => x"3d",
          4043 => x"08",
          4044 => x"b5",
          4045 => x"5c",
          4046 => x"06",
          4047 => x"b8",
          4048 => x"a8",
          4049 => x"85",
          4050 => x"18",
          4051 => x"83",
          4052 => x"11",
          4053 => x"84",
          4054 => x"0d",
          4055 => x"fd",
          4056 => x"08",
          4057 => x"b5",
          4058 => x"5c",
          4059 => x"06",
          4060 => x"b8",
          4061 => x"c0",
          4062 => x"85",
          4063 => x"18",
          4064 => x"2b",
          4065 => x"83",
          4066 => x"2b",
          4067 => x"70",
          4068 => x"80",
          4069 => x"ba",
          4070 => x"56",
          4071 => x"17",
          4072 => x"18",
          4073 => x"5a",
          4074 => x"81",
          4075 => x"08",
          4076 => x"18",
          4077 => x"5e",
          4078 => x"38",
          4079 => x"09",
          4080 => x"b4",
          4081 => x"7b",
          4082 => x"3f",
          4083 => x"b4",
          4084 => x"81",
          4085 => x"84",
          4086 => x"06",
          4087 => x"83",
          4088 => x"08",
          4089 => x"8b",
          4090 => x"2e",
          4091 => x"5b",
          4092 => x"08",
          4093 => x"33",
          4094 => x"84",
          4095 => x"06",
          4096 => x"83",
          4097 => x"08",
          4098 => x"7d",
          4099 => x"82",
          4100 => x"81",
          4101 => x"17",
          4102 => x"52",
          4103 => x"7a",
          4104 => x"17",
          4105 => x"18",
          4106 => x"5a",
          4107 => x"81",
          4108 => x"08",
          4109 => x"18",
          4110 => x"55",
          4111 => x"38",
          4112 => x"09",
          4113 => x"b4",
          4114 => x"7d",
          4115 => x"3f",
          4116 => x"b4",
          4117 => x"7b",
          4118 => x"3f",
          4119 => x"bb",
          4120 => x"60",
          4121 => x"81",
          4122 => x"08",
          4123 => x"78",
          4124 => x"80",
          4125 => x"77",
          4126 => x"04",
          4127 => x"58",
          4128 => x"76",
          4129 => x"33",
          4130 => x"81",
          4131 => x"53",
          4132 => x"f2",
          4133 => x"2e",
          4134 => x"b4",
          4135 => x"38",
          4136 => x"7b",
          4137 => x"b8",
          4138 => x"b9",
          4139 => x"77",
          4140 => x"04",
          4141 => x"ff",
          4142 => x"05",
          4143 => x"5c",
          4144 => x"19",
          4145 => x"09",
          4146 => x"77",
          4147 => x"51",
          4148 => x"80",
          4149 => x"77",
          4150 => x"b7",
          4151 => x"79",
          4152 => x"98",
          4153 => x"06",
          4154 => x"34",
          4155 => x"34",
          4156 => x"34",
          4157 => x"34",
          4158 => x"39",
          4159 => x"a8",
          4160 => x"59",
          4161 => x"0b",
          4162 => x"74",
          4163 => x"38",
          4164 => x"81",
          4165 => x"ba",
          4166 => x"58",
          4167 => x"58",
          4168 => x"06",
          4169 => x"06",
          4170 => x"2e",
          4171 => x"06",
          4172 => x"5a",
          4173 => x"34",
          4174 => x"56",
          4175 => x"74",
          4176 => x"74",
          4177 => x"33",
          4178 => x"84",
          4179 => x"06",
          4180 => x"83",
          4181 => x"1b",
          4182 => x"8c",
          4183 => x"27",
          4184 => x"82",
          4185 => x"53",
          4186 => x"d8",
          4187 => x"85",
          4188 => x"1a",
          4189 => x"ff",
          4190 => x"56",
          4191 => x"76",
          4192 => x"07",
          4193 => x"83",
          4194 => x"76",
          4195 => x"33",
          4196 => x"84",
          4197 => x"06",
          4198 => x"83",
          4199 => x"1b",
          4200 => x"8c",
          4201 => x"27",
          4202 => x"74",
          4203 => x"38",
          4204 => x"81",
          4205 => x"5a",
          4206 => x"b8",
          4207 => x"57",
          4208 => x"8c",
          4209 => x"ae",
          4210 => x"34",
          4211 => x"31",
          4212 => x"5f",
          4213 => x"f0",
          4214 => x"2e",
          4215 => x"54",
          4216 => x"33",
          4217 => x"d0",
          4218 => x"70",
          4219 => x"cf",
          4220 => x"7c",
          4221 => x"84",
          4222 => x"19",
          4223 => x"1b",
          4224 => x"40",
          4225 => x"82",
          4226 => x"81",
          4227 => x"1e",
          4228 => x"ed",
          4229 => x"81",
          4230 => x"19",
          4231 => x"fd",
          4232 => x"06",
          4233 => x"59",
          4234 => x"88",
          4235 => x"fa",
          4236 => x"76",
          4237 => x"b8",
          4238 => x"8f",
          4239 => x"42",
          4240 => x"7d",
          4241 => x"7d",
          4242 => x"7d",
          4243 => x"fa",
          4244 => x"71",
          4245 => x"38",
          4246 => x"80",
          4247 => x"80",
          4248 => x"54",
          4249 => x"7b",
          4250 => x"16",
          4251 => x"38",
          4252 => x"38",
          4253 => x"84",
          4254 => x"38",
          4255 => x"2e",
          4256 => x"70",
          4257 => x"7b",
          4258 => x"aa",
          4259 => x"ff",
          4260 => x"8c",
          4261 => x"ff",
          4262 => x"ca",
          4263 => x"3f",
          4264 => x"27",
          4265 => x"84",
          4266 => x"9c",
          4267 => x"c4",
          4268 => x"1b",
          4269 => x"38",
          4270 => x"eb",
          4271 => x"81",
          4272 => x"08",
          4273 => x"25",
          4274 => x"54",
          4275 => x"38",
          4276 => x"38",
          4277 => x"fe",
          4278 => x"fe",
          4279 => x"96",
          4280 => x"ff",
          4281 => x"3f",
          4282 => x"08",
          4283 => x"80",
          4284 => x"38",
          4285 => x"0c",
          4286 => x"08",
          4287 => x"ff",
          4288 => x"81",
          4289 => x"55",
          4290 => x"0d",
          4291 => x"8c",
          4292 => x"58",
          4293 => x"b8",
          4294 => x"f5",
          4295 => x"ff",
          4296 => x"ba",
          4297 => x"56",
          4298 => x"55",
          4299 => x"7c",
          4300 => x"80",
          4301 => x"06",
          4302 => x"19",
          4303 => x"df",
          4304 => x"80",
          4305 => x"0b",
          4306 => x"27",
          4307 => x"0c",
          4308 => x"53",
          4309 => x"73",
          4310 => x"83",
          4311 => x"0c",
          4312 => x"8a",
          4313 => x"8c",
          4314 => x"08",
          4315 => x"8a",
          4316 => x"73",
          4317 => x"53",
          4318 => x"59",
          4319 => x"22",
          4320 => x"5a",
          4321 => x"39",
          4322 => x"84",
          4323 => x"08",
          4324 => x"ba",
          4325 => x"17",
          4326 => x"27",
          4327 => x"73",
          4328 => x"81",
          4329 => x"0d",
          4330 => x"90",
          4331 => x"f0",
          4332 => x"0b",
          4333 => x"84",
          4334 => x"83",
          4335 => x"15",
          4336 => x"38",
          4337 => x"55",
          4338 => x"98",
          4339 => x"1b",
          4340 => x"75",
          4341 => x"04",
          4342 => x"ff",
          4343 => x"da",
          4344 => x"3f",
          4345 => x"81",
          4346 => x"38",
          4347 => x"2e",
          4348 => x"8c",
          4349 => x"2e",
          4350 => x"76",
          4351 => x"08",
          4352 => x"80",
          4353 => x"ba",
          4354 => x"81",
          4355 => x"ff",
          4356 => x"1a",
          4357 => x"fe",
          4358 => x"56",
          4359 => x"8a",
          4360 => x"08",
          4361 => x"b8",
          4362 => x"80",
          4363 => x"15",
          4364 => x"19",
          4365 => x"38",
          4366 => x"81",
          4367 => x"ba",
          4368 => x"56",
          4369 => x"0b",
          4370 => x"04",
          4371 => x"19",
          4372 => x"e4",
          4373 => x"f3",
          4374 => x"34",
          4375 => x"55",
          4376 => x"38",
          4377 => x"09",
          4378 => x"b4",
          4379 => x"75",
          4380 => x"3f",
          4381 => x"74",
          4382 => x"2e",
          4383 => x"18",
          4384 => x"05",
          4385 => x"fd",
          4386 => x"29",
          4387 => x"5c",
          4388 => x"8c",
          4389 => x"0d",
          4390 => x"5a",
          4391 => x"58",
          4392 => x"38",
          4393 => x"b4",
          4394 => x"83",
          4395 => x"2e",
          4396 => x"54",
          4397 => x"33",
          4398 => x"08",
          4399 => x"57",
          4400 => x"82",
          4401 => x"58",
          4402 => x"8b",
          4403 => x"06",
          4404 => x"81",
          4405 => x"70",
          4406 => x"07",
          4407 => x"38",
          4408 => x"88",
          4409 => x"81",
          4410 => x"7b",
          4411 => x"08",
          4412 => x"38",
          4413 => x"38",
          4414 => x"0d",
          4415 => x"7e",
          4416 => x"3f",
          4417 => x"2e",
          4418 => x"ba",
          4419 => x"08",
          4420 => x"08",
          4421 => x"fe",
          4422 => x"82",
          4423 => x"81",
          4424 => x"05",
          4425 => x"e0",
          4426 => x"79",
          4427 => x"38",
          4428 => x"80",
          4429 => x"81",
          4430 => x"ac",
          4431 => x"2e",
          4432 => x"fe",
          4433 => x"09",
          4434 => x"84",
          4435 => x"84",
          4436 => x"77",
          4437 => x"57",
          4438 => x"38",
          4439 => x"1a",
          4440 => x"41",
          4441 => x"81",
          4442 => x"5a",
          4443 => x"17",
          4444 => x"33",
          4445 => x"7a",
          4446 => x"fe",
          4447 => x"05",
          4448 => x"1a",
          4449 => x"cc",
          4450 => x"06",
          4451 => x"79",
          4452 => x"10",
          4453 => x"1d",
          4454 => x"9d",
          4455 => x"38",
          4456 => x"a8",
          4457 => x"2a",
          4458 => x"81",
          4459 => x"81",
          4460 => x"76",
          4461 => x"38",
          4462 => x"ba",
          4463 => x"3d",
          4464 => x"52",
          4465 => x"8c",
          4466 => x"80",
          4467 => x"0b",
          4468 => x"1c",
          4469 => x"76",
          4470 => x"78",
          4471 => x"06",
          4472 => x"b8",
          4473 => x"e0",
          4474 => x"85",
          4475 => x"1c",
          4476 => x"9c",
          4477 => x"80",
          4478 => x"bf",
          4479 => x"77",
          4480 => x"80",
          4481 => x"55",
          4482 => x"80",
          4483 => x"38",
          4484 => x"8b",
          4485 => x"29",
          4486 => x"57",
          4487 => x"19",
          4488 => x"7f",
          4489 => x"81",
          4490 => x"a0",
          4491 => x"5a",
          4492 => x"71",
          4493 => x"40",
          4494 => x"80",
          4495 => x"0b",
          4496 => x"f5",
          4497 => x"84",
          4498 => x"38",
          4499 => x"0d",
          4500 => x"7d",
          4501 => x"3f",
          4502 => x"2e",
          4503 => x"ba",
          4504 => x"08",
          4505 => x"08",
          4506 => x"fd",
          4507 => x"82",
          4508 => x"81",
          4509 => x"05",
          4510 => x"db",
          4511 => x"77",
          4512 => x"70",
          4513 => x"fe",
          4514 => x"5a",
          4515 => x"33",
          4516 => x"08",
          4517 => x"76",
          4518 => x"74",
          4519 => x"3f",
          4520 => x"8c",
          4521 => x"c8",
          4522 => x"81",
          4523 => x"fe",
          4524 => x"77",
          4525 => x"1b",
          4526 => x"71",
          4527 => x"ff",
          4528 => x"8d",
          4529 => x"59",
          4530 => x"05",
          4531 => x"2b",
          4532 => x"80",
          4533 => x"84",
          4534 => x"84",
          4535 => x"70",
          4536 => x"81",
          4537 => x"08",
          4538 => x"76",
          4539 => x"ff",
          4540 => x"81",
          4541 => x"38",
          4542 => x"60",
          4543 => x"b4",
          4544 => x"5e",
          4545 => x"ba",
          4546 => x"83",
          4547 => x"ff",
          4548 => x"68",
          4549 => x"a0",
          4550 => x"74",
          4551 => x"70",
          4552 => x"8e",
          4553 => x"22",
          4554 => x"3d",
          4555 => x"58",
          4556 => x"33",
          4557 => x"15",
          4558 => x"05",
          4559 => x"80",
          4560 => x"ab",
          4561 => x"5b",
          4562 => x"7a",
          4563 => x"05",
          4564 => x"34",
          4565 => x"7b",
          4566 => x"56",
          4567 => x"82",
          4568 => x"06",
          4569 => x"83",
          4570 => x"06",
          4571 => x"87",
          4572 => x"ff",
          4573 => x"78",
          4574 => x"84",
          4575 => x"b0",
          4576 => x"84",
          4577 => x"ff",
          4578 => x"59",
          4579 => x"80",
          4580 => x"80",
          4581 => x"74",
          4582 => x"75",
          4583 => x"70",
          4584 => x"81",
          4585 => x"55",
          4586 => x"78",
          4587 => x"57",
          4588 => x"27",
          4589 => x"3f",
          4590 => x"1b",
          4591 => x"38",
          4592 => x"e7",
          4593 => x"ba",
          4594 => x"82",
          4595 => x"ab",
          4596 => x"80",
          4597 => x"2a",
          4598 => x"2e",
          4599 => x"fe",
          4600 => x"1b",
          4601 => x"3f",
          4602 => x"8c",
          4603 => x"08",
          4604 => x"56",
          4605 => x"85",
          4606 => x"77",
          4607 => x"81",
          4608 => x"18",
          4609 => x"8c",
          4610 => x"81",
          4611 => x"76",
          4612 => x"56",
          4613 => x"38",
          4614 => x"56",
          4615 => x"81",
          4616 => x"38",
          4617 => x"84",
          4618 => x"08",
          4619 => x"75",
          4620 => x"75",
          4621 => x"81",
          4622 => x"1c",
          4623 => x"33",
          4624 => x"81",
          4625 => x"1c",
          4626 => x"8c",
          4627 => x"81",
          4628 => x"75",
          4629 => x"08",
          4630 => x"58",
          4631 => x"8b",
          4632 => x"55",
          4633 => x"70",
          4634 => x"74",
          4635 => x"33",
          4636 => x"34",
          4637 => x"75",
          4638 => x"04",
          4639 => x"07",
          4640 => x"74",
          4641 => x"3f",
          4642 => x"8c",
          4643 => x"bd",
          4644 => x"7c",
          4645 => x"3f",
          4646 => x"81",
          4647 => x"08",
          4648 => x"19",
          4649 => x"27",
          4650 => x"82",
          4651 => x"08",
          4652 => x"90",
          4653 => x"51",
          4654 => x"58",
          4655 => x"79",
          4656 => x"57",
          4657 => x"05",
          4658 => x"76",
          4659 => x"59",
          4660 => x"ff",
          4661 => x"08",
          4662 => x"2e",
          4663 => x"76",
          4664 => x"81",
          4665 => x"1c",
          4666 => x"8c",
          4667 => x"81",
          4668 => x"75",
          4669 => x"1f",
          4670 => x"5f",
          4671 => x"1c",
          4672 => x"1c",
          4673 => x"29",
          4674 => x"76",
          4675 => x"10",
          4676 => x"56",
          4677 => x"55",
          4678 => x"76",
          4679 => x"85",
          4680 => x"58",
          4681 => x"ff",
          4682 => x"1f",
          4683 => x"81",
          4684 => x"83",
          4685 => x"e1",
          4686 => x"ba",
          4687 => x"05",
          4688 => x"39",
          4689 => x"1c",
          4690 => x"d0",
          4691 => x"08",
          4692 => x"83",
          4693 => x"08",
          4694 => x"60",
          4695 => x"82",
          4696 => x"81",
          4697 => x"1c",
          4698 => x"52",
          4699 => x"77",
          4700 => x"08",
          4701 => x"e5",
          4702 => x"fb",
          4703 => x"80",
          4704 => x"7c",
          4705 => x"81",
          4706 => x"81",
          4707 => x"ba",
          4708 => x"bc",
          4709 => x"34",
          4710 => x"55",
          4711 => x"82",
          4712 => x"38",
          4713 => x"39",
          4714 => x"2e",
          4715 => x"1a",
          4716 => x"56",
          4717 => x"fd",
          4718 => x"1d",
          4719 => x"33",
          4720 => x"81",
          4721 => x"05",
          4722 => x"ce",
          4723 => x"0d",
          4724 => x"80",
          4725 => x"80",
          4726 => x"ff",
          4727 => x"60",
          4728 => x"5b",
          4729 => x"77",
          4730 => x"5b",
          4731 => x"d0",
          4732 => x"58",
          4733 => x"38",
          4734 => x"5d",
          4735 => x"30",
          4736 => x"5a",
          4737 => x"80",
          4738 => x"1f",
          4739 => x"70",
          4740 => x"a0",
          4741 => x"bc",
          4742 => x"72",
          4743 => x"8b",
          4744 => x"38",
          4745 => x"81",
          4746 => x"59",
          4747 => x"ff",
          4748 => x"80",
          4749 => x"53",
          4750 => x"bf",
          4751 => x"17",
          4752 => x"34",
          4753 => x"53",
          4754 => x"9c",
          4755 => x"1e",
          4756 => x"11",
          4757 => x"71",
          4758 => x"72",
          4759 => x"64",
          4760 => x"33",
          4761 => x"40",
          4762 => x"23",
          4763 => x"88",
          4764 => x"23",
          4765 => x"fe",
          4766 => x"ff",
          4767 => x"52",
          4768 => x"91",
          4769 => x"ff",
          4770 => x"ad",
          4771 => x"74",
          4772 => x"97",
          4773 => x"0b",
          4774 => x"75",
          4775 => x"fd",
          4776 => x"76",
          4777 => x"80",
          4778 => x"f9",
          4779 => x"58",
          4780 => x"cd",
          4781 => x"57",
          4782 => x"7c",
          4783 => x"14",
          4784 => x"99",
          4785 => x"11",
          4786 => x"38",
          4787 => x"5e",
          4788 => x"70",
          4789 => x"78",
          4790 => x"81",
          4791 => x"5e",
          4792 => x"38",
          4793 => x"cc",
          4794 => x"70",
          4795 => x"fc",
          4796 => x"08",
          4797 => x"33",
          4798 => x"38",
          4799 => x"df",
          4800 => x"98",
          4801 => x"96",
          4802 => x"75",
          4803 => x"16",
          4804 => x"81",
          4805 => x"df",
          4806 => x"81",
          4807 => x"8b",
          4808 => x"23",
          4809 => x"06",
          4810 => x"27",
          4811 => x"55",
          4812 => x"2e",
          4813 => x"b2",
          4814 => x"a8",
          4815 => x"56",
          4816 => x"75",
          4817 => x"70",
          4818 => x"ee",
          4819 => x"81",
          4820 => x"fd",
          4821 => x"23",
          4822 => x"52",
          4823 => x"fe",
          4824 => x"80",
          4825 => x"73",
          4826 => x"2e",
          4827 => x"80",
          4828 => x"dd",
          4829 => x"70",
          4830 => x"72",
          4831 => x"33",
          4832 => x"74",
          4833 => x"83",
          4834 => x"3f",
          4835 => x"06",
          4836 => x"73",
          4837 => x"04",
          4838 => x"06",
          4839 => x"38",
          4840 => x"34",
          4841 => x"84",
          4842 => x"93",
          4843 => x"32",
          4844 => x"41",
          4845 => x"38",
          4846 => x"55",
          4847 => x"72",
          4848 => x"25",
          4849 => x"38",
          4850 => x"2b",
          4851 => x"76",
          4852 => x"59",
          4853 => x"78",
          4854 => x"32",
          4855 => x"56",
          4856 => x"38",
          4857 => x"dd",
          4858 => x"76",
          4859 => x"80",
          4860 => x"72",
          4861 => x"82",
          4862 => x"53",
          4863 => x"80",
          4864 => x"70",
          4865 => x"38",
          4866 => x"17",
          4867 => x"14",
          4868 => x"09",
          4869 => x"1d",
          4870 => x"56",
          4871 => x"72",
          4872 => x"22",
          4873 => x"80",
          4874 => x"83",
          4875 => x"70",
          4876 => x"2e",
          4877 => x"72",
          4878 => x"59",
          4879 => x"07",
          4880 => x"54",
          4881 => x"7c",
          4882 => x"2e",
          4883 => x"77",
          4884 => x"8b",
          4885 => x"18",
          4886 => x"81",
          4887 => x"38",
          4888 => x"2e",
          4889 => x"e3",
          4890 => x"2e",
          4891 => x"74",
          4892 => x"2a",
          4893 => x"81",
          4894 => x"79",
          4895 => x"06",
          4896 => x"88",
          4897 => x"51",
          4898 => x"ab",
          4899 => x"08",
          4900 => x"8c",
          4901 => x"f7",
          4902 => x"79",
          4903 => x"2a",
          4904 => x"7b",
          4905 => x"16",
          4906 => x"81",
          4907 => x"40",
          4908 => x"38",
          4909 => x"83",
          4910 => x"22",
          4911 => x"fc",
          4912 => x"2e",
          4913 => x"10",
          4914 => x"a0",
          4915 => x"26",
          4916 => x"81",
          4917 => x"73",
          4918 => x"77",
          4919 => x"3f",
          4920 => x"56",
          4921 => x"38",
          4922 => x"fa",
          4923 => x"2a",
          4924 => x"83",
          4925 => x"06",
          4926 => x"d2",
          4927 => x"33",
          4928 => x"82",
          4929 => x"08",
          4930 => x"22",
          4931 => x"76",
          4932 => x"ab",
          4933 => x"5a",
          4934 => x"fc",
          4935 => x"8c",
          4936 => x"79",
          4937 => x"0b",
          4938 => x"81",
          4939 => x"80",
          4940 => x"ba",
          4941 => x"80",
          4942 => x"27",
          4943 => x"7b",
          4944 => x"7d",
          4945 => x"39",
          4946 => x"74",
          4947 => x"8c",
          4948 => x"2a",
          4949 => x"c4",
          4950 => x"9c",
          4951 => x"26",
          4952 => x"85",
          4953 => x"b4",
          4954 => x"59",
          4955 => x"75",
          4956 => x"70",
          4957 => x"ee",
          4958 => x"80",
          4959 => x"99",
          4960 => x"81",
          4961 => x"59",
          4962 => x"07",
          4963 => x"83",
          4964 => x"7b",
          4965 => x"81",
          4966 => x"39",
          4967 => x"b4",
          4968 => x"78",
          4969 => x"7a",
          4970 => x"5b",
          4971 => x"d2",
          4972 => x"15",
          4973 => x"07",
          4974 => x"fd",
          4975 => x"88",
          4976 => x"1b",
          4977 => x"79",
          4978 => x"79",
          4979 => x"76",
          4980 => x"a3",
          4981 => x"81",
          4982 => x"0b",
          4983 => x"04",
          4984 => x"05",
          4985 => x"80",
          4986 => x"5b",
          4987 => x"79",
          4988 => x"26",
          4989 => x"38",
          4990 => x"c7",
          4991 => x"76",
          4992 => x"84",
          4993 => x"8c",
          4994 => x"76",
          4995 => x"33",
          4996 => x"81",
          4997 => x"84",
          4998 => x"81",
          4999 => x"96",
          5000 => x"84",
          5001 => x"81",
          5002 => x"a4",
          5003 => x"06",
          5004 => x"7f",
          5005 => x"38",
          5006 => x"58",
          5007 => x"83",
          5008 => x"7a",
          5009 => x"b8",
          5010 => x"58",
          5011 => x"08",
          5012 => x"59",
          5013 => x"99",
          5014 => x"18",
          5015 => x"83",
          5016 => x"a5",
          5017 => x"ba",
          5018 => x"38",
          5019 => x"38",
          5020 => x"38",
          5021 => x"33",
          5022 => x"84",
          5023 => x"38",
          5024 => x"33",
          5025 => x"a4",
          5026 => x"82",
          5027 => x"2b",
          5028 => x"88",
          5029 => x"45",
          5030 => x"0c",
          5031 => x"80",
          5032 => x"ff",
          5033 => x"81",
          5034 => x"06",
          5035 => x"5a",
          5036 => x"59",
          5037 => x"18",
          5038 => x"80",
          5039 => x"71",
          5040 => x"18",
          5041 => x"8d",
          5042 => x"17",
          5043 => x"2b",
          5044 => x"d8",
          5045 => x"71",
          5046 => x"14",
          5047 => x"33",
          5048 => x"42",
          5049 => x"18",
          5050 => x"8d",
          5051 => x"7d",
          5052 => x"75",
          5053 => x"7a",
          5054 => x"ba",
          5055 => x"80",
          5056 => x"08",
          5057 => x"38",
          5058 => x"83",
          5059 => x"85",
          5060 => x"9c",
          5061 => x"1d",
          5062 => x"1a",
          5063 => x"87",
          5064 => x"7b",
          5065 => x"ac",
          5066 => x"2e",
          5067 => x"2a",
          5068 => x"ff",
          5069 => x"a0",
          5070 => x"94",
          5071 => x"ff",
          5072 => x"2e",
          5073 => x"d1",
          5074 => x"d1",
          5075 => x"d1",
          5076 => x"98",
          5077 => x"8c",
          5078 => x"84",
          5079 => x"76",
          5080 => x"57",
          5081 => x"82",
          5082 => x"5d",
          5083 => x"80",
          5084 => x"5c",
          5085 => x"81",
          5086 => x"5b",
          5087 => x"77",
          5088 => x"81",
          5089 => x"58",
          5090 => x"70",
          5091 => x"70",
          5092 => x"09",
          5093 => x"38",
          5094 => x"07",
          5095 => x"7a",
          5096 => x"84",
          5097 => x"98",
          5098 => x"80",
          5099 => x"81",
          5100 => x"38",
          5101 => x"33",
          5102 => x"81",
          5103 => x"eb",
          5104 => x"07",
          5105 => x"75",
          5106 => x"3d",
          5107 => x"16",
          5108 => x"a5",
          5109 => x"17",
          5110 => x"07",
          5111 => x"88",
          5112 => x"52",
          5113 => x"70",
          5114 => x"17",
          5115 => x"38",
          5116 => x"70",
          5117 => x"71",
          5118 => x"1c",
          5119 => x"08",
          5120 => x"fb",
          5121 => x"0b",
          5122 => x"7a",
          5123 => x"53",
          5124 => x"ff",
          5125 => x"76",
          5126 => x"74",
          5127 => x"38",
          5128 => x"2b",
          5129 => x"d4",
          5130 => x"80",
          5131 => x"81",
          5132 => x"eb",
          5133 => x"07",
          5134 => x"81",
          5135 => x"81",
          5136 => x"81",
          5137 => x"09",
          5138 => x"76",
          5139 => x"f8",
          5140 => x"5a",
          5141 => x"a8",
          5142 => x"e5",
          5143 => x"05",
          5144 => x"33",
          5145 => x"56",
          5146 => x"75",
          5147 => x"8a",
          5148 => x"7b",
          5149 => x"81",
          5150 => x"1b",
          5151 => x"85",
          5152 => x"82",
          5153 => x"fa",
          5154 => x"97",
          5155 => x"2e",
          5156 => x"18",
          5157 => x"b7",
          5158 => x"97",
          5159 => x"18",
          5160 => x"70",
          5161 => x"05",
          5162 => x"5b",
          5163 => x"d1",
          5164 => x"0b",
          5165 => x"5a",
          5166 => x"7a",
          5167 => x"31",
          5168 => x"80",
          5169 => x"e1",
          5170 => x"59",
          5171 => x"39",
          5172 => x"33",
          5173 => x"81",
          5174 => x"81",
          5175 => x"78",
          5176 => x"7a",
          5177 => x"38",
          5178 => x"81",
          5179 => x"84",
          5180 => x"ff",
          5181 => x"79",
          5182 => x"84",
          5183 => x"71",
          5184 => x"d4",
          5185 => x"38",
          5186 => x"33",
          5187 => x"81",
          5188 => x"75",
          5189 => x"42",
          5190 => x"d2",
          5191 => x"84",
          5192 => x"33",
          5193 => x"81",
          5194 => x"75",
          5195 => x"5c",
          5196 => x"f2",
          5197 => x"84",
          5198 => x"33",
          5199 => x"81",
          5200 => x"75",
          5201 => x"84",
          5202 => x"33",
          5203 => x"81",
          5204 => x"75",
          5205 => x"59",
          5206 => x"5b",
          5207 => x"e4",
          5208 => x"e4",
          5209 => x"ec",
          5210 => x"18",
          5211 => x"f8",
          5212 => x"f2",
          5213 => x"53",
          5214 => x"52",
          5215 => x"8c",
          5216 => x"a4",
          5217 => x"34",
          5218 => x"40",
          5219 => x"82",
          5220 => x"8d",
          5221 => x"a0",
          5222 => x"91",
          5223 => x"e5",
          5224 => x"80",
          5225 => x"71",
          5226 => x"7d",
          5227 => x"61",
          5228 => x"11",
          5229 => x"71",
          5230 => x"72",
          5231 => x"ac",
          5232 => x"43",
          5233 => x"75",
          5234 => x"82",
          5235 => x"f2",
          5236 => x"83",
          5237 => x"f5",
          5238 => x"b4",
          5239 => x"78",
          5240 => x"e7",
          5241 => x"02",
          5242 => x"93",
          5243 => x"40",
          5244 => x"70",
          5245 => x"55",
          5246 => x"73",
          5247 => x"38",
          5248 => x"24",
          5249 => x"d1",
          5250 => x"80",
          5251 => x"54",
          5252 => x"34",
          5253 => x"7c",
          5254 => x"3d",
          5255 => x"3f",
          5256 => x"ba",
          5257 => x"0b",
          5258 => x"04",
          5259 => x"06",
          5260 => x"38",
          5261 => x"05",
          5262 => x"38",
          5263 => x"5f",
          5264 => x"70",
          5265 => x"05",
          5266 => x"55",
          5267 => x"70",
          5268 => x"16",
          5269 => x"16",
          5270 => x"30",
          5271 => x"2e",
          5272 => x"be",
          5273 => x"72",
          5274 => x"54",
          5275 => x"84",
          5276 => x"99",
          5277 => x"83",
          5278 => x"54",
          5279 => x"02",
          5280 => x"59",
          5281 => x"74",
          5282 => x"05",
          5283 => x"ed",
          5284 => x"84",
          5285 => x"80",
          5286 => x"8c",
          5287 => x"6d",
          5288 => x"9a",
          5289 => x"ba",
          5290 => x"77",
          5291 => x"ca",
          5292 => x"76",
          5293 => x"07",
          5294 => x"2a",
          5295 => x"d1",
          5296 => x"33",
          5297 => x"42",
          5298 => x"84",
          5299 => x"80",
          5300 => x"17",
          5301 => x"66",
          5302 => x"67",
          5303 => x"80",
          5304 => x"7c",
          5305 => x"80",
          5306 => x"1c",
          5307 => x"0b",
          5308 => x"83",
          5309 => x"38",
          5310 => x"53",
          5311 => x"38",
          5312 => x"38",
          5313 => x"39",
          5314 => x"2b",
          5315 => x"38",
          5316 => x"fe",
          5317 => x"80",
          5318 => x"06",
          5319 => x"81",
          5320 => x"89",
          5321 => x"f6",
          5322 => x"75",
          5323 => x"07",
          5324 => x"0c",
          5325 => x"33",
          5326 => x"73",
          5327 => x"83",
          5328 => x"0c",
          5329 => x"33",
          5330 => x"81",
          5331 => x"75",
          5332 => x"0c",
          5333 => x"57",
          5334 => x"23",
          5335 => x"1a",
          5336 => x"85",
          5337 => x"84",
          5338 => x"38",
          5339 => x"70",
          5340 => x"30",
          5341 => x"79",
          5342 => x"76",
          5343 => x"86",
          5344 => x"db",
          5345 => x"ba",
          5346 => x"57",
          5347 => x"cb",
          5348 => x"02",
          5349 => x"7d",
          5350 => x"55",
          5351 => x"57",
          5352 => x"57",
          5353 => x"57",
          5354 => x"51",
          5355 => x"78",
          5356 => x"38",
          5357 => x"57",
          5358 => x"94",
          5359 => x"2b",
          5360 => x"fc",
          5361 => x"bd",
          5362 => x"cb",
          5363 => x"ba",
          5364 => x"84",
          5365 => x"38",
          5366 => x"99",
          5367 => x"ff",
          5368 => x"83",
          5369 => x"94",
          5370 => x"27",
          5371 => x"0c",
          5372 => x"84",
          5373 => x"ff",
          5374 => x"94",
          5375 => x"fb",
          5376 => x"33",
          5377 => x"7e",
          5378 => x"17",
          5379 => x"0b",
          5380 => x"17",
          5381 => x"34",
          5382 => x"17",
          5383 => x"33",
          5384 => x"fb",
          5385 => x"7f",
          5386 => x"08",
          5387 => x"5a",
          5388 => x"38",
          5389 => x"81",
          5390 => x"84",
          5391 => x"ff",
          5392 => x"7e",
          5393 => x"57",
          5394 => x"79",
          5395 => x"16",
          5396 => x"17",
          5397 => x"84",
          5398 => x"06",
          5399 => x"83",
          5400 => x"08",
          5401 => x"74",
          5402 => x"82",
          5403 => x"81",
          5404 => x"16",
          5405 => x"52",
          5406 => x"3f",
          5407 => x"1a",
          5408 => x"98",
          5409 => x"83",
          5410 => x"9a",
          5411 => x"fe",
          5412 => x"f9",
          5413 => x"29",
          5414 => x"80",
          5415 => x"15",
          5416 => x"39",
          5417 => x"e4",
          5418 => x"da",
          5419 => x"79",
          5420 => x"5b",
          5421 => x"65",
          5422 => x"7e",
          5423 => x"38",
          5424 => x"38",
          5425 => x"38",
          5426 => x"59",
          5427 => x"55",
          5428 => x"38",
          5429 => x"38",
          5430 => x"56",
          5431 => x"1a",
          5432 => x"56",
          5433 => x"80",
          5434 => x"83",
          5435 => x"8a",
          5436 => x"06",
          5437 => x"38",
          5438 => x"84",
          5439 => x"38",
          5440 => x"1a",
          5441 => x"05",
          5442 => x"38",
          5443 => x"1b",
          5444 => x"83",
          5445 => x"59",
          5446 => x"77",
          5447 => x"75",
          5448 => x"7c",
          5449 => x"e0",
          5450 => x"38",
          5451 => x"80",
          5452 => x"31",
          5453 => x"80",
          5454 => x"58",
          5455 => x"77",
          5456 => x"55",
          5457 => x"7b",
          5458 => x"78",
          5459 => x"94",
          5460 => x"38",
          5461 => x"92",
          5462 => x"0c",
          5463 => x"8e",
          5464 => x"ff",
          5465 => x"7b",
          5466 => x"56",
          5467 => x"80",
          5468 => x"5f",
          5469 => x"e4",
          5470 => x"52",
          5471 => x"3f",
          5472 => x"38",
          5473 => x"0c",
          5474 => x"08",
          5475 => x"58",
          5476 => x"fe",
          5477 => x"33",
          5478 => x"16",
          5479 => x"74",
          5480 => x"81",
          5481 => x"da",
          5482 => x"19",
          5483 => x"1a",
          5484 => x"81",
          5485 => x"09",
          5486 => x"8c",
          5487 => x"a8",
          5488 => x"5c",
          5489 => x"e1",
          5490 => x"2e",
          5491 => x"54",
          5492 => x"53",
          5493 => x"9d",
          5494 => x"76",
          5495 => x"fe",
          5496 => x"51",
          5497 => x"08",
          5498 => x"51",
          5499 => x"08",
          5500 => x"74",
          5501 => x"81",
          5502 => x"ba",
          5503 => x"0b",
          5504 => x"8c",
          5505 => x"0d",
          5506 => x"5a",
          5507 => x"2e",
          5508 => x"2e",
          5509 => x"2e",
          5510 => x"22",
          5511 => x"38",
          5512 => x"82",
          5513 => x"82",
          5514 => x"2a",
          5515 => x"80",
          5516 => x"7b",
          5517 => x"38",
          5518 => x"81",
          5519 => x"82",
          5520 => x"05",
          5521 => x"aa",
          5522 => x"08",
          5523 => x"74",
          5524 => x"2e",
          5525 => x"88",
          5526 => x"0c",
          5527 => x"08",
          5528 => x"fe",
          5529 => x"58",
          5530 => x"16",
          5531 => x"05",
          5532 => x"38",
          5533 => x"77",
          5534 => x"5f",
          5535 => x"31",
          5536 => x"81",
          5537 => x"84",
          5538 => x"b4",
          5539 => x"78",
          5540 => x"18",
          5541 => x"74",
          5542 => x"81",
          5543 => x"ef",
          5544 => x"77",
          5545 => x"08",
          5546 => x"08",
          5547 => x"1e",
          5548 => x"75",
          5549 => x"1b",
          5550 => x"33",
          5551 => x"90",
          5552 => x"8c",
          5553 => x"ba",
          5554 => x"16",
          5555 => x"56",
          5556 => x"59",
          5557 => x"71",
          5558 => x"38",
          5559 => x"78",
          5560 => x"33",
          5561 => x"09",
          5562 => x"77",
          5563 => x"51",
          5564 => x"08",
          5565 => x"5c",
          5566 => x"38",
          5567 => x"11",
          5568 => x"58",
          5569 => x"81",
          5570 => x"57",
          5571 => x"60",
          5572 => x"a3",
          5573 => x"b8",
          5574 => x"40",
          5575 => x"ba",
          5576 => x"ff",
          5577 => x"17",
          5578 => x"31",
          5579 => x"a0",
          5580 => x"16",
          5581 => x"06",
          5582 => x"08",
          5583 => x"81",
          5584 => x"7e",
          5585 => x"57",
          5586 => x"83",
          5587 => x"60",
          5588 => x"58",
          5589 => x"fd",
          5590 => x"51",
          5591 => x"08",
          5592 => x"38",
          5593 => x"76",
          5594 => x"84",
          5595 => x"08",
          5596 => x"b4",
          5597 => x"81",
          5598 => x"3f",
          5599 => x"84",
          5600 => x"16",
          5601 => x"a0",
          5602 => x"16",
          5603 => x"06",
          5604 => x"08",
          5605 => x"81",
          5606 => x"60",
          5607 => x"51",
          5608 => x"08",
          5609 => x"74",
          5610 => x"81",
          5611 => x"70",
          5612 => x"96",
          5613 => x"c6",
          5614 => x"34",
          5615 => x"55",
          5616 => x"38",
          5617 => x"09",
          5618 => x"b4",
          5619 => x"76",
          5620 => x"87",
          5621 => x"1b",
          5622 => x"0b",
          5623 => x"8c",
          5624 => x"91",
          5625 => x"0c",
          5626 => x"7d",
          5627 => x"38",
          5628 => x"38",
          5629 => x"38",
          5630 => x"59",
          5631 => x"55",
          5632 => x"38",
          5633 => x"06",
          5634 => x"38",
          5635 => x"17",
          5636 => x"33",
          5637 => x"78",
          5638 => x"51",
          5639 => x"08",
          5640 => x"56",
          5641 => x"38",
          5642 => x"07",
          5643 => x"08",
          5644 => x"06",
          5645 => x"7a",
          5646 => x"9c",
          5647 => x"5b",
          5648 => x"18",
          5649 => x"2a",
          5650 => x"2a",
          5651 => x"2a",
          5652 => x"34",
          5653 => x"98",
          5654 => x"34",
          5655 => x"93",
          5656 => x"1c",
          5657 => x"84",
          5658 => x"bf",
          5659 => x"75",
          5660 => x"04",
          5661 => x"17",
          5662 => x"ff",
          5663 => x"8c",
          5664 => x"08",
          5665 => x"18",
          5666 => x"55",
          5667 => x"38",
          5668 => x"09",
          5669 => x"b4",
          5670 => x"7a",
          5671 => x"ef",
          5672 => x"90",
          5673 => x"88",
          5674 => x"18",
          5675 => x"2a",
          5676 => x"2a",
          5677 => x"2a",
          5678 => x"34",
          5679 => x"98",
          5680 => x"34",
          5681 => x"93",
          5682 => x"1c",
          5683 => x"84",
          5684 => x"bf",
          5685 => x"fe",
          5686 => x"90",
          5687 => x"06",
          5688 => x"08",
          5689 => x"0d",
          5690 => x"84",
          5691 => x"08",
          5692 => x"9e",
          5693 => x"96",
          5694 => x"8e",
          5695 => x"58",
          5696 => x"52",
          5697 => x"75",
          5698 => x"89",
          5699 => x"ff",
          5700 => x"81",
          5701 => x"08",
          5702 => x"ff",
          5703 => x"2e",
          5704 => x"33",
          5705 => x"2e",
          5706 => x"2e",
          5707 => x"80",
          5708 => x"e8",
          5709 => x"8c",
          5710 => x"8c",
          5711 => x"d0",
          5712 => x"53",
          5713 => x"73",
          5714 => x"73",
          5715 => x"83",
          5716 => x"56",
          5717 => x"75",
          5718 => x"12",
          5719 => x"38",
          5720 => x"54",
          5721 => x"89",
          5722 => x"54",
          5723 => x"51",
          5724 => x"38",
          5725 => x"70",
          5726 => x"07",
          5727 => x"38",
          5728 => x"78",
          5729 => x"cf",
          5730 => x"76",
          5731 => x"0d",
          5732 => x"99",
          5733 => x"8c",
          5734 => x"2e",
          5735 => x"98",
          5736 => x"98",
          5737 => x"84",
          5738 => x"08",
          5739 => x"33",
          5740 => x"24",
          5741 => x"70",
          5742 => x"80",
          5743 => x"33",
          5744 => x"73",
          5745 => x"83",
          5746 => x"74",
          5747 => x"04",
          5748 => x"81",
          5749 => x"ba",
          5750 => x"16",
          5751 => x"71",
          5752 => x"0c",
          5753 => x"12",
          5754 => x"98",
          5755 => x"80",
          5756 => x"5d",
          5757 => x"e4",
          5758 => x"3d",
          5759 => x"08",
          5760 => x"38",
          5761 => x"98",
          5762 => x"80",
          5763 => x"2e",
          5764 => x"3d",
          5765 => x"a4",
          5766 => x"84",
          5767 => x"80",
          5768 => x"08",
          5769 => x"08",
          5770 => x"c7",
          5771 => x"52",
          5772 => x"3f",
          5773 => x"38",
          5774 => x"0c",
          5775 => x"08",
          5776 => x"88",
          5777 => x"59",
          5778 => x"38",
          5779 => x"7a",
          5780 => x"8c",
          5781 => x"9f",
          5782 => x"f5",
          5783 => x"ba",
          5784 => x"08",
          5785 => x"88",
          5786 => x"59",
          5787 => x"38",
          5788 => x"8c",
          5789 => x"3f",
          5790 => x"8c",
          5791 => x"84",
          5792 => x"38",
          5793 => x"7a",
          5794 => x"82",
          5795 => x"90",
          5796 => x"17",
          5797 => x"38",
          5798 => x"95",
          5799 => x"17",
          5800 => x"3d",
          5801 => x"59",
          5802 => x"eb",
          5803 => x"11",
          5804 => x"3d",
          5805 => x"60",
          5806 => x"d1",
          5807 => x"fc",
          5808 => x"59",
          5809 => x"81",
          5810 => x"5a",
          5811 => x"78",
          5812 => x"27",
          5813 => x"7c",
          5814 => x"57",
          5815 => x"70",
          5816 => x"09",
          5817 => x"80",
          5818 => x"80",
          5819 => x"94",
          5820 => x"2b",
          5821 => x"f0",
          5822 => x"71",
          5823 => x"07",
          5824 => x"52",
          5825 => x"ba",
          5826 => x"80",
          5827 => x"81",
          5828 => x"70",
          5829 => x"88",
          5830 => x"08",
          5831 => x"83",
          5832 => x"08",
          5833 => x"74",
          5834 => x"82",
          5835 => x"81",
          5836 => x"16",
          5837 => x"52",
          5838 => x"3f",
          5839 => x"80",
          5840 => x"7b",
          5841 => x"70",
          5842 => x"08",
          5843 => x"7e",
          5844 => x"38",
          5845 => x"18",
          5846 => x"70",
          5847 => x"fe",
          5848 => x"81",
          5849 => x"81",
          5850 => x"38",
          5851 => x"34",
          5852 => x"3d",
          5853 => x"58",
          5854 => x"38",
          5855 => x"38",
          5856 => x"38",
          5857 => x"59",
          5858 => x"53",
          5859 => x"38",
          5860 => x"38",
          5861 => x"81",
          5862 => x"58",
          5863 => x"8a",
          5864 => x"56",
          5865 => x"52",
          5866 => x"84",
          5867 => x"70",
          5868 => x"84",
          5869 => x"38",
          5870 => x"0c",
          5871 => x"58",
          5872 => x"75",
          5873 => x"31",
          5874 => x"90",
          5875 => x"51",
          5876 => x"38",
          5877 => x"3f",
          5878 => x"8c",
          5879 => x"ff",
          5880 => x"b4",
          5881 => x"27",
          5882 => x"ff",
          5883 => x"81",
          5884 => x"3d",
          5885 => x"2a",
          5886 => x"38",
          5887 => x"58",
          5888 => x"b6",
          5889 => x"08",
          5890 => x"8c",
          5891 => x"07",
          5892 => x"ff",
          5893 => x"9c",
          5894 => x"9c",
          5895 => x"0c",
          5896 => x"16",
          5897 => x"2e",
          5898 => x"73",
          5899 => x"39",
          5900 => x"08",
          5901 => x"06",
          5902 => x"fe",
          5903 => x"55",
          5904 => x"8a",
          5905 => x"08",
          5906 => x"53",
          5907 => x"15",
          5908 => x"74",
          5909 => x"8c",
          5910 => x"33",
          5911 => x"8c",
          5912 => x"38",
          5913 => x"39",
          5914 => x"3f",
          5915 => x"8c",
          5916 => x"8c",
          5917 => x"ba",
          5918 => x"16",
          5919 => x"16",
          5920 => x"8b",
          5921 => x"56",
          5922 => x"80",
          5923 => x"3d",
          5924 => x"ba",
          5925 => x"80",
          5926 => x"54",
          5927 => x"0d",
          5928 => x"51",
          5929 => x"08",
          5930 => x"38",
          5931 => x"59",
          5932 => x"33",
          5933 => x"79",
          5934 => x"08",
          5935 => x"88",
          5936 => x"5a",
          5937 => x"77",
          5938 => x"22",
          5939 => x"ff",
          5940 => x"55",
          5941 => x"2e",
          5942 => x"fe",
          5943 => x"f6",
          5944 => x"71",
          5945 => x"07",
          5946 => x"39",
          5947 => x"74",
          5948 => x"72",
          5949 => x"71",
          5950 => x"84",
          5951 => x"94",
          5952 => x"38",
          5953 => x"0c",
          5954 => x"51",
          5955 => x"08",
          5956 => x"75",
          5957 => x"0d",
          5958 => x"80",
          5959 => x"80",
          5960 => x"80",
          5961 => x"16",
          5962 => x"97",
          5963 => x"75",
          5964 => x"f3",
          5965 => x"bd",
          5966 => x"ba",
          5967 => x"ba",
          5968 => x"51",
          5969 => x"51",
          5970 => x"08",
          5971 => x"9f",
          5972 => x"57",
          5973 => x"3d",
          5974 => x"53",
          5975 => x"51",
          5976 => x"08",
          5977 => x"9f",
          5978 => x"57",
          5979 => x"ff",
          5980 => x"84",
          5981 => x"81",
          5982 => x"84",
          5983 => x"fe",
          5984 => x"fe",
          5985 => x"80",
          5986 => x"52",
          5987 => x"08",
          5988 => x"8a",
          5989 => x"3d",
          5990 => x"b5",
          5991 => x"84",
          5992 => x"cb",
          5993 => x"80",
          5994 => x"d1",
          5995 => x"bd",
          5996 => x"3d",
          5997 => x"0c",
          5998 => x"66",
          5999 => x"ec",
          6000 => x"3f",
          6001 => x"8c",
          6002 => x"08",
          6003 => x"08",
          6004 => x"8d",
          6005 => x"8c",
          6006 => x"8c",
          6007 => x"2e",
          6008 => x"84",
          6009 => x"80",
          6010 => x"5d",
          6011 => x"ef",
          6012 => x"7c",
          6013 => x"b8",
          6014 => x"fc",
          6015 => x"2e",
          6016 => x"b4",
          6017 => x"80",
          6018 => x"2e",
          6019 => x"83",
          6020 => x"2b",
          6021 => x"70",
          6022 => x"80",
          6023 => x"30",
          6024 => x"05",
          6025 => x"41",
          6026 => x"5e",
          6027 => x"0c",
          6028 => x"81",
          6029 => x"84",
          6030 => x"81",
          6031 => x"70",
          6032 => x"fc",
          6033 => x"08",
          6034 => x"83",
          6035 => x"08",
          6036 => x"74",
          6037 => x"82",
          6038 => x"81",
          6039 => x"17",
          6040 => x"52",
          6041 => x"3f",
          6042 => x"42",
          6043 => x"51",
          6044 => x"08",
          6045 => x"8c",
          6046 => x"ba",
          6047 => x"08",
          6048 => x"62",
          6049 => x"76",
          6050 => x"94",
          6051 => x"58",
          6052 => x"77",
          6053 => x"33",
          6054 => x"80",
          6055 => x"ff",
          6056 => x"55",
          6057 => x"77",
          6058 => x"5a",
          6059 => x"84",
          6060 => x"18",
          6061 => x"5a",
          6062 => x"89",
          6063 => x"08",
          6064 => x"33",
          6065 => x"15",
          6066 => x"78",
          6067 => x"5a",
          6068 => x"56",
          6069 => x"70",
          6070 => x"55",
          6071 => x"17",
          6072 => x"b7",
          6073 => x"08",
          6074 => x"88",
          6075 => x"38",
          6076 => x"94",
          6077 => x"c0",
          6078 => x"80",
          6079 => x"75",
          6080 => x"3d",
          6081 => x"80",
          6082 => x"fe",
          6083 => x"84",
          6084 => x"38",
          6085 => x"d8",
          6086 => x"82",
          6087 => x"51",
          6088 => x"08",
          6089 => x"11",
          6090 => x"74",
          6091 => x"17",
          6092 => x"73",
          6093 => x"26",
          6094 => x"33",
          6095 => x"8c",
          6096 => x"38",
          6097 => x"39",
          6098 => x"73",
          6099 => x"c7",
          6100 => x"fe",
          6101 => x"ff",
          6102 => x"08",
          6103 => x"ae",
          6104 => x"9c",
          6105 => x"ba",
          6106 => x"58",
          6107 => x"08",
          6108 => x"08",
          6109 => x"74",
          6110 => x"52",
          6111 => x"ba",
          6112 => x"80",
          6113 => x"fc",
          6114 => x"84",
          6115 => x"38",
          6116 => x"dc",
          6117 => x"80",
          6118 => x"51",
          6119 => x"08",
          6120 => x"11",
          6121 => x"74",
          6122 => x"0c",
          6123 => x"84",
          6124 => x"ff",
          6125 => x"17",
          6126 => x"fe",
          6127 => x"59",
          6128 => x"39",
          6129 => x"fe",
          6130 => x"18",
          6131 => x"0b",
          6132 => x"39",
          6133 => x"81",
          6134 => x"82",
          6135 => x"a8",
          6136 => x"ba",
          6137 => x"80",
          6138 => x"0c",
          6139 => x"3d",
          6140 => x"ff",
          6141 => x"56",
          6142 => x"81",
          6143 => x"06",
          6144 => x"76",
          6145 => x"38",
          6146 => x"06",
          6147 => x"38",
          6148 => x"9a",
          6149 => x"33",
          6150 => x"2e",
          6151 => x"06",
          6152 => x"87",
          6153 => x"83",
          6154 => x"8c",
          6155 => x"ff",
          6156 => x"56",
          6157 => x"84",
          6158 => x"91",
          6159 => x"84",
          6160 => x"84",
          6161 => x"95",
          6162 => x"2b",
          6163 => x"5d",
          6164 => x"08",
          6165 => x"08",
          6166 => x"3d",
          6167 => x"80",
          6168 => x"8b",
          6169 => x"84",
          6170 => x"75",
          6171 => x"5a",
          6172 => x"2e",
          6173 => x"81",
          6174 => x"7b",
          6175 => x"fd",
          6176 => x"3f",
          6177 => x"0c",
          6178 => x"98",
          6179 => x"08",
          6180 => x"33",
          6181 => x"81",
          6182 => x"53",
          6183 => x"fe",
          6184 => x"80",
          6185 => x"75",
          6186 => x"38",
          6187 => x"81",
          6188 => x"7c",
          6189 => x"51",
          6190 => x"08",
          6191 => x"ff",
          6192 => x"06",
          6193 => x"39",
          6194 => x"52",
          6195 => x"3f",
          6196 => x"2e",
          6197 => x"ba",
          6198 => x"08",
          6199 => x"08",
          6200 => x"fe",
          6201 => x"82",
          6202 => x"81",
          6203 => x"05",
          6204 => x"fe",
          6205 => x"39",
          6206 => x"38",
          6207 => x"3f",
          6208 => x"8c",
          6209 => x"ba",
          6210 => x"84",
          6211 => x"38",
          6212 => x"fd",
          6213 => x"38",
          6214 => x"08",
          6215 => x"b0",
          6216 => x"17",
          6217 => x"34",
          6218 => x"38",
          6219 => x"fd",
          6220 => x"fd",
          6221 => x"e3",
          6222 => x"bc",
          6223 => x"c0",
          6224 => x"ba",
          6225 => x"84",
          6226 => x"7d",
          6227 => x"5a",
          6228 => x"08",
          6229 => x"88",
          6230 => x"0d",
          6231 => x"09",
          6232 => x"05",
          6233 => x"58",
          6234 => x"5f",
          6235 => x"ff",
          6236 => x"75",
          6237 => x"38",
          6238 => x"2e",
          6239 => x"ff",
          6240 => x"38",
          6241 => x"33",
          6242 => x"fe",
          6243 => x"56",
          6244 => x"8a",
          6245 => x"08",
          6246 => x"b8",
          6247 => x"80",
          6248 => x"15",
          6249 => x"17",
          6250 => x"38",
          6251 => x"81",
          6252 => x"84",
          6253 => x"18",
          6254 => x"39",
          6255 => x"17",
          6256 => x"fe",
          6257 => x"8c",
          6258 => x"83",
          6259 => x"08",
          6260 => x"fe",
          6261 => x"82",
          6262 => x"75",
          6263 => x"05",
          6264 => x"fe",
          6265 => x"56",
          6266 => x"27",
          6267 => x"27",
          6268 => x"fe",
          6269 => x"5a",
          6270 => x"96",
          6271 => x"fd",
          6272 => x"2e",
          6273 => x"76",
          6274 => x"8c",
          6275 => x"fe",
          6276 => x"77",
          6277 => x"18",
          6278 => x"7b",
          6279 => x"26",
          6280 => x"0c",
          6281 => x"55",
          6282 => x"56",
          6283 => x"f0",
          6284 => x"a0",
          6285 => x"16",
          6286 => x"0b",
          6287 => x"80",
          6288 => x"ce",
          6289 => x"a1",
          6290 => x"0b",
          6291 => x"ff",
          6292 => x"17",
          6293 => x"d3",
          6294 => x"2e",
          6295 => x"80",
          6296 => x"74",
          6297 => x"81",
          6298 => x"ef",
          6299 => x"17",
          6300 => x"06",
          6301 => x"34",
          6302 => x"17",
          6303 => x"80",
          6304 => x"1c",
          6305 => x"84",
          6306 => x"08",
          6307 => x"8c",
          6308 => x"08",
          6309 => x"34",
          6310 => x"6a",
          6311 => x"88",
          6312 => x"33",
          6313 => x"69",
          6314 => x"57",
          6315 => x"fe",
          6316 => x"56",
          6317 => x"0d",
          6318 => x"ec",
          6319 => x"80",
          6320 => x"90",
          6321 => x"7a",
          6322 => x"34",
          6323 => x"b8",
          6324 => x"7b",
          6325 => x"77",
          6326 => x"69",
          6327 => x"57",
          6328 => x"fe",
          6329 => x"56",
          6330 => x"3d",
          6331 => x"79",
          6332 => x"05",
          6333 => x"75",
          6334 => x"38",
          6335 => x"53",
          6336 => x"3d",
          6337 => x"8c",
          6338 => x"2e",
          6339 => x"b1",
          6340 => x"b2",
          6341 => x"59",
          6342 => x"08",
          6343 => x"02",
          6344 => x"5d",
          6345 => x"92",
          6346 => x"75",
          6347 => x"81",
          6348 => x"ef",
          6349 => x"58",
          6350 => x"33",
          6351 => x"15",
          6352 => x"52",
          6353 => x"ba",
          6354 => x"85",
          6355 => x"81",
          6356 => x"0c",
          6357 => x"11",
          6358 => x"74",
          6359 => x"81",
          6360 => x"7a",
          6361 => x"83",
          6362 => x"5f",
          6363 => x"33",
          6364 => x"9f",
          6365 => x"89",
          6366 => x"57",
          6367 => x"26",
          6368 => x"06",
          6369 => x"59",
          6370 => x"85",
          6371 => x"32",
          6372 => x"7a",
          6373 => x"95",
          6374 => x"7b",
          6375 => x"7e",
          6376 => x"24",
          6377 => x"53",
          6378 => x"3d",
          6379 => x"8c",
          6380 => x"b2",
          6381 => x"08",
          6382 => x"77",
          6383 => x"8c",
          6384 => x"92",
          6385 => x"02",
          6386 => x"5a",
          6387 => x"70",
          6388 => x"79",
          6389 => x"8b",
          6390 => x"2a",
          6391 => x"75",
          6392 => x"7f",
          6393 => x"18",
          6394 => x"5c",
          6395 => x"3d",
          6396 => x"9b",
          6397 => x"2b",
          6398 => x"7d",
          6399 => x"9c",
          6400 => x"7d",
          6401 => x"76",
          6402 => x"5e",
          6403 => x"7a",
          6404 => x"aa",
          6405 => x"bc",
          6406 => x"52",
          6407 => x"3f",
          6408 => x"38",
          6409 => x"0c",
          6410 => x"56",
          6411 => x"5a",
          6412 => x"38",
          6413 => x"56",
          6414 => x"2a",
          6415 => x"33",
          6416 => x"93",
          6417 => x"ec",
          6418 => x"80",
          6419 => x"83",
          6420 => x"b2",
          6421 => x"2e",
          6422 => x"fb",
          6423 => x"84",
          6424 => x"16",
          6425 => x"b4",
          6426 => x"16",
          6427 => x"09",
          6428 => x"76",
          6429 => x"51",
          6430 => x"08",
          6431 => x"58",
          6432 => x"aa",
          6433 => x"34",
          6434 => x"08",
          6435 => x"51",
          6436 => x"08",
          6437 => x"ff",
          6438 => x"f9",
          6439 => x"38",
          6440 => x"ba",
          6441 => x"3d",
          6442 => x"0c",
          6443 => x"94",
          6444 => x"2b",
          6445 => x"8d",
          6446 => x"fb",
          6447 => x"2e",
          6448 => x"0c",
          6449 => x"16",
          6450 => x"51",
          6451 => x"ba",
          6452 => x"fe",
          6453 => x"17",
          6454 => x"31",
          6455 => x"a0",
          6456 => x"16",
          6457 => x"06",
          6458 => x"08",
          6459 => x"81",
          6460 => x"79",
          6461 => x"17",
          6462 => x"18",
          6463 => x"81",
          6464 => x"38",
          6465 => x"b4",
          6466 => x"ba",
          6467 => x"08",
          6468 => x"5d",
          6469 => x"81",
          6470 => x"18",
          6471 => x"33",
          6472 => x"fb",
          6473 => x"df",
          6474 => x"05",
          6475 => x"cc",
          6476 => x"d8",
          6477 => x"ba",
          6478 => x"84",
          6479 => x"78",
          6480 => x"51",
          6481 => x"08",
          6482 => x"02",
          6483 => x"54",
          6484 => x"06",
          6485 => x"06",
          6486 => x"55",
          6487 => x"0b",
          6488 => x"9a",
          6489 => x"8c",
          6490 => x"0d",
          6491 => x"05",
          6492 => x"3f",
          6493 => x"8c",
          6494 => x"ba",
          6495 => x"5a",
          6496 => x"ff",
          6497 => x"55",
          6498 => x"80",
          6499 => x"86",
          6500 => x"22",
          6501 => x"59",
          6502 => x"88",
          6503 => x"90",
          6504 => x"98",
          6505 => x"57",
          6506 => x"fe",
          6507 => x"84",
          6508 => x"e8",
          6509 => x"53",
          6510 => x"51",
          6511 => x"08",
          6512 => x"ba",
          6513 => x"57",
          6514 => x"76",
          6515 => x"76",
          6516 => x"5b",
          6517 => x"70",
          6518 => x"81",
          6519 => x"56",
          6520 => x"82",
          6521 => x"55",
          6522 => x"98",
          6523 => x"52",
          6524 => x"3f",
          6525 => x"38",
          6526 => x"0c",
          6527 => x"33",
          6528 => x"2e",
          6529 => x"2e",
          6530 => x"05",
          6531 => x"90",
          6532 => x"33",
          6533 => x"71",
          6534 => x"59",
          6535 => x"3d",
          6536 => x"52",
          6537 => x"8b",
          6538 => x"ba",
          6539 => x"76",
          6540 => x"38",
          6541 => x"39",
          6542 => x"16",
          6543 => x"fe",
          6544 => x"8c",
          6545 => x"e8",
          6546 => x"34",
          6547 => x"84",
          6548 => x"17",
          6549 => x"33",
          6550 => x"fe",
          6551 => x"a0",
          6552 => x"16",
          6553 => x"59",
          6554 => x"81",
          6555 => x"84",
          6556 => x"38",
          6557 => x"fe",
          6558 => x"57",
          6559 => x"84",
          6560 => x"66",
          6561 => x"7c",
          6562 => x"34",
          6563 => x"38",
          6564 => x"34",
          6565 => x"18",
          6566 => x"79",
          6567 => x"79",
          6568 => x"82",
          6569 => x"a2",
          6570 => x"ba",
          6571 => x"82",
          6572 => x"57",
          6573 => x"34",
          6574 => x"a3",
          6575 => x"06",
          6576 => x"81",
          6577 => x"5c",
          6578 => x"55",
          6579 => x"74",
          6580 => x"74",
          6581 => x"84",
          6582 => x"84",
          6583 => x"57",
          6584 => x"e7",
          6585 => x"81",
          6586 => x"2e",
          6587 => x"2e",
          6588 => x"81",
          6589 => x"2e",
          6590 => x"06",
          6591 => x"78",
          6592 => x"81",
          6593 => x"38",
          6594 => x"88",
          6595 => x"5d",
          6596 => x"81",
          6597 => x"08",
          6598 => x"58",
          6599 => x"38",
          6600 => x"81",
          6601 => x"99",
          6602 => x"70",
          6603 => x"81",
          6604 => x"ed",
          6605 => x"95",
          6606 => x"3f",
          6607 => x"8c",
          6608 => x"75",
          6609 => x"04",
          6610 => x"3f",
          6611 => x"06",
          6612 => x"75",
          6613 => x"04",
          6614 => x"39",
          6615 => x"3f",
          6616 => x"8c",
          6617 => x"82",
          6618 => x"55",
          6619 => x"70",
          6620 => x"74",
          6621 => x"1e",
          6622 => x"84",
          6623 => x"87",
          6624 => x"86",
          6625 => x"08",
          6626 => x"38",
          6627 => x"38",
          6628 => x"fe",
          6629 => x"57",
          6630 => x"81",
          6631 => x"08",
          6632 => x"57",
          6633 => x"b2",
          6634 => x"2e",
          6635 => x"54",
          6636 => x"33",
          6637 => x"8c",
          6638 => x"81",
          6639 => x"78",
          6640 => x"33",
          6641 => x"81",
          6642 => x"78",
          6643 => x"d7",
          6644 => x"a5",
          6645 => x"a1",
          6646 => x"ba",
          6647 => x"87",
          6648 => x"76",
          6649 => x"57",
          6650 => x"34",
          6651 => x"56",
          6652 => x"7e",
          6653 => x"58",
          6654 => x"ff",
          6655 => x"38",
          6656 => x"70",
          6657 => x"74",
          6658 => x"e5",
          6659 => x"1e",
          6660 => x"84",
          6661 => x"81",
          6662 => x"18",
          6663 => x"51",
          6664 => x"08",
          6665 => x"38",
          6666 => x"b4",
          6667 => x"7b",
          6668 => x"18",
          6669 => x"84",
          6670 => x"74",
          6671 => x"d1",
          6672 => x"ba",
          6673 => x"fe",
          6674 => x"80",
          6675 => x"81",
          6676 => x"05",
          6677 => x"fe",
          6678 => x"3d",
          6679 => x"cb",
          6680 => x"76",
          6681 => x"74",
          6682 => x"73",
          6683 => x"84",
          6684 => x"81",
          6685 => x"81",
          6686 => x"81",
          6687 => x"38",
          6688 => x"17",
          6689 => x"5d",
          6690 => x"8a",
          6691 => x"7c",
          6692 => x"3f",
          6693 => x"72",
          6694 => x"05",
          6695 => x"55",
          6696 => x"19",
          6697 => x"77",
          6698 => x"76",
          6699 => x"7f",
          6700 => x"83",
          6701 => x"81",
          6702 => x"08",
          6703 => x"8c",
          6704 => x"78",
          6705 => x"09",
          6706 => x"54",
          6707 => x"0d",
          6708 => x"90",
          6709 => x"fe",
          6710 => x"81",
          6711 => x"77",
          6712 => x"80",
          6713 => x"58",
          6714 => x"54",
          6715 => x"53",
          6716 => x"3f",
          6717 => x"8c",
          6718 => x"ff",
          6719 => x"7e",
          6720 => x"2e",
          6721 => x"79",
          6722 => x"c0",
          6723 => x"15",
          6724 => x"5a",
          6725 => x"7d",
          6726 => x"81",
          6727 => x"54",
          6728 => x"39",
          6729 => x"82",
          6730 => x"c0",
          6731 => x"84",
          6732 => x"3d",
          6733 => x"81",
          6734 => x"0b",
          6735 => x"79",
          6736 => x"81",
          6737 => x"56",
          6738 => x"ed",
          6739 => x"84",
          6740 => x"84",
          6741 => x"d4",
          6742 => x"2e",
          6743 => x"84",
          6744 => x"12",
          6745 => x"51",
          6746 => x"08",
          6747 => x"56",
          6748 => x"82",
          6749 => x"84",
          6750 => x"83",
          6751 => x"84",
          6752 => x"55",
          6753 => x"82",
          6754 => x"15",
          6755 => x"7e",
          6756 => x"26",
          6757 => x"26",
          6758 => x"55",
          6759 => x"a6",
          6760 => x"77",
          6761 => x"85",
          6762 => x"77",
          6763 => x"b0",
          6764 => x"81",
          6765 => x"fe",
          6766 => x"8c",
          6767 => x"05",
          6768 => x"88",
          6769 => x"82",
          6770 => x"f8",
          6771 => x"b2",
          6772 => x"82",
          6773 => x"33",
          6774 => x"88",
          6775 => x"07",
          6776 => x"ba",
          6777 => x"71",
          6778 => x"14",
          6779 => x"33",
          6780 => x"a3",
          6781 => x"54",
          6782 => x"4d",
          6783 => x"90",
          6784 => x"82",
          6785 => x"06",
          6786 => x"38",
          6787 => x"89",
          6788 => x"f4",
          6789 => x"43",
          6790 => x"38",
          6791 => x"81",
          6792 => x"74",
          6793 => x"98",
          6794 => x"82",
          6795 => x"80",
          6796 => x"38",
          6797 => x"3f",
          6798 => x"55",
          6799 => x"96",
          6800 => x"10",
          6801 => x"72",
          6802 => x"ff",
          6803 => x"47",
          6804 => x"11",
          6805 => x"58",
          6806 => x"b8",
          6807 => x"16",
          6808 => x"26",
          6809 => x"31",
          6810 => x"fc",
          6811 => x"40",
          6812 => x"82",
          6813 => x"83",
          6814 => x"27",
          6815 => x"77",
          6816 => x"ef",
          6817 => x"57",
          6818 => x"0d",
          6819 => x"fb",
          6820 => x"0c",
          6821 => x"04",
          6822 => x"06",
          6823 => x"38",
          6824 => x"05",
          6825 => x"38",
          6826 => x"7d",
          6827 => x"05",
          6828 => x"33",
          6829 => x"99",
          6830 => x"ff",
          6831 => x"64",
          6832 => x"81",
          6833 => x"9f",
          6834 => x"81",
          6835 => x"75",
          6836 => x"9f",
          6837 => x"80",
          6838 => x"1f",
          6839 => x"38",
          6840 => x"f8",
          6841 => x"ca",
          6842 => x"08",
          6843 => x"06",
          6844 => x"83",
          6845 => x"7e",
          6846 => x"31",
          6847 => x"d2",
          6848 => x"7b",
          6849 => x"39",
          6850 => x"80",
          6851 => x"30",
          6852 => x"ba",
          6853 => x"7a",
          6854 => x"7b",
          6855 => x"84",
          6856 => x"ba",
          6857 => x"2e",
          6858 => x"8b",
          6859 => x"7a",
          6860 => x"55",
          6861 => x"ff",
          6862 => x"83",
          6863 => x"81",
          6864 => x"58",
          6865 => x"60",
          6866 => x"61",
          6867 => x"34",
          6868 => x"61",
          6869 => x"7b",
          6870 => x"05",
          6871 => x"48",
          6872 => x"2a",
          6873 => x"34",
          6874 => x"86",
          6875 => x"55",
          6876 => x"2a",
          6877 => x"61",
          6878 => x"34",
          6879 => x"9a",
          6880 => x"7e",
          6881 => x"48",
          6882 => x"2a",
          6883 => x"98",
          6884 => x"98",
          6885 => x"2e",
          6886 => x"34",
          6887 => x"a9",
          6888 => x"34",
          6889 => x"61",
          6890 => x"6a",
          6891 => x"a4",
          6892 => x"93",
          6893 => x"57",
          6894 => x"76",
          6895 => x"55",
          6896 => x"49",
          6897 => x"05",
          6898 => x"7e",
          6899 => x"8f",
          6900 => x"fa",
          6901 => x"2e",
          6902 => x"80",
          6903 => x"15",
          6904 => x"5b",
          6905 => x"ff",
          6906 => x"38",
          6907 => x"2a",
          6908 => x"05",
          6909 => x"64",
          6910 => x"2a",
          6911 => x"59",
          6912 => x"78",
          6913 => x"fe",
          6914 => x"85",
          6915 => x"80",
          6916 => x"15",
          6917 => x"7a",
          6918 => x"81",
          6919 => x"38",
          6920 => x"66",
          6921 => x"38",
          6922 => x"52",
          6923 => x"ba",
          6924 => x"76",
          6925 => x"8c",
          6926 => x"58",
          6927 => x"84",
          6928 => x"58",
          6929 => x"81",
          6930 => x"80",
          6931 => x"05",
          6932 => x"38",
          6933 => x"34",
          6934 => x"34",
          6935 => x"82",
          6936 => x"77",
          6937 => x"fd",
          6938 => x"d1",
          6939 => x"ba",
          6940 => x"76",
          6941 => x"08",
          6942 => x"c6",
          6943 => x"34",
          6944 => x"ba",
          6945 => x"62",
          6946 => x"2a",
          6947 => x"62",
          6948 => x"05",
          6949 => x"83",
          6950 => x"60",
          6951 => x"81",
          6952 => x"38",
          6953 => x"c3",
          6954 => x"08",
          6955 => x"84",
          6956 => x"ba",
          6957 => x"39",
          6958 => x"c4",
          6959 => x"57",
          6960 => x"58",
          6961 => x"26",
          6962 => x"10",
          6963 => x"74",
          6964 => x"ee",
          6965 => x"f9",
          6966 => x"84",
          6967 => x"a0",
          6968 => x"fc",
          6969 => x"f0",
          6970 => x"57",
          6971 => x"83",
          6972 => x"f8",
          6973 => x"f4",
          6974 => x"68",
          6975 => x"af",
          6976 => x"61",
          6977 => x"68",
          6978 => x"5b",
          6979 => x"2a",
          6980 => x"c6",
          6981 => x"80",
          6982 => x"80",
          6983 => x"c6",
          6984 => x"7c",
          6985 => x"34",
          6986 => x"05",
          6987 => x"a7",
          6988 => x"80",
          6989 => x"05",
          6990 => x"61",
          6991 => x"34",
          6992 => x"b3",
          6993 => x"05",
          6994 => x"93",
          6995 => x"59",
          6996 => x"33",
          6997 => x"15",
          6998 => x"76",
          6999 => x"81",
          7000 => x"da",
          7001 => x"53",
          7002 => x"3f",
          7003 => x"b0",
          7004 => x"77",
          7005 => x"84",
          7006 => x"51",
          7007 => x"81",
          7008 => x"0d",
          7009 => x"34",
          7010 => x"4c",
          7011 => x"34",
          7012 => x"34",
          7013 => x"86",
          7014 => x"ff",
          7015 => x"05",
          7016 => x"65",
          7017 => x"54",
          7018 => x"fe",
          7019 => x"57",
          7020 => x"ff",
          7021 => x"80",
          7022 => x"7b",
          7023 => x"57",
          7024 => x"57",
          7025 => x"61",
          7026 => x"83",
          7027 => x"e6",
          7028 => x"05",
          7029 => x"83",
          7030 => x"78",
          7031 => x"2a",
          7032 => x"7a",
          7033 => x"05",
          7034 => x"76",
          7035 => x"83",
          7036 => x"05",
          7037 => x"6b",
          7038 => x"52",
          7039 => x"54",
          7040 => x"fe",
          7041 => x"f7",
          7042 => x"5b",
          7043 => x"57",
          7044 => x"3d",
          7045 => x"53",
          7046 => x"3f",
          7047 => x"38",
          7048 => x"90",
          7049 => x"34",
          7050 => x"38",
          7051 => x"34",
          7052 => x"74",
          7053 => x"04",
          7054 => x"b3",
          7055 => x"80",
          7056 => x"76",
          7057 => x"17",
          7058 => x"81",
          7059 => x"74",
          7060 => x"0c",
          7061 => x"05",
          7062 => x"08",
          7063 => x"32",
          7064 => x"70",
          7065 => x"1b",
          7066 => x"52",
          7067 => x"39",
          7068 => x"33",
          7069 => x"57",
          7070 => x"34",
          7071 => x"3d",
          7072 => x"f7",
          7073 => x"c0",
          7074 => x"59",
          7075 => x"bb",
          7076 => x"81",
          7077 => x"75",
          7078 => x"11",
          7079 => x"08",
          7080 => x"8c",
          7081 => x"38",
          7082 => x"3d",
          7083 => x"55",
          7084 => x"51",
          7085 => x"70",
          7086 => x"30",
          7087 => x"8d",
          7088 => x"81",
          7089 => x"3d",
          7090 => x"84",
          7091 => x"52",
          7092 => x"83",
          7093 => x"8c",
          7094 => x"ff",
          7095 => x"09",
          7096 => x"e4",
          7097 => x"71",
          7098 => x"ff",
          7099 => x"26",
          7100 => x"05",
          7101 => x"80",
          7102 => x"8c",
          7103 => x"3d",
          7104 => x"05",
          7105 => x"70",
          7106 => x"72",
          7107 => x"04",
          7108 => x"ef",
          7109 => x"70",
          7110 => x"84",
          7111 => x"04",
          7112 => x"ff",
          7113 => x"ff",
          7114 => x"75",
          7115 => x"70",
          7116 => x"70",
          7117 => x"56",
          7118 => x"82",
          7119 => x"54",
          7120 => x"54",
          7121 => x"38",
          7122 => x"52",
          7123 => x"75",
          7124 => x"80",
          7125 => x"ba",
          7126 => x"ed",
          7127 => x"26",
          7128 => x"a8",
          7129 => x"16",
          7130 => x"75",
          7131 => x"83",
          7132 => x"88",
          7133 => x"51",
          7134 => x"ff",
          7135 => x"70",
          7136 => x"39",
          7137 => x"57",
          7138 => x"ff",
          7139 => x"75",
          7140 => x"70",
          7141 => x"ff",
          7142 => x"05",
          7143 => x"00",
          7144 => x"ff",
          7145 => x"00",
          7146 => x"80",
          7147 => x"6a",
          7148 => x"54",
          7149 => x"3e",
          7150 => x"28",
          7151 => x"12",
          7152 => x"fc",
          7153 => x"e6",
          7154 => x"d0",
          7155 => x"ba",
          7156 => x"59",
          7157 => x"59",
          7158 => x"59",
          7159 => x"59",
          7160 => x"59",
          7161 => x"59",
          7162 => x"59",
          7163 => x"59",
          7164 => x"59",
          7165 => x"59",
          7166 => x"59",
          7167 => x"59",
          7168 => x"59",
          7169 => x"59",
          7170 => x"59",
          7171 => x"59",
          7172 => x"59",
          7173 => x"59",
          7174 => x"59",
          7175 => x"59",
          7176 => x"59",
          7177 => x"7b",
          7178 => x"59",
          7179 => x"59",
          7180 => x"59",
          7181 => x"59",
          7182 => x"59",
          7183 => x"59",
          7184 => x"59",
          7185 => x"59",
          7186 => x"10",
          7187 => x"94",
          7188 => x"71",
          7189 => x"d8",
          7190 => x"59",
          7191 => x"59",
          7192 => x"59",
          7193 => x"59",
          7194 => x"59",
          7195 => x"59",
          7196 => x"59",
          7197 => x"59",
          7198 => x"59",
          7199 => x"59",
          7200 => x"59",
          7201 => x"59",
          7202 => x"59",
          7203 => x"59",
          7204 => x"59",
          7205 => x"59",
          7206 => x"59",
          7207 => x"59",
          7208 => x"59",
          7209 => x"59",
          7210 => x"59",
          7211 => x"59",
          7212 => x"59",
          7213 => x"59",
          7214 => x"59",
          7215 => x"59",
          7216 => x"7a",
          7217 => x"59",
          7218 => x"59",
          7219 => x"59",
          7220 => x"59",
          7221 => x"62",
          7222 => x"4b",
          7223 => x"5b",
          7224 => x"44",
          7225 => x"34",
          7226 => x"4c",
          7227 => x"28",
          7228 => x"7f",
          7229 => x"49",
          7230 => x"d8",
          7231 => x"6e",
          7232 => x"9d",
          7233 => x"24",
          7234 => x"fb",
          7235 => x"95",
          7236 => x"d8",
          7237 => x"9d",
          7238 => x"49",
          7239 => x"8f",
          7240 => x"d5",
          7241 => x"fa",
          7242 => x"9f",
          7243 => x"5c",
          7244 => x"5c",
          7245 => x"5c",
          7246 => x"5c",
          7247 => x"5c",
          7248 => x"5c",
          7249 => x"5c",
          7250 => x"5c",
          7251 => x"5c",
          7252 => x"5c",
          7253 => x"5c",
          7254 => x"5c",
          7255 => x"5c",
          7256 => x"5c",
          7257 => x"74",
          7258 => x"4f",
          7259 => x"66",
          7260 => x"17",
          7261 => x"5c",
          7262 => x"07",
          7263 => x"b0",
          7264 => x"f5",
          7265 => x"d1",
          7266 => x"5c",
          7267 => x"02",
          7268 => x"43",
          7269 => x"77",
          7270 => x"2c",
          7271 => x"83",
          7272 => x"c5",
          7273 => x"83",
          7274 => x"83",
          7275 => x"83",
          7276 => x"ad",
          7277 => x"83",
          7278 => x"83",
          7279 => x"83",
          7280 => x"83",
          7281 => x"83",
          7282 => x"83",
          7283 => x"83",
          7284 => x"83",
          7285 => x"83",
          7286 => x"83",
          7287 => x"83",
          7288 => x"83",
          7289 => x"d3",
          7290 => x"83",
          7291 => x"83",
          7292 => x"5a",
          7293 => x"3d",
          7294 => x"1b",
          7295 => x"1b",
          7296 => x"1b",
          7297 => x"f6",
          7298 => x"1b",
          7299 => x"1b",
          7300 => x"1b",
          7301 => x"1b",
          7302 => x"1b",
          7303 => x"1b",
          7304 => x"1b",
          7305 => x"1b",
          7306 => x"1b",
          7307 => x"1b",
          7308 => x"1b",
          7309 => x"00",
          7310 => x"da",
          7311 => x"8b",
          7312 => x"68",
          7313 => x"58",
          7314 => x"36",
          7315 => x"12",
          7316 => x"72",
          7317 => x"4a",
          7318 => x"94",
          7319 => x"d1",
          7320 => x"d1",
          7321 => x"d1",
          7322 => x"d1",
          7323 => x"d1",
          7324 => x"d1",
          7325 => x"d1",
          7326 => x"d1",
          7327 => x"d1",
          7328 => x"d1",
          7329 => x"bf",
          7330 => x"d1",
          7331 => x"d1",
          7332 => x"d2",
          7333 => x"2e",
          7334 => x"0f",
          7335 => x"f9",
          7336 => x"e3",
          7337 => x"c9",
          7338 => x"fd",
          7339 => x"49",
          7340 => x"fd",
          7341 => x"fd",
          7342 => x"fd",
          7343 => x"fd",
          7344 => x"7f",
          7345 => x"fd",
          7346 => x"fd",
          7347 => x"fd",
          7348 => x"fd",
          7349 => x"fd",
          7350 => x"fd",
          7351 => x"fd",
          7352 => x"fd",
          7353 => x"fd",
          7354 => x"fd",
          7355 => x"fd",
          7356 => x"fd",
          7357 => x"fd",
          7358 => x"fd",
          7359 => x"fd",
          7360 => x"fd",
          7361 => x"fd",
          7362 => x"fd",
          7363 => x"1d",
          7364 => x"fd",
          7365 => x"fd",
          7366 => x"fd",
          7367 => x"fd",
          7368 => x"fd",
          7369 => x"fd",
          7370 => x"fd",
          7371 => x"2b",
          7372 => x"b8",
          7373 => x"b8",
          7374 => x"e1",
          7375 => x"fd",
          7376 => x"fd",
          7377 => x"16",
          7378 => x"fd",
          7379 => x"58",
          7380 => x"18",
          7381 => x"fd",
          7382 => x"69",
          7383 => x"63",
          7384 => x"69",
          7385 => x"61",
          7386 => x"65",
          7387 => x"65",
          7388 => x"70",
          7389 => x"66",
          7390 => x"6d",
          7391 => x"00",
          7392 => x"00",
          7393 => x"00",
          7394 => x"00",
          7395 => x"00",
          7396 => x"74",
          7397 => x"65",
          7398 => x"6f",
          7399 => x"74",
          7400 => x"00",
          7401 => x"73",
          7402 => x"73",
          7403 => x"6f",
          7404 => x"00",
          7405 => x"20",
          7406 => x"00",
          7407 => x"65",
          7408 => x"72",
          7409 => x"00",
          7410 => x"79",
          7411 => x"69",
          7412 => x"00",
          7413 => x"63",
          7414 => x"6d",
          7415 => x"00",
          7416 => x"20",
          7417 => x"00",
          7418 => x"2c",
          7419 => x"69",
          7420 => x"65",
          7421 => x"00",
          7422 => x"61",
          7423 => x"00",
          7424 => x"61",
          7425 => x"69",
          7426 => x"6d",
          7427 => x"6f",
          7428 => x"00",
          7429 => x"74",
          7430 => x"64",
          7431 => x"76",
          7432 => x"72",
          7433 => x"61",
          7434 => x"00",
          7435 => x"72",
          7436 => x"74",
          7437 => x"00",
          7438 => x"6e",
          7439 => x"61",
          7440 => x"00",
          7441 => x"72",
          7442 => x"69",
          7443 => x"00",
          7444 => x"64",
          7445 => x"00",
          7446 => x"20",
          7447 => x"65",
          7448 => x"70",
          7449 => x"6e",
          7450 => x"66",
          7451 => x"6e",
          7452 => x"6b",
          7453 => x"61",
          7454 => x"65",
          7455 => x"72",
          7456 => x"6b",
          7457 => x"00",
          7458 => x"2e",
          7459 => x"75",
          7460 => x"25",
          7461 => x"75",
          7462 => x"73",
          7463 => x"00",
          7464 => x"00",
          7465 => x"00",
          7466 => x"58",
          7467 => x"00",
          7468 => x"00",
          7469 => x"00",
          7470 => x"20",
          7471 => x"00",
          7472 => x"00",
          7473 => x"30",
          7474 => x"31",
          7475 => x"55",
          7476 => x"30",
          7477 => x"25",
          7478 => x"00",
          7479 => x"65",
          7480 => x"61",
          7481 => x"00",
          7482 => x"58",
          7483 => x"75",
          7484 => x"54",
          7485 => x"74",
          7486 => x"00",
          7487 => x"58",
          7488 => x"75",
          7489 => x"54",
          7490 => x"74",
          7491 => x"00",
          7492 => x"52",
          7493 => x"75",
          7494 => x"54",
          7495 => x"74",
          7496 => x"00",
          7497 => x"65",
          7498 => x"00",
          7499 => x"6e",
          7500 => x"00",
          7501 => x"20",
          7502 => x"72",
          7503 => x"62",
          7504 => x"6d",
          7505 => x"00",
          7506 => x"63",
          7507 => x"00",
          7508 => x"2e",
          7509 => x"6c",
          7510 => x"6e",
          7511 => x"65",
          7512 => x"64",
          7513 => x"61",
          7514 => x"20",
          7515 => x"79",
          7516 => x"00",
          7517 => x"00",
          7518 => x"69",
          7519 => x"64",
          7520 => x"00",
          7521 => x"6d",
          7522 => x"00",
          7523 => x"00",
          7524 => x"25",
          7525 => x"00",
          7526 => x"62",
          7527 => x"2e",
          7528 => x"74",
          7529 => x"61",
          7530 => x"69",
          7531 => x"00",
          7532 => x"20",
          7533 => x"25",
          7534 => x"2e",
          7535 => x"6c",
          7536 => x"65",
          7537 => x"28",
          7538 => x"00",
          7539 => x"6e",
          7540 => x"40",
          7541 => x"2e",
          7542 => x"6c",
          7543 => x"2d",
          7544 => x"6c",
          7545 => x"00",
          7546 => x"6e",
          7547 => x"00",
          7548 => x"30",
          7549 => x"38",
          7550 => x"29",
          7551 => x"79",
          7552 => x"00",
          7553 => x"30",
          7554 => x"61",
          7555 => x"2e",
          7556 => x"70",
          7557 => x"00",
          7558 => x"74",
          7559 => x"5c",
          7560 => x"00",
          7561 => x"65",
          7562 => x"64",
          7563 => x"74",
          7564 => x"73",
          7565 => x"64",
          7566 => x"00",
          7567 => x"64",
          7568 => x"25",
          7569 => x"00",
          7570 => x"66",
          7571 => x"6f",
          7572 => x"65",
          7573 => x"6d",
          7574 => x"65",
          7575 => x"72",
          7576 => x"00",
          7577 => x"20",
          7578 => x"65",
          7579 => x"64",
          7580 => x"25",
          7581 => x"00",
          7582 => x"20",
          7583 => x"53",
          7584 => x"64",
          7585 => x"25",
          7586 => x"00",
          7587 => x"63",
          7588 => x"20",
          7589 => x"20",
          7590 => x"25",
          7591 => x"00",
          7592 => x"00",
          7593 => x"20",
          7594 => x"20",
          7595 => x"20",
          7596 => x"25",
          7597 => x"00",
          7598 => x"74",
          7599 => x"6b",
          7600 => x"20",
          7601 => x"25",
          7602 => x"48",
          7603 => x"20",
          7604 => x"65",
          7605 => x"43",
          7606 => x"65",
          7607 => x"30",
          7608 => x"00",
          7609 => x"41",
          7610 => x"20",
          7611 => x"20",
          7612 => x"25",
          7613 => x"48",
          7614 => x"20",
          7615 => x"20",
          7616 => x"20",
          7617 => x"00",
          7618 => x"49",
          7619 => x"20",
          7620 => x"45",
          7621 => x"00",
          7622 => x"52",
          7623 => x"43",
          7624 => x"3d",
          7625 => x"00",
          7626 => x"45",
          7627 => x"54",
          7628 => x"3d",
          7629 => x"00",
          7630 => x"43",
          7631 => x"44",
          7632 => x"3d",
          7633 => x"00",
          7634 => x"20",
          7635 => x"25",
          7636 => x"58",
          7637 => x"20",
          7638 => x"20",
          7639 => x"3a",
          7640 => x"00",
          7641 => x"4e",
          7642 => x"25",
          7643 => x"58",
          7644 => x"20",
          7645 => x"20",
          7646 => x"3a",
          7647 => x"00",
          7648 => x"53",
          7649 => x"25",
          7650 => x"58",
          7651 => x"72",
          7652 => x"63",
          7653 => x"00",
          7654 => x"00",
          7655 => x"00",
          7656 => x"00",
          7657 => x"00",
          7658 => x"00",
          7659 => x"b4",
          7660 => x"02",
          7661 => x"00",
          7662 => x"ac",
          7663 => x"04",
          7664 => x"00",
          7665 => x"a4",
          7666 => x"06",
          7667 => x"00",
          7668 => x"9c",
          7669 => x"01",
          7670 => x"00",
          7671 => x"94",
          7672 => x"0b",
          7673 => x"00",
          7674 => x"8c",
          7675 => x"0a",
          7676 => x"00",
          7677 => x"84",
          7678 => x"0c",
          7679 => x"00",
          7680 => x"7c",
          7681 => x"0f",
          7682 => x"00",
          7683 => x"74",
          7684 => x"10",
          7685 => x"00",
          7686 => x"6c",
          7687 => x"12",
          7688 => x"00",
          7689 => x"64",
          7690 => x"14",
          7691 => x"00",
          7692 => x"00",
          7693 => x"00",
          7694 => x"7e",
          7695 => x"7e",
          7696 => x"7e",
          7697 => x"7e",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"00",
          7703 => x"6e",
          7704 => x"2f",
          7705 => x"68",
          7706 => x"66",
          7707 => x"73",
          7708 => x"00",
          7709 => x"00",
          7710 => x"00",
          7711 => x"6c",
          7712 => x"00",
          7713 => x"74",
          7714 => x"20",
          7715 => x"74",
          7716 => x"65",
          7717 => x"2e",
          7718 => x"0a",
          7719 => x"7e",
          7720 => x"00",
          7721 => x"00",
          7722 => x"30",
          7723 => x"31",
          7724 => x"32",
          7725 => x"33",
          7726 => x"34",
          7727 => x"35",
          7728 => x"37",
          7729 => x"38",
          7730 => x"39",
          7731 => x"30",
          7732 => x"7e",
          7733 => x"7e",
          7734 => x"00",
          7735 => x"00",
          7736 => x"00",
          7737 => x"2c",
          7738 => x"64",
          7739 => x"78",
          7740 => x"64",
          7741 => x"25",
          7742 => x"2c",
          7743 => x"00",
          7744 => x"00",
          7745 => x"00",
          7746 => x"64",
          7747 => x"6f",
          7748 => x"6f",
          7749 => x"25",
          7750 => x"78",
          7751 => x"25",
          7752 => x"78",
          7753 => x"25",
          7754 => x"00",
          7755 => x"74",
          7756 => x"69",
          7757 => x"20",
          7758 => x"44",
          7759 => x"00",
          7760 => x"74",
          7761 => x"69",
          7762 => x"74",
          7763 => x"69",
          7764 => x"00",
          7765 => x"3c",
          7766 => x"00",
          7767 => x"00",
          7768 => x"33",
          7769 => x"4d",
          7770 => x"00",
          7771 => x"20",
          7772 => x"20",
          7773 => x"4e",
          7774 => x"46",
          7775 => x"00",
          7776 => x"00",
          7777 => x"00",
          7778 => x"12",
          7779 => x"00",
          7780 => x"80",
          7781 => x"8f",
          7782 => x"55",
          7783 => x"9f",
          7784 => x"a7",
          7785 => x"af",
          7786 => x"b7",
          7787 => x"bf",
          7788 => x"c7",
          7789 => x"cf",
          7790 => x"d7",
          7791 => x"df",
          7792 => x"e7",
          7793 => x"ef",
          7794 => x"f7",
          7795 => x"ff",
          7796 => x"2f",
          7797 => x"7c",
          7798 => x"04",
          7799 => x"00",
          7800 => x"02",
          7801 => x"20",
          7802 => x"fc",
          7803 => x"e0",
          7804 => x"eb",
          7805 => x"ec",
          7806 => x"e6",
          7807 => x"f2",
          7808 => x"d6",
          7809 => x"a5",
          7810 => x"ed",
          7811 => x"d1",
          7812 => x"10",
          7813 => x"a1",
          7814 => x"92",
          7815 => x"61",
          7816 => x"63",
          7817 => x"5c",
          7818 => x"34",
          7819 => x"3c",
          7820 => x"54",
          7821 => x"50",
          7822 => x"64",
          7823 => x"52",
          7824 => x"18",
          7825 => x"8c",
          7826 => x"df",
          7827 => x"c3",
          7828 => x"98",
          7829 => x"c6",
          7830 => x"b1",
          7831 => x"21",
          7832 => x"19",
          7833 => x"b2",
          7834 => x"1a",
          7835 => x"07",
          7836 => x"00",
          7837 => x"39",
          7838 => x"79",
          7839 => x"43",
          7840 => x"84",
          7841 => x"87",
          7842 => x"8b",
          7843 => x"90",
          7844 => x"94",
          7845 => x"98",
          7846 => x"9c",
          7847 => x"a0",
          7848 => x"a4",
          7849 => x"a7",
          7850 => x"ac",
          7851 => x"af",
          7852 => x"b3",
          7853 => x"b8",
          7854 => x"bc",
          7855 => x"c0",
          7856 => x"c4",
          7857 => x"c8",
          7858 => x"ca",
          7859 => x"01",
          7860 => x"f3",
          7861 => x"f4",
          7862 => x"12",
          7863 => x"3b",
          7864 => x"3f",
          7865 => x"46",
          7866 => x"81",
          7867 => x"8a",
          7868 => x"90",
          7869 => x"5f",
          7870 => x"94",
          7871 => x"67",
          7872 => x"62",
          7873 => x"9c",
          7874 => x"73",
          7875 => x"77",
          7876 => x"7b",
          7877 => x"7f",
          7878 => x"a9",
          7879 => x"87",
          7880 => x"b2",
          7881 => x"8f",
          7882 => x"7b",
          7883 => x"ff",
          7884 => x"88",
          7885 => x"11",
          7886 => x"a3",
          7887 => x"03",
          7888 => x"d8",
          7889 => x"f9",
          7890 => x"f6",
          7891 => x"fa",
          7892 => x"50",
          7893 => x"8a",
          7894 => x"cf",
          7895 => x"44",
          7896 => x"00",
          7897 => x"00",
          7898 => x"00",
          7899 => x"20",
          7900 => x"40",
          7901 => x"59",
          7902 => x"5d",
          7903 => x"08",
          7904 => x"bb",
          7905 => x"cb",
          7906 => x"f9",
          7907 => x"fb",
          7908 => x"08",
          7909 => x"04",
          7910 => x"bc",
          7911 => x"d0",
          7912 => x"e5",
          7913 => x"01",
          7914 => x"32",
          7915 => x"01",
          7916 => x"30",
          7917 => x"67",
          7918 => x"80",
          7919 => x"41",
          7920 => x"00",
          7921 => x"00",
          7922 => x"00",
          7923 => x"00",
          7924 => x"00",
          7925 => x"00",
          7926 => x"00",
          7927 => x"00",
          7928 => x"00",
          7929 => x"00",
          7930 => x"00",
          7931 => x"00",
          7932 => x"00",
          7933 => x"00",
          7934 => x"00",
          7935 => x"00",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"00",
          7940 => x"00",
          7941 => x"00",
          7942 => x"00",
          7943 => x"00",
          7944 => x"00",
          7945 => x"00",
          7946 => x"00",
          7947 => x"00",
          7948 => x"00",
          7949 => x"00",
          7950 => x"00",
          7951 => x"00",
          7952 => x"00",
          7953 => x"00",
          7954 => x"00",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"00",
          7959 => x"00",
          7960 => x"00",
          7961 => x"00",
          7962 => x"00",
          7963 => x"00",
          7964 => x"00",
          7965 => x"00",
          7966 => x"00",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"00",
          7983 => x"00",
          7984 => x"00",
          7985 => x"00",
          7986 => x"01",
          7987 => x"01",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"00",
          7996 => x"00",
          7997 => x"00",
          7998 => x"00",
          7999 => x"00",
          8000 => x"e4",
          8001 => x"ec",
          8002 => x"f4",
          8003 => x"80",
          8004 => x"0d",
          8005 => x"f0",
          8006 => x"78",
          8007 => x"70",
          8008 => x"68",
          8009 => x"38",
          8010 => x"2e",
          8011 => x"2f",
          8012 => x"f0",
          8013 => x"f0",
          8014 => x"0d",
          8015 => x"f0",
          8016 => x"58",
          8017 => x"50",
          8018 => x"48",
          8019 => x"38",
          8020 => x"2e",
          8021 => x"2f",
          8022 => x"f0",
          8023 => x"f0",
          8024 => x"0d",
          8025 => x"f0",
          8026 => x"58",
          8027 => x"50",
          8028 => x"48",
          8029 => x"28",
          8030 => x"3e",
          8031 => x"2f",
          8032 => x"f0",
          8033 => x"f0",
          8034 => x"f0",
          8035 => x"f0",
          8036 => x"18",
          8037 => x"10",
          8038 => x"08",
          8039 => x"f0",
          8040 => x"f0",
          8041 => x"1c",
          8042 => x"f0",
          8043 => x"f0",
          8044 => x"cd",
          8045 => x"f0",
          8046 => x"dd",
          8047 => x"b1",
          8048 => x"73",
          8049 => x"a2",
          8050 => x"b9",
          8051 => x"be",
          8052 => x"f0",
          8053 => x"f0",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"01",
          9089 => x"f3",
          9090 => x"fb",
          9091 => x"c3",
          9092 => x"e6",
          9093 => x"63",
          9094 => x"6a",
          9095 => x"23",
          9096 => x"2c",
          9097 => x"03",
          9098 => x"0b",
          9099 => x"13",
          9100 => x"52",
          9101 => x"83",
          9102 => x"8b",
          9103 => x"93",
          9104 => x"bc",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"00",
          9113 => x"00",
          9114 => x"00",
          9115 => x"00",
          9116 => x"00",
          9117 => x"00",
          9118 => x"00",
          9119 => x"00",
          9120 => x"03",
          9121 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"87",
             1 => x"e9",
             2 => x"00",
             3 => x"00",
             4 => x"8c",
             5 => x"90",
             6 => x"00",
             7 => x"00",
             8 => x"06",
             9 => x"82",
            10 => x"06",
            11 => x"00",
            12 => x"06",
            13 => x"09",
            14 => x"09",
            15 => x"0b",
            16 => x"81",
            17 => x"09",
            18 => x"81",
            19 => x"00",
            20 => x"24",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"05",
            26 => x"0a",
            27 => x"53",
            28 => x"26",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"9f",
            45 => x"93",
            46 => x"00",
            47 => x"00",
            48 => x"2a",
            49 => x"09",
            50 => x"53",
            51 => x"00",
            52 => x"53",
            53 => x"81",
            54 => x"07",
            55 => x"00",
            56 => x"81",
            57 => x"09",
            58 => x"00",
            59 => x"00",
            60 => x"81",
            61 => x"09",
            62 => x"04",
            63 => x"00",
            64 => x"81",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"09",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"72",
            73 => x"51",
            74 => x"00",
            75 => x"00",
            76 => x"06",
            77 => x"83",
            78 => x"06",
            79 => x"00",
            80 => x"06",
            81 => x"83",
            82 => x"0b",
            83 => x"00",
            84 => x"8c",
            85 => x"0b",
            86 => x"56",
            87 => x"04",
            88 => x"8c",
            89 => x"0b",
            90 => x"56",
            91 => x"04",
            92 => x"70",
            93 => x"ff",
            94 => x"72",
            95 => x"51",
            96 => x"70",
            97 => x"06",
            98 => x"09",
            99 => x"51",
           100 => x"05",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"05",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"05",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"05",
           125 => x"04",
           126 => x"ff",
           127 => x"ff",
           128 => x"06",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"85",
           134 => x"0b",
           135 => x"0b",
           136 => x"c6",
           137 => x"0b",
           138 => x"0b",
           139 => x"86",
           140 => x"0b",
           141 => x"0b",
           142 => x"c6",
           143 => x"0b",
           144 => x"0b",
           145 => x"8a",
           146 => x"0b",
           147 => x"0b",
           148 => x"ce",
           149 => x"0b",
           150 => x"0b",
           151 => x"92",
           152 => x"0b",
           153 => x"0b",
           154 => x"d6",
           155 => x"0b",
           156 => x"0b",
           157 => x"9a",
           158 => x"0b",
           159 => x"0b",
           160 => x"de",
           161 => x"0b",
           162 => x"0b",
           163 => x"a2",
           164 => x"0b",
           165 => x"0b",
           166 => x"e6",
           167 => x"0b",
           168 => x"0b",
           169 => x"aa",
           170 => x"0b",
           171 => x"0b",
           172 => x"ed",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"8c",
           193 => x"d5",
           194 => x"c0",
           195 => x"a2",
           196 => x"c0",
           197 => x"a0",
           198 => x"c0",
           199 => x"a0",
           200 => x"c0",
           201 => x"94",
           202 => x"c0",
           203 => x"a1",
           204 => x"c0",
           205 => x"af",
           206 => x"c0",
           207 => x"ad",
           208 => x"c0",
           209 => x"94",
           210 => x"c0",
           211 => x"95",
           212 => x"c0",
           213 => x"95",
           214 => x"c0",
           215 => x"b1",
           216 => x"c0",
           217 => x"80",
           218 => x"80",
           219 => x"0c",
           220 => x"08",
           221 => x"98",
           222 => x"98",
           223 => x"ba",
           224 => x"ba",
           225 => x"84",
           226 => x"84",
           227 => x"04",
           228 => x"2d",
           229 => x"90",
           230 => x"e7",
           231 => x"80",
           232 => x"d8",
           233 => x"c0",
           234 => x"82",
           235 => x"80",
           236 => x"0c",
           237 => x"08",
           238 => x"98",
           239 => x"98",
           240 => x"ba",
           241 => x"ba",
           242 => x"84",
           243 => x"84",
           244 => x"04",
           245 => x"2d",
           246 => x"90",
           247 => x"eb",
           248 => x"80",
           249 => x"ff",
           250 => x"c0",
           251 => x"83",
           252 => x"80",
           253 => x"0c",
           254 => x"08",
           255 => x"98",
           256 => x"98",
           257 => x"ba",
           258 => x"ba",
           259 => x"84",
           260 => x"84",
           261 => x"04",
           262 => x"2d",
           263 => x"90",
           264 => x"d7",
           265 => x"80",
           266 => x"f6",
           267 => x"c0",
           268 => x"83",
           269 => x"80",
           270 => x"0c",
           271 => x"08",
           272 => x"98",
           273 => x"98",
           274 => x"ba",
           275 => x"ba",
           276 => x"84",
           277 => x"84",
           278 => x"04",
           279 => x"2d",
           280 => x"90",
           281 => x"8e",
           282 => x"80",
           283 => x"f4",
           284 => x"c0",
           285 => x"81",
           286 => x"80",
           287 => x"0c",
           288 => x"08",
           289 => x"98",
           290 => x"98",
           291 => x"ba",
           292 => x"ba",
           293 => x"84",
           294 => x"84",
           295 => x"04",
           296 => x"84",
           297 => x"04",
           298 => x"2d",
           299 => x"90",
           300 => x"85",
           301 => x"80",
           302 => x"f2",
           303 => x"c0",
           304 => x"81",
           305 => x"80",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"04",
           311 => x"83",
           312 => x"10",
           313 => x"51",
           314 => x"06",
           315 => x"10",
           316 => x"ed",
           317 => x"ba",
           318 => x"38",
           319 => x"0b",
           320 => x"51",
           321 => x"0d",
           322 => x"08",
           323 => x"08",
           324 => x"04",
           325 => x"11",
           326 => x"25",
           327 => x"72",
           328 => x"38",
           329 => x"30",
           330 => x"55",
           331 => x"71",
           332 => x"fa",
           333 => x"ba",
           334 => x"ba",
           335 => x"34",
           336 => x"70",
           337 => x"54",
           338 => x"34",
           339 => x"88",
           340 => x"8c",
           341 => x"0d",
           342 => x"05",
           343 => x"3d",
           344 => x"e4",
           345 => x"80",
           346 => x"3d",
           347 => x"52",
           348 => x"04",
           349 => x"5d",
           350 => x"1e",
           351 => x"06",
           352 => x"2e",
           353 => x"33",
           354 => x"81",
           355 => x"80",
           356 => x"7e",
           357 => x"32",
           358 => x"55",
           359 => x"38",
           360 => x"06",
           361 => x"7a",
           362 => x"76",
           363 => x"73",
           364 => x"04",
           365 => x"10",
           366 => x"98",
           367 => x"8b",
           368 => x"5b",
           369 => x"38",
           370 => x"38",
           371 => x"f7",
           372 => x"09",
           373 => x"5a",
           374 => x"76",
           375 => x"52",
           376 => x"57",
           377 => x"7a",
           378 => x"78",
           379 => x"54",
           380 => x"80",
           381 => x"83",
           382 => x"73",
           383 => x"27",
           384 => x"eb",
           385 => x"fe",
           386 => x"59",
           387 => x"84",
           388 => x"06",
           389 => x"5e",
           390 => x"84",
           391 => x"ba",
           392 => x"72",
           393 => x"08",
           394 => x"05",
           395 => x"ca",
           396 => x"ba",
           397 => x"9c",
           398 => x"56",
           399 => x"80",
           400 => x"90",
           401 => x"81",
           402 => x"38",
           403 => x"80",
           404 => x"77",
           405 => x"05",
           406 => x"2a",
           407 => x"2e",
           408 => x"ff",
           409 => x"cc",
           410 => x"83",
           411 => x"74",
           412 => x"f0",
           413 => x"90",
           414 => x"53",
           415 => x"81",
           416 => x"38",
           417 => x"86",
           418 => x"54",
           419 => x"54",
           420 => x"81",
           421 => x"77",
           422 => x"80",
           423 => x"80",
           424 => x"51",
           425 => x"80",
           426 => x"2c",
           427 => x"38",
           428 => x"b2",
           429 => x"81",
           430 => x"55",
           431 => x"52",
           432 => x"81",
           433 => x"70",
           434 => x"24",
           435 => x"06",
           436 => x"38",
           437 => x"76",
           438 => x"80",
           439 => x"ba",
           440 => x"1e",
           441 => x"7d",
           442 => x"ec",
           443 => x"2e",
           444 => x"80",
           445 => x"2c",
           446 => x"91",
           447 => x"3f",
           448 => x"a0",
           449 => x"87",
           450 => x"07",
           451 => x"84",
           452 => x"06",
           453 => x"39",
           454 => x"0a",
           455 => x"72",
           456 => x"80",
           457 => x"5a",
           458 => x"70",
           459 => x"38",
           460 => x"80",
           461 => x"5f",
           462 => x"52",
           463 => x"ff",
           464 => x"57",
           465 => x"38",
           466 => x"33",
           467 => x"1a",
           468 => x"79",
           469 => x"7c",
           470 => x"51",
           471 => x"0a",
           472 => x"80",
           473 => x"90",
           474 => x"87",
           475 => x"7a",
           476 => x"60",
           477 => x"41",
           478 => x"7a",
           479 => x"9c",
           480 => x"7c",
           481 => x"f8",
           482 => x"7c",
           483 => x"f8",
           484 => x"08",
           485 => x"72",
           486 => x"3f",
           487 => x"06",
           488 => x"72",
           489 => x"80",
           490 => x"f7",
           491 => x"84",
           492 => x"58",
           493 => x"51",
           494 => x"83",
           495 => x"2b",
           496 => x"07",
           497 => x"38",
           498 => x"80",
           499 => x"2c",
           500 => x"d6",
           501 => x"3f",
           502 => x"bb",
           503 => x"fa",
           504 => x"ab",
           505 => x"7e",
           506 => x"39",
           507 => x"2b",
           508 => x"57",
           509 => x"ff",
           510 => x"fb",
           511 => x"2e",
           512 => x"52",
           513 => x"74",
           514 => x"f1",
           515 => x"98",
           516 => x"b7",
           517 => x"3f",
           518 => x"bb",
           519 => x"51",
           520 => x"83",
           521 => x"2b",
           522 => x"07",
           523 => x"52",
           524 => x"0d",
           525 => x"74",
           526 => x"04",
           527 => x"84",
           528 => x"81",
           529 => x"56",
           530 => x"2e",
           531 => x"70",
           532 => x"2e",
           533 => x"72",
           534 => x"84",
           535 => x"ff",
           536 => x"53",
           537 => x"f0",
           538 => x"08",
           539 => x"51",
           540 => x"ba",
           541 => x"57",
           542 => x"88",
           543 => x"7a",
           544 => x"70",
           545 => x"51",
           546 => x"2e",
           547 => x"81",
           548 => x"09",
           549 => x"84",
           550 => x"73",
           551 => x"80",
           552 => x"90",
           553 => x"8c",
           554 => x"70",
           555 => x"e3",
           556 => x"d5",
           557 => x"83",
           558 => x"7a",
           559 => x"32",
           560 => x"56",
           561 => x"06",
           562 => x"15",
           563 => x"91",
           564 => x"74",
           565 => x"08",
           566 => x"56",
           567 => x"0d",
           568 => x"51",
           569 => x"56",
           570 => x"15",
           571 => x"56",
           572 => x"11",
           573 => x"32",
           574 => x"54",
           575 => x"06",
           576 => x"81",
           577 => x"38",
           578 => x"80",
           579 => x"0c",
           580 => x"0c",
           581 => x"ba",
           582 => x"ff",
           583 => x"8c",
           584 => x"84",
           585 => x"3d",
           586 => x"55",
           587 => x"84",
           588 => x"38",
           589 => x"52",
           590 => x"38",
           591 => x"34",
           592 => x"87",
           593 => x"72",
           594 => x"fd",
           595 => x"54",
           596 => x"70",
           597 => x"81",
           598 => x"81",
           599 => x"84",
           600 => x"fc",
           601 => x"55",
           602 => x"73",
           603 => x"93",
           604 => x"73",
           605 => x"51",
           606 => x"0c",
           607 => x"73",
           608 => x"53",
           609 => x"71",
           610 => x"80",
           611 => x"53",
           612 => x"51",
           613 => x"0d",
           614 => x"05",
           615 => x"12",
           616 => x"51",
           617 => x"75",
           618 => x"81",
           619 => x"81",
           620 => x"84",
           621 => x"fd",
           622 => x"55",
           623 => x"71",
           624 => x"81",
           625 => x"ef",
           626 => x"3d",
           627 => x"7a",
           628 => x"38",
           629 => x"33",
           630 => x"06",
           631 => x"2e",
           632 => x"38",
           633 => x"86",
           634 => x"38",
           635 => x"2e",
           636 => x"51",
           637 => x"31",
           638 => x"04",
           639 => x"0d",
           640 => x"70",
           641 => x"8c",
           642 => x"52",
           643 => x"8c",
           644 => x"2e",
           645 => x"54",
           646 => x"84",
           647 => x"84",
           648 => x"8c",
           649 => x"0d",
           650 => x"54",
           651 => x"81",
           652 => x"8c",
           653 => x"09",
           654 => x"75",
           655 => x"0c",
           656 => x"75",
           657 => x"70",
           658 => x"81",
           659 => x"f4",
           660 => x"3d",
           661 => x"58",
           662 => x"38",
           663 => x"8c",
           664 => x"2e",
           665 => x"71",
           666 => x"52",
           667 => x"52",
           668 => x"13",
           669 => x"71",
           670 => x"74",
           671 => x"9f",
           672 => x"72",
           673 => x"06",
           674 => x"1c",
           675 => x"53",
           676 => x"52",
           677 => x"0d",
           678 => x"80",
           679 => x"80",
           680 => x"75",
           681 => x"70",
           682 => x"71",
           683 => x"06",
           684 => x"84",
           685 => x"75",
           686 => x"70",
           687 => x"71",
           688 => x"81",
           689 => x"75",
           690 => x"52",
           691 => x"55",
           692 => x"51",
           693 => x"04",
           694 => x"71",
           695 => x"ba",
           696 => x"84",
           697 => x"04",
           698 => x"a0",
           699 => x"51",
           700 => x"53",
           701 => x"38",
           702 => x"ba",
           703 => x"9f",
           704 => x"9f",
           705 => x"2a",
           706 => x"54",
           707 => x"a8",
           708 => x"74",
           709 => x"11",
           710 => x"06",
           711 => x"52",
           712 => x"38",
           713 => x"0d",
           714 => x"7a",
           715 => x"7c",
           716 => x"71",
           717 => x"59",
           718 => x"84",
           719 => x"84",
           720 => x"f7",
           721 => x"70",
           722 => x"56",
           723 => x"8f",
           724 => x"33",
           725 => x"73",
           726 => x"2e",
           727 => x"56",
           728 => x"58",
           729 => x"38",
           730 => x"14",
           731 => x"14",
           732 => x"73",
           733 => x"ff",
           734 => x"89",
           735 => x"77",
           736 => x"0c",
           737 => x"26",
           738 => x"38",
           739 => x"56",
           740 => x"0d",
           741 => x"70",
           742 => x"09",
           743 => x"70",
           744 => x"80",
           745 => x"80",
           746 => x"74",
           747 => x"56",
           748 => x"38",
           749 => x"0d",
           750 => x"0c",
           751 => x"ca",
           752 => x"8b",
           753 => x"7d",
           754 => x"08",
           755 => x"2e",
           756 => x"70",
           757 => x"a0",
           758 => x"f5",
           759 => x"d0",
           760 => x"80",
           761 => x"74",
           762 => x"27",
           763 => x"06",
           764 => x"06",
           765 => x"f9",
           766 => x"89",
           767 => x"27",
           768 => x"81",
           769 => x"56",
           770 => x"78",
           771 => x"75",
           772 => x"8c",
           773 => x"16",
           774 => x"59",
           775 => x"ff",
           776 => x"33",
           777 => x"38",
           778 => x"38",
           779 => x"d0",
           780 => x"73",
           781 => x"8c",
           782 => x"81",
           783 => x"55",
           784 => x"84",
           785 => x"80",
           786 => x"81",
           787 => x"ff",
           788 => x"8c",
           789 => x"05",
           790 => x"51",
           791 => x"83",
           792 => x"3d",
           793 => x"a8",
           794 => x"a4",
           795 => x"04",
           796 => x"83",
           797 => x"ef",
           798 => x"cf",
           799 => x"0d",
           800 => x"3f",
           801 => x"51",
           802 => x"83",
           803 => x"3d",
           804 => x"d0",
           805 => x"ec",
           806 => x"04",
           807 => x"83",
           808 => x"ee",
           809 => x"d1",
           810 => x"0d",
           811 => x"3f",
           812 => x"51",
           813 => x"83",
           814 => x"3d",
           815 => x"f8",
           816 => x"80",
           817 => x"04",
           818 => x"83",
           819 => x"02",
           820 => x"58",
           821 => x"73",
           822 => x"75",
           823 => x"74",
           824 => x"55",
           825 => x"53",
           826 => x"82",
           827 => x"57",
           828 => x"d0",
           829 => x"76",
           830 => x"30",
           831 => x"57",
           832 => x"c0",
           833 => x"26",
           834 => x"e8",
           835 => x"8c",
           836 => x"52",
           837 => x"76",
           838 => x"04",
           839 => x"88",
           840 => x"3d",
           841 => x"52",
           842 => x"ba",
           843 => x"ff",
           844 => x"ff",
           845 => x"59",
           846 => x"f4",
           847 => x"78",
           848 => x"08",
           849 => x"83",
           850 => x"97",
           851 => x"05",
           852 => x"80",
           853 => x"3f",
           854 => x"80",
           855 => x"38",
           856 => x"0d",
           857 => x"61",
           858 => x"7f",
           859 => x"8c",
           860 => x"0d",
           861 => x"02",
           862 => x"73",
           863 => x"5d",
           864 => x"7a",
           865 => x"3f",
           866 => x"80",
           867 => x"90",
           868 => x"82",
           869 => x"27",
           870 => x"d2",
           871 => x"84",
           872 => x"ec",
           873 => x"83",
           874 => x"56",
           875 => x"18",
           876 => x"7a",
           877 => x"9f",
           878 => x"73",
           879 => x"74",
           880 => x"27",
           881 => x"52",
           882 => x"56",
           883 => x"dc",
           884 => x"1c",
           885 => x"84",
           886 => x"2c",
           887 => x"38",
           888 => x"1e",
           889 => x"ff",
           890 => x"0d",
           891 => x"3f",
           892 => x"54",
           893 => x"26",
           894 => x"d2",
           895 => x"84",
           896 => x"ea",
           897 => x"38",
           898 => x"38",
           899 => x"db",
           900 => x"08",
           901 => x"78",
           902 => x"83",
           903 => x"14",
           904 => x"51",
           905 => x"ff",
           906 => x"df",
           907 => x"51",
           908 => x"f0",
           909 => x"3f",
           910 => x"39",
           911 => x"e9",
           912 => x"39",
           913 => x"08",
           914 => x"a8",
           915 => x"80",
           916 => x"38",
           917 => x"9b",
           918 => x"2b",
           919 => x"30",
           920 => x"07",
           921 => x"59",
           922 => x"e8",
           923 => x"ba",
           924 => x"70",
           925 => x"70",
           926 => x"06",
           927 => x"80",
           928 => x"39",
           929 => x"3d",
           930 => x"96",
           931 => x"51",
           932 => x"9d",
           933 => x"72",
           934 => x"71",
           935 => x"81",
           936 => x"72",
           937 => x"71",
           938 => x"81",
           939 => x"72",
           940 => x"71",
           941 => x"81",
           942 => x"72",
           943 => x"71",
           944 => x"53",
           945 => x"3d",
           946 => x"83",
           947 => x"51",
           948 => x"3d",
           949 => x"83",
           950 => x"51",
           951 => x"06",
           952 => x"39",
           953 => x"f4",
           954 => x"c1",
           955 => x"51",
           956 => x"c2",
           957 => x"d4",
           958 => x"9b",
           959 => x"06",
           960 => x"38",
           961 => x"3f",
           962 => x"80",
           963 => x"70",
           964 => x"fe",
           965 => x"9a",
           966 => x"f9",
           967 => x"84",
           968 => x"80",
           969 => x"81",
           970 => x"51",
           971 => x"3f",
           972 => x"52",
           973 => x"bd",
           974 => x"d4",
           975 => x"9a",
           976 => x"06",
           977 => x"38",
           978 => x"70",
           979 => x"0c",
           980 => x"d5",
           981 => x"06",
           982 => x"84",
           983 => x"b8",
           984 => x"51",
           985 => x"53",
           986 => x"0b",
           987 => x"ff",
           988 => x"f1",
           989 => x"78",
           990 => x"83",
           991 => x"80",
           992 => x"7b",
           993 => x"81",
           994 => x"2e",
           995 => x"be",
           996 => x"05",
           997 => x"84",
           998 => x"54",
           999 => x"da",
          1000 => x"84",
          1001 => x"80",
          1002 => x"5d",
          1003 => x"3d",
          1004 => x"38",
          1005 => x"3f",
          1006 => x"8c",
          1007 => x"ba",
          1008 => x"05",
          1009 => x"08",
          1010 => x"2e",
          1011 => x"51",
          1012 => x"8f",
          1013 => x"3d",
          1014 => x"38",
          1015 => x"81",
          1016 => x"53",
          1017 => x"dd",
          1018 => x"bc",
          1019 => x"90",
          1020 => x"7c",
          1021 => x"08",
          1022 => x"70",
          1023 => x"42",
          1024 => x"81",
          1025 => x"2e",
          1026 => x"06",
          1027 => x"81",
          1028 => x"81",
          1029 => x"38",
          1030 => x"d5",
          1031 => x"80",
          1032 => x"bc",
          1033 => x"70",
          1034 => x"91",
          1035 => x"84",
          1036 => x"84",
          1037 => x"0b",
          1038 => x"d1",
          1039 => x"82",
          1040 => x"80",
          1041 => x"51",
          1042 => x"80",
          1043 => x"7d",
          1044 => x"38",
          1045 => x"a2",
          1046 => x"ef",
          1047 => x"f8",
          1048 => x"70",
          1049 => x"39",
          1050 => x"59",
          1051 => x"78",
          1052 => x"79",
          1053 => x"88",
          1054 => x"d6",
          1055 => x"60",
          1056 => x"82",
          1057 => x"61",
          1058 => x"81",
          1059 => x"a4",
          1060 => x"3f",
          1061 => x"86",
          1062 => x"83",
          1063 => x"9c",
          1064 => x"89",
          1065 => x"39",
          1066 => x"52",
          1067 => x"39",
          1068 => x"83",
          1069 => x"59",
          1070 => x"80",
          1071 => x"b8",
          1072 => x"05",
          1073 => x"08",
          1074 => x"83",
          1075 => x"5a",
          1076 => x"2e",
          1077 => x"52",
          1078 => x"fa",
          1079 => x"53",
          1080 => x"84",
          1081 => x"38",
          1082 => x"b5",
          1083 => x"fe",
          1084 => x"e9",
          1085 => x"2e",
          1086 => x"11",
          1087 => x"3f",
          1088 => x"64",
          1089 => x"d7",
          1090 => x"ec",
          1091 => x"d0",
          1092 => x"78",
          1093 => x"26",
          1094 => x"46",
          1095 => x"11",
          1096 => x"3f",
          1097 => x"f4",
          1098 => x"ff",
          1099 => x"ba",
          1100 => x"78",
          1101 => x"51",
          1102 => x"53",
          1103 => x"3f",
          1104 => x"2e",
          1105 => x"ca",
          1106 => x"cf",
          1107 => x"ff",
          1108 => x"ba",
          1109 => x"b8",
          1110 => x"05",
          1111 => x"08",
          1112 => x"fe",
          1113 => x"e9",
          1114 => x"2e",
          1115 => x"ce",
          1116 => x"7c",
          1117 => x"7a",
          1118 => x"95",
          1119 => x"53",
          1120 => x"85",
          1121 => x"81",
          1122 => x"ff",
          1123 => x"e8",
          1124 => x"2e",
          1125 => x"11",
          1126 => x"3f",
          1127 => x"84",
          1128 => x"ff",
          1129 => x"ba",
          1130 => x"83",
          1131 => x"5a",
          1132 => x"5c",
          1133 => x"34",
          1134 => x"3d",
          1135 => x"51",
          1136 => x"80",
          1137 => x"fc",
          1138 => x"f3",
          1139 => x"68",
          1140 => x"51",
          1141 => x"53",
          1142 => x"3f",
          1143 => x"2e",
          1144 => x"97",
          1145 => x"68",
          1146 => x"34",
          1147 => x"fc",
          1148 => x"a3",
          1149 => x"f5",
          1150 => x"05",
          1151 => x"b8",
          1152 => x"05",
          1153 => x"08",
          1154 => x"3d",
          1155 => x"51",
          1156 => x"80",
          1157 => x"fc",
          1158 => x"d3",
          1159 => x"f5",
          1160 => x"53",
          1161 => x"84",
          1162 => x"8c",
          1163 => x"ad",
          1164 => x"27",
          1165 => x"84",
          1166 => x"38",
          1167 => x"39",
          1168 => x"96",
          1169 => x"ff",
          1170 => x"81",
          1171 => x"51",
          1172 => x"80",
          1173 => x"08",
          1174 => x"b8",
          1175 => x"05",
          1176 => x"08",
          1177 => x"79",
          1178 => x"c8",
          1179 => x"53",
          1180 => x"84",
          1181 => x"90",
          1182 => x"38",
          1183 => x"fe",
          1184 => x"e5",
          1185 => x"2e",
          1186 => x"88",
          1187 => x"32",
          1188 => x"7e",
          1189 => x"88",
          1190 => x"46",
          1191 => x"80",
          1192 => x"68",
          1193 => x"51",
          1194 => x"64",
          1195 => x"b8",
          1196 => x"05",
          1197 => x"08",
          1198 => x"71",
          1199 => x"3d",
          1200 => x"51",
          1201 => x"c6",
          1202 => x"80",
          1203 => x"40",
          1204 => x"11",
          1205 => x"3f",
          1206 => x"8c",
          1207 => x"22",
          1208 => x"45",
          1209 => x"80",
          1210 => x"8c",
          1211 => x"b8",
          1212 => x"05",
          1213 => x"08",
          1214 => x"02",
          1215 => x"81",
          1216 => x"fe",
          1217 => x"e0",
          1218 => x"2e",
          1219 => x"5d",
          1220 => x"e1",
          1221 => x"f3",
          1222 => x"54",
          1223 => x"51",
          1224 => x"52",
          1225 => x"39",
          1226 => x"f0",
          1227 => x"53",
          1228 => x"84",
          1229 => x"64",
          1230 => x"70",
          1231 => x"e7",
          1232 => x"80",
          1233 => x"08",
          1234 => x"33",
          1235 => x"f2",
          1236 => x"d8",
          1237 => x"f7",
          1238 => x"c0",
          1239 => x"f3",
          1240 => x"38",
          1241 => x"39",
          1242 => x"f9",
          1243 => x"78",
          1244 => x"08",
          1245 => x"33",
          1246 => x"f2",
          1247 => x"f3",
          1248 => x"38",
          1249 => x"39",
          1250 => x"2e",
          1251 => x"fb",
          1252 => x"7c",
          1253 => x"08",
          1254 => x"08",
          1255 => x"83",
          1256 => x"b5",
          1257 => x"ba",
          1258 => x"08",
          1259 => x"51",
          1260 => x"90",
          1261 => x"80",
          1262 => x"84",
          1263 => x"c0",
          1264 => x"84",
          1265 => x"84",
          1266 => x"57",
          1267 => x"da",
          1268 => x"07",
          1269 => x"c0",
          1270 => x"87",
          1271 => x"5c",
          1272 => x"05",
          1273 => x"ec",
          1274 => x"70",
          1275 => x"b6",
          1276 => x"3f",
          1277 => x"d2",
          1278 => x"95",
          1279 => x"55",
          1280 => x"83",
          1281 => x"83",
          1282 => x"97",
          1283 => x"3d",
          1284 => x"75",
          1285 => x"38",
          1286 => x"52",
          1287 => x"38",
          1288 => x"06",
          1289 => x"38",
          1290 => x"2e",
          1291 => x"2e",
          1292 => x"81",
          1293 => x"2e",
          1294 => x"8b",
          1295 => x"12",
          1296 => x"06",
          1297 => x"06",
          1298 => x"70",
          1299 => x"52",
          1300 => x"72",
          1301 => x"0c",
          1302 => x"87",
          1303 => x"38",
          1304 => x"12",
          1305 => x"06",
          1306 => x"38",
          1307 => x"81",
          1308 => x"81",
          1309 => x"3d",
          1310 => x"80",
          1311 => x"0d",
          1312 => x"51",
          1313 => x"80",
          1314 => x"0c",
          1315 => x"76",
          1316 => x"81",
          1317 => x"83",
          1318 => x"73",
          1319 => x"33",
          1320 => x"fe",
          1321 => x"73",
          1322 => x"33",
          1323 => x"e6",
          1324 => x"74",
          1325 => x"13",
          1326 => x"26",
          1327 => x"98",
          1328 => x"bc",
          1329 => x"b8",
          1330 => x"b4",
          1331 => x"b0",
          1332 => x"ac",
          1333 => x"a8",
          1334 => x"73",
          1335 => x"87",
          1336 => x"84",
          1337 => x"f3",
          1338 => x"9c",
          1339 => x"bc",
          1340 => x"98",
          1341 => x"87",
          1342 => x"1c",
          1343 => x"7b",
          1344 => x"08",
          1345 => x"98",
          1346 => x"87",
          1347 => x"1c",
          1348 => x"79",
          1349 => x"83",
          1350 => x"ff",
          1351 => x"1b",
          1352 => x"1b",
          1353 => x"83",
          1354 => x"51",
          1355 => x"04",
          1356 => x"53",
          1357 => x"80",
          1358 => x"98",
          1359 => x"ff",
          1360 => x"83",
          1361 => x"0c",
          1362 => x"e8",
          1363 => x"2b",
          1364 => x"2e",
          1365 => x"80",
          1366 => x"98",
          1367 => x"ff",
          1368 => x"0d",
          1369 => x"54",
          1370 => x"ba",
          1371 => x"51",
          1372 => x"72",
          1373 => x"25",
          1374 => x"85",
          1375 => x"9b",
          1376 => x"81",
          1377 => x"2e",
          1378 => x"08",
          1379 => x"54",
          1380 => x"91",
          1381 => x"e3",
          1382 => x"72",
          1383 => x"81",
          1384 => x"ff",
          1385 => x"70",
          1386 => x"90",
          1387 => x"8c",
          1388 => x"2a",
          1389 => x"38",
          1390 => x"80",
          1391 => x"06",
          1392 => x"c0",
          1393 => x"81",
          1394 => x"d8",
          1395 => x"33",
          1396 => x"52",
          1397 => x"0d",
          1398 => x"75",
          1399 => x"2e",
          1400 => x"c4",
          1401 => x"55",
          1402 => x"c0",
          1403 => x"81",
          1404 => x"8c",
          1405 => x"51",
          1406 => x"81",
          1407 => x"71",
          1408 => x"38",
          1409 => x"94",
          1410 => x"87",
          1411 => x"81",
          1412 => x"9b",
          1413 => x"3d",
          1414 => x"06",
          1415 => x"32",
          1416 => x"38",
          1417 => x"80",
          1418 => x"84",
          1419 => x"53",
          1420 => x"ff",
          1421 => x"70",
          1422 => x"80",
          1423 => x"a4",
          1424 => x"9e",
          1425 => x"c0",
          1426 => x"87",
          1427 => x"0c",
          1428 => x"d8",
          1429 => x"f2",
          1430 => x"83",
          1431 => x"08",
          1432 => x"b4",
          1433 => x"9e",
          1434 => x"c0",
          1435 => x"87",
          1436 => x"0c",
          1437 => x"f8",
          1438 => x"71",
          1439 => x"84",
          1440 => x"9e",
          1441 => x"c0",
          1442 => x"81",
          1443 => x"87",
          1444 => x"0a",
          1445 => x"38",
          1446 => x"87",
          1447 => x"0a",
          1448 => x"83",
          1449 => x"34",
          1450 => x"70",
          1451 => x"70",
          1452 => x"83",
          1453 => x"9e",
          1454 => x"51",
          1455 => x"81",
          1456 => x"0b",
          1457 => x"80",
          1458 => x"2e",
          1459 => x"91",
          1460 => x"08",
          1461 => x"52",
          1462 => x"71",
          1463 => x"c0",
          1464 => x"06",
          1465 => x"38",
          1466 => x"80",
          1467 => x"82",
          1468 => x"80",
          1469 => x"f3",
          1470 => x"90",
          1471 => x"52",
          1472 => x"52",
          1473 => x"87",
          1474 => x"80",
          1475 => x"83",
          1476 => x"34",
          1477 => x"70",
          1478 => x"80",
          1479 => x"f3",
          1480 => x"98",
          1481 => x"71",
          1482 => x"c0",
          1483 => x"51",
          1484 => x"81",
          1485 => x"c0",
          1486 => x"84",
          1487 => x"34",
          1488 => x"70",
          1489 => x"2e",
          1490 => x"9b",
          1491 => x"06",
          1492 => x"3d",
          1493 => x"fb",
          1494 => x"b6",
          1495 => x"73",
          1496 => x"c3",
          1497 => x"74",
          1498 => x"54",
          1499 => x"33",
          1500 => x"91",
          1501 => x"f3",
          1502 => x"83",
          1503 => x"38",
          1504 => x"90",
          1505 => x"83",
          1506 => x"75",
          1507 => x"54",
          1508 => x"33",
          1509 => x"95",
          1510 => x"f3",
          1511 => x"83",
          1512 => x"f2",
          1513 => x"ff",
          1514 => x"52",
          1515 => x"3f",
          1516 => x"94",
          1517 => x"bc",
          1518 => x"22",
          1519 => x"8d",
          1520 => x"84",
          1521 => x"84",
          1522 => x"76",
          1523 => x"08",
          1524 => x"e5",
          1525 => x"80",
          1526 => x"74",
          1527 => x"87",
          1528 => x"56",
          1529 => x"da",
          1530 => x"c0",
          1531 => x"ba",
          1532 => x"ff",
          1533 => x"3f",
          1534 => x"08",
          1535 => x"c9",
          1536 => x"84",
          1537 => x"84",
          1538 => x"51",
          1539 => x"33",
          1540 => x"ff",
          1541 => x"c8",
          1542 => x"3f",
          1543 => x"c4",
          1544 => x"f4",
          1545 => x"b3",
          1546 => x"83",
          1547 => x"83",
          1548 => x"f2",
          1549 => x"ff",
          1550 => x"56",
          1551 => x"aa",
          1552 => x"c0",
          1553 => x"ba",
          1554 => x"ff",
          1555 => x"55",
          1556 => x"cc",
          1557 => x"c8",
          1558 => x"80",
          1559 => x"83",
          1560 => x"83",
          1561 => x"fc",
          1562 => x"51",
          1563 => x"33",
          1564 => x"d7",
          1565 => x"88",
          1566 => x"80",
          1567 => x"f3",
          1568 => x"ff",
          1569 => x"56",
          1570 => x"39",
          1571 => x"cc",
          1572 => x"99",
          1573 => x"38",
          1574 => x"83",
          1575 => x"83",
          1576 => x"fb",
          1577 => x"08",
          1578 => x"83",
          1579 => x"83",
          1580 => x"fb",
          1581 => x"08",
          1582 => x"83",
          1583 => x"83",
          1584 => x"fa",
          1585 => x"08",
          1586 => x"83",
          1587 => x"83",
          1588 => x"fa",
          1589 => x"08",
          1590 => x"83",
          1591 => x"83",
          1592 => x"fa",
          1593 => x"08",
          1594 => x"83",
          1595 => x"83",
          1596 => x"f9",
          1597 => x"51",
          1598 => x"51",
          1599 => x"33",
          1600 => x"c4",
          1601 => x"33",
          1602 => x"10",
          1603 => x"08",
          1604 => x"e5",
          1605 => x"b4",
          1606 => x"0d",
          1607 => x"cd",
          1608 => x"c4",
          1609 => x"0d",
          1610 => x"b5",
          1611 => x"d4",
          1612 => x"0d",
          1613 => x"0b",
          1614 => x"f3",
          1615 => x"04",
          1616 => x"3d",
          1617 => x"80",
          1618 => x"88",
          1619 => x"ed",
          1620 => x"f3",
          1621 => x"76",
          1622 => x"8c",
          1623 => x"c0",
          1624 => x"17",
          1625 => x"08",
          1626 => x"ff",
          1627 => x"34",
          1628 => x"9f",
          1629 => x"85",
          1630 => x"f8",
          1631 => x"87",
          1632 => x"38",
          1633 => x"ba",
          1634 => x"e2",
          1635 => x"76",
          1636 => x"52",
          1637 => x"ff",
          1638 => x"84",
          1639 => x"83",
          1640 => x"80",
          1641 => x"0d",
          1642 => x"ad",
          1643 => x"57",
          1644 => x"91",
          1645 => x"75",
          1646 => x"70",
          1647 => x"84",
          1648 => x"08",
          1649 => x"08",
          1650 => x"81",
          1651 => x"99",
          1652 => x"57",
          1653 => x"54",
          1654 => x"0d",
          1655 => x"84",
          1656 => x"c3",
          1657 => x"d1",
          1658 => x"51",
          1659 => x"81",
          1660 => x"38",
          1661 => x"54",
          1662 => x"b6",
          1663 => x"76",
          1664 => x"5b",
          1665 => x"09",
          1666 => x"26",
          1667 => x"56",
          1668 => x"08",
          1669 => x"82",
          1670 => x"80",
          1671 => x"80",
          1672 => x"3f",
          1673 => x"38",
          1674 => x"ba",
          1675 => x"8c",
          1676 => x"08",
          1677 => x"77",
          1678 => x"83",
          1679 => x"3f",
          1680 => x"b2",
          1681 => x"aa",
          1682 => x"3d",
          1683 => x"5a",
          1684 => x"83",
          1685 => x"56",
          1686 => x"f4",
          1687 => x"cb",
          1688 => x"81",
          1689 => x"a0",
          1690 => x"93",
          1691 => x"ea",
          1692 => x"2b",
          1693 => x"2e",
          1694 => x"d1",
          1695 => x"2c",
          1696 => x"70",
          1697 => x"10",
          1698 => x"15",
          1699 => x"52",
          1700 => x"79",
          1701 => x"81",
          1702 => x"81",
          1703 => x"55",
          1704 => x"10",
          1705 => x"0b",
          1706 => x"77",
          1707 => x"15",
          1708 => x"75",
          1709 => x"c2",
          1710 => x"57",
          1711 => x"1b",
          1712 => x"d1",
          1713 => x"2c",
          1714 => x"83",
          1715 => x"5d",
          1716 => x"81",
          1717 => x"fe",
          1718 => x"38",
          1719 => x"0a",
          1720 => x"06",
          1721 => x"c0",
          1722 => x"51",
          1723 => x"33",
          1724 => x"83",
          1725 => x"42",
          1726 => x"76",
          1727 => x"39",
          1728 => x"38",
          1729 => x"39",
          1730 => x"84",
          1731 => x"34",
          1732 => x"55",
          1733 => x"10",
          1734 => x"08",
          1735 => x"0c",
          1736 => x"0b",
          1737 => x"d1",
          1738 => x"85",
          1739 => x"51",
          1740 => x"33",
          1741 => x"34",
          1742 => x"70",
          1743 => x"5b",
          1744 => x"38",
          1745 => x"58",
          1746 => x"70",
          1747 => x"fc",
          1748 => x"38",
          1749 => x"70",
          1750 => x"75",
          1751 => x"84",
          1752 => x"56",
          1753 => x"d5",
          1754 => x"9b",
          1755 => x"51",
          1756 => x"08",
          1757 => x"84",
          1758 => x"84",
          1759 => x"55",
          1760 => x"85",
          1761 => x"cd",
          1762 => x"08",
          1763 => x"10",
          1764 => x"57",
          1765 => x"56",
          1766 => x"51",
          1767 => x"08",
          1768 => x"08",
          1769 => x"52",
          1770 => x"d1",
          1771 => x"56",
          1772 => x"d5",
          1773 => x"83",
          1774 => x"51",
          1775 => x"08",
          1776 => x"84",
          1777 => x"84",
          1778 => x"55",
          1779 => x"81",
          1780 => x"57",
          1781 => x"84",
          1782 => x"76",
          1783 => x"33",
          1784 => x"d1",
          1785 => x"d1",
          1786 => x"27",
          1787 => x"52",
          1788 => x"34",
          1789 => x"b3",
          1790 => x"81",
          1791 => x"57",
          1792 => x"f9",
          1793 => x"d1",
          1794 => x"f9",
          1795 => x"d1",
          1796 => x"2c",
          1797 => x"60",
          1798 => x"f0",
          1799 => x"3f",
          1800 => x"70",
          1801 => x"57",
          1802 => x"38",
          1803 => x"ff",
          1804 => x"29",
          1805 => x"84",
          1806 => x"7b",
          1807 => x"08",
          1808 => x"74",
          1809 => x"05",
          1810 => x"5d",
          1811 => x"38",
          1812 => x"18",
          1813 => x"52",
          1814 => x"75",
          1815 => x"05",
          1816 => x"5b",
          1817 => x"38",
          1818 => x"34",
          1819 => x"51",
          1820 => x"0a",
          1821 => x"2c",
          1822 => x"78",
          1823 => x"39",
          1824 => x"2e",
          1825 => x"52",
          1826 => x"d1",
          1827 => x"d1",
          1828 => x"dd",
          1829 => x"5f",
          1830 => x"52",
          1831 => x"d1",
          1832 => x"84",
          1833 => x"77",
          1834 => x"57",
          1835 => x"f3",
          1836 => x"a4",
          1837 => x"8b",
          1838 => x"06",
          1839 => x"53",
          1840 => x"ba",
          1841 => x"33",
          1842 => x"70",
          1843 => x"38",
          1844 => x"2e",
          1845 => x"77",
          1846 => x"84",
          1847 => x"cc",
          1848 => x"3d",
          1849 => x"74",
          1850 => x"08",
          1851 => x"84",
          1852 => x"af",
          1853 => x"88",
          1854 => x"d0",
          1855 => x"d0",
          1856 => x"cc",
          1857 => x"fd",
          1858 => x"80",
          1859 => x"39",
          1860 => x"34",
          1861 => x"2e",
          1862 => x"88",
          1863 => x"f0",
          1864 => x"3f",
          1865 => x"ff",
          1866 => x"ff",
          1867 => x"7c",
          1868 => x"83",
          1869 => x"80",
          1870 => x"84",
          1871 => x"0c",
          1872 => x"33",
          1873 => x"80",
          1874 => x"33",
          1875 => x"34",
          1876 => x"34",
          1877 => x"ff",
          1878 => x"70",
          1879 => x"cc",
          1880 => x"24",
          1881 => x"52",
          1882 => x"d1",
          1883 => x"2c",
          1884 => x"56",
          1885 => x"d5",
          1886 => x"fb",
          1887 => x"80",
          1888 => x"cc",
          1889 => x"f3",
          1890 => x"88",
          1891 => x"80",
          1892 => x"98",
          1893 => x"55",
          1894 => x"a5",
          1895 => x"77",
          1896 => x"33",
          1897 => x"80",
          1898 => x"98",
          1899 => x"5b",
          1900 => x"16",
          1901 => x"d5",
          1902 => x"ab",
          1903 => x"81",
          1904 => x"d1",
          1905 => x"24",
          1906 => x"d1",
          1907 => x"58",
          1908 => x"d1",
          1909 => x"38",
          1910 => x"41",
          1911 => x"5b",
          1912 => x"80",
          1913 => x"98",
          1914 => x"58",
          1915 => x"55",
          1916 => x"ff",
          1917 => x"7a",
          1918 => x"60",
          1919 => x"84",
          1920 => x"d0",
          1921 => x"ff",
          1922 => x"ff",
          1923 => x"24",
          1924 => x"98",
          1925 => x"59",
          1926 => x"d5",
          1927 => x"b3",
          1928 => x"80",
          1929 => x"cc",
          1930 => x"f1",
          1931 => x"88",
          1932 => x"80",
          1933 => x"98",
          1934 => x"41",
          1935 => x"dd",
          1936 => x"80",
          1937 => x"ad",
          1938 => x"d1",
          1939 => x"ff",
          1940 => x"51",
          1941 => x"33",
          1942 => x"80",
          1943 => x"08",
          1944 => x"84",
          1945 => x"a9",
          1946 => x"88",
          1947 => x"d0",
          1948 => x"d0",
          1949 => x"39",
          1950 => x"ba",
          1951 => x"ba",
          1952 => x"f3",
          1953 => x"c3",
          1954 => x"16",
          1955 => x"3f",
          1956 => x"0a",
          1957 => x"33",
          1958 => x"38",
          1959 => x"70",
          1960 => x"58",
          1961 => x"38",
          1962 => x"80",
          1963 => x"57",
          1964 => x"38",
          1965 => x"80",
          1966 => x"fc",
          1967 => x"80",
          1968 => x"e8",
          1969 => x"80",
          1970 => x"f8",
          1971 => x"ee",
          1972 => x"3f",
          1973 => x"58",
          1974 => x"ff",
          1975 => x"3f",
          1976 => x"34",
          1977 => x"81",
          1978 => x"ab",
          1979 => x"33",
          1980 => x"74",
          1981 => x"f0",
          1982 => x"3f",
          1983 => x"ff",
          1984 => x"52",
          1985 => x"d1",
          1986 => x"d1",
          1987 => x"c7",
          1988 => x"d1",
          1989 => x"34",
          1990 => x"0d",
          1991 => x"84",
          1992 => x"84",
          1993 => x"05",
          1994 => x"97",
          1995 => x"84",
          1996 => x"58",
          1997 => x"93",
          1998 => x"51",
          1999 => x"08",
          2000 => x"84",
          2001 => x"a5",
          2002 => x"05",
          2003 => x"81",
          2004 => x"ff",
          2005 => x"84",
          2006 => x"81",
          2007 => x"7b",
          2008 => x"70",
          2009 => x"84",
          2010 => x"74",
          2011 => x"f0",
          2012 => x"3f",
          2013 => x"ff",
          2014 => x"52",
          2015 => x"d1",
          2016 => x"d1",
          2017 => x"c7",
          2018 => x"83",
          2019 => x"fc",
          2020 => x"70",
          2021 => x"3f",
          2022 => x"f3",
          2023 => x"a4",
          2024 => x"80",
          2025 => x"52",
          2026 => x"f3",
          2027 => x"06",
          2028 => x"38",
          2029 => x"39",
          2030 => x"53",
          2031 => x"3f",
          2032 => x"82",
          2033 => x"51",
          2034 => x"d1",
          2035 => x"34",
          2036 => x"0d",
          2037 => x"8c",
          2038 => x"ba",
          2039 => x"8c",
          2040 => x"f8",
          2041 => x"82",
          2042 => x"5a",
          2043 => x"81",
          2044 => x"08",
          2045 => x"8c",
          2046 => x"08",
          2047 => x"08",
          2048 => x"77",
          2049 => x"fc",
          2050 => x"05",
          2051 => x"80",
          2052 => x"06",
          2053 => x"53",
          2054 => x"ba",
          2055 => x"33",
          2056 => x"70",
          2057 => x"81",
          2058 => x"93",
          2059 => x"ff",
          2060 => x"77",
          2061 => x"53",
          2062 => x"3f",
          2063 => x"81",
          2064 => x"80",
          2065 => x"34",
          2066 => x"c7",
          2067 => x"2b",
          2068 => x"81",
          2069 => x"da",
          2070 => x"0c",
          2071 => x"83",
          2072 => x"41",
          2073 => x"9e",
          2074 => x"f7",
          2075 => x"c0",
          2076 => x"90",
          2077 => x"39",
          2078 => x"33",
          2079 => x"5b",
          2080 => x"72",
          2081 => x"25",
          2082 => x"a8",
          2083 => x"a3",
          2084 => x"9f",
          2085 => x"75",
          2086 => x"bd",
          2087 => x"f9",
          2088 => x"2b",
          2089 => x"7a",
          2090 => x"27",
          2091 => x"56",
          2092 => x"0c",
          2093 => x"27",
          2094 => x"98",
          2095 => x"55",
          2096 => x"74",
          2097 => x"53",
          2098 => x"87",
          2099 => x"33",
          2100 => x"33",
          2101 => x"41",
          2102 => x"0b",
          2103 => x"06",
          2104 => x"06",
          2105 => x"ff",
          2106 => x"58",
          2107 => x"87",
          2108 => x"79",
          2109 => x"7c",
          2110 => x"06",
          2111 => x"14",
          2112 => x"74",
          2113 => x"74",
          2114 => x"59",
          2115 => x"2e",
          2116 => x"72",
          2117 => x"70",
          2118 => x"33",
          2119 => x"39",
          2120 => x"b0",
          2121 => x"81",
          2122 => x"81",
          2123 => x"74",
          2124 => x"5e",
          2125 => x"73",
          2126 => x"71",
          2127 => x"80",
          2128 => x"f9",
          2129 => x"34",
          2130 => x"71",
          2131 => x"71",
          2132 => x"76",
          2133 => x"39",
          2134 => x"33",
          2135 => x"11",
          2136 => x"11",
          2137 => x"5b",
          2138 => x"70",
          2139 => x"ff",
          2140 => x"ff",
          2141 => x"ff",
          2142 => x"5e",
          2143 => x"57",
          2144 => x"31",
          2145 => x"7d",
          2146 => x"71",
          2147 => x"62",
          2148 => x"5f",
          2149 => x"85",
          2150 => x"31",
          2151 => x"fd",
          2152 => x"fd",
          2153 => x"31",
          2154 => x"3d",
          2155 => x"f4",
          2156 => x"ee",
          2157 => x"73",
          2158 => x"76",
          2159 => x"34",
          2160 => x"75",
          2161 => x"81",
          2162 => x"d8",
          2163 => x"54",
          2164 => x"f8",
          2165 => x"72",
          2166 => x"06",
          2167 => x"34",
          2168 => x"06",
          2169 => x"81",
          2170 => x"88",
          2171 => x"0b",
          2172 => x"ba",
          2173 => x"b8",
          2174 => x"f7",
          2175 => x"84",
          2176 => x"33",
          2177 => x"26",
          2178 => x"83",
          2179 => x"72",
          2180 => x"11",
          2181 => x"59",
          2182 => x"ff",
          2183 => x"58",
          2184 => x"83",
          2185 => x"83",
          2186 => x"76",
          2187 => x"ff",
          2188 => x"82",
          2189 => x"f9",
          2190 => x"83",
          2191 => x"5c",
          2192 => x"38",
          2193 => x"54",
          2194 => x"ac",
          2195 => x"55",
          2196 => x"34",
          2197 => x"70",
          2198 => x"84",
          2199 => x"9f",
          2200 => x"33",
          2201 => x"0b",
          2202 => x"81",
          2203 => x"9f",
          2204 => x"33",
          2205 => x"23",
          2206 => x"83",
          2207 => x"26",
          2208 => x"05",
          2209 => x"58",
          2210 => x"80",
          2211 => x"ff",
          2212 => x"29",
          2213 => x"27",
          2214 => x"e0",
          2215 => x"13",
          2216 => x"73",
          2217 => x"81",
          2218 => x"80",
          2219 => x"29",
          2220 => x"26",
          2221 => x"8c",
          2222 => x"f9",
          2223 => x"83",
          2224 => x"5c",
          2225 => x"38",
          2226 => x"81",
          2227 => x"33",
          2228 => x"06",
          2229 => x"05",
          2230 => x"78",
          2231 => x"73",
          2232 => x"b8",
          2233 => x"31",
          2234 => x"16",
          2235 => x"34",
          2236 => x"8a",
          2237 => x"75",
          2238 => x"13",
          2239 => x"80",
          2240 => x"fe",
          2241 => x"59",
          2242 => x"84",
          2243 => x"fc",
          2244 => x"05",
          2245 => x"38",
          2246 => x"51",
          2247 => x"51",
          2248 => x"f9",
          2249 => x"0c",
          2250 => x"f9",
          2251 => x"81",
          2252 => x"e2",
          2253 => x"bc",
          2254 => x"86",
          2255 => x"70",
          2256 => x"72",
          2257 => x"f9",
          2258 => x"33",
          2259 => x"11",
          2260 => x"38",
          2261 => x"80",
          2262 => x"0d",
          2263 => x"31",
          2264 => x"54",
          2265 => x"34",
          2266 => x"3d",
          2267 => x"05",
          2268 => x"55",
          2269 => x"53",
          2270 => x"84",
          2271 => x"80",
          2272 => x"bc",
          2273 => x"56",
          2274 => x"81",
          2275 => x"fe",
          2276 => x"05",
          2277 => x"70",
          2278 => x"70",
          2279 => x"80",
          2280 => x"06",
          2281 => x"53",
          2282 => x"06",
          2283 => x"b8",
          2284 => x"83",
          2285 => x"81",
          2286 => x"f9",
          2287 => x"0c",
          2288 => x"33",
          2289 => x"b8",
          2290 => x"81",
          2291 => x"f9",
          2292 => x"83",
          2293 => x"8c",
          2294 => x"b8",
          2295 => x"70",
          2296 => x"83",
          2297 => x"83",
          2298 => x"f9",
          2299 => x"51",
          2300 => x"39",
          2301 => x"83",
          2302 => x"ff",
          2303 => x"f9",
          2304 => x"b8",
          2305 => x"33",
          2306 => x"b8",
          2307 => x"33",
          2308 => x"70",
          2309 => x"83",
          2310 => x"07",
          2311 => x"ba",
          2312 => x"06",
          2313 => x"b8",
          2314 => x"33",
          2315 => x"70",
          2316 => x"83",
          2317 => x"07",
          2318 => x"82",
          2319 => x"06",
          2320 => x"f2",
          2321 => x"06",
          2322 => x"34",
          2323 => x"bf",
          2324 => x"05",
          2325 => x"bb",
          2326 => x"82",
          2327 => x"78",
          2328 => x"24",
          2329 => x"38",
          2330 => x"84",
          2331 => x"34",
          2332 => x"f9",
          2333 => x"83",
          2334 => x"0b",
          2335 => x"b8",
          2336 => x"34",
          2337 => x"0b",
          2338 => x"b8",
          2339 => x"56",
          2340 => x"7c",
          2341 => x"ff",
          2342 => x"34",
          2343 => x"83",
          2344 => x"23",
          2345 => x"0d",
          2346 => x"81",
          2347 => x"83",
          2348 => x"bd",
          2349 => x"84",
          2350 => x"33",
          2351 => x"55",
          2352 => x"e3",
          2353 => x"0b",
          2354 => x"79",
          2355 => x"e0",
          2356 => x"f8",
          2357 => x"70",
          2358 => x"52",
          2359 => x"83",
          2360 => x"7d",
          2361 => x"b8",
          2362 => x"7b",
          2363 => x"bd",
          2364 => x"84",
          2365 => x"84",
          2366 => x"a8",
          2367 => x"83",
          2368 => x"ff",
          2369 => x"52",
          2370 => x"3f",
          2371 => x"92",
          2372 => x"27",
          2373 => x"33",
          2374 => x"d5",
          2375 => x"5a",
          2376 => x"02",
          2377 => x"80",
          2378 => x"bc",
          2379 => x"a0",
          2380 => x"51",
          2381 => x"83",
          2382 => x"52",
          2383 => x"2e",
          2384 => x"f9",
          2385 => x"75",
          2386 => x"2e",
          2387 => x"83",
          2388 => x"72",
          2389 => x"b8",
          2390 => x"14",
          2391 => x"bd",
          2392 => x"29",
          2393 => x"f9",
          2394 => x"73",
          2395 => x"b8",
          2396 => x"84",
          2397 => x"83",
          2398 => x"72",
          2399 => x"57",
          2400 => x"14",
          2401 => x"59",
          2402 => x"84",
          2403 => x"38",
          2404 => x"34",
          2405 => x"2e",
          2406 => x"76",
          2407 => x"84",
          2408 => x"75",
          2409 => x"80",
          2410 => x"06",
          2411 => x"f1",
          2412 => x"34",
          2413 => x"33",
          2414 => x"34",
          2415 => x"89",
          2416 => x"fd",
          2417 => x"06",
          2418 => x"38",
          2419 => x"81",
          2420 => x"83",
          2421 => x"74",
          2422 => x"75",
          2423 => x"0b",
          2424 => x"04",
          2425 => x"fd",
          2426 => x"81",
          2427 => x"83",
          2428 => x"34",
          2429 => x"83",
          2430 => x"55",
          2431 => x"73",
          2432 => x"a0",
          2433 => x"81",
          2434 => x"90",
          2435 => x"3f",
          2436 => x"80",
          2437 => x"57",
          2438 => x"75",
          2439 => x"2e",
          2440 => x"d1",
          2441 => x"78",
          2442 => x"80",
          2443 => x"bd",
          2444 => x"5c",
          2445 => x"a0",
          2446 => x"83",
          2447 => x"72",
          2448 => x"78",
          2449 => x"bc",
          2450 => x"5a",
          2451 => x"b0",
          2452 => x"70",
          2453 => x"83",
          2454 => x"42",
          2455 => x"33",
          2456 => x"70",
          2457 => x"26",
          2458 => x"5a",
          2459 => x"75",
          2460 => x"ba",
          2461 => x"b7",
          2462 => x"81",
          2463 => x"38",
          2464 => x"80",
          2465 => x"80",
          2466 => x"bd",
          2467 => x"40",
          2468 => x"a0",
          2469 => x"83",
          2470 => x"72",
          2471 => x"78",
          2472 => x"bc",
          2473 => x"83",
          2474 => x"1b",
          2475 => x"ff",
          2476 => x"bd",
          2477 => x"43",
          2478 => x"84",
          2479 => x"77",
          2480 => x"fe",
          2481 => x"80",
          2482 => x"0d",
          2483 => x"78",
          2484 => x"2e",
          2485 => x"0b",
          2486 => x"ba",
          2487 => x"9b",
          2488 => x"75",
          2489 => x"8c",
          2490 => x"b9",
          2491 => x"34",
          2492 => x"84",
          2493 => x"ba",
          2494 => x"9b",
          2495 => x"b9",
          2496 => x"f9",
          2497 => x"72",
          2498 => x"88",
          2499 => x"34",
          2500 => x"33",
          2501 => x"12",
          2502 => x"be",
          2503 => x"71",
          2504 => x"33",
          2505 => x"b8",
          2506 => x"f9",
          2507 => x"72",
          2508 => x"83",
          2509 => x"05",
          2510 => x"81",
          2511 => x"0b",
          2512 => x"84",
          2513 => x"70",
          2514 => x"73",
          2515 => x"05",
          2516 => x"72",
          2517 => x"06",
          2518 => x"5a",
          2519 => x"78",
          2520 => x"76",
          2521 => x"f9",
          2522 => x"84",
          2523 => x"8d",
          2524 => x"80",
          2525 => x"84",
          2526 => x"8c",
          2527 => x"bc",
          2528 => x"bd",
          2529 => x"bb",
          2530 => x"84",
          2531 => x"8c",
          2532 => x"ff",
          2533 => x"83",
          2534 => x"70",
          2535 => x"70",
          2536 => x"87",
          2537 => x"22",
          2538 => x"83",
          2539 => x"44",
          2540 => x"81",
          2541 => x"06",
          2542 => x"75",
          2543 => x"81",
          2544 => x"81",
          2545 => x"40",
          2546 => x"a0",
          2547 => x"83",
          2548 => x"72",
          2549 => x"a0",
          2550 => x"f9",
          2551 => x"5a",
          2552 => x"b0",
          2553 => x"70",
          2554 => x"83",
          2555 => x"43",
          2556 => x"33",
          2557 => x"1a",
          2558 => x"7b",
          2559 => x"33",
          2560 => x"58",
          2561 => x"bd",
          2562 => x"05",
          2563 => x"95",
          2564 => x"38",
          2565 => x"b9",
          2566 => x"ff",
          2567 => x"c8",
          2568 => x"05",
          2569 => x"f9",
          2570 => x"9f",
          2571 => x"9c",
          2572 => x"84",
          2573 => x"83",
          2574 => x"72",
          2575 => x"05",
          2576 => x"7b",
          2577 => x"83",
          2578 => x"59",
          2579 => x"38",
          2580 => x"81",
          2581 => x"72",
          2582 => x"a8",
          2583 => x"84",
          2584 => x"83",
          2585 => x"5e",
          2586 => x"be",
          2587 => x"71",
          2588 => x"33",
          2589 => x"b8",
          2590 => x"f9",
          2591 => x"72",
          2592 => x"83",
          2593 => x"34",
          2594 => x"5b",
          2595 => x"84",
          2596 => x"38",
          2597 => x"34",
          2598 => x"59",
          2599 => x"f9",
          2600 => x"f9",
          2601 => x"81",
          2602 => x"72",
          2603 => x"5b",
          2604 => x"80",
          2605 => x"f9",
          2606 => x"71",
          2607 => x"0b",
          2608 => x"bc",
          2609 => x"83",
          2610 => x"1a",
          2611 => x"ff",
          2612 => x"bd",
          2613 => x"5a",
          2614 => x"98",
          2615 => x"81",
          2616 => x"fe",
          2617 => x"fe",
          2618 => x"0c",
          2619 => x"3d",
          2620 => x"59",
          2621 => x"83",
          2622 => x"58",
          2623 => x"0b",
          2624 => x"ba",
          2625 => x"f9",
          2626 => x"1b",
          2627 => x"84",
          2628 => x"5b",
          2629 => x"84",
          2630 => x"53",
          2631 => x"84",
          2632 => x"38",
          2633 => x"5a",
          2634 => x"83",
          2635 => x"22",
          2636 => x"cf",
          2637 => x"84",
          2638 => x"f9",
          2639 => x"f9",
          2640 => x"39",
          2641 => x"33",
          2642 => x"05",
          2643 => x"33",
          2644 => x"84",
          2645 => x"83",
          2646 => x"5a",
          2647 => x"18",
          2648 => x"29",
          2649 => x"60",
          2650 => x"b8",
          2651 => x"f9",
          2652 => x"72",
          2653 => x"83",
          2654 => x"34",
          2655 => x"58",
          2656 => x"b8",
          2657 => x"ff",
          2658 => x"80",
          2659 => x"83",
          2660 => x"38",
          2661 => x"b4",
          2662 => x"3f",
          2663 => x"3d",
          2664 => x"f9",
          2665 => x"f9",
          2666 => x"76",
          2667 => x"83",
          2668 => x"83",
          2669 => x"83",
          2670 => x"ff",
          2671 => x"7a",
          2672 => x"e0",
          2673 => x"06",
          2674 => x"81",
          2675 => x"05",
          2676 => x"94",
          2677 => x"3f",
          2678 => x"ba",
          2679 => x"90",
          2680 => x"24",
          2681 => x"f0",
          2682 => x"39",
          2683 => x"58",
          2684 => x"27",
          2685 => x"e0",
          2686 => x"b1",
          2687 => x"83",
          2688 => x"84",
          2689 => x"8f",
          2690 => x"b9",
          2691 => x"70",
          2692 => x"5e",
          2693 => x"e7",
          2694 => x"80",
          2695 => x"33",
          2696 => x"b8",
          2697 => x"27",
          2698 => x"34",
          2699 => x"bd",
          2700 => x"ff",
          2701 => x"a7",
          2702 => x"bc",
          2703 => x"f9",
          2704 => x"b7",
          2705 => x"76",
          2706 => x"75",
          2707 => x"84",
          2708 => x"8d",
          2709 => x"b9",
          2710 => x"70",
          2711 => x"42",
          2712 => x"cf",
          2713 => x"80",
          2714 => x"22",
          2715 => x"fc",
          2716 => x"f9",
          2717 => x"71",
          2718 => x"83",
          2719 => x"71",
          2720 => x"06",
          2721 => x"80",
          2722 => x"82",
          2723 => x"83",
          2724 => x"b9",
          2725 => x"e7",
          2726 => x"99",
          2727 => x"81",
          2728 => x"39",
          2729 => x"2e",
          2730 => x"83",
          2731 => x"b8",
          2732 => x"75",
          2733 => x"83",
          2734 => x"b9",
          2735 => x"c8",
          2736 => x"bc",
          2737 => x"33",
          2738 => x"25",
          2739 => x"bc",
          2740 => x"51",
          2741 => x"b9",
          2742 => x"8b",
          2743 => x"05",
          2744 => x"51",
          2745 => x"81",
          2746 => x"58",
          2747 => x"8d",
          2748 => x"38",
          2749 => x"26",
          2750 => x"81",
          2751 => x"97",
          2752 => x"77",
          2753 => x"33",
          2754 => x"b9",
          2755 => x"06",
          2756 => x"06",
          2757 => x"5c",
          2758 => x"5a",
          2759 => x"ff",
          2760 => x"27",
          2761 => x"bc",
          2762 => x"57",
          2763 => x"7a",
          2764 => x"af",
          2765 => x"80",
          2766 => x"33",
          2767 => x"7f",
          2768 => x"33",
          2769 => x"06",
          2770 => x"11",
          2771 => x"ba",
          2772 => x"70",
          2773 => x"33",
          2774 => x"81",
          2775 => x"ff",
          2776 => x"7c",
          2777 => x"33",
          2778 => x"ff",
          2779 => x"7c",
          2780 => x"57",
          2781 => x"b7",
          2782 => x"ee",
          2783 => x"bc",
          2784 => x"ba",
          2785 => x"26",
          2786 => x"7e",
          2787 => x"5e",
          2788 => x"5b",
          2789 => x"06",
          2790 => x"1d",
          2791 => x"f7",
          2792 => x"e0",
          2793 => x"1f",
          2794 => x"76",
          2795 => x"81",
          2796 => x"80",
          2797 => x"29",
          2798 => x"27",
          2799 => x"5f",
          2800 => x"81",
          2801 => x"58",
          2802 => x"81",
          2803 => x"ff",
          2804 => x"5e",
          2805 => x"f6",
          2806 => x"75",
          2807 => x"84",
          2808 => x"f6",
          2809 => x"33",
          2810 => x"59",
          2811 => x"84",
          2812 => x"09",
          2813 => x"bd",
          2814 => x"f9",
          2815 => x"ff",
          2816 => x"33",
          2817 => x"7e",
          2818 => x"f5",
          2819 => x"27",
          2820 => x"10",
          2821 => x"87",
          2822 => x"5a",
          2823 => x"06",
          2824 => x"79",
          2825 => x"83",
          2826 => x"90",
          2827 => x"07",
          2828 => x"7a",
          2829 => x"05",
          2830 => x"58",
          2831 => x"b8",
          2832 => x"5f",
          2833 => x"06",
          2834 => x"64",
          2835 => x"26",
          2836 => x"7b",
          2837 => x"1d",
          2838 => x"38",
          2839 => x"18",
          2840 => x"34",
          2841 => x"81",
          2842 => x"38",
          2843 => x"78",
          2844 => x"57",
          2845 => x"39",
          2846 => x"58",
          2847 => x"70",
          2848 => x"f0",
          2849 => x"57",
          2850 => x"be",
          2851 => x"34",
          2852 => x"56",
          2853 => x"33",
          2854 => x"34",
          2855 => x"33",
          2856 => x"33",
          2857 => x"83",
          2858 => x"83",
          2859 => x"ff",
          2860 => x"f9",
          2861 => x"56",
          2862 => x"83",
          2863 => x"07",
          2864 => x"39",
          2865 => x"81",
          2866 => x"c3",
          2867 => x"06",
          2868 => x"34",
          2869 => x"f9",
          2870 => x"06",
          2871 => x"b8",
          2872 => x"f9",
          2873 => x"b8",
          2874 => x"75",
          2875 => x"83",
          2876 => x"e0",
          2877 => x"fe",
          2878 => x"cf",
          2879 => x"f9",
          2880 => x"b8",
          2881 => x"75",
          2882 => x"83",
          2883 => x"07",
          2884 => x"b3",
          2885 => x"06",
          2886 => x"34",
          2887 => x"81",
          2888 => x"f9",
          2889 => x"b8",
          2890 => x"f9",
          2891 => x"b8",
          2892 => x"f9",
          2893 => x"b8",
          2894 => x"f9",
          2895 => x"b8",
          2896 => x"56",
          2897 => x"39",
          2898 => x"b0",
          2899 => x"fd",
          2900 => x"34",
          2901 => x"ec",
          2902 => x"f9",
          2903 => x"f9",
          2904 => x"78",
          2905 => x"b9",
          2906 => x"84",
          2907 => x"8c",
          2908 => x"f9",
          2909 => x"81",
          2910 => x"cf",
          2911 => x"dc",
          2912 => x"83",
          2913 => x"84",
          2914 => x"80",
          2915 => x"84",
          2916 => x"77",
          2917 => x"84",
          2918 => x"7a",
          2919 => x"fe",
          2920 => x"84",
          2921 => x"b9",
          2922 => x"f9",
          2923 => x"97",
          2924 => x"ff",
          2925 => x"39",
          2926 => x"52",
          2927 => x"39",
          2928 => x"8f",
          2929 => x"70",
          2930 => x"5f",
          2931 => x"51",
          2932 => x"75",
          2933 => x"f9",
          2934 => x"bc",
          2935 => x"2c",
          2936 => x"39",
          2937 => x"b7",
          2938 => x"75",
          2939 => x"f3",
          2940 => x"81",
          2941 => x"ee",
          2942 => x"b8",
          2943 => x"f9",
          2944 => x"a3",
          2945 => x"5f",
          2946 => x"ff",
          2947 => x"5b",
          2948 => x"81",
          2949 => x"ff",
          2950 => x"89",
          2951 => x"76",
          2952 => x"75",
          2953 => x"06",
          2954 => x"83",
          2955 => x"76",
          2956 => x"56",
          2957 => x"ff",
          2958 => x"80",
          2959 => x"77",
          2960 => x"71",
          2961 => x"87",
          2962 => x"80",
          2963 => x"06",
          2964 => x"5d",
          2965 => x"98",
          2966 => x"5e",
          2967 => x"81",
          2968 => x"58",
          2969 => x"81",
          2970 => x"ff",
          2971 => x"5d",
          2972 => x"e0",
          2973 => x"1e",
          2974 => x"76",
          2975 => x"81",
          2976 => x"80",
          2977 => x"29",
          2978 => x"26",
          2979 => x"f9",
          2980 => x"1c",
          2981 => x"84",
          2982 => x"84",
          2983 => x"fd",
          2984 => x"b7",
          2985 => x"11",
          2986 => x"38",
          2987 => x"77",
          2988 => x"80",
          2989 => x"83",
          2990 => x"70",
          2991 => x"56",
          2992 => x"56",
          2993 => x"39",
          2994 => x"b8",
          2995 => x"75",
          2996 => x"ef",
          2997 => x"06",
          2998 => x"70",
          2999 => x"7a",
          3000 => x"09",
          3001 => x"39",
          3002 => x"34",
          3003 => x"83",
          3004 => x"7b",
          3005 => x"f2",
          3006 => x"7a",
          3007 => x"81",
          3008 => x"77",
          3009 => x"26",
          3010 => x"05",
          3011 => x"70",
          3012 => x"d4",
          3013 => x"56",
          3014 => x"39",
          3015 => x"ad",
          3016 => x"84",
          3017 => x"f1",
          3018 => x"34",
          3019 => x"33",
          3020 => x"34",
          3021 => x"a7",
          3022 => x"33",
          3023 => x"80",
          3024 => x"3f",
          3025 => x"3d",
          3026 => x"ab",
          3027 => x"85",
          3028 => x"bf",
          3029 => x"90",
          3030 => x"f0",
          3031 => x"80",
          3032 => x"75",
          3033 => x"84",
          3034 => x"83",
          3035 => x"80",
          3036 => x"30",
          3037 => x"56",
          3038 => x"0c",
          3039 => x"09",
          3040 => x"83",
          3041 => x"07",
          3042 => x"c4",
          3043 => x"bd",
          3044 => x"29",
          3045 => x"f9",
          3046 => x"29",
          3047 => x"f8",
          3048 => x"81",
          3049 => x"73",
          3050 => x"87",
          3051 => x"88",
          3052 => x"86",
          3053 => x"f5",
          3054 => x"ff",
          3055 => x"cf",
          3056 => x"33",
          3057 => x"16",
          3058 => x"85",
          3059 => x"b4",
          3060 => x"75",
          3061 => x"2e",
          3062 => x"15",
          3063 => x"f7",
          3064 => x"ff",
          3065 => x"b3",
          3066 => x"2b",
          3067 => x"83",
          3068 => x"70",
          3069 => x"51",
          3070 => x"38",
          3071 => x"09",
          3072 => x"e4",
          3073 => x"80",
          3074 => x"ec",
          3075 => x"f7",
          3076 => x"5d",
          3077 => x"c0",
          3078 => x"8d",
          3079 => x"73",
          3080 => x"ca",
          3081 => x"8b",
          3082 => x"73",
          3083 => x"54",
          3084 => x"f7",
          3085 => x"81",
          3086 => x"72",
          3087 => x"f7",
          3088 => x"84",
          3089 => x"e8",
          3090 => x"54",
          3091 => x"0b",
          3092 => x"e0",
          3093 => x"06",
          3094 => x"38",
          3095 => x"f7",
          3096 => x"9c",
          3097 => x"83",
          3098 => x"83",
          3099 => x"91",
          3100 => x"9c",
          3101 => x"dc",
          3102 => x"54",
          3103 => x"54",
          3104 => x"98",
          3105 => x"81",
          3106 => x"38",
          3107 => x"b8",
          3108 => x"54",
          3109 => x"53",
          3110 => x"81",
          3111 => x"34",
          3112 => x"58",
          3113 => x"83",
          3114 => x"77",
          3115 => x"7d",
          3116 => x"2e",
          3117 => x"59",
          3118 => x"54",
          3119 => x"2e",
          3120 => x"06",
          3121 => x"27",
          3122 => x"54",
          3123 => x"10",
          3124 => x"2b",
          3125 => x"33",
          3126 => x"9c",
          3127 => x"ea",
          3128 => x"a8",
          3129 => x"a0",
          3130 => x"ff",
          3131 => x"b8",
          3132 => x"83",
          3133 => x"70",
          3134 => x"7d",
          3135 => x"06",
          3136 => x"c6",
          3137 => x"83",
          3138 => x"78",
          3139 => x"70",
          3140 => x"27",
          3141 => x"72",
          3142 => x"84",
          3143 => x"81",
          3144 => x"3f",
          3145 => x"0d",
          3146 => x"f9",
          3147 => x"38",
          3148 => x"5b",
          3149 => x"c9",
          3150 => x"34",
          3151 => x"ff",
          3152 => x"b1",
          3153 => x"81",
          3154 => x"d4",
          3155 => x"8a",
          3156 => x"81",
          3157 => x"83",
          3158 => x"c0",
          3159 => x"27",
          3160 => x"08",
          3161 => x"06",
          3162 => x"f7",
          3163 => x"83",
          3164 => x"53",
          3165 => x"e6",
          3166 => x"83",
          3167 => x"70",
          3168 => x"33",
          3169 => x"fa",
          3170 => x"06",
          3171 => x"2e",
          3172 => x"81",
          3173 => x"ef",
          3174 => x"39",
          3175 => x"54",
          3176 => x"b8",
          3177 => x"80",
          3178 => x"76",
          3179 => x"82",
          3180 => x"53",
          3181 => x"83",
          3182 => x"f6",
          3183 => x"81",
          3184 => x"80",
          3185 => x"83",
          3186 => x"ff",
          3187 => x"38",
          3188 => x"84",
          3189 => x"56",
          3190 => x"38",
          3191 => x"ff",
          3192 => x"51",
          3193 => x"aa",
          3194 => x"14",
          3195 => x"de",
          3196 => x"34",
          3197 => x"39",
          3198 => x"3f",
          3199 => x"80",
          3200 => x"02",
          3201 => x"f4",
          3202 => x"85",
          3203 => x"fe",
          3204 => x"f0",
          3205 => x"08",
          3206 => x"90",
          3207 => x"53",
          3208 => x"73",
          3209 => x"c0",
          3210 => x"27",
          3211 => x"38",
          3212 => x"56",
          3213 => x"56",
          3214 => x"c0",
          3215 => x"54",
          3216 => x"c0",
          3217 => x"f6",
          3218 => x"9c",
          3219 => x"38",
          3220 => x"c0",
          3221 => x"74",
          3222 => x"2e",
          3223 => x"75",
          3224 => x"38",
          3225 => x"ba",
          3226 => x"17",
          3227 => x"df",
          3228 => x"58",
          3229 => x"8c",
          3230 => x"0d",
          3231 => x"57",
          3232 => x"74",
          3233 => x"70",
          3234 => x"58",
          3235 => x"52",
          3236 => x"57",
          3237 => x"34",
          3238 => x"14",
          3239 => x"e1",
          3240 => x"08",
          3241 => x"80",
          3242 => x"c0",
          3243 => x"56",
          3244 => x"98",
          3245 => x"08",
          3246 => x"15",
          3247 => x"53",
          3248 => x"fe",
          3249 => x"08",
          3250 => x"cf",
          3251 => x"c7",
          3252 => x"ce",
          3253 => x"08",
          3254 => x"75",
          3255 => x"87",
          3256 => x"74",
          3257 => x"db",
          3258 => x"ff",
          3259 => x"72",
          3260 => x"76",
          3261 => x"ff",
          3262 => x"52",
          3263 => x"38",
          3264 => x"56",
          3265 => x"72",
          3266 => x"81",
          3267 => x"38",
          3268 => x"0d",
          3269 => x"58",
          3270 => x"8c",
          3271 => x"70",
          3272 => x"a5",
          3273 => x"3d",
          3274 => x"33",
          3275 => x"08",
          3276 => x"06",
          3277 => x"56",
          3278 => x"2a",
          3279 => x"2a",
          3280 => x"16",
          3281 => x"c6",
          3282 => x"52",
          3283 => x"81",
          3284 => x"55",
          3285 => x"f4",
          3286 => x"83",
          3287 => x"34",
          3288 => x"57",
          3289 => x"86",
          3290 => x"9c",
          3291 => x"ce",
          3292 => x"08",
          3293 => x"71",
          3294 => x"87",
          3295 => x"74",
          3296 => x"db",
          3297 => x"ff",
          3298 => x"72",
          3299 => x"87",
          3300 => x"05",
          3301 => x"87",
          3302 => x"2e",
          3303 => x"98",
          3304 => x"87",
          3305 => x"87",
          3306 => x"71",
          3307 => x"ff",
          3308 => x"38",
          3309 => x"d8",
          3310 => x"52",
          3311 => x"0c",
          3312 => x"81",
          3313 => x"ff",
          3314 => x"80",
          3315 => x"fc",
          3316 => x"84",
          3317 => x"fb",
          3318 => x"80",
          3319 => x"98",
          3320 => x"34",
          3321 => x"87",
          3322 => x"08",
          3323 => x"c0",
          3324 => x"9c",
          3325 => x"81",
          3326 => x"52",
          3327 => x"81",
          3328 => x"a4",
          3329 => x"80",
          3330 => x"80",
          3331 => x"80",
          3332 => x"9c",
          3333 => x"53",
          3334 => x"33",
          3335 => x"70",
          3336 => x"2e",
          3337 => x"51",
          3338 => x"71",
          3339 => x"80",
          3340 => x"52",
          3341 => x"16",
          3342 => x"39",
          3343 => x"fe",
          3344 => x"f9",
          3345 => x"71",
          3346 => x"06",
          3347 => x"81",
          3348 => x"2b",
          3349 => x"33",
          3350 => x"5c",
          3351 => x"52",
          3352 => x"af",
          3353 => x"12",
          3354 => x"07",
          3355 => x"71",
          3356 => x"53",
          3357 => x"24",
          3358 => x"14",
          3359 => x"07",
          3360 => x"56",
          3361 => x"ff",
          3362 => x"b9",
          3363 => x"85",
          3364 => x"88",
          3365 => x"84",
          3366 => x"b9",
          3367 => x"13",
          3368 => x"b9",
          3369 => x"73",
          3370 => x"16",
          3371 => x"2b",
          3372 => x"2a",
          3373 => x"75",
          3374 => x"86",
          3375 => x"2b",
          3376 => x"16",
          3377 => x"07",
          3378 => x"53",
          3379 => x"85",
          3380 => x"16",
          3381 => x"8b",
          3382 => x"5a",
          3383 => x"13",
          3384 => x"2a",
          3385 => x"34",
          3386 => x"08",
          3387 => x"88",
          3388 => x"88",
          3389 => x"34",
          3390 => x"08",
          3391 => x"71",
          3392 => x"05",
          3393 => x"2b",
          3394 => x"06",
          3395 => x"53",
          3396 => x"82",
          3397 => x"b9",
          3398 => x"12",
          3399 => x"07",
          3400 => x"71",
          3401 => x"70",
          3402 => x"57",
          3403 => x"14",
          3404 => x"82",
          3405 => x"2b",
          3406 => x"33",
          3407 => x"90",
          3408 => x"57",
          3409 => x"38",
          3410 => x"2b",
          3411 => x"2a",
          3412 => x"81",
          3413 => x"17",
          3414 => x"2b",
          3415 => x"14",
          3416 => x"07",
          3417 => x"58",
          3418 => x"75",
          3419 => x"f9",
          3420 => x"58",
          3421 => x"80",
          3422 => x"3f",
          3423 => x"0b",
          3424 => x"84",
          3425 => x"76",
          3426 => x"ec",
          3427 => x"75",
          3428 => x"b9",
          3429 => x"81",
          3430 => x"08",
          3431 => x"87",
          3432 => x"b9",
          3433 => x"07",
          3434 => x"2a",
          3435 => x"34",
          3436 => x"22",
          3437 => x"08",
          3438 => x"15",
          3439 => x"ee",
          3440 => x"53",
          3441 => x"fb",
          3442 => x"ff",
          3443 => x"ff",
          3444 => x"33",
          3445 => x"70",
          3446 => x"ff",
          3447 => x"75",
          3448 => x"12",
          3449 => x"ff",
          3450 => x"ff",
          3451 => x"5c",
          3452 => x"70",
          3453 => x"58",
          3454 => x"88",
          3455 => x"73",
          3456 => x"74",
          3457 => x"11",
          3458 => x"2b",
          3459 => x"56",
          3460 => x"83",
          3461 => x"26",
          3462 => x"2e",
          3463 => x"88",
          3464 => x"11",
          3465 => x"2a",
          3466 => x"34",
          3467 => x"08",
          3468 => x"82",
          3469 => x"b9",
          3470 => x"12",
          3471 => x"2b",
          3472 => x"83",
          3473 => x"58",
          3474 => x"12",
          3475 => x"83",
          3476 => x"54",
          3477 => x"84",
          3478 => x"33",
          3479 => x"83",
          3480 => x"53",
          3481 => x"15",
          3482 => x"55",
          3483 => x"33",
          3484 => x"54",
          3485 => x"71",
          3486 => x"70",
          3487 => x"71",
          3488 => x"05",
          3489 => x"15",
          3490 => x"fc",
          3491 => x"11",
          3492 => x"07",
          3493 => x"70",
          3494 => x"84",
          3495 => x"70",
          3496 => x"04",
          3497 => x"8b",
          3498 => x"84",
          3499 => x"2b",
          3500 => x"53",
          3501 => x"85",
          3502 => x"19",
          3503 => x"8b",
          3504 => x"86",
          3505 => x"2b",
          3506 => x"52",
          3507 => x"34",
          3508 => x"08",
          3509 => x"88",
          3510 => x"88",
          3511 => x"34",
          3512 => x"08",
          3513 => x"f9",
          3514 => x"58",
          3515 => x"54",
          3516 => x"0c",
          3517 => x"91",
          3518 => x"8c",
          3519 => x"f4",
          3520 => x"0b",
          3521 => x"53",
          3522 => x"cc",
          3523 => x"76",
          3524 => x"84",
          3525 => x"34",
          3526 => x"fc",
          3527 => x"0b",
          3528 => x"84",
          3529 => x"80",
          3530 => x"88",
          3531 => x"17",
          3532 => x"f8",
          3533 => x"fc",
          3534 => x"82",
          3535 => x"77",
          3536 => x"fe",
          3537 => x"41",
          3538 => x"59",
          3539 => x"38",
          3540 => x"80",
          3541 => x"60",
          3542 => x"2a",
          3543 => x"55",
          3544 => x"78",
          3545 => x"06",
          3546 => x"81",
          3547 => x"75",
          3548 => x"10",
          3549 => x"61",
          3550 => x"88",
          3551 => x"2c",
          3552 => x"43",
          3553 => x"42",
          3554 => x"15",
          3555 => x"07",
          3556 => x"81",
          3557 => x"2b",
          3558 => x"80",
          3559 => x"27",
          3560 => x"62",
          3561 => x"85",
          3562 => x"25",
          3563 => x"79",
          3564 => x"33",
          3565 => x"83",
          3566 => x"12",
          3567 => x"07",
          3568 => x"58",
          3569 => x"1e",
          3570 => x"8b",
          3571 => x"86",
          3572 => x"2b",
          3573 => x"14",
          3574 => x"07",
          3575 => x"5b",
          3576 => x"84",
          3577 => x"b9",
          3578 => x"85",
          3579 => x"2b",
          3580 => x"15",
          3581 => x"2a",
          3582 => x"57",
          3583 => x"34",
          3584 => x"81",
          3585 => x"ff",
          3586 => x"5e",
          3587 => x"34",
          3588 => x"11",
          3589 => x"71",
          3590 => x"81",
          3591 => x"88",
          3592 => x"55",
          3593 => x"34",
          3594 => x"33",
          3595 => x"83",
          3596 => x"83",
          3597 => x"88",
          3598 => x"55",
          3599 => x"1a",
          3600 => x"82",
          3601 => x"2b",
          3602 => x"2b",
          3603 => x"05",
          3604 => x"fc",
          3605 => x"1c",
          3606 => x"5f",
          3607 => x"54",
          3608 => x"0d",
          3609 => x"fc",
          3610 => x"23",
          3611 => x"ff",
          3612 => x"b9",
          3613 => x"0b",
          3614 => x"5d",
          3615 => x"1e",
          3616 => x"86",
          3617 => x"84",
          3618 => x"ff",
          3619 => x"ff",
          3620 => x"5b",
          3621 => x"18",
          3622 => x"10",
          3623 => x"05",
          3624 => x"0b",
          3625 => x"57",
          3626 => x"82",
          3627 => x"fe",
          3628 => x"84",
          3629 => x"95",
          3630 => x"fc",
          3631 => x"44",
          3632 => x"71",
          3633 => x"70",
          3634 => x"63",
          3635 => x"84",
          3636 => x"57",
          3637 => x"19",
          3638 => x"70",
          3639 => x"07",
          3640 => x"74",
          3641 => x"88",
          3642 => x"5d",
          3643 => x"ff",
          3644 => x"84",
          3645 => x"34",
          3646 => x"fc",
          3647 => x"3f",
          3648 => x"31",
          3649 => x"fa",
          3650 => x"76",
          3651 => x"17",
          3652 => x"07",
          3653 => x"81",
          3654 => x"2b",
          3655 => x"45",
          3656 => x"ff",
          3657 => x"38",
          3658 => x"83",
          3659 => x"fc",
          3660 => x"f4",
          3661 => x"0b",
          3662 => x"53",
          3663 => x"c4",
          3664 => x"7e",
          3665 => x"84",
          3666 => x"34",
          3667 => x"fc",
          3668 => x"0b",
          3669 => x"84",
          3670 => x"80",
          3671 => x"88",
          3672 => x"88",
          3673 => x"84",
          3674 => x"84",
          3675 => x"43",
          3676 => x"83",
          3677 => x"24",
          3678 => x"06",
          3679 => x"fc",
          3680 => x"38",
          3681 => x"73",
          3682 => x"04",
          3683 => x"33",
          3684 => x"7a",
          3685 => x"71",
          3686 => x"05",
          3687 => x"88",
          3688 => x"45",
          3689 => x"56",
          3690 => x"85",
          3691 => x"17",
          3692 => x"8b",
          3693 => x"86",
          3694 => x"2b",
          3695 => x"48",
          3696 => x"05",
          3697 => x"b9",
          3698 => x"33",
          3699 => x"06",
          3700 => x"7b",
          3701 => x"b9",
          3702 => x"83",
          3703 => x"2b",
          3704 => x"33",
          3705 => x"5e",
          3706 => x"76",
          3707 => x"b9",
          3708 => x"12",
          3709 => x"07",
          3710 => x"33",
          3711 => x"40",
          3712 => x"78",
          3713 => x"84",
          3714 => x"33",
          3715 => x"66",
          3716 => x"52",
          3717 => x"fe",
          3718 => x"1e",
          3719 => x"5c",
          3720 => x"0b",
          3721 => x"84",
          3722 => x"7f",
          3723 => x"a4",
          3724 => x"76",
          3725 => x"b9",
          3726 => x"81",
          3727 => x"08",
          3728 => x"87",
          3729 => x"b9",
          3730 => x"07",
          3731 => x"2a",
          3732 => x"34",
          3733 => x"22",
          3734 => x"08",
          3735 => x"1c",
          3736 => x"51",
          3737 => x"39",
          3738 => x"8b",
          3739 => x"84",
          3740 => x"2b",
          3741 => x"43",
          3742 => x"63",
          3743 => x"08",
          3744 => x"33",
          3745 => x"74",
          3746 => x"71",
          3747 => x"5f",
          3748 => x"64",
          3749 => x"34",
          3750 => x"81",
          3751 => x"ff",
          3752 => x"58",
          3753 => x"34",
          3754 => x"33",
          3755 => x"83",
          3756 => x"12",
          3757 => x"2b",
          3758 => x"88",
          3759 => x"5d",
          3760 => x"83",
          3761 => x"1f",
          3762 => x"2b",
          3763 => x"33",
          3764 => x"81",
          3765 => x"5d",
          3766 => x"60",
          3767 => x"83",
          3768 => x"86",
          3769 => x"2b",
          3770 => x"18",
          3771 => x"07",
          3772 => x"41",
          3773 => x"1e",
          3774 => x"84",
          3775 => x"2b",
          3776 => x"14",
          3777 => x"07",
          3778 => x"5a",
          3779 => x"34",
          3780 => x"fc",
          3781 => x"71",
          3782 => x"70",
          3783 => x"75",
          3784 => x"fc",
          3785 => x"33",
          3786 => x"74",
          3787 => x"88",
          3788 => x"f8",
          3789 => x"54",
          3790 => x"7f",
          3791 => x"84",
          3792 => x"81",
          3793 => x"2b",
          3794 => x"33",
          3795 => x"06",
          3796 => x"5b",
          3797 => x"81",
          3798 => x"1f",
          3799 => x"8b",
          3800 => x"86",
          3801 => x"2b",
          3802 => x"14",
          3803 => x"07",
          3804 => x"5c",
          3805 => x"77",
          3806 => x"84",
          3807 => x"33",
          3808 => x"83",
          3809 => x"87",
          3810 => x"88",
          3811 => x"41",
          3812 => x"16",
          3813 => x"33",
          3814 => x"81",
          3815 => x"5c",
          3816 => x"1a",
          3817 => x"82",
          3818 => x"2b",
          3819 => x"33",
          3820 => x"70",
          3821 => x"5a",
          3822 => x"1a",
          3823 => x"70",
          3824 => x"71",
          3825 => x"33",
          3826 => x"70",
          3827 => x"5a",
          3828 => x"83",
          3829 => x"1f",
          3830 => x"88",
          3831 => x"83",
          3832 => x"84",
          3833 => x"b9",
          3834 => x"05",
          3835 => x"44",
          3836 => x"87",
          3837 => x"2b",
          3838 => x"1d",
          3839 => x"2a",
          3840 => x"61",
          3841 => x"34",
          3842 => x"11",
          3843 => x"71",
          3844 => x"33",
          3845 => x"70",
          3846 => x"59",
          3847 => x"7a",
          3848 => x"08",
          3849 => x"88",
          3850 => x"88",
          3851 => x"34",
          3852 => x"08",
          3853 => x"71",
          3854 => x"05",
          3855 => x"2b",
          3856 => x"06",
          3857 => x"5c",
          3858 => x"82",
          3859 => x"b9",
          3860 => x"12",
          3861 => x"07",
          3862 => x"71",
          3863 => x"70",
          3864 => x"59",
          3865 => x"1e",
          3866 => x"f3",
          3867 => x"a1",
          3868 => x"ba",
          3869 => x"53",
          3870 => x"fe",
          3871 => x"3f",
          3872 => x"38",
          3873 => x"7a",
          3874 => x"76",
          3875 => x"8a",
          3876 => x"3d",
          3877 => x"84",
          3878 => x"08",
          3879 => x"52",
          3880 => x"bc",
          3881 => x"3d",
          3882 => x"b9",
          3883 => x"f8",
          3884 => x"84",
          3885 => x"84",
          3886 => x"81",
          3887 => x"08",
          3888 => x"85",
          3889 => x"76",
          3890 => x"34",
          3891 => x"22",
          3892 => x"83",
          3893 => x"51",
          3894 => x"89",
          3895 => x"10",
          3896 => x"f8",
          3897 => x"81",
          3898 => x"80",
          3899 => x"ff",
          3900 => x"81",
          3901 => x"ba",
          3902 => x"8c",
          3903 => x"0d",
          3904 => x"71",
          3905 => x"ec",
          3906 => x"06",
          3907 => x"88",
          3908 => x"53",
          3909 => x"0d",
          3910 => x"02",
          3911 => x"57",
          3912 => x"38",
          3913 => x"81",
          3914 => x"73",
          3915 => x"0c",
          3916 => x"8d",
          3917 => x"06",
          3918 => x"c0",
          3919 => x"79",
          3920 => x"80",
          3921 => x"81",
          3922 => x"0c",
          3923 => x"81",
          3924 => x"56",
          3925 => x"39",
          3926 => x"8c",
          3927 => x"59",
          3928 => x"84",
          3929 => x"06",
          3930 => x"58",
          3931 => x"78",
          3932 => x"3f",
          3933 => x"55",
          3934 => x"98",
          3935 => x"78",
          3936 => x"06",
          3937 => x"54",
          3938 => x"8b",
          3939 => x"19",
          3940 => x"79",
          3941 => x"fc",
          3942 => x"05",
          3943 => x"53",
          3944 => x"87",
          3945 => x"72",
          3946 => x"38",
          3947 => x"81",
          3948 => x"71",
          3949 => x"38",
          3950 => x"86",
          3951 => x"0c",
          3952 => x"0d",
          3953 => x"84",
          3954 => x"71",
          3955 => x"53",
          3956 => x"81",
          3957 => x"2e",
          3958 => x"55",
          3959 => x"08",
          3960 => x"87",
          3961 => x"82",
          3962 => x"38",
          3963 => x"38",
          3964 => x"58",
          3965 => x"56",
          3966 => x"a8",
          3967 => x"81",
          3968 => x"18",
          3969 => x"8c",
          3970 => x"78",
          3971 => x"04",
          3972 => x"18",
          3973 => x"fc",
          3974 => x"08",
          3975 => x"84",
          3976 => x"18",
          3977 => x"1a",
          3978 => x"56",
          3979 => x"82",
          3980 => x"81",
          3981 => x"1b",
          3982 => x"fc",
          3983 => x"75",
          3984 => x"38",
          3985 => x"09",
          3986 => x"5a",
          3987 => x"70",
          3988 => x"76",
          3989 => x"19",
          3990 => x"34",
          3991 => x"b9",
          3992 => x"34",
          3993 => x"f2",
          3994 => x"0b",
          3995 => x"84",
          3996 => x"9f",
          3997 => x"84",
          3998 => x"7a",
          3999 => x"56",
          4000 => x"2a",
          4001 => x"18",
          4002 => x"7a",
          4003 => x"34",
          4004 => x"19",
          4005 => x"a7",
          4006 => x"70",
          4007 => x"53",
          4008 => x"e8",
          4009 => x"80",
          4010 => x"3f",
          4011 => x"b7",
          4012 => x"60",
          4013 => x"76",
          4014 => x"26",
          4015 => x"8c",
          4016 => x"33",
          4017 => x"38",
          4018 => x"81",
          4019 => x"81",
          4020 => x"08",
          4021 => x"08",
          4022 => x"5c",
          4023 => x"de",
          4024 => x"52",
          4025 => x"84",
          4026 => x"ff",
          4027 => x"7a",
          4028 => x"17",
          4029 => x"2a",
          4030 => x"59",
          4031 => x"80",
          4032 => x"5d",
          4033 => x"b5",
          4034 => x"52",
          4035 => x"84",
          4036 => x"ff",
          4037 => x"79",
          4038 => x"17",
          4039 => x"07",
          4040 => x"5d",
          4041 => x"76",
          4042 => x"8f",
          4043 => x"18",
          4044 => x"2e",
          4045 => x"71",
          4046 => x"81",
          4047 => x"53",
          4048 => x"f7",
          4049 => x"2e",
          4050 => x"b4",
          4051 => x"10",
          4052 => x"81",
          4053 => x"07",
          4054 => x"3d",
          4055 => x"06",
          4056 => x"18",
          4057 => x"2e",
          4058 => x"71",
          4059 => x"81",
          4060 => x"53",
          4061 => x"f6",
          4062 => x"2e",
          4063 => x"b4",
          4064 => x"82",
          4065 => x"05",
          4066 => x"90",
          4067 => x"33",
          4068 => x"71",
          4069 => x"84",
          4070 => x"5a",
          4071 => x"b4",
          4072 => x"81",
          4073 => x"81",
          4074 => x"09",
          4075 => x"8c",
          4076 => x"a8",
          4077 => x"5b",
          4078 => x"84",
          4079 => x"2e",
          4080 => x"54",
          4081 => x"53",
          4082 => x"98",
          4083 => x"54",
          4084 => x"53",
          4085 => x"3f",
          4086 => x"81",
          4087 => x"08",
          4088 => x"18",
          4089 => x"27",
          4090 => x"82",
          4091 => x"08",
          4092 => x"17",
          4093 => x"18",
          4094 => x"5a",
          4095 => x"81",
          4096 => x"08",
          4097 => x"18",
          4098 => x"5e",
          4099 => x"38",
          4100 => x"09",
          4101 => x"b4",
          4102 => x"7b",
          4103 => x"3f",
          4104 => x"b4",
          4105 => x"81",
          4106 => x"81",
          4107 => x"09",
          4108 => x"8c",
          4109 => x"a8",
          4110 => x"5b",
          4111 => x"91",
          4112 => x"2e",
          4113 => x"54",
          4114 => x"53",
          4115 => x"90",
          4116 => x"54",
          4117 => x"53",
          4118 => x"f8",
          4119 => x"f9",
          4120 => x"0d",
          4121 => x"58",
          4122 => x"1a",
          4123 => x"74",
          4124 => x"81",
          4125 => x"38",
          4126 => x"0d",
          4127 => x"05",
          4128 => x"5c",
          4129 => x"19",
          4130 => x"09",
          4131 => x"77",
          4132 => x"51",
          4133 => x"80",
          4134 => x"77",
          4135 => x"b0",
          4136 => x"05",
          4137 => x"76",
          4138 => x"79",
          4139 => x"34",
          4140 => x"0d",
          4141 => x"fe",
          4142 => x"08",
          4143 => x"58",
          4144 => x"83",
          4145 => x"2e",
          4146 => x"54",
          4147 => x"33",
          4148 => x"08",
          4149 => x"5a",
          4150 => x"fe",
          4151 => x"06",
          4152 => x"70",
          4153 => x"0a",
          4154 => x"7d",
          4155 => x"1d",
          4156 => x"1d",
          4157 => x"1d",
          4158 => x"e8",
          4159 => x"2a",
          4160 => x"59",
          4161 => x"80",
          4162 => x"5d",
          4163 => x"d4",
          4164 => x"52",
          4165 => x"84",
          4166 => x"ff",
          4167 => x"7b",
          4168 => x"ff",
          4169 => x"81",
          4170 => x"80",
          4171 => x"f0",
          4172 => x"56",
          4173 => x"1a",
          4174 => x"05",
          4175 => x"5f",
          4176 => x"54",
          4177 => x"1a",
          4178 => x"58",
          4179 => x"81",
          4180 => x"08",
          4181 => x"a8",
          4182 => x"ba",
          4183 => x"7a",
          4184 => x"74",
          4185 => x"75",
          4186 => x"ee",
          4187 => x"2e",
          4188 => x"b4",
          4189 => x"83",
          4190 => x"2a",
          4191 => x"2a",
          4192 => x"06",
          4193 => x"0b",
          4194 => x"54",
          4195 => x"1a",
          4196 => x"5a",
          4197 => x"81",
          4198 => x"08",
          4199 => x"a8",
          4200 => x"ba",
          4201 => x"77",
          4202 => x"55",
          4203 => x"bd",
          4204 => x"52",
          4205 => x"7b",
          4206 => x"53",
          4207 => x"52",
          4208 => x"ba",
          4209 => x"fd",
          4210 => x"1a",
          4211 => x"08",
          4212 => x"08",
          4213 => x"fc",
          4214 => x"82",
          4215 => x"81",
          4216 => x"19",
          4217 => x"fc",
          4218 => x"19",
          4219 => x"ed",
          4220 => x"08",
          4221 => x"38",
          4222 => x"b4",
          4223 => x"a0",
          4224 => x"5f",
          4225 => x"38",
          4226 => x"09",
          4227 => x"7c",
          4228 => x"51",
          4229 => x"39",
          4230 => x"81",
          4231 => x"58",
          4232 => x"fe",
          4233 => x"06",
          4234 => x"76",
          4235 => x"f9",
          4236 => x"7b",
          4237 => x"05",
          4238 => x"2b",
          4239 => x"07",
          4240 => x"34",
          4241 => x"34",
          4242 => x"34",
          4243 => x"34",
          4244 => x"7e",
          4245 => x"8a",
          4246 => x"2e",
          4247 => x"27",
          4248 => x"56",
          4249 => x"76",
          4250 => x"81",
          4251 => x"89",
          4252 => x"b2",
          4253 => x"3f",
          4254 => x"d0",
          4255 => x"81",
          4256 => x"09",
          4257 => x"70",
          4258 => x"82",
          4259 => x"06",
          4260 => x"ba",
          4261 => x"57",
          4262 => x"58",
          4263 => x"a4",
          4264 => x"08",
          4265 => x"55",
          4266 => x"38",
          4267 => x"26",
          4268 => x"81",
          4269 => x"83",
          4270 => x"ef",
          4271 => x"08",
          4272 => x"8c",
          4273 => x"80",
          4274 => x"08",
          4275 => x"85",
          4276 => x"9a",
          4277 => x"27",
          4278 => x"27",
          4279 => x"fe",
          4280 => x"38",
          4281 => x"f5",
          4282 => x"8c",
          4283 => x"07",
          4284 => x"c4",
          4285 => x"1a",
          4286 => x"1a",
          4287 => x"38",
          4288 => x"33",
          4289 => x"75",
          4290 => x"3d",
          4291 => x"0c",
          4292 => x"08",
          4293 => x"ff",
          4294 => x"51",
          4295 => x"55",
          4296 => x"84",
          4297 => x"ff",
          4298 => x"81",
          4299 => x"7a",
          4300 => x"f0",
          4301 => x"9f",
          4302 => x"90",
          4303 => x"80",
          4304 => x"26",
          4305 => x"82",
          4306 => x"79",
          4307 => x"19",
          4308 => x"08",
          4309 => x"38",
          4310 => x"73",
          4311 => x"19",
          4312 => x"0c",
          4313 => x"ba",
          4314 => x"17",
          4315 => x"38",
          4316 => x"59",
          4317 => x"08",
          4318 => x"80",
          4319 => x"17",
          4320 => x"05",
          4321 => x"91",
          4322 => x"3f",
          4323 => x"8c",
          4324 => x"84",
          4325 => x"9c",
          4326 => x"73",
          4327 => x"54",
          4328 => x"39",
          4329 => x"3d",
          4330 => x"08",
          4331 => x"57",
          4332 => x"80",
          4333 => x"55",
          4334 => x"79",
          4335 => x"81",
          4336 => x"a9",
          4337 => x"57",
          4338 => x"77",
          4339 => x"78",
          4340 => x"56",
          4341 => x"0d",
          4342 => x"22",
          4343 => x"7b",
          4344 => x"9c",
          4345 => x"56",
          4346 => x"d0",
          4347 => x"ff",
          4348 => x"ba",
          4349 => x"80",
          4350 => x"52",
          4351 => x"8c",
          4352 => x"08",
          4353 => x"84",
          4354 => x"38",
          4355 => x"2e",
          4356 => x"83",
          4357 => x"38",
          4358 => x"59",
          4359 => x"38",
          4360 => x"1b",
          4361 => x"0c",
          4362 => x"55",
          4363 => x"ff",
          4364 => x"8a",
          4365 => x"80",
          4366 => x"52",
          4367 => x"84",
          4368 => x"16",
          4369 => x"84",
          4370 => x"0d",
          4371 => x"b8",
          4372 => x"56",
          4373 => x"80",
          4374 => x"1a",
          4375 => x"31",
          4376 => x"e8",
          4377 => x"2e",
          4378 => x"54",
          4379 => x"53",
          4380 => x"c8",
          4381 => x"55",
          4382 => x"76",
          4383 => x"94",
          4384 => x"fe",
          4385 => x"27",
          4386 => x"71",
          4387 => x"0c",
          4388 => x"ba",
          4389 => x"3d",
          4390 => x"08",
          4391 => x"08",
          4392 => x"d2",
          4393 => x"58",
          4394 => x"38",
          4395 => x"78",
          4396 => x"81",
          4397 => x"19",
          4398 => x"8c",
          4399 => x"81",
          4400 => x"76",
          4401 => x"33",
          4402 => x"38",
          4403 => x"ff",
          4404 => x"76",
          4405 => x"32",
          4406 => x"25",
          4407 => x"93",
          4408 => x"61",
          4409 => x"2e",
          4410 => x"52",
          4411 => x"8c",
          4412 => x"b2",
          4413 => x"dc",
          4414 => x"3d",
          4415 => x"53",
          4416 => x"a8",
          4417 => x"78",
          4418 => x"84",
          4419 => x"19",
          4420 => x"8c",
          4421 => x"27",
          4422 => x"60",
          4423 => x"38",
          4424 => x"08",
          4425 => x"51",
          4426 => x"39",
          4427 => x"e7",
          4428 => x"7a",
          4429 => x"77",
          4430 => x"7f",
          4431 => x"7d",
          4432 => x"5d",
          4433 => x"2e",
          4434 => x"39",
          4435 => x"7a",
          4436 => x"04",
          4437 => x"33",
          4438 => x"cb",
          4439 => x"9a",
          4440 => x"56",
          4441 => x"70",
          4442 => x"51",
          4443 => x"8c",
          4444 => x"71",
          4445 => x"56",
          4446 => x"81",
          4447 => x"61",
          4448 => x"81",
          4449 => x"27",
          4450 => x"81",
          4451 => x"38",
          4452 => x"79",
          4453 => x"ff",
          4454 => x"fd",
          4455 => x"ca",
          4456 => x"7c",
          4457 => x"81",
          4458 => x"70",
          4459 => x"70",
          4460 => x"59",
          4461 => x"81",
          4462 => x"84",
          4463 => x"ef",
          4464 => x"80",
          4465 => x"ba",
          4466 => x"82",
          4467 => x"ff",
          4468 => x"98",
          4469 => x"08",
          4470 => x"33",
          4471 => x"81",
          4472 => x"53",
          4473 => x"dc",
          4474 => x"2e",
          4475 => x"b4",
          4476 => x"38",
          4477 => x"76",
          4478 => x"33",
          4479 => x"58",
          4480 => x"2e",
          4481 => x"06",
          4482 => x"74",
          4483 => x"e5",
          4484 => x"58",
          4485 => x"80",
          4486 => x"33",
          4487 => x"ff",
          4488 => x"74",
          4489 => x"33",
          4490 => x"0b",
          4491 => x"05",
          4492 => x"33",
          4493 => x"42",
          4494 => x"75",
          4495 => x"ff",
          4496 => x"51",
          4497 => x"5a",
          4498 => x"8f",
          4499 => x"3d",
          4500 => x"53",
          4501 => x"80",
          4502 => x"78",
          4503 => x"84",
          4504 => x"1b",
          4505 => x"8c",
          4506 => x"27",
          4507 => x"79",
          4508 => x"38",
          4509 => x"08",
          4510 => x"51",
          4511 => x"39",
          4512 => x"33",
          4513 => x"60",
          4514 => x"06",
          4515 => x"19",
          4516 => x"1f",
          4517 => x"5f",
          4518 => x"55",
          4519 => x"92",
          4520 => x"ba",
          4521 => x"fe",
          4522 => x"38",
          4523 => x"0c",
          4524 => x"7e",
          4525 => x"8c",
          4526 => x"33",
          4527 => x"76",
          4528 => x"06",
          4529 => x"77",
          4530 => x"79",
          4531 => x"88",
          4532 => x"2e",
          4533 => x"ff",
          4534 => x"3f",
          4535 => x"05",
          4536 => x"56",
          4537 => x"8c",
          4538 => x"38",
          4539 => x"27",
          4540 => x"2a",
          4541 => x"92",
          4542 => x"10",
          4543 => x"fe",
          4544 => x"06",
          4545 => x"84",
          4546 => x"76",
          4547 => x"81",
          4548 => x"0d",
          4549 => x"81",
          4550 => x"56",
          4551 => x"08",
          4552 => x"2e",
          4553 => x"70",
          4554 => x"95",
          4555 => x"7b",
          4556 => x"57",
          4557 => x"ff",
          4558 => x"db",
          4559 => x"76",
          4560 => x"0b",
          4561 => x"40",
          4562 => x"8b",
          4563 => x"81",
          4564 => x"58",
          4565 => x"85",
          4566 => x"22",
          4567 => x"74",
          4568 => x"81",
          4569 => x"70",
          4570 => x"81",
          4571 => x"2e",
          4572 => x"57",
          4573 => x"38",
          4574 => x"02",
          4575 => x"76",
          4576 => x"27",
          4577 => x"34",
          4578 => x"59",
          4579 => x"59",
          4580 => x"56",
          4581 => x"55",
          4582 => x"56",
          4583 => x"1a",
          4584 => x"09",
          4585 => x"a0",
          4586 => x"3d",
          4587 => x"33",
          4588 => x"76",
          4589 => x"8f",
          4590 => x"81",
          4591 => x"91",
          4592 => x"82",
          4593 => x"84",
          4594 => x"06",
          4595 => x"33",
          4596 => x"05",
          4597 => x"81",
          4598 => x"80",
          4599 => x"51",
          4600 => x"08",
          4601 => x"8c",
          4602 => x"ba",
          4603 => x"8c",
          4604 => x"08",
          4605 => x"2e",
          4606 => x"7f",
          4607 => x"38",
          4608 => x"81",
          4609 => x"ba",
          4610 => x"56",
          4611 => x"56",
          4612 => x"33",
          4613 => x"c9",
          4614 => x"07",
          4615 => x"38",
          4616 => x"89",
          4617 => x"3f",
          4618 => x"8c",
          4619 => x"58",
          4620 => x"58",
          4621 => x"7f",
          4622 => x"b4",
          4623 => x"1c",
          4624 => x"38",
          4625 => x"81",
          4626 => x"ba",
          4627 => x"57",
          4628 => x"58",
          4629 => x"1f",
          4630 => x"05",
          4631 => x"38",
          4632 => x"58",
          4633 => x"77",
          4634 => x"55",
          4635 => x"1f",
          4636 => x"1b",
          4637 => x"56",
          4638 => x"0d",
          4639 => x"72",
          4640 => x"38",
          4641 => x"c2",
          4642 => x"ba",
          4643 => x"fe",
          4644 => x"53",
          4645 => x"80",
          4646 => x"09",
          4647 => x"8c",
          4648 => x"a8",
          4649 => x"08",
          4650 => x"60",
          4651 => x"8c",
          4652 => x"2b",
          4653 => x"7d",
          4654 => x"08",
          4655 => x"38",
          4656 => x"8b",
          4657 => x"29",
          4658 => x"57",
          4659 => x"19",
          4660 => x"81",
          4661 => x"1e",
          4662 => x"77",
          4663 => x"7a",
          4664 => x"38",
          4665 => x"81",
          4666 => x"ba",
          4667 => x"57",
          4668 => x"58",
          4669 => x"9c",
          4670 => x"5c",
          4671 => x"8b",
          4672 => x"9a",
          4673 => x"8d",
          4674 => x"59",
          4675 => x"78",
          4676 => x"58",
          4677 => x"05",
          4678 => x"34",
          4679 => x"76",
          4680 => x"18",
          4681 => x"83",
          4682 => x"10",
          4683 => x"2e",
          4684 => x"0b",
          4685 => x"e9",
          4686 => x"84",
          4687 => x"ff",
          4688 => x"eb",
          4689 => x"b8",
          4690 => x"59",
          4691 => x"8c",
          4692 => x"08",
          4693 => x"1d",
          4694 => x"41",
          4695 => x"38",
          4696 => x"09",
          4697 => x"b4",
          4698 => x"78",
          4699 => x"3f",
          4700 => x"1f",
          4701 => x"81",
          4702 => x"38",
          4703 => x"76",
          4704 => x"39",
          4705 => x"39",
          4706 => x"52",
          4707 => x"84",
          4708 => x"06",
          4709 => x"1d",
          4710 => x"31",
          4711 => x"38",
          4712 => x"aa",
          4713 => x"f8",
          4714 => x"80",
          4715 => x"75",
          4716 => x"59",
          4717 => x"fa",
          4718 => x"a0",
          4719 => x"1c",
          4720 => x"39",
          4721 => x"08",
          4722 => x"51",
          4723 => x"3d",
          4724 => x"5c",
          4725 => x"08",
          4726 => x"08",
          4727 => x"71",
          4728 => x"58",
          4729 => x"38",
          4730 => x"1b",
          4731 => x"80",
          4732 => x"06",
          4733 => x"83",
          4734 => x"22",
          4735 => x"7a",
          4736 => x"06",
          4737 => x"57",
          4738 => x"89",
          4739 => x"16",
          4740 => x"74",
          4741 => x"81",
          4742 => x"70",
          4743 => x"77",
          4744 => x"8b",
          4745 => x"34",
          4746 => x"05",
          4747 => x"27",
          4748 => x"55",
          4749 => x"33",
          4750 => x"38",
          4751 => x"7c",
          4752 => x"17",
          4753 => x"55",
          4754 => x"34",
          4755 => x"88",
          4756 => x"83",
          4757 => x"2b",
          4758 => x"70",
          4759 => x"07",
          4760 => x"17",
          4761 => x"5b",
          4762 => x"1e",
          4763 => x"71",
          4764 => x"1e",
          4765 => x"55",
          4766 => x"81",
          4767 => x"b5",
          4768 => x"81",
          4769 => x"83",
          4770 => x"27",
          4771 => x"38",
          4772 => x"74",
          4773 => x"80",
          4774 => x"19",
          4775 => x"79",
          4776 => x"30",
          4777 => x"72",
          4778 => x"80",
          4779 => x"05",
          4780 => x"5b",
          4781 => x"5a",
          4782 => x"38",
          4783 => x"89",
          4784 => x"78",
          4785 => x"8c",
          4786 => x"b4",
          4787 => x"06",
          4788 => x"14",
          4789 => x"73",
          4790 => x"16",
          4791 => x"33",
          4792 => x"b7",
          4793 => x"53",
          4794 => x"25",
          4795 => x"58",
          4796 => x"70",
          4797 => x"70",
          4798 => x"83",
          4799 => x"81",
          4800 => x"38",
          4801 => x"33",
          4802 => x"9f",
          4803 => x"8c",
          4804 => x"70",
          4805 => x"81",
          4806 => x"2e",
          4807 => x"27",
          4808 => x"76",
          4809 => x"ff",
          4810 => x"73",
          4811 => x"5b",
          4812 => x"dc",
          4813 => x"26",
          4814 => x"e5",
          4815 => x"54",
          4816 => x"73",
          4817 => x"33",
          4818 => x"73",
          4819 => x"7a",
          4820 => x"80",
          4821 => x"7d",
          4822 => x"05",
          4823 => x"2e",
          4824 => x"73",
          4825 => x"25",
          4826 => x"80",
          4827 => x"54",
          4828 => x"2e",
          4829 => x"30",
          4830 => x"57",
          4831 => x"73",
          4832 => x"55",
          4833 => x"39",
          4834 => x"e7",
          4835 => x"ff",
          4836 => x"54",
          4837 => x"0d",
          4838 => x"ff",
          4839 => x"e3",
          4840 => x"1d",
          4841 => x"3f",
          4842 => x"0c",
          4843 => x"dc",
          4844 => x"07",
          4845 => x"a1",
          4846 => x"33",
          4847 => x"38",
          4848 => x"80",
          4849 => x"e1",
          4850 => x"82",
          4851 => x"38",
          4852 => x"17",
          4853 => x"17",
          4854 => x"a0",
          4855 => x"42",
          4856 => x"84",
          4857 => x"76",
          4858 => x"80",
          4859 => x"38",
          4860 => x"06",
          4861 => x"2e",
          4862 => x"06",
          4863 => x"76",
          4864 => x"05",
          4865 => x"9d",
          4866 => x"ff",
          4867 => x"fe",
          4868 => x"2e",
          4869 => x"a0",
          4870 => x"05",
          4871 => x"38",
          4872 => x"70",
          4873 => x"74",
          4874 => x"2e",
          4875 => x"30",
          4876 => x"77",
          4877 => x"38",
          4878 => x"81",
          4879 => x"72",
          4880 => x"51",
          4881 => x"38",
          4882 => x"77",
          4883 => x"75",
          4884 => x"5b",
          4885 => x"77",
          4886 => x"22",
          4887 => x"95",
          4888 => x"e5",
          4889 => x"82",
          4890 => x"8c",
          4891 => x"55",
          4892 => x"81",
          4893 => x"7d",
          4894 => x"38",
          4895 => x"81",
          4896 => x"79",
          4897 => x"7b",
          4898 => x"08",
          4899 => x"8c",
          4900 => x"ba",
          4901 => x"fb",
          4902 => x"5a",
          4903 => x"82",
          4904 => x"38",
          4905 => x"8c",
          4906 => x"39",
          4907 => x"22",
          4908 => x"f0",
          4909 => x"79",
          4910 => x"18",
          4911 => x"06",
          4912 => x"ae",
          4913 => x"76",
          4914 => x"0b",
          4915 => x"73",
          4916 => x"70",
          4917 => x"8a",
          4918 => x"58",
          4919 => x"bf",
          4920 => x"33",
          4921 => x"d6",
          4922 => x"77",
          4923 => x"84",
          4924 => x"2e",
          4925 => x"ff",
          4926 => x"80",
          4927 => x"62",
          4928 => x"2e",
          4929 => x"7b",
          4930 => x"77",
          4931 => x"38",
          4932 => x"fb",
          4933 => x"56",
          4934 => x"81",
          4935 => x"77",
          4936 => x"38",
          4937 => x"85",
          4938 => x"09",
          4939 => x"ff",
          4940 => x"84",
          4941 => x"74",
          4942 => x"75",
          4943 => x"78",
          4944 => x"07",
          4945 => x"a4",
          4946 => x"52",
          4947 => x"ba",
          4948 => x"87",
          4949 => x"2e",
          4950 => x"e6",
          4951 => x"ff",
          4952 => x"81",
          4953 => x"e5",
          4954 => x"54",
          4955 => x"73",
          4956 => x"33",
          4957 => x"73",
          4958 => x"78",
          4959 => x"73",
          4960 => x"70",
          4961 => x"15",
          4962 => x"81",
          4963 => x"70",
          4964 => x"53",
          4965 => x"34",
          4966 => x"fc",
          4967 => x"e5",
          4968 => x"53",
          4969 => x"df",
          4970 => x"5b",
          4971 => x"5b",
          4972 => x"cc",
          4973 => x"2b",
          4974 => x"57",
          4975 => x"75",
          4976 => x"81",
          4977 => x"74",
          4978 => x"39",
          4979 => x"5a",
          4980 => x"fa",
          4981 => x"2a",
          4982 => x"85",
          4983 => x"0d",
          4984 => x"88",
          4985 => x"5e",
          4986 => x"59",
          4987 => x"38",
          4988 => x"9f",
          4989 => x"d0",
          4990 => x"85",
          4991 => x"80",
          4992 => x"10",
          4993 => x"5a",
          4994 => x"38",
          4995 => x"77",
          4996 => x"38",
          4997 => x"3f",
          4998 => x"70",
          4999 => x"86",
          5000 => x"5d",
          5001 => x"34",
          5002 => x"bb",
          5003 => x"ff",
          5004 => x"58",
          5005 => x"8d",
          5006 => x"8a",
          5007 => x"7a",
          5008 => x"0c",
          5009 => x"53",
          5010 => x"52",
          5011 => x"8c",
          5012 => x"81",
          5013 => x"78",
          5014 => x"b6",
          5015 => x"56",
          5016 => x"85",
          5017 => x"84",
          5018 => x"bf",
          5019 => x"cd",
          5020 => x"c5",
          5021 => x"18",
          5022 => x"7c",
          5023 => x"ad",
          5024 => x"18",
          5025 => x"75",
          5026 => x"33",
          5027 => x"88",
          5028 => x"07",
          5029 => x"5a",
          5030 => x"18",
          5031 => x"34",
          5032 => x"81",
          5033 => x"7c",
          5034 => x"ff",
          5035 => x"33",
          5036 => x"77",
          5037 => x"ff",
          5038 => x"38",
          5039 => x"33",
          5040 => x"88",
          5041 => x"5a",
          5042 => x"cc",
          5043 => x"88",
          5044 => x"80",
          5045 => x"33",
          5046 => x"81",
          5047 => x"75",
          5048 => x"42",
          5049 => x"c6",
          5050 => x"58",
          5051 => x"38",
          5052 => x"79",
          5053 => x"74",
          5054 => x"84",
          5055 => x"08",
          5056 => x"8c",
          5057 => x"83",
          5058 => x"26",
          5059 => x"26",
          5060 => x"70",
          5061 => x"7b",
          5062 => x"b0",
          5063 => x"8a",
          5064 => x"58",
          5065 => x"16",
          5066 => x"82",
          5067 => x"81",
          5068 => x"83",
          5069 => x"78",
          5070 => x"0b",
          5071 => x"0c",
          5072 => x"83",
          5073 => x"84",
          5074 => x"84",
          5075 => x"84",
          5076 => x"0b",
          5077 => x"ba",
          5078 => x"0b",
          5079 => x"04",
          5080 => x"06",
          5081 => x"38",
          5082 => x"05",
          5083 => x"38",
          5084 => x"40",
          5085 => x"70",
          5086 => x"05",
          5087 => x"56",
          5088 => x"70",
          5089 => x"17",
          5090 => x"17",
          5091 => x"30",
          5092 => x"2e",
          5093 => x"be",
          5094 => x"72",
          5095 => x"55",
          5096 => x"1c",
          5097 => x"ff",
          5098 => x"78",
          5099 => x"2a",
          5100 => x"c5",
          5101 => x"78",
          5102 => x"09",
          5103 => x"81",
          5104 => x"7b",
          5105 => x"38",
          5106 => x"93",
          5107 => x"fa",
          5108 => x"2e",
          5109 => x"80",
          5110 => x"2b",
          5111 => x"07",
          5112 => x"07",
          5113 => x"7a",
          5114 => x"90",
          5115 => x"be",
          5116 => x"30",
          5117 => x"3d",
          5118 => x"b6",
          5119 => x"78",
          5120 => x"80",
          5121 => x"ff",
          5122 => x"56",
          5123 => x"7a",
          5124 => x"51",
          5125 => x"08",
          5126 => x"56",
          5127 => x"bf",
          5128 => x"88",
          5129 => x"82",
          5130 => x"38",
          5131 => x"75",
          5132 => x"81",
          5133 => x"7a",
          5134 => x"75",
          5135 => x"77",
          5136 => x"ba",
          5137 => x"2e",
          5138 => x"81",
          5139 => x"2e",
          5140 => x"5a",
          5141 => x"f8",
          5142 => x"83",
          5143 => x"81",
          5144 => x"40",
          5145 => x"52",
          5146 => x"38",
          5147 => x"81",
          5148 => x"58",
          5149 => x"70",
          5150 => x"ff",
          5151 => x"2e",
          5152 => x"38",
          5153 => x"7c",
          5154 => x"0c",
          5155 => x"80",
          5156 => x"8a",
          5157 => x"ff",
          5158 => x"0c",
          5159 => x"ee",
          5160 => x"78",
          5161 => x"81",
          5162 => x"1b",
          5163 => x"83",
          5164 => x"85",
          5165 => x"5c",
          5166 => x"33",
          5167 => x"71",
          5168 => x"77",
          5169 => x"2e",
          5170 => x"83",
          5171 => x"c6",
          5172 => x"18",
          5173 => x"75",
          5174 => x"38",
          5175 => x"08",
          5176 => x"5b",
          5177 => x"9b",
          5178 => x"52",
          5179 => x"3f",
          5180 => x"38",
          5181 => x"0c",
          5182 => x"34",
          5183 => x"33",
          5184 => x"82",
          5185 => x"fc",
          5186 => x"12",
          5187 => x"07",
          5188 => x"2b",
          5189 => x"45",
          5190 => x"a4",
          5191 => x"38",
          5192 => x"12",
          5193 => x"07",
          5194 => x"2b",
          5195 => x"5b",
          5196 => x"e4",
          5197 => x"38",
          5198 => x"12",
          5199 => x"07",
          5200 => x"2b",
          5201 => x"5d",
          5202 => x"12",
          5203 => x"07",
          5204 => x"2b",
          5205 => x"0c",
          5206 => x"45",
          5207 => x"d1",
          5208 => x"d1",
          5209 => x"d1",
          5210 => x"98",
          5211 => x"24",
          5212 => x"56",
          5213 => x"08",
          5214 => x"33",
          5215 => x"ba",
          5216 => x"81",
          5217 => x"18",
          5218 => x"31",
          5219 => x"38",
          5220 => x"81",
          5221 => x"fd",
          5222 => x"f3",
          5223 => x"83",
          5224 => x"39",
          5225 => x"33",
          5226 => x"58",
          5227 => x"42",
          5228 => x"83",
          5229 => x"2b",
          5230 => x"70",
          5231 => x"07",
          5232 => x"5a",
          5233 => x"39",
          5234 => x"38",
          5235 => x"2e",
          5236 => x"5a",
          5237 => x"79",
          5238 => x"54",
          5239 => x"53",
          5240 => x"ad",
          5241 => x"0d",
          5242 => x"43",
          5243 => x"5a",
          5244 => x"78",
          5245 => x"26",
          5246 => x"38",
          5247 => x"d9",
          5248 => x"74",
          5249 => x"84",
          5250 => x"73",
          5251 => x"62",
          5252 => x"74",
          5253 => x"54",
          5254 => x"93",
          5255 => x"81",
          5256 => x"84",
          5257 => x"8b",
          5258 => x"0d",
          5259 => x"ff",
          5260 => x"91",
          5261 => x"d0",
          5262 => x"f7",
          5263 => x"5e",
          5264 => x"79",
          5265 => x"81",
          5266 => x"57",
          5267 => x"15",
          5268 => x"9f",
          5269 => x"e0",
          5270 => x"74",
          5271 => x"76",
          5272 => x"ff",
          5273 => x"70",
          5274 => x"57",
          5275 => x"1b",
          5276 => x"ff",
          5277 => x"7a",
          5278 => x"0c",
          5279 => x"6c",
          5280 => x"56",
          5281 => x"38",
          5282 => x"cc",
          5283 => x"58",
          5284 => x"57",
          5285 => x"38",
          5286 => x"ba",
          5287 => x"40",
          5288 => x"e1",
          5289 => x"84",
          5290 => x"38",
          5291 => x"81",
          5292 => x"38",
          5293 => x"88",
          5294 => x"83",
          5295 => x"81",
          5296 => x"12",
          5297 => x"33",
          5298 => x"2e",
          5299 => x"34",
          5300 => x"90",
          5301 => x"34",
          5302 => x"7e",
          5303 => x"34",
          5304 => x"5d",
          5305 => x"5b",
          5306 => x"9d",
          5307 => x"80",
          5308 => x"0b",
          5309 => x"e2",
          5310 => x"08",
          5311 => x"89",
          5312 => x"8a",
          5313 => x"a3",
          5314 => x"98",
          5315 => x"b8",
          5316 => x"7c",
          5317 => x"02",
          5318 => x"81",
          5319 => x"77",
          5320 => x"2e",
          5321 => x"81",
          5322 => x"56",
          5323 => x"c0",
          5324 => x"1b",
          5325 => x"11",
          5326 => x"07",
          5327 => x"7b",
          5328 => x"1a",
          5329 => x"12",
          5330 => x"07",
          5331 => x"2b",
          5332 => x"05",
          5333 => x"59",
          5334 => x"1a",
          5335 => x"91",
          5336 => x"77",
          5337 => x"2e",
          5338 => x"f1",
          5339 => x"22",
          5340 => x"76",
          5341 => x"5b",
          5342 => x"70",
          5343 => x"84",
          5344 => x"ac",
          5345 => x"84",
          5346 => x"82",
          5347 => x"80",
          5348 => x"39",
          5349 => x"5e",
          5350 => x"06",
          5351 => x"88",
          5352 => x"87",
          5353 => x"84",
          5354 => x"79",
          5355 => x"08",
          5356 => x"c8",
          5357 => x"31",
          5358 => x"33",
          5359 => x"90",
          5360 => x"fd",
          5361 => x"81",
          5362 => x"ab",
          5363 => x"84",
          5364 => x"38",
          5365 => x"d9",
          5366 => x"83",
          5367 => x"51",
          5368 => x"08",
          5369 => x"11",
          5370 => x"75",
          5371 => x"18",
          5372 => x"74",
          5373 => x"26",
          5374 => x"0b",
          5375 => x"34",
          5376 => x"17",
          5377 => x"07",
          5378 => x"8e",
          5379 => x"a1",
          5380 => x"91",
          5381 => x"17",
          5382 => x"9a",
          5383 => x"7d",
          5384 => x"06",
          5385 => x"7f",
          5386 => x"16",
          5387 => x"33",
          5388 => x"b5",
          5389 => x"52",
          5390 => x"3f",
          5391 => x"38",
          5392 => x"0c",
          5393 => x"0c",
          5394 => x"80",
          5395 => x"b4",
          5396 => x"81",
          5397 => x"3f",
          5398 => x"81",
          5399 => x"08",
          5400 => x"17",
          5401 => x"55",
          5402 => x"38",
          5403 => x"09",
          5404 => x"b4",
          5405 => x"79",
          5406 => x"b8",
          5407 => x"94",
          5408 => x"77",
          5409 => x"75",
          5410 => x"f8",
          5411 => x"08",
          5412 => x"27",
          5413 => x"71",
          5414 => x"74",
          5415 => x"2a",
          5416 => x"ed",
          5417 => x"f7",
          5418 => x"f7",
          5419 => x"80",
          5420 => x"57",
          5421 => x"62",
          5422 => x"80",
          5423 => x"9f",
          5424 => x"97",
          5425 => x"8f",
          5426 => x"59",
          5427 => x"80",
          5428 => x"8c",
          5429 => x"84",
          5430 => x"87",
          5431 => x"94",
          5432 => x"56",
          5433 => x"7b",
          5434 => x"75",
          5435 => x"38",
          5436 => x"2a",
          5437 => x"d3",
          5438 => x"27",
          5439 => x"f0",
          5440 => x"98",
          5441 => x"fe",
          5442 => x"e7",
          5443 => x"b0",
          5444 => x"2e",
          5445 => x"2a",
          5446 => x"38",
          5447 => x"38",
          5448 => x"53",
          5449 => x"9f",
          5450 => x"98",
          5451 => x"75",
          5452 => x"77",
          5453 => x"84",
          5454 => x"58",
          5455 => x"33",
          5456 => x"15",
          5457 => x"58",
          5458 => x"0c",
          5459 => x"59",
          5460 => x"af",
          5461 => x"0c",
          5462 => x"8c",
          5463 => x"fe",
          5464 => x"83",
          5465 => x"5b",
          5466 => x"76",
          5467 => x"38",
          5468 => x"41",
          5469 => x"80",
          5470 => x"19",
          5471 => x"b1",
          5472 => x"85",
          5473 => x"1a",
          5474 => x"1b",
          5475 => x"5a",
          5476 => x"2e",
          5477 => x"56",
          5478 => x"ff",
          5479 => x"38",
          5480 => x"70",
          5481 => x"75",
          5482 => x"b4",
          5483 => x"81",
          5484 => x"3f",
          5485 => x"2e",
          5486 => x"ba",
          5487 => x"08",
          5488 => x"08",
          5489 => x"fe",
          5490 => x"82",
          5491 => x"81",
          5492 => x"05",
          5493 => x"ff",
          5494 => x"39",
          5495 => x"56",
          5496 => x"79",
          5497 => x"8c",
          5498 => x"33",
          5499 => x"8c",
          5500 => x"38",
          5501 => x"39",
          5502 => x"84",
          5503 => x"82",
          5504 => x"ba",
          5505 => x"3d",
          5506 => x"5c",
          5507 => x"80",
          5508 => x"80",
          5509 => x"80",
          5510 => x"1b",
          5511 => x"fd",
          5512 => x"76",
          5513 => x"74",
          5514 => x"81",
          5515 => x"76",
          5516 => x"08",
          5517 => x"84",
          5518 => x"82",
          5519 => x"7e",
          5520 => x"ff",
          5521 => x"78",
          5522 => x"1a",
          5523 => x"38",
          5524 => x"ff",
          5525 => x"0c",
          5526 => x"1b",
          5527 => x"1b",
          5528 => x"08",
          5529 => x"58",
          5530 => x"8a",
          5531 => x"08",
          5532 => x"de",
          5533 => x"5c",
          5534 => x"19",
          5535 => x"79",
          5536 => x"52",
          5537 => x"3f",
          5538 => x"60",
          5539 => x"74",
          5540 => x"b8",
          5541 => x"56",
          5542 => x"70",
          5543 => x"75",
          5544 => x"34",
          5545 => x"7e",
          5546 => x"1c",
          5547 => x"8c",
          5548 => x"75",
          5549 => x"8c",
          5550 => x"1a",
          5551 => x"7a",
          5552 => x"ba",
          5553 => x"84",
          5554 => x"83",
          5555 => x"60",
          5556 => x"08",
          5557 => x"80",
          5558 => x"83",
          5559 => x"08",
          5560 => x"17",
          5561 => x"2e",
          5562 => x"54",
          5563 => x"33",
          5564 => x"8c",
          5565 => x"81",
          5566 => x"bf",
          5567 => x"06",
          5568 => x"56",
          5569 => x"70",
          5570 => x"05",
          5571 => x"38",
          5572 => x"fe",
          5573 => x"53",
          5574 => x"52",
          5575 => x"84",
          5576 => x"06",
          5577 => x"83",
          5578 => x"08",
          5579 => x"74",
          5580 => x"82",
          5581 => x"81",
          5582 => x"16",
          5583 => x"52",
          5584 => x"3f",
          5585 => x"08",
          5586 => x"38",
          5587 => x"38",
          5588 => x"08",
          5589 => x"58",
          5590 => x"79",
          5591 => x"8c",
          5592 => x"d8",
          5593 => x"39",
          5594 => x"3f",
          5595 => x"8c",
          5596 => x"54",
          5597 => x"53",
          5598 => x"b8",
          5599 => x"38",
          5600 => x"b4",
          5601 => x"77",
          5602 => x"82",
          5603 => x"81",
          5604 => x"16",
          5605 => x"52",
          5606 => x"3f",
          5607 => x"33",
          5608 => x"8c",
          5609 => x"38",
          5610 => x"39",
          5611 => x"16",
          5612 => x"ff",
          5613 => x"80",
          5614 => x"17",
          5615 => x"31",
          5616 => x"98",
          5617 => x"2e",
          5618 => x"54",
          5619 => x"53",
          5620 => x"96",
          5621 => x"94",
          5622 => x"81",
          5623 => x"ba",
          5624 => x"0b",
          5625 => x"8c",
          5626 => x"0d",
          5627 => x"9f",
          5628 => x"97",
          5629 => x"8f",
          5630 => x"58",
          5631 => x"80",
          5632 => x"d8",
          5633 => x"81",
          5634 => x"c8",
          5635 => x"b4",
          5636 => x"17",
          5637 => x"54",
          5638 => x"33",
          5639 => x"8c",
          5640 => x"81",
          5641 => x"90",
          5642 => x"a0",
          5643 => x"77",
          5644 => x"ff",
          5645 => x"34",
          5646 => x"34",
          5647 => x"56",
          5648 => x"8c",
          5649 => x"88",
          5650 => x"90",
          5651 => x"98",
          5652 => x"7a",
          5653 => x"0b",
          5654 => x"18",
          5655 => x"0b",
          5656 => x"83",
          5657 => x"3f",
          5658 => x"81",
          5659 => x"34",
          5660 => x"0d",
          5661 => x"b8",
          5662 => x"5b",
          5663 => x"ba",
          5664 => x"8c",
          5665 => x"a8",
          5666 => x"57",
          5667 => x"8e",
          5668 => x"2e",
          5669 => x"54",
          5670 => x"53",
          5671 => x"92",
          5672 => x"78",
          5673 => x"74",
          5674 => x"8c",
          5675 => x"88",
          5676 => x"90",
          5677 => x"98",
          5678 => x"7a",
          5679 => x"0b",
          5680 => x"18",
          5681 => x"0b",
          5682 => x"83",
          5683 => x"3f",
          5684 => x"81",
          5685 => x"34",
          5686 => x"ff",
          5687 => x"81",
          5688 => x"78",
          5689 => x"3d",
          5690 => x"3f",
          5691 => x"8c",
          5692 => x"2e",
          5693 => x"2e",
          5694 => x"2e",
          5695 => x"22",
          5696 => x"80",
          5697 => x"38",
          5698 => x"0c",
          5699 => x"51",
          5700 => x"08",
          5701 => x"75",
          5702 => x"0d",
          5703 => x"80",
          5704 => x"57",
          5705 => x"ba",
          5706 => x"ba",
          5707 => x"51",
          5708 => x"d1",
          5709 => x"0c",
          5710 => x"ba",
          5711 => x"33",
          5712 => x"53",
          5713 => x"19",
          5714 => x"54",
          5715 => x"0b",
          5716 => x"79",
          5717 => x"33",
          5718 => x"9f",
          5719 => x"89",
          5720 => x"53",
          5721 => x"26",
          5722 => x"06",
          5723 => x"55",
          5724 => x"85",
          5725 => x"32",
          5726 => x"76",
          5727 => x"92",
          5728 => x"83",
          5729 => x"fe",
          5730 => x"77",
          5731 => x"3d",
          5732 => x"52",
          5733 => x"ba",
          5734 => x"80",
          5735 => x"0c",
          5736 => x"52",
          5737 => x"3f",
          5738 => x"8c",
          5739 => x"05",
          5740 => x"77",
          5741 => x"33",
          5742 => x"75",
          5743 => x"11",
          5744 => x"07",
          5745 => x"79",
          5746 => x"0c",
          5747 => x"0d",
          5748 => x"09",
          5749 => x"84",
          5750 => x"95",
          5751 => x"2b",
          5752 => x"1b",
          5753 => x"98",
          5754 => x"0c",
          5755 => x"0d",
          5756 => x"08",
          5757 => x"80",
          5758 => x"e5",
          5759 => x"8c",
          5760 => x"c8",
          5761 => x"61",
          5762 => x"58",
          5763 => x"80",
          5764 => x"98",
          5765 => x"ff",
          5766 => x"59",
          5767 => x"60",
          5768 => x"16",
          5769 => x"8c",
          5770 => x"83",
          5771 => x"16",
          5772 => x"c9",
          5773 => x"85",
          5774 => x"17",
          5775 => x"3d",
          5776 => x"71",
          5777 => x"40",
          5778 => x"da",
          5779 => x"52",
          5780 => x"ba",
          5781 => x"82",
          5782 => x"a8",
          5783 => x"84",
          5784 => x"3d",
          5785 => x"71",
          5786 => x"58",
          5787 => x"fd",
          5788 => x"ba",
          5789 => x"e2",
          5790 => x"ba",
          5791 => x"78",
          5792 => x"c8",
          5793 => x"52",
          5794 => x"7f",
          5795 => x"2e",
          5796 => x"81",
          5797 => x"f5",
          5798 => x"81",
          5799 => x"7e",
          5800 => x"e6",
          5801 => x"59",
          5802 => x"76",
          5803 => x"08",
          5804 => x"da",
          5805 => x"77",
          5806 => x"84",
          5807 => x"e5",
          5808 => x"59",
          5809 => x"38",
          5810 => x"5f",
          5811 => x"7a",
          5812 => x"7a",
          5813 => x"33",
          5814 => x"17",
          5815 => x"7c",
          5816 => x"2e",
          5817 => x"59",
          5818 => x"0c",
          5819 => x"33",
          5820 => x"90",
          5821 => x"fd",
          5822 => x"33",
          5823 => x"79",
          5824 => x"80",
          5825 => x"84",
          5826 => x"08",
          5827 => x"39",
          5828 => x"16",
          5829 => x"ff",
          5830 => x"8c",
          5831 => x"08",
          5832 => x"17",
          5833 => x"55",
          5834 => x"38",
          5835 => x"09",
          5836 => x"b4",
          5837 => x"7d",
          5838 => x"b8",
          5839 => x"18",
          5840 => x"af",
          5841 => x"33",
          5842 => x"70",
          5843 => x"5a",
          5844 => x"e8",
          5845 => x"08",
          5846 => x"7c",
          5847 => x"27",
          5848 => x"18",
          5849 => x"70",
          5850 => x"d4",
          5851 => x"7c",
          5852 => x"e4",
          5853 => x"7d",
          5854 => x"9f",
          5855 => x"97",
          5856 => x"8f",
          5857 => x"59",
          5858 => x"80",
          5859 => x"c2",
          5860 => x"ba",
          5861 => x"26",
          5862 => x"80",
          5863 => x"79",
          5864 => x"5a",
          5865 => x"75",
          5866 => x"3f",
          5867 => x"54",
          5868 => x"3f",
          5869 => x"d5",
          5870 => x"17",
          5871 => x"56",
          5872 => x"38",
          5873 => x"76",
          5874 => x"0c",
          5875 => x"06",
          5876 => x"fe",
          5877 => x"f3",
          5878 => x"ba",
          5879 => x"73",
          5880 => x"82",
          5881 => x"08",
          5882 => x"0c",
          5883 => x"34",
          5884 => x"8b",
          5885 => x"81",
          5886 => x"bb",
          5887 => x"80",
          5888 => x"fe",
          5889 => x"15",
          5890 => x"73",
          5891 => x"c0",
          5892 => x"83",
          5893 => x"38",
          5894 => x"77",
          5895 => x"8c",
          5896 => x"94",
          5897 => x"80",
          5898 => x"0c",
          5899 => x"a8",
          5900 => x"15",
          5901 => x"ff",
          5902 => x"79",
          5903 => x"5a",
          5904 => x"38",
          5905 => x"18",
          5906 => x"5a",
          5907 => x"8c",
          5908 => x"52",
          5909 => x"ba",
          5910 => x"14",
          5911 => x"ba",
          5912 => x"cf",
          5913 => x"c9",
          5914 => x"cb",
          5915 => x"ba",
          5916 => x"ba",
          5917 => x"84",
          5918 => x"98",
          5919 => x"91",
          5920 => x"0c",
          5921 => x"7c",
          5922 => x"38",
          5923 => x"8d",
          5924 => x"84",
          5925 => x"08",
          5926 => x"74",
          5927 => x"3d",
          5928 => x"75",
          5929 => x"8c",
          5930 => x"d1",
          5931 => x"59",
          5932 => x"16",
          5933 => x"54",
          5934 => x"16",
          5935 => x"71",
          5936 => x"5d",
          5937 => x"38",
          5938 => x"18",
          5939 => x"51",
          5940 => x"08",
          5941 => x"80",
          5942 => x"fe",
          5943 => x"fe",
          5944 => x"33",
          5945 => x"7a",
          5946 => x"bc",
          5947 => x"54",
          5948 => x"53",
          5949 => x"52",
          5950 => x"22",
          5951 => x"2e",
          5952 => x"84",
          5953 => x"8c",
          5954 => x"33",
          5955 => x"8c",
          5956 => x"71",
          5957 => x"3d",
          5958 => x"74",
          5959 => x"73",
          5960 => x"72",
          5961 => x"84",
          5962 => x"81",
          5963 => x"53",
          5964 => x"80",
          5965 => x"9d",
          5966 => x"84",
          5967 => x"84",
          5968 => x"74",
          5969 => x"74",
          5970 => x"8c",
          5971 => x"07",
          5972 => x"55",
          5973 => x"8a",
          5974 => x"52",
          5975 => x"74",
          5976 => x"8c",
          5977 => x"07",
          5978 => x"55",
          5979 => x"51",
          5980 => x"08",
          5981 => x"04",
          5982 => x"3f",
          5983 => x"72",
          5984 => x"56",
          5985 => x"57",
          5986 => x"3d",
          5987 => x"8c",
          5988 => x"2e",
          5989 => x"95",
          5990 => x"ff",
          5991 => x"55",
          5992 => x"80",
          5993 => x"58",
          5994 => x"2e",
          5995 => x"b0",
          5996 => x"95",
          5997 => x"8c",
          5998 => x"0d",
          5999 => x"3d",
          6000 => x"b9",
          6001 => x"ba",
          6002 => x"74",
          6003 => x"13",
          6004 => x"26",
          6005 => x"ba",
          6006 => x"ba",
          6007 => x"81",
          6008 => x"08",
          6009 => x"77",
          6010 => x"5c",
          6011 => x"82",
          6012 => x"5d",
          6013 => x"53",
          6014 => x"fe",
          6015 => x"80",
          6016 => x"79",
          6017 => x"7d",
          6018 => x"82",
          6019 => x"05",
          6020 => x"90",
          6021 => x"33",
          6022 => x"71",
          6023 => x"70",
          6024 => x"84",
          6025 => x"43",
          6026 => x"40",
          6027 => x"7f",
          6028 => x"33",
          6029 => x"79",
          6030 => x"04",
          6031 => x"17",
          6032 => x"fe",
          6033 => x"8c",
          6034 => x"08",
          6035 => x"18",
          6036 => x"55",
          6037 => x"38",
          6038 => x"09",
          6039 => x"b4",
          6040 => x"7c",
          6041 => x"e0",
          6042 => x"77",
          6043 => x"77",
          6044 => x"8c",
          6045 => x"ba",
          6046 => x"84",
          6047 => x"8c",
          6048 => x"18",
          6049 => x"08",
          6050 => x"7a",
          6051 => x"07",
          6052 => x"39",
          6053 => x"71",
          6054 => x"70",
          6055 => x"06",
          6056 => x"5f",
          6057 => x"39",
          6058 => x"58",
          6059 => x"0c",
          6060 => x"84",
          6061 => x"58",
          6062 => x"57",
          6063 => x"76",
          6064 => x"74",
          6065 => x"86",
          6066 => x"78",
          6067 => x"73",
          6068 => x"33",
          6069 => x"33",
          6070 => x"87",
          6071 => x"94",
          6072 => x"27",
          6073 => x"17",
          6074 => x"27",
          6075 => x"b3",
          6076 => x"0c",
          6077 => x"80",
          6078 => x"75",
          6079 => x"34",
          6080 => x"8b",
          6081 => x"27",
          6082 => x"fe",
          6083 => x"59",
          6084 => x"e9",
          6085 => x"82",
          6086 => x"2e",
          6087 => x"75",
          6088 => x"8c",
          6089 => x"fe",
          6090 => x"74",
          6091 => x"94",
          6092 => x"54",
          6093 => x"79",
          6094 => x"15",
          6095 => x"ba",
          6096 => x"95",
          6097 => x"8f",
          6098 => x"54",
          6099 => x"fe",
          6100 => x"51",
          6101 => x"08",
          6102 => x"8c",
          6103 => x"81",
          6104 => x"08",
          6105 => x"84",
          6106 => x"08",
          6107 => x"8c",
          6108 => x"8c",
          6109 => x"38",
          6110 => x"74",
          6111 => x"84",
          6112 => x"08",
          6113 => x"fe",
          6114 => x"59",
          6115 => x"cb",
          6116 => x"80",
          6117 => x"2e",
          6118 => x"75",
          6119 => x"8c",
          6120 => x"fe",
          6121 => x"74",
          6122 => x"17",
          6123 => x"73",
          6124 => x"26",
          6125 => x"90",
          6126 => x"56",
          6127 => x"33",
          6128 => x"e7",
          6129 => x"54",
          6130 => x"90",
          6131 => x"81",
          6132 => x"f0",
          6133 => x"39",
          6134 => x"0d",
          6135 => x"52",
          6136 => x"84",
          6137 => x"08",
          6138 => x"8c",
          6139 => x"a8",
          6140 => x"59",
          6141 => x"08",
          6142 => x"02",
          6143 => x"81",
          6144 => x"38",
          6145 => x"c4",
          6146 => x"81",
          6147 => x"b4",
          6148 => x"33",
          6149 => x"73",
          6150 => x"83",
          6151 => x"81",
          6152 => x"38",
          6153 => x"ff",
          6154 => x"ba",
          6155 => x"55",
          6156 => x"08",
          6157 => x"38",
          6158 => x"ff",
          6159 => x"56",
          6160 => x"0b",
          6161 => x"04",
          6162 => x"98",
          6163 => x"5d",
          6164 => x"8c",
          6165 => x"8c",
          6166 => x"a8",
          6167 => x"2e",
          6168 => x"ff",
          6169 => x"56",
          6170 => x"38",
          6171 => x"56",
          6172 => x"80",
          6173 => x"55",
          6174 => x"08",
          6175 => x"75",
          6176 => x"db",
          6177 => x"8c",
          6178 => x"5d",
          6179 => x"17",
          6180 => x"17",
          6181 => x"09",
          6182 => x"75",
          6183 => x"51",
          6184 => x"08",
          6185 => x"58",
          6186 => x"ab",
          6187 => x"34",
          6188 => x"08",
          6189 => x"78",
          6190 => x"8c",
          6191 => x"2e",
          6192 => x"81",
          6193 => x"c8",
          6194 => x"7c",
          6195 => x"90",
          6196 => x"7a",
          6197 => x"84",
          6198 => x"17",
          6199 => x"8c",
          6200 => x"27",
          6201 => x"74",
          6202 => x"38",
          6203 => x"08",
          6204 => x"51",
          6205 => x"c5",
          6206 => x"e1",
          6207 => x"e4",
          6208 => x"ba",
          6209 => x"84",
          6210 => x"38",
          6211 => x"cb",
          6212 => x"fe",
          6213 => x"b3",
          6214 => x"19",
          6215 => x"ff",
          6216 => x"84",
          6217 => x"18",
          6218 => x"a1",
          6219 => x"56",
          6220 => x"56",
          6221 => x"39",
          6222 => x"ff",
          6223 => x"b2",
          6224 => x"84",
          6225 => x"75",
          6226 => x"04",
          6227 => x"52",
          6228 => x"8c",
          6229 => x"38",
          6230 => x"3d",
          6231 => x"2e",
          6232 => x"f3",
          6233 => x"56",
          6234 => x"7d",
          6235 => x"5d",
          6236 => x"08",
          6237 => x"83",
          6238 => x"81",
          6239 => x"08",
          6240 => x"c9",
          6241 => x"12",
          6242 => x"38",
          6243 => x"5a",
          6244 => x"38",
          6245 => x"19",
          6246 => x"0c",
          6247 => x"55",
          6248 => x"ff",
          6249 => x"8a",
          6250 => x"f9",
          6251 => x"52",
          6252 => x"3f",
          6253 => x"81",
          6254 => x"84",
          6255 => x"b8",
          6256 => x"58",
          6257 => x"ba",
          6258 => x"08",
          6259 => x"18",
          6260 => x"27",
          6261 => x"7a",
          6262 => x"38",
          6263 => x"08",
          6264 => x"51",
          6265 => x"81",
          6266 => x"7c",
          6267 => x"08",
          6268 => x"51",
          6269 => x"08",
          6270 => x"fd",
          6271 => x"2e",
          6272 => x"ff",
          6273 => x"52",
          6274 => x"ba",
          6275 => x"08",
          6276 => x"59",
          6277 => x"94",
          6278 => x"5c",
          6279 => x"7a",
          6280 => x"8c",
          6281 => x"22",
          6282 => x"81",
          6283 => x"fe",
          6284 => x"56",
          6285 => x"ff",
          6286 => x"ae",
          6287 => x"0b",
          6288 => x"80",
          6289 => x"34",
          6290 => x"cc",
          6291 => x"83",
          6292 => x"d2",
          6293 => x"80",
          6294 => x"83",
          6295 => x"0b",
          6296 => x"56",
          6297 => x"70",
          6298 => x"75",
          6299 => x"d9",
          6300 => x"ff",
          6301 => x"17",
          6302 => x"f3",
          6303 => x"2e",
          6304 => x"83",
          6305 => x"3f",
          6306 => x"8c",
          6307 => x"ba",
          6308 => x"8c",
          6309 => x"17",
          6310 => x"7d",
          6311 => x"77",
          6312 => x"7c",
          6313 => x"38",
          6314 => x"7d",
          6315 => x"51",
          6316 => x"08",
          6317 => x"3d",
          6318 => x"80",
          6319 => x"76",
          6320 => x"7b",
          6321 => x"34",
          6322 => x"17",
          6323 => x"1a",
          6324 => x"39",
          6325 => x"34",
          6326 => x"34",
          6327 => x"7d",
          6328 => x"51",
          6329 => x"08",
          6330 => x"b3",
          6331 => x"5f",
          6332 => x"81",
          6333 => x"56",
          6334 => x"ed",
          6335 => x"82",
          6336 => x"b2",
          6337 => x"ba",
          6338 => x"80",
          6339 => x"0c",
          6340 => x"0c",
          6341 => x"52",
          6342 => x"8c",
          6343 => x"38",
          6344 => x"06",
          6345 => x"0b",
          6346 => x"55",
          6347 => x"70",
          6348 => x"74",
          6349 => x"7a",
          6350 => x"57",
          6351 => x"ff",
          6352 => x"08",
          6353 => x"84",
          6354 => x"08",
          6355 => x"2e",
          6356 => x"8c",
          6357 => x"d0",
          6358 => x"58",
          6359 => x"78",
          6360 => x"78",
          6361 => x"08",
          6362 => x"5e",
          6363 => x"5c",
          6364 => x"ff",
          6365 => x"26",
          6366 => x"06",
          6367 => x"99",
          6368 => x"ff",
          6369 => x"2a",
          6370 => x"06",
          6371 => x"7a",
          6372 => x"2a",
          6373 => x"2e",
          6374 => x"5c",
          6375 => x"08",
          6376 => x"83",
          6377 => x"82",
          6378 => x"b2",
          6379 => x"ba",
          6380 => x"fd",
          6381 => x"3d",
          6382 => x"38",
          6383 => x"ba",
          6384 => x"fd",
          6385 => x"19",
          6386 => x"56",
          6387 => x"75",
          6388 => x"5a",
          6389 => x"33",
          6390 => x"84",
          6391 => x"38",
          6392 => x"34",
          6393 => x"8b",
          6394 => x"57",
          6395 => x"a7",
          6396 => x"7f",
          6397 => x"88",
          6398 => x"57",
          6399 => x"16",
          6400 => x"75",
          6401 => x"22",
          6402 => x"57",
          6403 => x"75",
          6404 => x"2e",
          6405 => x"83",
          6406 => x"17",
          6407 => x"f1",
          6408 => x"85",
          6409 => x"18",
          6410 => x"56",
          6411 => x"33",
          6412 => x"bb",
          6413 => x"5d",
          6414 => x"88",
          6415 => x"76",
          6416 => x"06",
          6417 => x"80",
          6418 => x"75",
          6419 => x"0b",
          6420 => x"08",
          6421 => x"ff",
          6422 => x"fe",
          6423 => x"55",
          6424 => x"b8",
          6425 => x"5a",
          6426 => x"83",
          6427 => x"2e",
          6428 => x"54",
          6429 => x"33",
          6430 => x"8c",
          6431 => x"81",
          6432 => x"77",
          6433 => x"7a",
          6434 => x"19",
          6435 => x"78",
          6436 => x"8c",
          6437 => x"2e",
          6438 => x"2e",
          6439 => x"db",
          6440 => x"84",
          6441 => x"b1",
          6442 => x"8c",
          6443 => x"33",
          6444 => x"90",
          6445 => x"fd",
          6446 => x"2e",
          6447 => x"80",
          6448 => x"8c",
          6449 => x"b4",
          6450 => x"33",
          6451 => x"84",
          6452 => x"06",
          6453 => x"83",
          6454 => x"08",
          6455 => x"74",
          6456 => x"82",
          6457 => x"81",
          6458 => x"16",
          6459 => x"52",
          6460 => x"3f",
          6461 => x"b4",
          6462 => x"81",
          6463 => x"3f",
          6464 => x"c9",
          6465 => x"34",
          6466 => x"84",
          6467 => x"18",
          6468 => x"33",
          6469 => x"fc",
          6470 => x"a0",
          6471 => x"17",
          6472 => x"5c",
          6473 => x"80",
          6474 => x"e3",
          6475 => x"3d",
          6476 => x"a2",
          6477 => x"84",
          6478 => x"75",
          6479 => x"04",
          6480 => x"05",
          6481 => x"8c",
          6482 => x"38",
          6483 => x"06",
          6484 => x"a7",
          6485 => x"71",
          6486 => x"57",
          6487 => x"81",
          6488 => x"e2",
          6489 => x"ba",
          6490 => x"3d",
          6491 => x"cc",
          6492 => x"d9",
          6493 => x"ba",
          6494 => x"84",
          6495 => x"78",
          6496 => x"51",
          6497 => x"08",
          6498 => x"02",
          6499 => x"56",
          6500 => x"18",
          6501 => x"07",
          6502 => x"76",
          6503 => x"76",
          6504 => x"76",
          6505 => x"78",
          6506 => x"51",
          6507 => x"08",
          6508 => x"04",
          6509 => x"80",
          6510 => x"3d",
          6511 => x"8c",
          6512 => x"84",
          6513 => x"56",
          6514 => x"70",
          6515 => x"38",
          6516 => x"56",
          6517 => x"81",
          6518 => x"2e",
          6519 => x"58",
          6520 => x"2e",
          6521 => x"5a",
          6522 => x"81",
          6523 => x"16",
          6524 => x"c9",
          6525 => x"85",
          6526 => x"17",
          6527 => x"70",
          6528 => x"83",
          6529 => x"84",
          6530 => x"b8",
          6531 => x"71",
          6532 => x"14",
          6533 => x"33",
          6534 => x"57",
          6535 => x"9a",
          6536 => x"80",
          6537 => x"f4",
          6538 => x"84",
          6539 => x"38",
          6540 => x"b8",
          6541 => x"b0",
          6542 => x"b8",
          6543 => x"5b",
          6544 => x"ba",
          6545 => x"fe",
          6546 => x"17",
          6547 => x"31",
          6548 => x"a0",
          6549 => x"16",
          6550 => x"06",
          6551 => x"08",
          6552 => x"81",
          6553 => x"79",
          6554 => x"52",
          6555 => x"3f",
          6556 => x"8d",
          6557 => x"51",
          6558 => x"08",
          6559 => x"38",
          6560 => x"08",
          6561 => x"19",
          6562 => x"75",
          6563 => x"ec",
          6564 => x"76",
          6565 => x"ff",
          6566 => x"58",
          6567 => x"39",
          6568 => x"0d",
          6569 => x"52",
          6570 => x"84",
          6571 => x"08",
          6572 => x"7d",
          6573 => x"58",
          6574 => x"74",
          6575 => x"ff",
          6576 => x"27",
          6577 => x"5c",
          6578 => x"57",
          6579 => x"0c",
          6580 => x"38",
          6581 => x"52",
          6582 => x"3f",
          6583 => x"06",
          6584 => x"83",
          6585 => x"70",
          6586 => x"80",
          6587 => x"77",
          6588 => x"70",
          6589 => x"80",
          6590 => x"81",
          6591 => x"59",
          6592 => x"27",
          6593 => x"96",
          6594 => x"76",
          6595 => x"05",
          6596 => x"70",
          6597 => x"3d",
          6598 => x"5b",
          6599 => x"d1",
          6600 => x"76",
          6601 => x"2e",
          6602 => x"16",
          6603 => x"09",
          6604 => x"79",
          6605 => x"52",
          6606 => x"e4",
          6607 => x"ba",
          6608 => x"56",
          6609 => x"0d",
          6610 => x"e7",
          6611 => x"ff",
          6612 => x"56",
          6613 => x"0d",
          6614 => x"c3",
          6615 => x"ee",
          6616 => x"ba",
          6617 => x"2e",
          6618 => x"57",
          6619 => x"76",
          6620 => x"55",
          6621 => x"83",
          6622 => x"3f",
          6623 => x"ff",
          6624 => x"38",
          6625 => x"8c",
          6626 => x"ee",
          6627 => x"e6",
          6628 => x"58",
          6629 => x"08",
          6630 => x"09",
          6631 => x"8c",
          6632 => x"08",
          6633 => x"2e",
          6634 => x"79",
          6635 => x"81",
          6636 => x"18",
          6637 => x"ba",
          6638 => x"57",
          6639 => x"57",
          6640 => x"70",
          6641 => x"2e",
          6642 => x"25",
          6643 => x"81",
          6644 => x"2e",
          6645 => x"ef",
          6646 => x"84",
          6647 => x"38",
          6648 => x"38",
          6649 => x"6c",
          6650 => x"58",
          6651 => x"6b",
          6652 => x"6c",
          6653 => x"05",
          6654 => x"34",
          6655 => x"eb",
          6656 => x"76",
          6657 => x"55",
          6658 => x"5a",
          6659 => x"83",
          6660 => x"3f",
          6661 => x"39",
          6662 => x"b4",
          6663 => x"33",
          6664 => x"8c",
          6665 => x"c3",
          6666 => x"34",
          6667 => x"5c",
          6668 => x"82",
          6669 => x"38",
          6670 => x"39",
          6671 => x"ed",
          6672 => x"84",
          6673 => x"38",
          6674 => x"78",
          6675 => x"39",
          6676 => x"08",
          6677 => x"51",
          6678 => x"f2",
          6679 => x"80",
          6680 => x"56",
          6681 => x"55",
          6682 => x"54",
          6683 => x"22",
          6684 => x"2e",
          6685 => x"75",
          6686 => x"75",
          6687 => x"a2",
          6688 => x"90",
          6689 => x"56",
          6690 => x"7e",
          6691 => x"55",
          6692 => x"82",
          6693 => x"70",
          6694 => x"08",
          6695 => x"5f",
          6696 => x"9c",
          6697 => x"58",
          6698 => x"52",
          6699 => x"15",
          6700 => x"26",
          6701 => x"08",
          6702 => x"8c",
          6703 => x"ba",
          6704 => x"59",
          6705 => x"2e",
          6706 => x"75",
          6707 => x"3d",
          6708 => x"0c",
          6709 => x"51",
          6710 => x"08",
          6711 => x"73",
          6712 => x"7b",
          6713 => x"56",
          6714 => x"18",
          6715 => x"73",
          6716 => x"dd",
          6717 => x"ba",
          6718 => x"19",
          6719 => x"38",
          6720 => x"80",
          6721 => x"0c",
          6722 => x"80",
          6723 => x"9c",
          6724 => x"58",
          6725 => x"76",
          6726 => x"33",
          6727 => x"75",
          6728 => x"97",
          6729 => x"39",
          6730 => x"fe",
          6731 => x"39",
          6732 => x"a3",
          6733 => x"05",
          6734 => x"ff",
          6735 => x"40",
          6736 => x"70",
          6737 => x"56",
          6738 => x"74",
          6739 => x"38",
          6740 => x"24",
          6741 => x"d1",
          6742 => x"80",
          6743 => x"16",
          6744 => x"81",
          6745 => x"79",
          6746 => x"8c",
          6747 => x"5d",
          6748 => x"75",
          6749 => x"7f",
          6750 => x"53",
          6751 => x"3f",
          6752 => x"6d",
          6753 => x"74",
          6754 => x"ff",
          6755 => x"38",
          6756 => x"7f",
          6757 => x"0a",
          6758 => x"06",
          6759 => x"2a",
          6760 => x"2b",
          6761 => x"2e",
          6762 => x"25",
          6763 => x"83",
          6764 => x"38",
          6765 => x"51",
          6766 => x"ba",
          6767 => x"ff",
          6768 => x"71",
          6769 => x"77",
          6770 => x"82",
          6771 => x"83",
          6772 => x"2e",
          6773 => x"11",
          6774 => x"71",
          6775 => x"72",
          6776 => x"83",
          6777 => x"33",
          6778 => x"81",
          6779 => x"75",
          6780 => x"42",
          6781 => x"4e",
          6782 => x"78",
          6783 => x"82",
          6784 => x"26",
          6785 => x"81",
          6786 => x"f9",
          6787 => x"2e",
          6788 => x"83",
          6789 => x"46",
          6790 => x"c2",
          6791 => x"57",
          6792 => x"58",
          6793 => x"26",
          6794 => x"10",
          6795 => x"74",
          6796 => x"ee",
          6797 => x"ba",
          6798 => x"05",
          6799 => x"26",
          6800 => x"08",
          6801 => x"11",
          6802 => x"83",
          6803 => x"a0",
          6804 => x"66",
          6805 => x"31",
          6806 => x"89",
          6807 => x"29",
          6808 => x"79",
          6809 => x"7d",
          6810 => x"56",
          6811 => x"08",
          6812 => x"62",
          6813 => x"38",
          6814 => x"08",
          6815 => x"38",
          6816 => x"89",
          6817 => x"8b",
          6818 => x"3d",
          6819 => x"4e",
          6820 => x"8c",
          6821 => x"0c",
          6822 => x"ff",
          6823 => x"91",
          6824 => x"d0",
          6825 => x"b2",
          6826 => x"5c",
          6827 => x"81",
          6828 => x"58",
          6829 => x"62",
          6830 => x"81",
          6831 => x"45",
          6832 => x"70",
          6833 => x"70",
          6834 => x"09",
          6835 => x"38",
          6836 => x"07",
          6837 => x"7a",
          6838 => x"84",
          6839 => x"98",
          6840 => x"3d",
          6841 => x"fe",
          6842 => x"8c",
          6843 => x"77",
          6844 => x"75",
          6845 => x"57",
          6846 => x"7f",
          6847 => x"fa",
          6848 => x"38",
          6849 => x"95",
          6850 => x"67",
          6851 => x"70",
          6852 => x"84",
          6853 => x"38",
          6854 => x"80",
          6855 => x"76",
          6856 => x"84",
          6857 => x"81",
          6858 => x"27",
          6859 => x"57",
          6860 => x"57",
          6861 => x"34",
          6862 => x"61",
          6863 => x"70",
          6864 => x"05",
          6865 => x"38",
          6866 => x"82",
          6867 => x"05",
          6868 => x"6a",
          6869 => x"5c",
          6870 => x"90",
          6871 => x"5a",
          6872 => x"9e",
          6873 => x"05",
          6874 => x"26",
          6875 => x"06",
          6876 => x"88",
          6877 => x"f8",
          6878 => x"05",
          6879 => x"61",
          6880 => x"34",
          6881 => x"2a",
          6882 => x"90",
          6883 => x"7e",
          6884 => x"ba",
          6885 => x"83",
          6886 => x"05",
          6887 => x"61",
          6888 => x"05",
          6889 => x"74",
          6890 => x"4b",
          6891 => x"61",
          6892 => x"34",
          6893 => x"59",
          6894 => x"33",
          6895 => x"15",
          6896 => x"05",
          6897 => x"ff",
          6898 => x"54",
          6899 => x"c6",
          6900 => x"08",
          6901 => x"83",
          6902 => x"55",
          6903 => x"ff",
          6904 => x"41",
          6905 => x"87",
          6906 => x"83",
          6907 => x"88",
          6908 => x"81",
          6909 => x"78",
          6910 => x"98",
          6911 => x"65",
          6912 => x"59",
          6913 => x"51",
          6914 => x"08",
          6915 => x"55",
          6916 => x"ff",
          6917 => x"77",
          6918 => x"7f",
          6919 => x"89",
          6920 => x"38",
          6921 => x"83",
          6922 => x"60",
          6923 => x"84",
          6924 => x"1b",
          6925 => x"38",
          6926 => x"86",
          6927 => x"38",
          6928 => x"81",
          6929 => x"2a",
          6930 => x"84",
          6931 => x"81",
          6932 => x"f4",
          6933 => x"6b",
          6934 => x"67",
          6935 => x"67",
          6936 => x"34",
          6937 => x"80",
          6938 => x"f7",
          6939 => x"84",
          6940 => x"57",
          6941 => x"8c",
          6942 => x"83",
          6943 => x"05",
          6944 => x"84",
          6945 => x"34",
          6946 => x"88",
          6947 => x"34",
          6948 => x"cc",
          6949 => x"61",
          6950 => x"53",
          6951 => x"3f",
          6952 => x"c9",
          6953 => x"fe",
          6954 => x"8c",
          6955 => x"08",
          6956 => x"84",
          6957 => x"e4",
          6958 => x"f6",
          6959 => x"2a",
          6960 => x"56",
          6961 => x"77",
          6962 => x"77",
          6963 => x"58",
          6964 => x"27",
          6965 => x"f5",
          6966 => x"10",
          6967 => x"5c",
          6968 => x"08",
          6969 => x"ff",
          6970 => x"8e",
          6971 => x"08",
          6972 => x"7a",
          6973 => x"7a",
          6974 => x"39",
          6975 => x"f8",
          6976 => x"75",
          6977 => x"49",
          6978 => x"2a",
          6979 => x"98",
          6980 => x"f9",
          6981 => x"34",
          6982 => x"61",
          6983 => x"80",
          6984 => x"34",
          6985 => x"05",
          6986 => x"a6",
          6987 => x"61",
          6988 => x"34",
          6989 => x"ae",
          6990 => x"81",
          6991 => x"05",
          6992 => x"61",
          6993 => x"c0",
          6994 => x"34",
          6995 => x"e8",
          6996 => x"58",
          6997 => x"ff",
          6998 => x"38",
          6999 => x"70",
          7000 => x"74",
          7001 => x"80",
          7002 => x"d9",
          7003 => x"f4",
          7004 => x"42",
          7005 => x"54",
          7006 => x"79",
          7007 => x"39",
          7008 => x"3d",
          7009 => x"61",
          7010 => x"05",
          7011 => x"4c",
          7012 => x"05",
          7013 => x"61",
          7014 => x"34",
          7015 => x"89",
          7016 => x"8f",
          7017 => x"76",
          7018 => x"51",
          7019 => x"56",
          7020 => x"34",
          7021 => x"5c",
          7022 => x"34",
          7023 => x"05",
          7024 => x"05",
          7025 => x"f2",
          7026 => x"61",
          7027 => x"83",
          7028 => x"e7",
          7029 => x"61",
          7030 => x"59",
          7031 => x"90",
          7032 => x"34",
          7033 => x"eb",
          7034 => x"34",
          7035 => x"61",
          7036 => x"ef",
          7037 => x"aa",
          7038 => x"60",
          7039 => x"81",
          7040 => x"51",
          7041 => x"55",
          7042 => x"61",
          7043 => x"5a",
          7044 => x"8d",
          7045 => x"81",
          7046 => x"b4",
          7047 => x"9e",
          7048 => x"2e",
          7049 => x"58",
          7050 => x"86",
          7051 => x"76",
          7052 => x"55",
          7053 => x"0d",
          7054 => x"05",
          7055 => x"2e",
          7056 => x"80",
          7057 => x"77",
          7058 => x"34",
          7059 => x"38",
          7060 => x"18",
          7061 => x"fc",
          7062 => x"76",
          7063 => x"7a",
          7064 => x"2a",
          7065 => x"88",
          7066 => x"8d",
          7067 => x"a3",
          7068 => x"05",
          7069 => x"77",
          7070 => x"58",
          7071 => x"a1",
          7072 => x"80",
          7073 => x"80",
          7074 => x"56",
          7075 => x"74",
          7076 => x"0c",
          7077 => x"80",
          7078 => x"ac",
          7079 => x"76",
          7080 => x"ba",
          7081 => x"ba",
          7082 => x"9f",
          7083 => x"11",
          7084 => x"08",
          7085 => x"32",
          7086 => x"70",
          7087 => x"39",
          7088 => x"ff",
          7089 => x"9f",
          7090 => x"02",
          7091 => x"80",
          7092 => x"72",
          7093 => x"ba",
          7094 => x"ff",
          7095 => x"2e",
          7096 => x"2e",
          7097 => x"72",
          7098 => x"83",
          7099 => x"ff",
          7100 => x"d0",
          7101 => x"81",
          7102 => x"ba",
          7103 => x"fe",
          7104 => x"84",
          7105 => x"53",
          7106 => x"53",
          7107 => x"0d",
          7108 => x"06",
          7109 => x"38",
          7110 => x"22",
          7111 => x"0d",
          7112 => x"83",
          7113 => x"83",
          7114 => x"56",
          7115 => x"74",
          7116 => x"30",
          7117 => x"54",
          7118 => x"70",
          7119 => x"2a",
          7120 => x"52",
          7121 => x"cf",
          7122 => x"05",
          7123 => x"25",
          7124 => x"70",
          7125 => x"84",
          7126 => x"83",
          7127 => x"88",
          7128 => x"ca",
          7129 => x"a0",
          7130 => x"51",
          7131 => x"70",
          7132 => x"39",
          7133 => x"57",
          7134 => x"ff",
          7135 => x"16",
          7136 => x"d0",
          7137 => x"06",
          7138 => x"83",
          7139 => x"39",
          7140 => x"31",
          7141 => x"55",
          7142 => x"75",
          7143 => x"39",
          7144 => x"ff",
          7145 => x"ff",
          7146 => x"19",
          7147 => x"19",
          7148 => x"19",
          7149 => x"19",
          7150 => x"19",
          7151 => x"19",
          7152 => x"18",
          7153 => x"18",
          7154 => x"18",
          7155 => x"18",
          7156 => x"1f",
          7157 => x"1f",
          7158 => x"1f",
          7159 => x"1f",
          7160 => x"1f",
          7161 => x"1f",
          7162 => x"1f",
          7163 => x"1f",
          7164 => x"1f",
          7165 => x"1f",
          7166 => x"1f",
          7167 => x"1f",
          7168 => x"1f",
          7169 => x"1f",
          7170 => x"1f",
          7171 => x"1f",
          7172 => x"1f",
          7173 => x"1f",
          7174 => x"1f",
          7175 => x"1f",
          7176 => x"1f",
          7177 => x"24",
          7178 => x"1f",
          7179 => x"1f",
          7180 => x"1f",
          7181 => x"1f",
          7182 => x"1f",
          7183 => x"1f",
          7184 => x"1f",
          7185 => x"1f",
          7186 => x"23",
          7187 => x"22",
          7188 => x"23",
          7189 => x"21",
          7190 => x"1f",
          7191 => x"1f",
          7192 => x"1f",
          7193 => x"1f",
          7194 => x"1f",
          7195 => x"1f",
          7196 => x"1f",
          7197 => x"1f",
          7198 => x"1f",
          7199 => x"1f",
          7200 => x"1f",
          7201 => x"1f",
          7202 => x"1f",
          7203 => x"1f",
          7204 => x"1f",
          7205 => x"1f",
          7206 => x"1f",
          7207 => x"1f",
          7208 => x"1f",
          7209 => x"1f",
          7210 => x"1f",
          7211 => x"1f",
          7212 => x"1f",
          7213 => x"1f",
          7214 => x"1f",
          7215 => x"1f",
          7216 => x"21",
          7217 => x"1f",
          7218 => x"1f",
          7219 => x"1f",
          7220 => x"1f",
          7221 => x"21",
          7222 => x"21",
          7223 => x"21",
          7224 => x"21",
          7225 => x"32",
          7226 => x"32",
          7227 => x"32",
          7228 => x"3a",
          7229 => x"36",
          7230 => x"34",
          7231 => x"36",
          7232 => x"36",
          7233 => x"39",
          7234 => x"38",
          7235 => x"37",
          7236 => x"34",
          7237 => x"36",
          7238 => x"36",
          7239 => x"46",
          7240 => x"46",
          7241 => x"46",
          7242 => x"47",
          7243 => x"47",
          7244 => x"47",
          7245 => x"47",
          7246 => x"47",
          7247 => x"47",
          7248 => x"47",
          7249 => x"47",
          7250 => x"47",
          7251 => x"47",
          7252 => x"47",
          7253 => x"47",
          7254 => x"47",
          7255 => x"47",
          7256 => x"47",
          7257 => x"48",
          7258 => x"48",
          7259 => x"47",
          7260 => x"48",
          7261 => x"47",
          7262 => x"48",
          7263 => x"47",
          7264 => x"47",
          7265 => x"47",
          7266 => x"47",
          7267 => x"54",
          7268 => x"55",
          7269 => x"54",
          7270 => x"54",
          7271 => x"52",
          7272 => x"57",
          7273 => x"52",
          7274 => x"52",
          7275 => x"52",
          7276 => x"57",
          7277 => x"52",
          7278 => x"52",
          7279 => x"52",
          7280 => x"52",
          7281 => x"52",
          7282 => x"52",
          7283 => x"52",
          7284 => x"52",
          7285 => x"52",
          7286 => x"52",
          7287 => x"52",
          7288 => x"52",
          7289 => x"53",
          7290 => x"52",
          7291 => x"52",
          7292 => x"53",
          7293 => x"53",
          7294 => x"59",
          7295 => x"59",
          7296 => x"59",
          7297 => x"58",
          7298 => x"59",
          7299 => x"59",
          7300 => x"59",
          7301 => x"59",
          7302 => x"59",
          7303 => x"59",
          7304 => x"59",
          7305 => x"59",
          7306 => x"59",
          7307 => x"59",
          7308 => x"59",
          7309 => x"5a",
          7310 => x"59",
          7311 => x"5a",
          7312 => x"5a",
          7313 => x"5a",
          7314 => x"5a",
          7315 => x"5a",
          7316 => x"59",
          7317 => x"59",
          7318 => x"59",
          7319 => x"61",
          7320 => x"61",
          7321 => x"61",
          7322 => x"61",
          7323 => x"61",
          7324 => x"61",
          7325 => x"61",
          7326 => x"61",
          7327 => x"61",
          7328 => x"61",
          7329 => x"63",
          7330 => x"61",
          7331 => x"61",
          7332 => x"5e",
          7333 => x"df",
          7334 => x"df",
          7335 => x"de",
          7336 => x"de",
          7337 => x"de",
          7338 => x"0b",
          7339 => x"0f",
          7340 => x"0b",
          7341 => x"0b",
          7342 => x"0b",
          7343 => x"0d",
          7344 => x"0f",
          7345 => x"0b",
          7346 => x"0b",
          7347 => x"0b",
          7348 => x"0b",
          7349 => x"0b",
          7350 => x"0b",
          7351 => x"0b",
          7352 => x"0b",
          7353 => x"0b",
          7354 => x"0b",
          7355 => x"0b",
          7356 => x"0b",
          7357 => x"0b",
          7358 => x"0b",
          7359 => x"0b",
          7360 => x"0b",
          7361 => x"0b",
          7362 => x"0b",
          7363 => x"0f",
          7364 => x"0b",
          7365 => x"0b",
          7366 => x"0b",
          7367 => x"0b",
          7368 => x"0b",
          7369 => x"0b",
          7370 => x"0b",
          7371 => x"0e",
          7372 => x"0e",
          7373 => x"0e",
          7374 => x"0e",
          7375 => x"0b",
          7376 => x"0b",
          7377 => x"0c",
          7378 => x"0b",
          7379 => x"0f",
          7380 => x"0c",
          7381 => x"0b",
          7382 => x"6e",
          7383 => x"6f",
          7384 => x"6e",
          7385 => x"6f",
          7386 => x"78",
          7387 => x"6c",
          7388 => x"6f",
          7389 => x"69",
          7390 => x"75",
          7391 => x"62",
          7392 => x"77",
          7393 => x"65",
          7394 => x"65",
          7395 => x"00",
          7396 => x"73",
          7397 => x"73",
          7398 => x"66",
          7399 => x"73",
          7400 => x"73",
          7401 => x"61",
          7402 => x"61",
          7403 => x"6c",
          7404 => x"00",
          7405 => x"6e",
          7406 => x"00",
          7407 => x"74",
          7408 => x"6f",
          7409 => x"00",
          7410 => x"6e",
          7411 => x"66",
          7412 => x"00",
          7413 => x"69",
          7414 => x"65",
          7415 => x"00",
          7416 => x"73",
          7417 => x"2e",
          7418 => x"74",
          7419 => x"74",
          7420 => x"63",
          7421 => x"00",
          7422 => x"20",
          7423 => x"2e",
          7424 => x"70",
          7425 => x"66",
          7426 => x"65",
          7427 => x"20",
          7428 => x"2e",
          7429 => x"6f",
          7430 => x"65",
          7431 => x"69",
          7432 => x"65",
          7433 => x"76",
          7434 => x"00",
          7435 => x"77",
          7436 => x"6f",
          7437 => x"00",
          7438 => x"61",
          7439 => x"76",
          7440 => x"00",
          7441 => x"6c",
          7442 => x"78",
          7443 => x"00",
          7444 => x"20",
          7445 => x"00",
          7446 => x"64",
          7447 => x"6d",
          7448 => x"20",
          7449 => x"75",
          7450 => x"20",
          7451 => x"75",
          7452 => x"73",
          7453 => x"65",
          7454 => x"74",
          7455 => x"72",
          7456 => x"73",
          7457 => x"00",
          7458 => x"73",
          7459 => x"6c",
          7460 => x"20",
          7461 => x"6c",
          7462 => x"2f",
          7463 => x"00",
          7464 => x"00",
          7465 => x"00",
          7466 => x"32",
          7467 => x"00",
          7468 => x"00",
          7469 => x"00",
          7470 => x"20",
          7471 => x"53",
          7472 => x"28",
          7473 => x"32",
          7474 => x"2e",
          7475 => x"50",
          7476 => x"25",
          7477 => x"20",
          7478 => x"00",
          7479 => x"74",
          7480 => x"48",
          7481 => x"00",
          7482 => x"54",
          7483 => x"72",
          7484 => x"52",
          7485 => x"6e",
          7486 => x"00",
          7487 => x"54",
          7488 => x"72",
          7489 => x"52",
          7490 => x"6e",
          7491 => x"00",
          7492 => x"57",
          7493 => x"72",
          7494 => x"43",
          7495 => x"6e",
          7496 => x"00",
          7497 => x"74",
          7498 => x"00",
          7499 => x"69",
          7500 => x"74",
          7501 => x"67",
          7502 => x"65",
          7503 => x"61",
          7504 => x"69",
          7505 => x"00",
          7506 => x"65",
          7507 => x"00",
          7508 => x"75",
          7509 => x"69",
          7510 => x"69",
          7511 => x"73",
          7512 => x"72",
          7513 => x"65",
          7514 => x"74",
          7515 => x"6c",
          7516 => x"00",
          7517 => x"00",
          7518 => x"6e",
          7519 => x"65",
          7520 => x"00",
          7521 => x"6d",
          7522 => x"00",
          7523 => x"6e",
          7524 => x"5c",
          7525 => x"00",
          7526 => x"65",
          7527 => x"2e",
          7528 => x"73",
          7529 => x"20",
          7530 => x"74",
          7531 => x"00",
          7532 => x"67",
          7533 => x"20",
          7534 => x"2e",
          7535 => x"6c",
          7536 => x"6e",
          7537 => x"20",
          7538 => x"00",
          7539 => x"69",
          7540 => x"20",
          7541 => x"20",
          7542 => x"38",
          7543 => x"58",
          7544 => x"38",
          7545 => x"2d",
          7546 => x"69",
          7547 => x"00",
          7548 => x"25",
          7549 => x"30",
          7550 => x"78",
          7551 => x"70",
          7552 => x"00",
          7553 => x"25",
          7554 => x"65",
          7555 => x"2e",
          7556 => x"6d",
          7557 => x"79",
          7558 => x"65",
          7559 => x"3a",
          7560 => x"00",
          7561 => x"20",
          7562 => x"65",
          7563 => x"6f",
          7564 => x"73",
          7565 => x"6e",
          7566 => x"3f",
          7567 => x"25",
          7568 => x"3a",
          7569 => x"0a",
          7570 => x"6e",
          7571 => x"69",
          7572 => x"44",
          7573 => x"69",
          7574 => x"74",
          7575 => x"64",
          7576 => x"00",
          7577 => x"55",
          7578 => x"56",
          7579 => x"64",
          7580 => x"20",
          7581 => x"00",
          7582 => x"55",
          7583 => x"20",
          7584 => x"64",
          7585 => x"20",
          7586 => x"00",
          7587 => x"61",
          7588 => x"74",
          7589 => x"73",
          7590 => x"20",
          7591 => x"00",
          7592 => x"00",
          7593 => x"55",
          7594 => x"20",
          7595 => x"20",
          7596 => x"20",
          7597 => x"00",
          7598 => x"73",
          7599 => x"63",
          7600 => x"20",
          7601 => x"20",
          7602 => x"4d",
          7603 => x"20",
          7604 => x"6e",
          7605 => x"20",
          7606 => x"72",
          7607 => x"25",
          7608 => x"00",
          7609 => x"52",
          7610 => x"6b",
          7611 => x"20",
          7612 => x"20",
          7613 => x"4d",
          7614 => x"20",
          7615 => x"20",
          7616 => x"20",
          7617 => x"00",
          7618 => x"20",
          7619 => x"20",
          7620 => x"4e",
          7621 => x"00",
          7622 => x"54",
          7623 => x"28",
          7624 => x"73",
          7625 => x"0a",
          7626 => x"4d",
          7627 => x"28",
          7628 => x"20",
          7629 => x"0a",
          7630 => x"20",
          7631 => x"28",
          7632 => x"20",
          7633 => x"0a",
          7634 => x"4d",
          7635 => x"28",
          7636 => x"38",
          7637 => x"20",
          7638 => x"20",
          7639 => x"58",
          7640 => x"0a",
          7641 => x"53",
          7642 => x"28",
          7643 => x"38",
          7644 => x"20",
          7645 => x"20",
          7646 => x"58",
          7647 => x"0a",
          7648 => x"20",
          7649 => x"28",
          7650 => x"38",
          7651 => x"66",
          7652 => x"20",
          7653 => x"00",
          7654 => x"6e",
          7655 => x"00",
          7656 => x"00",
          7657 => x"00",
          7658 => x"00",
          7659 => x"f0",
          7660 => x"00",
          7661 => x"00",
          7662 => x"f0",
          7663 => x"00",
          7664 => x"00",
          7665 => x"f0",
          7666 => x"00",
          7667 => x"00",
          7668 => x"f0",
          7669 => x"00",
          7670 => x"00",
          7671 => x"f0",
          7672 => x"00",
          7673 => x"00",
          7674 => x"f0",
          7675 => x"00",
          7676 => x"00",
          7677 => x"f0",
          7678 => x"00",
          7679 => x"00",
          7680 => x"f0",
          7681 => x"00",
          7682 => x"00",
          7683 => x"f0",
          7684 => x"00",
          7685 => x"00",
          7686 => x"f0",
          7687 => x"00",
          7688 => x"00",
          7689 => x"f0",
          7690 => x"00",
          7691 => x"00",
          7692 => x"44",
          7693 => x"42",
          7694 => x"36",
          7695 => x"34",
          7696 => x"33",
          7697 => x"31",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"00",
          7703 => x"6e",
          7704 => x"6e",
          7705 => x"20",
          7706 => x"20",
          7707 => x"69",
          7708 => x"2e",
          7709 => x"79",
          7710 => x"00",
          7711 => x"36",
          7712 => x"00",
          7713 => x"20",
          7714 => x"74",
          7715 => x"73",
          7716 => x"6c",
          7717 => x"46",
          7718 => x"73",
          7719 => x"31",
          7720 => x"41",
          7721 => x"43",
          7722 => x"31",
          7723 => x"31",
          7724 => x"31",
          7725 => x"31",
          7726 => x"31",
          7727 => x"31",
          7728 => x"31",
          7729 => x"31",
          7730 => x"31",
          7731 => x"32",
          7732 => x"32",
          7733 => x"33",
          7734 => x"46",
          7735 => x"00",
          7736 => x"00",
          7737 => x"64",
          7738 => x"25",
          7739 => x"32",
          7740 => x"25",
          7741 => x"3a",
          7742 => x"64",
          7743 => x"2c",
          7744 => x"00",
          7745 => x"00",
          7746 => x"25",
          7747 => x"70",
          7748 => x"73",
          7749 => x"3a",
          7750 => x"32",
          7751 => x"3a",
          7752 => x"32",
          7753 => x"3a",
          7754 => x"00",
          7755 => x"69",
          7756 => x"6e",
          7757 => x"64",
          7758 => x"53",
          7759 => x"00",
          7760 => x"69",
          7761 => x"72",
          7762 => x"20",
          7763 => x"66",
          7764 => x"00",
          7765 => x"3a",
          7766 => x"00",
          7767 => x"00",
          7768 => x"54",
          7769 => x"90",
          7770 => x"30",
          7771 => x"45",
          7772 => x"20",
          7773 => x"20",
          7774 => x"20",
          7775 => x"20",
          7776 => x"00",
          7777 => x"00",
          7778 => x"10",
          7779 => x"00",
          7780 => x"8f",
          7781 => x"8e",
          7782 => x"55",
          7783 => x"9e",
          7784 => x"a6",
          7785 => x"ae",
          7786 => x"b6",
          7787 => x"be",
          7788 => x"c6",
          7789 => x"ce",
          7790 => x"d6",
          7791 => x"de",
          7792 => x"e6",
          7793 => x"ee",
          7794 => x"f6",
          7795 => x"fe",
          7796 => x"5d",
          7797 => x"3f",
          7798 => x"00",
          7799 => x"02",
          7800 => x"00",
          7801 => x"00",
          7802 => x"00",
          7803 => x"00",
          7804 => x"00",
          7805 => x"00",
          7806 => x"00",
          7807 => x"00",
          7808 => x"00",
          7809 => x"00",
          7810 => x"00",
          7811 => x"00",
          7812 => x"23",
          7813 => x"00",
          7814 => x"25",
          7815 => x"25",
          7816 => x"25",
          7817 => x"25",
          7818 => x"25",
          7819 => x"25",
          7820 => x"25",
          7821 => x"25",
          7822 => x"25",
          7823 => x"25",
          7824 => x"25",
          7825 => x"25",
          7826 => x"00",
          7827 => x"03",
          7828 => x"03",
          7829 => x"03",
          7830 => x"00",
          7831 => x"23",
          7832 => x"22",
          7833 => x"00",
          7834 => x"03",
          7835 => x"03",
          7836 => x"01",
          7837 => x"01",
          7838 => x"01",
          7839 => x"02",
          7840 => x"01",
          7841 => x"01",
          7842 => x"01",
          7843 => x"01",
          7844 => x"01",
          7845 => x"01",
          7846 => x"01",
          7847 => x"01",
          7848 => x"01",
          7849 => x"01",
          7850 => x"01",
          7851 => x"01",
          7852 => x"01",
          7853 => x"01",
          7854 => x"01",
          7855 => x"01",
          7856 => x"01",
          7857 => x"01",
          7858 => x"01",
          7859 => x"00",
          7860 => x"01",
          7861 => x"01",
          7862 => x"01",
          7863 => x"02",
          7864 => x"02",
          7865 => x"02",
          7866 => x"01",
          7867 => x"01",
          7868 => x"01",
          7869 => x"02",
          7870 => x"01",
          7871 => x"02",
          7872 => x"2c",
          7873 => x"01",
          7874 => x"02",
          7875 => x"02",
          7876 => x"02",
          7877 => x"02",
          7878 => x"01",
          7879 => x"02",
          7880 => x"01",
          7881 => x"02",
          7882 => x"03",
          7883 => x"03",
          7884 => x"03",
          7885 => x"03",
          7886 => x"03",
          7887 => x"00",
          7888 => x"03",
          7889 => x"03",
          7890 => x"03",
          7891 => x"03",
          7892 => x"04",
          7893 => x"04",
          7894 => x"04",
          7895 => x"01",
          7896 => x"00",
          7897 => x"1e",
          7898 => x"1f",
          7899 => x"1f",
          7900 => x"1f",
          7901 => x"1f",
          7902 => x"1f",
          7903 => x"06",
          7904 => x"1f",
          7905 => x"1f",
          7906 => x"1f",
          7907 => x"1f",
          7908 => x"06",
          7909 => x"00",
          7910 => x"1f",
          7911 => x"1f",
          7912 => x"1f",
          7913 => x"00",
          7914 => x"21",
          7915 => x"00",
          7916 => x"2c",
          7917 => x"2c",
          7918 => x"2c",
          7919 => x"ff",
          7920 => x"00",
          7921 => x"01",
          7922 => x"00",
          7923 => x"01",
          7924 => x"00",
          7925 => x"03",
          7926 => x"00",
          7927 => x"03",
          7928 => x"00",
          7929 => x"03",
          7930 => x"00",
          7931 => x"04",
          7932 => x"00",
          7933 => x"04",
          7934 => x"00",
          7935 => x"04",
          7936 => x"00",
          7937 => x"04",
          7938 => x"00",
          7939 => x"04",
          7940 => x"00",
          7941 => x"04",
          7942 => x"00",
          7943 => x"04",
          7944 => x"00",
          7945 => x"05",
          7946 => x"00",
          7947 => x"05",
          7948 => x"00",
          7949 => x"05",
          7950 => x"00",
          7951 => x"05",
          7952 => x"00",
          7953 => x"07",
          7954 => x"00",
          7955 => x"07",
          7956 => x"00",
          7957 => x"08",
          7958 => x"00",
          7959 => x"08",
          7960 => x"00",
          7961 => x"08",
          7962 => x"00",
          7963 => x"08",
          7964 => x"00",
          7965 => x"08",
          7966 => x"00",
          7967 => x"08",
          7968 => x"00",
          7969 => x"09",
          7970 => x"00",
          7971 => x"09",
          7972 => x"00",
          7973 => x"09",
          7974 => x"00",
          7975 => x"09",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"00",
          7983 => x"78",
          7984 => x"e1",
          7985 => x"e1",
          7986 => x"01",
          7987 => x"10",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"00",
          7996 => x"00",
          7997 => x"00",
          7998 => x"00",
          7999 => x"00",
          8000 => x"f0",
          8001 => x"f0",
          8002 => x"f0",
          8003 => x"fd",
          8004 => x"3a",
          8005 => x"f0",
          8006 => x"77",
          8007 => x"6f",
          8008 => x"67",
          8009 => x"37",
          8010 => x"2c",
          8011 => x"3f",
          8012 => x"f0",
          8013 => x"f0",
          8014 => x"3b",
          8015 => x"f0",
          8016 => x"57",
          8017 => x"4f",
          8018 => x"47",
          8019 => x"37",
          8020 => x"2c",
          8021 => x"3f",
          8022 => x"f0",
          8023 => x"f0",
          8024 => x"2a",
          8025 => x"f0",
          8026 => x"57",
          8027 => x"4f",
          8028 => x"47",
          8029 => x"27",
          8030 => x"3c",
          8031 => x"3f",
          8032 => x"f0",
          8033 => x"f0",
          8034 => x"f0",
          8035 => x"f0",
          8036 => x"17",
          8037 => x"0f",
          8038 => x"07",
          8039 => x"f0",
          8040 => x"f0",
          8041 => x"f0",
          8042 => x"f0",
          8043 => x"f0",
          8044 => x"4d",
          8045 => x"f0",
          8046 => x"78",
          8047 => x"d5",
          8048 => x"4c",
          8049 => x"5f",
          8050 => x"d0",
          8051 => x"bb",
          8052 => x"f0",
          8053 => x"f0",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"01",
          9089 => x"f2",
          9090 => x"fa",
          9091 => x"c2",
          9092 => x"e5",
          9093 => x"62",
          9094 => x"6b",
          9095 => x"22",
          9096 => x"4f",
          9097 => x"02",
          9098 => x"0a",
          9099 => x"12",
          9100 => x"1a",
          9101 => x"82",
          9102 => x"8a",
          9103 => x"92",
          9104 => x"9a",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"00",
          9113 => x"00",
          9114 => x"00",
          9115 => x"00",
          9116 => x"00",
          9117 => x"00",
          9118 => x"00",
          9119 => x"00",
          9120 => x"00",
          9121 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"93",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"2d",
             6 => x"00",
             7 => x"00",
             8 => x"fd",
             9 => x"05",
            10 => x"ff",
            11 => x"00",
            12 => x"fd",
            13 => x"06",
            14 => x"2b",
            15 => x"0b",
            16 => x"09",
            17 => x"06",
            18 => x"0a",
            19 => x"00",
            20 => x"72",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"73",
            25 => x"81",
            26 => x"10",
            27 => x"51",
            28 => x"72",
            29 => x"04",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"0a",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"72",
            45 => x"0b",
            46 => x"00",
            47 => x"00",
            48 => x"72",
            49 => x"74",
            50 => x"07",
            51 => x"00",
            52 => x"71",
            53 => x"09",
            54 => x"2b",
            55 => x"04",
            56 => x"09",
            57 => x"05",
            58 => x"04",
            59 => x"00",
            60 => x"09",
            61 => x"05",
            62 => x"51",
            63 => x"00",
            64 => x"09",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"72",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"09",
            73 => x"53",
            74 => x"00",
            75 => x"00",
            76 => x"fc",
            77 => x"05",
            78 => x"ff",
            79 => x"00",
            80 => x"fc",
            81 => x"73",
            82 => x"0b",
            83 => x"00",
            84 => x"08",
            85 => x"0b",
            86 => x"08",
            87 => x"51",
            88 => x"08",
            89 => x"0b",
            90 => x"08",
            91 => x"51",
            92 => x"09",
            93 => x"06",
            94 => x"09",
            95 => x"51",
            96 => x"09",
            97 => x"81",
            98 => x"73",
            99 => x"07",
           100 => x"ff",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"81",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"84",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"0d",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"8c",
           134 => x"04",
           135 => x"0b",
           136 => x"8c",
           137 => x"04",
           138 => x"0b",
           139 => x"8d",
           140 => x"04",
           141 => x"0b",
           142 => x"8d",
           143 => x"04",
           144 => x"0b",
           145 => x"8e",
           146 => x"04",
           147 => x"0b",
           148 => x"8e",
           149 => x"04",
           150 => x"0b",
           151 => x"8f",
           152 => x"04",
           153 => x"0b",
           154 => x"8f",
           155 => x"04",
           156 => x"0b",
           157 => x"90",
           158 => x"04",
           159 => x"0b",
           160 => x"90",
           161 => x"04",
           162 => x"0b",
           163 => x"91",
           164 => x"04",
           165 => x"0b",
           166 => x"91",
           167 => x"04",
           168 => x"0b",
           169 => x"92",
           170 => x"04",
           171 => x"0b",
           172 => x"92",
           173 => x"04",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"00",
           193 => x"80",
           194 => x"80",
           195 => x"0c",
           196 => x"80",
           197 => x"0c",
           198 => x"80",
           199 => x"0c",
           200 => x"80",
           201 => x"0c",
           202 => x"80",
           203 => x"0c",
           204 => x"80",
           205 => x"0c",
           206 => x"80",
           207 => x"0c",
           208 => x"80",
           209 => x"0c",
           210 => x"80",
           211 => x"0c",
           212 => x"80",
           213 => x"0c",
           214 => x"80",
           215 => x"0c",
           216 => x"80",
           217 => x"0c",
           218 => x"08",
           219 => x"98",
           220 => x"98",
           221 => x"ba",
           222 => x"ba",
           223 => x"84",
           224 => x"84",
           225 => x"04",
           226 => x"2d",
           227 => x"90",
           228 => x"c9",
           229 => x"80",
           230 => x"d2",
           231 => x"c0",
           232 => x"82",
           233 => x"80",
           234 => x"0c",
           235 => x"08",
           236 => x"98",
           237 => x"98",
           238 => x"ba",
           239 => x"ba",
           240 => x"84",
           241 => x"84",
           242 => x"04",
           243 => x"2d",
           244 => x"90",
           245 => x"a9",
           246 => x"80",
           247 => x"84",
           248 => x"c0",
           249 => x"82",
           250 => x"80",
           251 => x"0c",
           252 => x"08",
           253 => x"98",
           254 => x"98",
           255 => x"ba",
           256 => x"ba",
           257 => x"84",
           258 => x"84",
           259 => x"04",
           260 => x"2d",
           261 => x"90",
           262 => x"b0",
           263 => x"80",
           264 => x"e7",
           265 => x"c0",
           266 => x"82",
           267 => x"80",
           268 => x"0c",
           269 => x"08",
           270 => x"98",
           271 => x"98",
           272 => x"ba",
           273 => x"ba",
           274 => x"84",
           275 => x"84",
           276 => x"04",
           277 => x"2d",
           278 => x"90",
           279 => x"dc",
           280 => x"80",
           281 => x"b8",
           282 => x"c0",
           283 => x"81",
           284 => x"80",
           285 => x"0c",
           286 => x"08",
           287 => x"98",
           288 => x"98",
           289 => x"ba",
           290 => x"ba",
           291 => x"84",
           292 => x"84",
           293 => x"04",
           294 => x"2d",
           295 => x"90",
           296 => x"2d",
           297 => x"90",
           298 => x"ca",
           299 => x"80",
           300 => x"dd",
           301 => x"c0",
           302 => x"81",
           303 => x"80",
           304 => x"0c",
           305 => x"08",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"51",
           311 => x"73",
           312 => x"10",
           313 => x"0c",
           314 => x"81",
           315 => x"71",
           316 => x"72",
           317 => x"84",
           318 => x"8e",
           319 => x"0c",
           320 => x"81",
           321 => x"3d",
           322 => x"52",
           323 => x"f0",
           324 => x"0d",
           325 => x"85",
           326 => x"73",
           327 => x"52",
           328 => x"d3",
           329 => x"70",
           330 => x"55",
           331 => x"38",
           332 => x"8e",
           333 => x"84",
           334 => x"84",
           335 => x"57",
           336 => x"30",
           337 => x"54",
           338 => x"75",
           339 => x"0c",
           340 => x"ba",
           341 => x"3d",
           342 => x"99",
           343 => x"8e",
           344 => x"3d",
           345 => x"54",
           346 => x"fd",
           347 => x"76",
           348 => x"0d",
           349 => x"42",
           350 => x"85",
           351 => x"81",
           352 => x"7b",
           353 => x"7b",
           354 => x"38",
           355 => x"72",
           356 => x"5f",
           357 => x"b0",
           358 => x"54",
           359 => x"a9",
           360 => x"81",
           361 => x"38",
           362 => x"57",
           363 => x"54",
           364 => x"0d",
           365 => x"10",
           366 => x"70",
           367 => x"29",
           368 => x"5a",
           369 => x"86",
           370 => x"bd",
           371 => x"fe",
           372 => x"2e",
           373 => x"74",
           374 => x"5a",
           375 => x"7c",
           376 => x"33",
           377 => x"39",
           378 => x"55",
           379 => x"40",
           380 => x"72",
           381 => x"10",
           382 => x"04",
           383 => x"73",
           384 => x"8a",
           385 => x"76",
           386 => x"ff",
           387 => x"60",
           388 => x"cf",
           389 => x"9c",
           390 => x"3f",
           391 => x"84",
           392 => x"53",
           393 => x"8c",
           394 => x"81",
           395 => x"90",
           396 => x"84",
           397 => x"ba",
           398 => x"40",
           399 => x"84",
           400 => x"70",
           401 => x"70",
           402 => x"9e",
           403 => x"80",
           404 => x"38",
           405 => x"80",
           406 => x"83",
           407 => x"80",
           408 => x"81",
           409 => x"86",
           410 => x"70",
           411 => x"5b",
           412 => x"85",
           413 => x"70",
           414 => x"59",
           415 => x"7a",
           416 => x"eb",
           417 => x"73",
           418 => x"06",
           419 => x"06",
           420 => x"2a",
           421 => x"38",
           422 => x"80",
           423 => x"54",
           424 => x"b0",
           425 => x"80",
           426 => x"90",
           427 => x"e5",
           428 => x"2e",
           429 => x"29",
           430 => x"5b",
           431 => x"7c",
           432 => x"79",
           433 => x"05",
           434 => x"80",
           435 => x"81",
           436 => x"b9",
           437 => x"38",
           438 => x"76",
           439 => x"84",
           440 => x"ff",
           441 => x"3f",
           442 => x"06",
           443 => x"80",
           444 => x"80",
           445 => x"90",
           446 => x"fc",
           447 => x"f4",
           448 => x"7a",
           449 => x"fa",
           450 => x"c0",
           451 => x"61",
           452 => x"cf",
           453 => x"fd",
           454 => x"80",
           455 => x"2b",
           456 => x"fc",
           457 => x"52",
           458 => x"2a",
           459 => x"c9",
           460 => x"fc",
           461 => x"54",
           462 => x"7c",
           463 => x"39",
           464 => x"5b",
           465 => x"ca",
           466 => x"57",
           467 => x"ff",
           468 => x"54",
           469 => x"38",
           470 => x"33",
           471 => x"fc",
           472 => x"84",
           473 => x"70",
           474 => x"7b",
           475 => x"57",
           476 => x"7f",
           477 => x"40",
           478 => x"38",
           479 => x"ba",
           480 => x"07",
           481 => x"38",
           482 => x"80",
           483 => x"38",
           484 => x"71",
           485 => x"5f",
           486 => x"f6",
           487 => x"ff",
           488 => x"5a",
           489 => x"7a",
           490 => x"76",
           491 => x"60",
           492 => x"5d",
           493 => x"75",
           494 => x"08",
           495 => x"90",
           496 => x"80",
           497 => x"88",
           498 => x"80",
           499 => x"90",
           500 => x"fa",
           501 => x"c4",
           502 => x"83",
           503 => x"06",
           504 => x"83",
           505 => x"5f",
           506 => x"d8",
           507 => x"90",
           508 => x"06",
           509 => x"38",
           510 => x"82",
           511 => x"80",
           512 => x"7c",
           513 => x"3f",
           514 => x"f7",
           515 => x"31",
           516 => x"f9",
           517 => x"c4",
           518 => x"82",
           519 => x"75",
           520 => x"08",
           521 => x"90",
           522 => x"82",
           523 => x"06",
           524 => x"3d",
           525 => x"52",
           526 => x"0d",
           527 => x"0b",
           528 => x"70",
           529 => x"51",
           530 => x"77",
           531 => x"74",
           532 => x"77",
           533 => x"52",
           534 => x"2d",
           535 => x"38",
           536 => x"33",
           537 => x"d5",
           538 => x"f0",
           539 => x"8a",
           540 => x"84",
           541 => x"ff",
           542 => x"0c",
           543 => x"78",
           544 => x"33",
           545 => x"06",
           546 => x"77",
           547 => x"70",
           548 => x"2e",
           549 => x"75",
           550 => x"04",
           551 => x"72",
           552 => x"51",
           553 => x"ba",
           554 => x"74",
           555 => x"72",
           556 => x"84",
           557 => x"3f",
           558 => x"78",
           559 => x"81",
           560 => x"ff",
           561 => x"81",
           562 => x"8c",
           563 => x"25",
           564 => x"34",
           565 => x"15",
           566 => x"76",
           567 => x"3d",
           568 => x"06",
           569 => x"ff",
           570 => x"8c",
           571 => x"76",
           572 => x"85",
           573 => x"81",
           574 => x"ff",
           575 => x"81",
           576 => x"2a",
           577 => x"c3",
           578 => x"71",
           579 => x"76",
           580 => x"17",
           581 => x"84",
           582 => x"74",
           583 => x"34",
           584 => x"0c",
           585 => x"87",
           586 => x"08",
           587 => x"52",
           588 => x"b9",
           589 => x"54",
           590 => x"85",
           591 => x"17",
           592 => x"0c",
           593 => x"53",
           594 => x"39",
           595 => x"54",
           596 => x"51",
           597 => x"70",
           598 => x"70",
           599 => x"73",
           600 => x"04",
           601 => x"55",
           602 => x"38",
           603 => x"2e",
           604 => x"33",
           605 => x"11",
           606 => x"8c",
           607 => x"55",
           608 => x"75",
           609 => x"53",
           610 => x"70",
           611 => x"13",
           612 => x"11",
           613 => x"3d",
           614 => x"81",
           615 => x"ff",
           616 => x"0c",
           617 => x"0d",
           618 => x"70",
           619 => x"70",
           620 => x"73",
           621 => x"04",
           622 => x"55",
           623 => x"38",
           624 => x"70",
           625 => x"70",
           626 => x"85",
           627 => x"78",
           628 => x"a1",
           629 => x"57",
           630 => x"81",
           631 => x"80",
           632 => x"e1",
           633 => x"0c",
           634 => x"f1",
           635 => x"80",
           636 => x"81",
           637 => x"72",
           638 => x"0d",
           639 => x"3d",
           640 => x"53",
           641 => x"ba",
           642 => x"05",
           643 => x"ba",
           644 => x"80",
           645 => x"15",
           646 => x"52",
           647 => x"3f",
           648 => x"ba",
           649 => x"3d",
           650 => x"53",
           651 => x"70",
           652 => x"2e",
           653 => x"2e",
           654 => x"70",
           655 => x"8c",
           656 => x"0d",
           657 => x"54",
           658 => x"70",
           659 => x"70",
           660 => x"85",
           661 => x"7a",
           662 => x"8b",
           663 => x"ba",
           664 => x"80",
           665 => x"3f",
           666 => x"80",
           667 => x"73",
           668 => x"81",
           669 => x"76",
           670 => x"56",
           671 => x"74",
           672 => x"78",
           673 => x"81",
           674 => x"ff",
           675 => x"55",
           676 => x"07",
           677 => x"3d",
           678 => x"fc",
           679 => x"07",
           680 => x"31",
           681 => x"06",
           682 => x"88",
           683 => x"f0",
           684 => x"2b",
           685 => x"53",
           686 => x"30",
           687 => x"77",
           688 => x"70",
           689 => x"06",
           690 => x"51",
           691 => x"53",
           692 => x"56",
           693 => x"0d",
           694 => x"54",
           695 => x"84",
           696 => x"31",
           697 => x"0d",
           698 => x"54",
           699 => x"76",
           700 => x"08",
           701 => x"8d",
           702 => x"84",
           703 => x"71",
           704 => x"71",
           705 => x"71",
           706 => x"57",
           707 => x"2e",
           708 => x"07",
           709 => x"ff",
           710 => x"72",
           711 => x"56",
           712 => x"da",
           713 => x"3d",
           714 => x"2c",
           715 => x"32",
           716 => x"32",
           717 => x"56",
           718 => x"3f",
           719 => x"31",
           720 => x"04",
           721 => x"80",
           722 => x"56",
           723 => x"06",
           724 => x"70",
           725 => x"38",
           726 => x"b0",
           727 => x"80",
           728 => x"8a",
           729 => x"c4",
           730 => x"e0",
           731 => x"d0",
           732 => x"90",
           733 => x"81",
           734 => x"81",
           735 => x"38",
           736 => x"79",
           737 => x"a0",
           738 => x"84",
           739 => x"81",
           740 => x"3d",
           741 => x"0c",
           742 => x"2e",
           743 => x"15",
           744 => x"73",
           745 => x"73",
           746 => x"a0",
           747 => x"80",
           748 => x"e1",
           749 => x"3d",
           750 => x"78",
           751 => x"fe",
           752 => x"0c",
           753 => x"7b",
           754 => x"77",
           755 => x"a0",
           756 => x"15",
           757 => x"73",
           758 => x"80",
           759 => x"38",
           760 => x"26",
           761 => x"a0",
           762 => x"74",
           763 => x"ff",
           764 => x"ff",
           765 => x"38",
           766 => x"54",
           767 => x"78",
           768 => x"13",
           769 => x"56",
           770 => x"38",
           771 => x"56",
           772 => x"ba",
           773 => x"70",
           774 => x"56",
           775 => x"fe",
           776 => x"70",
           777 => x"a6",
           778 => x"a0",
           779 => x"38",
           780 => x"89",
           781 => x"ba",
           782 => x"58",
           783 => x"55",
           784 => x"0b",
           785 => x"04",
           786 => x"08",
           787 => x"04",
           788 => x"26",
           789 => x"cc",
           790 => x"e4",
           791 => x"04",
           792 => x"83",
           793 => x"ef",
           794 => x"cf",
           795 => x"0d",
           796 => x"3f",
           797 => x"51",
           798 => x"83",
           799 => x"3d",
           800 => x"f1",
           801 => x"a4",
           802 => x"04",
           803 => x"83",
           804 => x"ee",
           805 => x"d0",
           806 => x"0d",
           807 => x"3f",
           808 => x"51",
           809 => x"83",
           810 => x"3d",
           811 => x"99",
           812 => x"d0",
           813 => x"04",
           814 => x"83",
           815 => x"ed",
           816 => x"d2",
           817 => x"0d",
           818 => x"3f",
           819 => x"66",
           820 => x"5b",
           821 => x"07",
           822 => x"57",
           823 => x"57",
           824 => x"51",
           825 => x"81",
           826 => x"58",
           827 => x"08",
           828 => x"80",
           829 => x"3f",
           830 => x"7b",
           831 => x"57",
           832 => x"87",
           833 => x"e7",
           834 => x"87",
           835 => x"ba",
           836 => x"78",
           837 => x"3f",
           838 => x"0d",
           839 => x"98",
           840 => x"96",
           841 => x"75",
           842 => x"84",
           843 => x"08",
           844 => x"2e",
           845 => x"57",
           846 => x"51",
           847 => x"52",
           848 => x"8c",
           849 => x"52",
           850 => x"ff",
           851 => x"84",
           852 => x"58",
           853 => x"ec",
           854 => x"76",
           855 => x"8a",
           856 => x"3d",
           857 => x"56",
           858 => x"53",
           859 => x"ba",
           860 => x"3d",
           861 => x"63",
           862 => x"73",
           863 => x"5f",
           864 => x"38",
           865 => x"fe",
           866 => x"3f",
           867 => x"7c",
           868 => x"2e",
           869 => x"7a",
           870 => x"83",
           871 => x"14",
           872 => x"51",
           873 => x"38",
           874 => x"80",
           875 => x"75",
           876 => x"72",
           877 => x"53",
           878 => x"74",
           879 => x"57",
           880 => x"74",
           881 => x"08",
           882 => x"16",
           883 => x"d2",
           884 => x"79",
           885 => x"3f",
           886 => x"98",
           887 => x"ee",
           888 => x"7b",
           889 => x"38",
           890 => x"3d",
           891 => x"ae",
           892 => x"53",
           893 => x"74",
           894 => x"83",
           895 => x"14",
           896 => x"51",
           897 => x"c0",
           898 => x"df",
           899 => x"51",
           900 => x"f0",
           901 => x"3f",
           902 => x"39",
           903 => x"84",
           904 => x"a0",
           905 => x"fd",
           906 => x"27",
           907 => x"c4",
           908 => x"d5",
           909 => x"84",
           910 => x"d8",
           911 => x"51",
           912 => x"91",
           913 => x"8c",
           914 => x"72",
           915 => x"72",
           916 => x"e0",
           917 => x"51",
           918 => x"98",
           919 => x"70",
           920 => x"72",
           921 => x"58",
           922 => x"fd",
           923 => x"84",
           924 => x"2c",
           925 => x"32",
           926 => x"07",
           927 => x"53",
           928 => x"b9",
           929 => x"8f",
           930 => x"c0",
           931 => x"81",
           932 => x"51",
           933 => x"3f",
           934 => x"52",
           935 => x"70",
           936 => x"38",
           937 => x"52",
           938 => x"70",
           939 => x"38",
           940 => x"52",
           941 => x"70",
           942 => x"38",
           943 => x"52",
           944 => x"06",
           945 => x"84",
           946 => x"3f",
           947 => x"80",
           948 => x"84",
           949 => x"3f",
           950 => x"80",
           951 => x"81",
           952 => x"cb",
           953 => x"d3",
           954 => x"9b",
           955 => x"06",
           956 => x"38",
           957 => x"83",
           958 => x"51",
           959 => x"81",
           960 => x"f0",
           961 => x"8a",
           962 => x"3f",
           963 => x"2a",
           964 => x"2e",
           965 => x"51",
           966 => x"9a",
           967 => x"72",
           968 => x"71",
           969 => x"39",
           970 => x"c4",
           971 => x"ba",
           972 => x"51",
           973 => x"ff",
           974 => x"83",
           975 => x"51",
           976 => x"81",
           977 => x"b8",
           978 => x"80",
           979 => x"98",
           980 => x"b6",
           981 => x"ff",
           982 => x"2e",
           983 => x"e3",
           984 => x"e0",
           985 => x"f8",
           986 => x"3f",
           987 => x"81",
           988 => x"82",
           989 => x"38",
           990 => x"2e",
           991 => x"79",
           992 => x"5c",
           993 => x"38",
           994 => x"a0",
           995 => x"26",
           996 => x"84",
           997 => x"3f",
           998 => x"08",
           999 => x"e8",
          1000 => x"38",
          1001 => x"83",
          1002 => x"06",
          1003 => x"9a",
          1004 => x"dd",
          1005 => x"92",
          1006 => x"ba",
          1007 => x"84",
          1008 => x"80",
          1009 => x"8c",
          1010 => x"80",
          1011 => x"08",
          1012 => x"08",
          1013 => x"a5",
          1014 => x"8f",
          1015 => x"7a",
          1016 => x"80",
          1017 => x"d5",
          1018 => x"ba",
          1019 => x"54",
          1020 => x"52",
          1021 => x"8c",
          1022 => x"30",
          1023 => x"5b",
          1024 => x"38",
          1025 => x"80",
          1026 => x"ff",
          1027 => x"7f",
          1028 => x"7c",
          1029 => x"f2",
          1030 => x"83",
          1031 => x"48",
          1032 => x"e8",
          1033 => x"33",
          1034 => x"fd",
          1035 => x"52",
          1036 => x"3f",
          1037 => x"81",
          1038 => x"84",
          1039 => x"51",
          1040 => x"08",
          1041 => x"08",
          1042 => x"ef",
          1043 => x"59",
          1044 => x"d3",
          1045 => x"82",
          1046 => x"83",
          1047 => x"80",
          1048 => x"67",
          1049 => x"90",
          1050 => x"33",
          1051 => x"38",
          1052 => x"5a",
          1053 => x"df",
          1054 => x"83",
          1055 => x"3f",
          1056 => x"51",
          1057 => x"08",
          1058 => x"38",
          1059 => x"fb",
          1060 => x"d1",
          1061 => x"fe",
          1062 => x"55",
          1063 => x"d6",
          1064 => x"fd",
          1065 => x"f5",
          1066 => x"81",
          1067 => x"e5",
          1068 => x"39",
          1069 => x"80",
          1070 => x"de",
          1071 => x"39",
          1072 => x"80",
          1073 => x"8c",
          1074 => x"52",
          1075 => x"68",
          1076 => x"80",
          1077 => x"08",
          1078 => x"3f",
          1079 => x"11",
          1080 => x"3f",
          1081 => x"f5",
          1082 => x"d0",
          1083 => x"3d",
          1084 => x"51",
          1085 => x"80",
          1086 => x"f0",
          1087 => x"88",
          1088 => x"38",
          1089 => x"83",
          1090 => x"d5",
          1091 => x"51",
          1092 => x"59",
          1093 => x"9f",
          1094 => x"70",
          1095 => x"f4",
          1096 => x"c0",
          1097 => x"f8",
          1098 => x"53",
          1099 => x"84",
          1100 => x"59",
          1101 => x"c0",
          1102 => x"08",
          1103 => x"a9",
          1104 => x"ae",
          1105 => x"87",
          1106 => x"59",
          1107 => x"53",
          1108 => x"84",
          1109 => x"38",
          1110 => x"80",
          1111 => x"8c",
          1112 => x"3d",
          1113 => x"51",
          1114 => x"80",
          1115 => x"51",
          1116 => x"78",
          1117 => x"33",
          1118 => x"2e",
          1119 => x"33",
          1120 => x"ce",
          1121 => x"19",
          1122 => x"3d",
          1123 => x"51",
          1124 => x"80",
          1125 => x"fc",
          1126 => x"d4",
          1127 => x"f7",
          1128 => x"53",
          1129 => x"84",
          1130 => x"38",
          1131 => x"68",
          1132 => x"65",
          1133 => x"7c",
          1134 => x"b8",
          1135 => x"05",
          1136 => x"08",
          1137 => x"fe",
          1138 => x"e7",
          1139 => x"38",
          1140 => x"84",
          1141 => x"08",
          1142 => x"f1",
          1143 => x"ae",
          1144 => x"84",
          1145 => x"39",
          1146 => x"79",
          1147 => x"fe",
          1148 => x"e7",
          1149 => x"2e",
          1150 => x"db",
          1151 => x"49",
          1152 => x"80",
          1153 => x"8c",
          1154 => x"b8",
          1155 => x"05",
          1156 => x"08",
          1157 => x"fe",
          1158 => x"e6",
          1159 => x"2e",
          1160 => x"11",
          1161 => x"3f",
          1162 => x"ba",
          1163 => x"cb",
          1164 => x"7a",
          1165 => x"70",
          1166 => x"f5",
          1167 => x"c5",
          1168 => x"87",
          1169 => x"3d",
          1170 => x"3f",
          1171 => x"78",
          1172 => x"08",
          1173 => x"8c",
          1174 => x"39",
          1175 => x"80",
          1176 => x"8c",
          1177 => x"5a",
          1178 => x"f2",
          1179 => x"11",
          1180 => x"3f",
          1181 => x"f3",
          1182 => x"8a",
          1183 => x"3d",
          1184 => x"51",
          1185 => x"80",
          1186 => x"7a",
          1187 => x"90",
          1188 => x"2a",
          1189 => x"2e",
          1190 => x"88",
          1191 => x"3f",
          1192 => x"52",
          1193 => x"ac",
          1194 => x"64",
          1195 => x"45",
          1196 => x"80",
          1197 => x"8c",
          1198 => x"64",
          1199 => x"b8",
          1200 => x"05",
          1201 => x"08",
          1202 => x"02",
          1203 => x"05",
          1204 => x"f0",
          1205 => x"d8",
          1206 => x"f2",
          1207 => x"05",
          1208 => x"7d",
          1209 => x"ff",
          1210 => x"ba",
          1211 => x"39",
          1212 => x"80",
          1213 => x"8c",
          1214 => x"5c",
          1215 => x"68",
          1216 => x"3d",
          1217 => x"51",
          1218 => x"80",
          1219 => x"0c",
          1220 => x"f7",
          1221 => x"06",
          1222 => x"98",
          1223 => x"7c",
          1224 => x"7b",
          1225 => x"82",
          1226 => x"3f",
          1227 => x"11",
          1228 => x"3f",
          1229 => x"38",
          1230 => x"79",
          1231 => x"f7",
          1232 => x"7b",
          1233 => x"d4",
          1234 => x"91",
          1235 => x"83",
          1236 => x"83",
          1237 => x"59",
          1238 => x"d3",
          1239 => x"83",
          1240 => x"a5",
          1241 => x"8b",
          1242 => x"3f",
          1243 => x"59",
          1244 => x"dc",
          1245 => x"93",
          1246 => x"83",
          1247 => x"83",
          1248 => x"9b",
          1249 => x"ee",
          1250 => x"80",
          1251 => x"49",
          1252 => x"5d",
          1253 => x"ec",
          1254 => x"f8",
          1255 => x"39",
          1256 => x"fb",
          1257 => x"84",
          1258 => x"70",
          1259 => x"74",
          1260 => x"08",
          1261 => x"84",
          1262 => x"74",
          1263 => x"87",
          1264 => x"87",
          1265 => x"3f",
          1266 => x"08",
          1267 => x"51",
          1268 => x"08",
          1269 => x"87",
          1270 => x"0b",
          1271 => x"ec",
          1272 => x"84",
          1273 => x"d5",
          1274 => x"0c",
          1275 => x"56",
          1276 => x"87",
          1277 => x"83",
          1278 => x"c4",
          1279 => x"52",
          1280 => x"54",
          1281 => x"52",
          1282 => x"8d",
          1283 => x"fb",
          1284 => x"80",
          1285 => x"83",
          1286 => x"52",
          1287 => x"91",
          1288 => x"ff",
          1289 => x"f1",
          1290 => x"a2",
          1291 => x"81",
          1292 => x"70",
          1293 => x"a0",
          1294 => x"2e",
          1295 => x"81",
          1296 => x"ff",
          1297 => x"81",
          1298 => x"32",
          1299 => x"52",
          1300 => x"80",
          1301 => x"76",
          1302 => x"0c",
          1303 => x"c4",
          1304 => x"81",
          1305 => x"ff",
          1306 => x"e4",
          1307 => x"55",
          1308 => x"09",
          1309 => x"fc",
          1310 => x"38",
          1311 => x"3d",
          1312 => x"72",
          1313 => x"08",
          1314 => x"8c",
          1315 => x"0d",
          1316 => x"53",
          1317 => x"38",
          1318 => x"52",
          1319 => x"13",
          1320 => x"80",
          1321 => x"52",
          1322 => x"13",
          1323 => x"80",
          1324 => x"52",
          1325 => x"8a",
          1326 => x"e7",
          1327 => x"c0",
          1328 => x"98",
          1329 => x"98",
          1330 => x"98",
          1331 => x"98",
          1332 => x"98",
          1333 => x"98",
          1334 => x"0c",
          1335 => x"0b",
          1336 => x"71",
          1337 => x"04",
          1338 => x"98",
          1339 => x"98",
          1340 => x"c0",
          1341 => x"34",
          1342 => x"83",
          1343 => x"5c",
          1344 => x"ac",
          1345 => x"c0",
          1346 => x"34",
          1347 => x"88",
          1348 => x"5a",
          1349 => x"79",
          1350 => x"ff",
          1351 => x"85",
          1352 => x"83",
          1353 => x"7d",
          1354 => x"f4",
          1355 => x"0d",
          1356 => x"33",
          1357 => x"51",
          1358 => x"08",
          1359 => x"71",
          1360 => x"72",
          1361 => x"8c",
          1362 => x"80",
          1363 => x"98",
          1364 => x"ff",
          1365 => x"51",
          1366 => x"08",
          1367 => x"71",
          1368 => x"3d",
          1369 => x"2b",
          1370 => x"84",
          1371 => x"2c",
          1372 => x"73",
          1373 => x"73",
          1374 => x"0c",
          1375 => x"02",
          1376 => x"70",
          1377 => x"80",
          1378 => x"94",
          1379 => x"53",
          1380 => x"71",
          1381 => x"70",
          1382 => x"53",
          1383 => x"2a",
          1384 => x"81",
          1385 => x"52",
          1386 => x"94",
          1387 => x"ba",
          1388 => x"91",
          1389 => x"97",
          1390 => x"72",
          1391 => x"81",
          1392 => x"87",
          1393 => x"70",
          1394 => x"38",
          1395 => x"05",
          1396 => x"52",
          1397 => x"3d",
          1398 => x"80",
          1399 => x"77",
          1400 => x"f2",
          1401 => x"57",
          1402 => x"87",
          1403 => x"70",
          1404 => x"2e",
          1405 => x"06",
          1406 => x"32",
          1407 => x"38",
          1408 => x"cf",
          1409 => x"c0",
          1410 => x"38",
          1411 => x"0c",
          1412 => x"ff",
          1413 => x"88",
          1414 => x"81",
          1415 => x"81",
          1416 => x"c1",
          1417 => x"71",
          1418 => x"94",
          1419 => x"06",
          1420 => x"39",
          1421 => x"08",
          1422 => x"70",
          1423 => x"9e",
          1424 => x"c0",
          1425 => x"87",
          1426 => x"0c",
          1427 => x"d4",
          1428 => x"f2",
          1429 => x"83",
          1430 => x"08",
          1431 => x"b0",
          1432 => x"9e",
          1433 => x"c0",
          1434 => x"87",
          1435 => x"0c",
          1436 => x"f4",
          1437 => x"f2",
          1438 => x"52",
          1439 => x"9e",
          1440 => x"c0",
          1441 => x"87",
          1442 => x"0c",
          1443 => x"0b",
          1444 => x"80",
          1445 => x"fb",
          1446 => x"0b",
          1447 => x"80",
          1448 => x"2e",
          1449 => x"8e",
          1450 => x"08",
          1451 => x"52",
          1452 => x"71",
          1453 => x"c0",
          1454 => x"06",
          1455 => x"38",
          1456 => x"80",
          1457 => x"a0",
          1458 => x"80",
          1459 => x"f3",
          1460 => x"90",
          1461 => x"52",
          1462 => x"52",
          1463 => x"87",
          1464 => x"80",
          1465 => x"83",
          1466 => x"34",
          1467 => x"70",
          1468 => x"70",
          1469 => x"83",
          1470 => x"9e",
          1471 => x"51",
          1472 => x"81",
          1473 => x"0b",
          1474 => x"c0",
          1475 => x"2e",
          1476 => x"96",
          1477 => x"08",
          1478 => x"70",
          1479 => x"83",
          1480 => x"08",
          1481 => x"51",
          1482 => x"87",
          1483 => x"06",
          1484 => x"38",
          1485 => x"87",
          1486 => x"70",
          1487 => x"9a",
          1488 => x"08",
          1489 => x"80",
          1490 => x"f3",
          1491 => x"87",
          1492 => x"83",
          1493 => x"39",
          1494 => x"ff",
          1495 => x"54",
          1496 => x"51",
          1497 => x"55",
          1498 => x"33",
          1499 => x"90",
          1500 => x"f3",
          1501 => x"83",
          1502 => x"38",
          1503 => x"b3",
          1504 => x"84",
          1505 => x"74",
          1506 => x"56",
          1507 => x"33",
          1508 => x"94",
          1509 => x"f3",
          1510 => x"83",
          1511 => x"38",
          1512 => x"83",
          1513 => x"51",
          1514 => x"08",
          1515 => x"ae",
          1516 => x"da",
          1517 => x"da",
          1518 => x"fc",
          1519 => x"b5",
          1520 => x"bd",
          1521 => x"3f",
          1522 => x"29",
          1523 => x"8c",
          1524 => x"b4",
          1525 => x"74",
          1526 => x"55",
          1527 => x"3f",
          1528 => x"08",
          1529 => x"c9",
          1530 => x"84",
          1531 => x"84",
          1532 => x"51",
          1533 => x"f4",
          1534 => x"84",
          1535 => x"51",
          1536 => x"bd",
          1537 => x"54",
          1538 => x"c4",
          1539 => x"8e",
          1540 => x"38",
          1541 => x"c0",
          1542 => x"c1",
          1543 => x"d9",
          1544 => x"f2",
          1545 => x"ff",
          1546 => x"52",
          1547 => x"3f",
          1548 => x"83",
          1549 => x"51",
          1550 => x"08",
          1551 => x"c8",
          1552 => x"84",
          1553 => x"84",
          1554 => x"51",
          1555 => x"33",
          1556 => x"fe",
          1557 => x"bf",
          1558 => x"73",
          1559 => x"39",
          1560 => x"3f",
          1561 => x"2e",
          1562 => x"8c",
          1563 => x"94",
          1564 => x"38",
          1565 => x"bf",
          1566 => x"73",
          1567 => x"83",
          1568 => x"51",
          1569 => x"33",
          1570 => x"d2",
          1571 => x"dc",
          1572 => x"f3",
          1573 => x"e3",
          1574 => x"52",
          1575 => x"3f",
          1576 => x"2e",
          1577 => x"d8",
          1578 => x"52",
          1579 => x"3f",
          1580 => x"2e",
          1581 => x"d0",
          1582 => x"52",
          1583 => x"3f",
          1584 => x"2e",
          1585 => x"c8",
          1586 => x"52",
          1587 => x"3f",
          1588 => x"2e",
          1589 => x"e0",
          1590 => x"52",
          1591 => x"3f",
          1592 => x"2e",
          1593 => x"e8",
          1594 => x"52",
          1595 => x"3f",
          1596 => x"2e",
          1597 => x"98",
          1598 => x"a0",
          1599 => x"8e",
          1600 => x"38",
          1601 => x"05",
          1602 => x"71",
          1603 => x"71",
          1604 => x"af",
          1605 => x"de",
          1606 => x"3d",
          1607 => x"af",
          1608 => x"de",
          1609 => x"3d",
          1610 => x"af",
          1611 => x"de",
          1612 => x"3d",
          1613 => x"80",
          1614 => x"83",
          1615 => x"0c",
          1616 => x"ad",
          1617 => x"58",
          1618 => x"82",
          1619 => x"80",
          1620 => x"83",
          1621 => x"52",
          1622 => x"ba",
          1623 => x"51",
          1624 => x"81",
          1625 => x"8c",
          1626 => x"08",
          1627 => x"74",
          1628 => x"07",
          1629 => x"2e",
          1630 => x"f3",
          1631 => x"82",
          1632 => x"8f",
          1633 => x"84",
          1634 => x"83",
          1635 => x"78",
          1636 => x"76",
          1637 => x"51",
          1638 => x"56",
          1639 => x"52",
          1640 => x"3f",
          1641 => x"3d",
          1642 => x"08",
          1643 => x"33",
          1644 => x"81",
          1645 => x"56",
          1646 => x"05",
          1647 => x"3f",
          1648 => x"73",
          1649 => x"8c",
          1650 => x"73",
          1651 => x"2e",
          1652 => x"06",
          1653 => x"80",
          1654 => x"3d",
          1655 => x"ff",
          1656 => x"c7",
          1657 => x"2e",
          1658 => x"76",
          1659 => x"08",
          1660 => x"c9",
          1661 => x"57",
          1662 => x"ff",
          1663 => x"76",
          1664 => x"70",
          1665 => x"2e",
          1666 => x"75",
          1667 => x"59",
          1668 => x"8c",
          1669 => x"56",
          1670 => x"08",
          1671 => x"53",
          1672 => x"cc",
          1673 => x"ba",
          1674 => x"84",
          1675 => x"ba",
          1676 => x"8c",
          1677 => x"80",
          1678 => x"16",
          1679 => x"8e",
          1680 => x"ff",
          1681 => x"0c",
          1682 => x"b5",
          1683 => x"08",
          1684 => x"34",
          1685 => x"08",
          1686 => x"f3",
          1687 => x"82",
          1688 => x"38",
          1689 => x"90",
          1690 => x"38",
          1691 => x"51",
          1692 => x"98",
          1693 => x"ff",
          1694 => x"84",
          1695 => x"98",
          1696 => x"2b",
          1697 => x"70",
          1698 => x"08",
          1699 => x"46",
          1700 => x"74",
          1701 => x"27",
          1702 => x"29",
          1703 => x"57",
          1704 => x"75",
          1705 => x"80",
          1706 => x"57",
          1707 => x"d8",
          1708 => x"78",
          1709 => x"2e",
          1710 => x"81",
          1711 => x"81",
          1712 => x"84",
          1713 => x"97",
          1714 => x"2b",
          1715 => x"5f",
          1716 => x"2e",
          1717 => x"34",
          1718 => x"ba",
          1719 => x"80",
          1720 => x"ff",
          1721 => x"80",
          1722 => x"2b",
          1723 => x"16",
          1724 => x"38",
          1725 => x"33",
          1726 => x"38",
          1727 => x"f2",
          1728 => x"ab",
          1729 => x"b2",
          1730 => x"76",
          1731 => x"c4",
          1732 => x"62",
          1733 => x"74",
          1734 => x"76",
          1735 => x"7f",
          1736 => x"80",
          1737 => x"84",
          1738 => x"fd",
          1739 => x"88",
          1740 => x"d0",
          1741 => x"d0",
          1742 => x"33",
          1743 => x"33",
          1744 => x"d6",
          1745 => x"15",
          1746 => x"16",
          1747 => x"3f",
          1748 => x"da",
          1749 => x"05",
          1750 => x"38",
          1751 => x"34",
          1752 => x"33",
          1753 => x"84",
          1754 => x"b5",
          1755 => x"a0",
          1756 => x"f0",
          1757 => x"3f",
          1758 => x"7a",
          1759 => x"06",
          1760 => x"a6",
          1761 => x"fb",
          1762 => x"f0",
          1763 => x"10",
          1764 => x"08",
          1765 => x"08",
          1766 => x"75",
          1767 => x"8c",
          1768 => x"8c",
          1769 => x"75",
          1770 => x"84",
          1771 => x"56",
          1772 => x"84",
          1773 => x"b4",
          1774 => x"a0",
          1775 => x"f0",
          1776 => x"3f",
          1777 => x"74",
          1778 => x"06",
          1779 => x"70",
          1780 => x"5b",
          1781 => x"38",
          1782 => x"57",
          1783 => x"70",
          1784 => x"84",
          1785 => x"84",
          1786 => x"78",
          1787 => x"08",
          1788 => x"d0",
          1789 => x"ff",
          1790 => x"70",
          1791 => x"5a",
          1792 => x"38",
          1793 => x"84",
          1794 => x"2e",
          1795 => x"84",
          1796 => x"98",
          1797 => x"5a",
          1798 => x"d5",
          1799 => x"b4",
          1800 => x"2b",
          1801 => x"5a",
          1802 => x"86",
          1803 => x"51",
          1804 => x"0a",
          1805 => x"2c",
          1806 => x"74",
          1807 => x"f0",
          1808 => x"3f",
          1809 => x"0a",
          1810 => x"33",
          1811 => x"b9",
          1812 => x"81",
          1813 => x"08",
          1814 => x"3f",
          1815 => x"0a",
          1816 => x"33",
          1817 => x"e6",
          1818 => x"78",
          1819 => x"33",
          1820 => x"80",
          1821 => x"98",
          1822 => x"55",
          1823 => x"b6",
          1824 => x"80",
          1825 => x"08",
          1826 => x"84",
          1827 => x"84",
          1828 => x"55",
          1829 => x"05",
          1830 => x"08",
          1831 => x"84",
          1832 => x"3f",
          1833 => x"58",
          1834 => x"33",
          1835 => x"83",
          1836 => x"f3",
          1837 => x"74",
          1838 => x"fc",
          1839 => x"70",
          1840 => x"84",
          1841 => x"fc",
          1842 => x"05",
          1843 => x"ad",
          1844 => x"80",
          1845 => x"58",
          1846 => x"0b",
          1847 => x"d1",
          1848 => x"b4",
          1849 => x"55",
          1850 => x"f0",
          1851 => x"3f",
          1852 => x"ff",
          1853 => x"52",
          1854 => x"d1",
          1855 => x"d1",
          1856 => x"74",
          1857 => x"9f",
          1858 => x"34",
          1859 => x"be",
          1860 => x"1d",
          1861 => x"80",
          1862 => x"52",
          1863 => x"d5",
          1864 => x"ac",
          1865 => x"51",
          1866 => x"33",
          1867 => x"34",
          1868 => x"38",
          1869 => x"3f",
          1870 => x"0b",
          1871 => x"8c",
          1872 => x"d0",
          1873 => x"7a",
          1874 => x"cc",
          1875 => x"cc",
          1876 => x"d0",
          1877 => x"51",
          1878 => x"33",
          1879 => x"d1",
          1880 => x"76",
          1881 => x"08",
          1882 => x"84",
          1883 => x"98",
          1884 => x"59",
          1885 => x"84",
          1886 => x"ac",
          1887 => x"81",
          1888 => x"d1",
          1889 => x"24",
          1890 => x"52",
          1891 => x"81",
          1892 => x"70",
          1893 => x"51",
          1894 => x"f3",
          1895 => x"33",
          1896 => x"76",
          1897 => x"81",
          1898 => x"70",
          1899 => x"57",
          1900 => x"7b",
          1901 => x"84",
          1902 => x"ff",
          1903 => x"29",
          1904 => x"84",
          1905 => x"76",
          1906 => x"84",
          1907 => x"58",
          1908 => x"84",
          1909 => x"ae",
          1910 => x"57",
          1911 => x"16",
          1912 => x"81",
          1913 => x"70",
          1914 => x"57",
          1915 => x"18",
          1916 => x"81",
          1917 => x"33",
          1918 => x"76",
          1919 => x"75",
          1920 => x"d1",
          1921 => x"81",
          1922 => x"81",
          1923 => x"76",
          1924 => x"70",
          1925 => x"57",
          1926 => x"84",
          1927 => x"aa",
          1928 => x"81",
          1929 => x"d1",
          1930 => x"25",
          1931 => x"52",
          1932 => x"81",
          1933 => x"70",
          1934 => x"57",
          1935 => x"f0",
          1936 => x"75",
          1937 => x"ff",
          1938 => x"84",
          1939 => x"81",
          1940 => x"7b",
          1941 => x"cc",
          1942 => x"74",
          1943 => x"f0",
          1944 => x"3f",
          1945 => x"ff",
          1946 => x"52",
          1947 => x"d1",
          1948 => x"d1",
          1949 => x"c7",
          1950 => x"84",
          1951 => x"84",
          1952 => x"83",
          1953 => x"80",
          1954 => x"7b",
          1955 => x"d4",
          1956 => x"80",
          1957 => x"cc",
          1958 => x"da",
          1959 => x"2b",
          1960 => x"5d",
          1961 => x"8e",
          1962 => x"08",
          1963 => x"a4",
          1964 => x"bb",
          1965 => x"75",
          1966 => x"f3",
          1967 => x"74",
          1968 => x"81",
          1969 => x"51",
          1970 => x"f3",
          1971 => x"5f",
          1972 => x"b8",
          1973 => x"18",
          1974 => x"38",
          1975 => x"ee",
          1976 => x"cc",
          1977 => x"06",
          1978 => x"ff",
          1979 => x"cc",
          1980 => x"5d",
          1981 => x"d5",
          1982 => x"fc",
          1983 => x"51",
          1984 => x"08",
          1985 => x"84",
          1986 => x"84",
          1987 => x"55",
          1988 => x"84",
          1989 => x"cc",
          1990 => x"3d",
          1991 => x"3f",
          1992 => x"34",
          1993 => x"81",
          1994 => x"aa",
          1995 => x"06",
          1996 => x"33",
          1997 => x"f1",
          1998 => x"88",
          1999 => x"f0",
          2000 => x"3f",
          2001 => x"ff",
          2002 => x"ff",
          2003 => x"76",
          2004 => x"51",
          2005 => x"08",
          2006 => x"08",
          2007 => x"52",
          2008 => x"1d",
          2009 => x"33",
          2010 => x"58",
          2011 => x"d5",
          2012 => x"8c",
          2013 => x"51",
          2014 => x"08",
          2015 => x"84",
          2016 => x"84",
          2017 => x"55",
          2018 => x"3f",
          2019 => x"87",
          2020 => x"19",
          2021 => x"a0",
          2022 => x"83",
          2023 => x"f3",
          2024 => x"74",
          2025 => x"7b",
          2026 => x"83",
          2027 => x"ff",
          2028 => x"f2",
          2029 => x"b1",
          2030 => x"76",
          2031 => x"8f",
          2032 => x"51",
          2033 => x"08",
          2034 => x"84",
          2035 => x"cc",
          2036 => x"3d",
          2037 => x"ba",
          2038 => x"84",
          2039 => x"ba",
          2040 => x"f3",
          2041 => x"51",
          2042 => x"08",
          2043 => x"09",
          2044 => x"8c",
          2045 => x"ba",
          2046 => x"8c",
          2047 => x"8c",
          2048 => x"80",
          2049 => x"f3",
          2050 => x"a4",
          2051 => x"74",
          2052 => x"fc",
          2053 => x"70",
          2054 => x"84",
          2055 => x"fc",
          2056 => x"05",
          2057 => x"38",
          2058 => x"57",
          2059 => x"75",
          2060 => x"38",
          2061 => x"76",
          2062 => x"f8",
          2063 => x"70",
          2064 => x"27",
          2065 => x"fc",
          2066 => x"d4",
          2067 => x"82",
          2068 => x"05",
          2069 => x"80",
          2070 => x"75",
          2071 => x"10",
          2072 => x"40",
          2073 => x"ff",
          2074 => x"fe",
          2075 => x"f1",
          2076 => x"9f",
          2077 => x"e4",
          2078 => x"05",
          2079 => x"33",
          2080 => x"38",
          2081 => x"73",
          2082 => x"82",
          2083 => x"87",
          2084 => x"56",
          2085 => x"38",
          2086 => x"f9",
          2087 => x"83",
          2088 => x"90",
          2089 => x"07",
          2090 => x"77",
          2091 => x"05",
          2092 => x"55",
          2093 => x"78",
          2094 => x"84",
          2095 => x"55",
          2096 => x"74",
          2097 => x"13",
          2098 => x"04",
          2099 => x"bc",
          2100 => x"bd",
          2101 => x"5b",
          2102 => x"80",
          2103 => x"ff",
          2104 => x"ff",
          2105 => x"ff",
          2106 => x"5d",
          2107 => x"26",
          2108 => x"56",
          2109 => x"06",
          2110 => x"ff",
          2111 => x"29",
          2112 => x"74",
          2113 => x"33",
          2114 => x"1b",
          2115 => x"80",
          2116 => x"53",
          2117 => x"73",
          2118 => x"b8",
          2119 => x"e8",
          2120 => x"a3",
          2121 => x"70",
          2122 => x"70",
          2123 => x"70",
          2124 => x"56",
          2125 => x"38",
          2126 => x"06",
          2127 => x"79",
          2128 => x"83",
          2129 => x"bd",
          2130 => x"2b",
          2131 => x"07",
          2132 => x"5b",
          2133 => x"be",
          2134 => x"bc",
          2135 => x"10",
          2136 => x"29",
          2137 => x"57",
          2138 => x"80",
          2139 => x"81",
          2140 => x"81",
          2141 => x"83",
          2142 => x"05",
          2143 => x"5e",
          2144 => x"7a",
          2145 => x"53",
          2146 => x"06",
          2147 => x"06",
          2148 => x"58",
          2149 => x"26",
          2150 => x"73",
          2151 => x"79",
          2152 => x"7b",
          2153 => x"78",
          2154 => x"fb",
          2155 => x"80",
          2156 => x"86",
          2157 => x"80",
          2158 => x"8a",
          2159 => x"74",
          2160 => x"8a",
          2161 => x"34",
          2162 => x"fa",
          2163 => x"08",
          2164 => x"81",
          2165 => x"55",
          2166 => x"ff",
          2167 => x"75",
          2168 => x"77",
          2169 => x"8c",
          2170 => x"06",
          2171 => x"d0",
          2172 => x"84",
          2173 => x"84",
          2174 => x"04",
          2175 => x"02",
          2176 => x"ff",
          2177 => x"79",
          2178 => x"33",
          2179 => x"33",
          2180 => x"80",
          2181 => x"57",
          2182 => x"ff",
          2183 => x"57",
          2184 => x"38",
          2185 => x"74",
          2186 => x"33",
          2187 => x"81",
          2188 => x"26",
          2189 => x"83",
          2190 => x"70",
          2191 => x"33",
          2192 => x"89",
          2193 => x"29",
          2194 => x"26",
          2195 => x"54",
          2196 => x"16",
          2197 => x"75",
          2198 => x"54",
          2199 => x"73",
          2200 => x"b8",
          2201 => x"a0",
          2202 => x"70",
          2203 => x"9f",
          2204 => x"fe",
          2205 => x"ba",
          2206 => x"77",
          2207 => x"73",
          2208 => x"81",
          2209 => x"29",
          2210 => x"a0",
          2211 => x"81",
          2212 => x"71",
          2213 => x"79",
          2214 => x"54",
          2215 => x"88",
          2216 => x"34",
          2217 => x"70",
          2218 => x"b8",
          2219 => x"71",
          2220 => x"75",
          2221 => x"ba",
          2222 => x"83",
          2223 => x"70",
          2224 => x"33",
          2225 => x"f9",
          2226 => x"78",
          2227 => x"bc",
          2228 => x"81",
          2229 => x"81",
          2230 => x"29",
          2231 => x"54",
          2232 => x"f9",
          2233 => x"76",
          2234 => x"e0",
          2235 => x"57",
          2236 => x"fe",
          2237 => x"34",
          2238 => x"ff",
          2239 => x"39",
          2240 => x"56",
          2241 => x"33",
          2242 => x"34",
          2243 => x"39",
          2244 => x"9f",
          2245 => x"9b",
          2246 => x"05",
          2247 => x"33",
          2248 => x"83",
          2249 => x"8c",
          2250 => x"83",
          2251 => x"70",
          2252 => x"2e",
          2253 => x"f9",
          2254 => x"0c",
          2255 => x"33",
          2256 => x"2c",
          2257 => x"83",
          2258 => x"bc",
          2259 => x"ff",
          2260 => x"83",
          2261 => x"34",
          2262 => x"3d",
          2263 => x"73",
          2264 => x"06",
          2265 => x"bd",
          2266 => x"86",
          2267 => x"72",
          2268 => x"55",
          2269 => x"70",
          2270 => x"0b",
          2271 => x"04",
          2272 => x"f9",
          2273 => x"05",
          2274 => x"38",
          2275 => x"34",
          2276 => x"8f",
          2277 => x"38",
          2278 => x"51",
          2279 => x"70",
          2280 => x"f0",
          2281 => x"52",
          2282 => x"81",
          2283 => x"f9",
          2284 => x"0c",
          2285 => x"33",
          2286 => x"83",
          2287 => x"8c",
          2288 => x"b8",
          2289 => x"f9",
          2290 => x"33",
          2291 => x"83",
          2292 => x"0b",
          2293 => x"ba",
          2294 => x"f9",
          2295 => x"51",
          2296 => x"39",
          2297 => x"70",
          2298 => x"83",
          2299 => x"07",
          2300 => x"93",
          2301 => x"06",
          2302 => x"34",
          2303 => x"81",
          2304 => x"f9",
          2305 => x"b8",
          2306 => x"f9",
          2307 => x"b8",
          2308 => x"51",
          2309 => x"39",
          2310 => x"b0",
          2311 => x"fe",
          2312 => x"ef",
          2313 => x"f9",
          2314 => x"b8",
          2315 => x"51",
          2316 => x"39",
          2317 => x"a0",
          2318 => x"fe",
          2319 => x"8f",
          2320 => x"fd",
          2321 => x"fa",
          2322 => x"b8",
          2323 => x"02",
          2324 => x"c3",
          2325 => x"f9",
          2326 => x"b8",
          2327 => x"59",
          2328 => x"82",
          2329 => x"82",
          2330 => x"0b",
          2331 => x"bc",
          2332 => x"83",
          2333 => x"78",
          2334 => x"80",
          2335 => x"84",
          2336 => x"bc",
          2337 => x"82",
          2338 => x"84",
          2339 => x"33",
          2340 => x"54",
          2341 => x"51",
          2342 => x"82",
          2343 => x"7a",
          2344 => x"ba",
          2345 => x"3d",
          2346 => x"34",
          2347 => x"0b",
          2348 => x"f9",
          2349 => x"23",
          2350 => x"8e",
          2351 => x"79",
          2352 => x"83",
          2353 => x"80",
          2354 => x"79",
          2355 => x"b9",
          2356 => x"e3",
          2357 => x"1a",
          2358 => x"33",
          2359 => x"38",
          2360 => x"3f",
          2361 => x"84",
          2362 => x"34",
          2363 => x"f9",
          2364 => x"0b",
          2365 => x"b8",
          2366 => x"34",
          2367 => x"0b",
          2368 => x"51",
          2369 => x"08",
          2370 => x"f6",
          2371 => x"ff",
          2372 => x"08",
          2373 => x"19",
          2374 => x"ff",
          2375 => x"06",
          2376 => x"7a",
          2377 => x"b8",
          2378 => x"f9",
          2379 => x"a3",
          2380 => x"53",
          2381 => x"70",
          2382 => x"33",
          2383 => x"81",
          2384 => x"81",
          2385 => x"38",
          2386 => x"88",
          2387 => x"33",
          2388 => x"33",
          2389 => x"84",
          2390 => x"80",
          2391 => x"f9",
          2392 => x"71",
          2393 => x"83",
          2394 => x"33",
          2395 => x"f9",
          2396 => x"34",
          2397 => x"06",
          2398 => x"33",
          2399 => x"55",
          2400 => x"de",
          2401 => x"06",
          2402 => x"38",
          2403 => x"ea",
          2404 => x"bd",
          2405 => x"80",
          2406 => x"57",
          2407 => x"0b",
          2408 => x"04",
          2409 => x"24",
          2410 => x"81",
          2411 => x"51",
          2412 => x"bd",
          2413 => x"15",
          2414 => x"74",
          2415 => x"fe",
          2416 => x"51",
          2417 => x"ff",
          2418 => x"91",
          2419 => x"3f",
          2420 => x"54",
          2421 => x"39",
          2422 => x"39",
          2423 => x"80",
          2424 => x"0d",
          2425 => x"06",
          2426 => x"70",
          2427 => x"73",
          2428 => x"bd",
          2429 => x"3f",
          2430 => x"06",
          2431 => x"38",
          2432 => x"fe",
          2433 => x"34",
          2434 => x"fe",
          2435 => x"d8",
          2436 => x"02",
          2437 => x"08",
          2438 => x"38",
          2439 => x"8a",
          2440 => x"82",
          2441 => x"38",
          2442 => x"b8",
          2443 => x"f9",
          2444 => x"5e",
          2445 => x"a3",
          2446 => x"33",
          2447 => x"22",
          2448 => x"40",
          2449 => x"f9",
          2450 => x"40",
          2451 => x"a3",
          2452 => x"33",
          2453 => x"22",
          2454 => x"11",
          2455 => x"b8",
          2456 => x"1d",
          2457 => x"61",
          2458 => x"33",
          2459 => x"56",
          2460 => x"84",
          2461 => x"78",
          2462 => x"25",
          2463 => x"b3",
          2464 => x"38",
          2465 => x"b8",
          2466 => x"f9",
          2467 => x"40",
          2468 => x"a3",
          2469 => x"33",
          2470 => x"22",
          2471 => x"56",
          2472 => x"f9",
          2473 => x"57",
          2474 => x"80",
          2475 => x"81",
          2476 => x"f9",
          2477 => x"42",
          2478 => x"60",
          2479 => x"58",
          2480 => x"27",
          2481 => x"34",
          2482 => x"3d",
          2483 => x"38",
          2484 => x"8d",
          2485 => x"80",
          2486 => x"84",
          2487 => x"78",
          2488 => x"56",
          2489 => x"b9",
          2490 => x"84",
          2491 => x"18",
          2492 => x"0b",
          2493 => x"84",
          2494 => x"78",
          2495 => x"84",
          2496 => x"83",
          2497 => x"72",
          2498 => x"b8",
          2499 => x"1d",
          2500 => x"bd",
          2501 => x"29",
          2502 => x"f9",
          2503 => x"76",
          2504 => x"b8",
          2505 => x"84",
          2506 => x"83",
          2507 => x"72",
          2508 => x"59",
          2509 => x"de",
          2510 => x"39",
          2511 => x"80",
          2512 => x"39",
          2513 => x"33",
          2514 => x"33",
          2515 => x"80",
          2516 => x"5d",
          2517 => x"ff",
          2518 => x"59",
          2519 => x"38",
          2520 => x"57",
          2521 => x"83",
          2522 => x"0b",
          2523 => x"b9",
          2524 => x"34",
          2525 => x"0b",
          2526 => x"ba",
          2527 => x"f9",
          2528 => x"f9",
          2529 => x"f9",
          2530 => x"0b",
          2531 => x"ba",
          2532 => x"80",
          2533 => x"38",
          2534 => x"33",
          2535 => x"33",
          2536 => x"11",
          2537 => x"ba",
          2538 => x"70",
          2539 => x"33",
          2540 => x"7d",
          2541 => x"ff",
          2542 => x"38",
          2543 => x"7b",
          2544 => x"78",
          2545 => x"5f",
          2546 => x"a3",
          2547 => x"33",
          2548 => x"22",
          2549 => x"40",
          2550 => x"83",
          2551 => x"05",
          2552 => x"a3",
          2553 => x"33",
          2554 => x"22",
          2555 => x"11",
          2556 => x"b8",
          2557 => x"81",
          2558 => x"7c",
          2559 => x"81",
          2560 => x"19",
          2561 => x"f9",
          2562 => x"ff",
          2563 => x"2e",
          2564 => x"d7",
          2565 => x"84",
          2566 => x"38",
          2567 => x"84",
          2568 => x"98",
          2569 => x"83",
          2570 => x"e7",
          2571 => x"0c",
          2572 => x"33",
          2573 => x"06",
          2574 => x"06",
          2575 => x"80",
          2576 => x"72",
          2577 => x"06",
          2578 => x"5c",
          2579 => x"ef",
          2580 => x"7a",
          2581 => x"72",
          2582 => x"b8",
          2583 => x"34",
          2584 => x"33",
          2585 => x"12",
          2586 => x"f9",
          2587 => x"76",
          2588 => x"b8",
          2589 => x"84",
          2590 => x"83",
          2591 => x"72",
          2592 => x"59",
          2593 => x"18",
          2594 => x"06",
          2595 => x"38",
          2596 => x"fb",
          2597 => x"bd",
          2598 => x"5d",
          2599 => x"83",
          2600 => x"83",
          2601 => x"72",
          2602 => x"72",
          2603 => x"5b",
          2604 => x"a0",
          2605 => x"83",
          2606 => x"72",
          2607 => x"a0",
          2608 => x"f9",
          2609 => x"5e",
          2610 => x"80",
          2611 => x"81",
          2612 => x"f9",
          2613 => x"44",
          2614 => x"84",
          2615 => x"70",
          2616 => x"27",
          2617 => x"34",
          2618 => x"88",
          2619 => x"9c",
          2620 => x"33",
          2621 => x"34",
          2622 => x"06",
          2623 => x"81",
          2624 => x"84",
          2625 => x"83",
          2626 => x"88",
          2627 => x"33",
          2628 => x"33",
          2629 => x"39",
          2630 => x"11",
          2631 => x"3f",
          2632 => x"f0",
          2633 => x"57",
          2634 => x"10",
          2635 => x"05",
          2636 => x"fb",
          2637 => x"5c",
          2638 => x"83",
          2639 => x"83",
          2640 => x"e5",
          2641 => x"bc",
          2642 => x"29",
          2643 => x"19",
          2644 => x"34",
          2645 => x"33",
          2646 => x"12",
          2647 => x"be",
          2648 => x"71",
          2649 => x"33",
          2650 => x"84",
          2651 => x"83",
          2652 => x"72",
          2653 => x"5a",
          2654 => x"1e",
          2655 => x"5c",
          2656 => x"84",
          2657 => x"38",
          2658 => x"34",
          2659 => x"b8",
          2660 => x"bd",
          2661 => x"f3",
          2662 => x"e4",
          2663 => x"9c",
          2664 => x"83",
          2665 => x"83",
          2666 => x"57",
          2667 => x"39",
          2668 => x"34",
          2669 => x"34",
          2670 => x"34",
          2671 => x"5b",
          2672 => x"b9",
          2673 => x"81",
          2674 => x"33",
          2675 => x"81",
          2676 => x"52",
          2677 => x"fe",
          2678 => x"84",
          2679 => x"f8",
          2680 => x"a0",
          2681 => x"f7",
          2682 => x"c0",
          2683 => x"5b",
          2684 => x"7b",
          2685 => x"b9",
          2686 => x"75",
          2687 => x"10",
          2688 => x"04",
          2689 => x"2e",
          2690 => x"84",
          2691 => x"09",
          2692 => x"59",
          2693 => x"fd",
          2694 => x"75",
          2695 => x"e1",
          2696 => x"84",
          2697 => x"7b",
          2698 => x"bd",
          2699 => x"f9",
          2700 => x"81",
          2701 => x"fd",
          2702 => x"f9",
          2703 => x"83",
          2704 => x"84",
          2705 => x"76",
          2706 => x"56",
          2707 => x"39",
          2708 => x"2e",
          2709 => x"84",
          2710 => x"09",
          2711 => x"59",
          2712 => x"fc",
          2713 => x"7a",
          2714 => x"e0",
          2715 => x"06",
          2716 => x"83",
          2717 => x"72",
          2718 => x"11",
          2719 => x"58",
          2720 => x"ff",
          2721 => x"fe",
          2722 => x"84",
          2723 => x"0b",
          2724 => x"84",
          2725 => x"fb",
          2726 => x"77",
          2727 => x"38",
          2728 => x"d0",
          2729 => x"80",
          2730 => x"33",
          2731 => x"84",
          2732 => x"56",
          2733 => x"76",
          2734 => x"84",
          2735 => x"8c",
          2736 => x"f9",
          2737 => x"ff",
          2738 => x"60",
          2739 => x"f9",
          2740 => x"98",
          2741 => x"84",
          2742 => x"27",
          2743 => x"e0",
          2744 => x"f8",
          2745 => x"70",
          2746 => x"58",
          2747 => x"b9",
          2748 => x"8d",
          2749 => x"83",
          2750 => x"76",
          2751 => x"fa",
          2752 => x"81",
          2753 => x"e3",
          2754 => x"84",
          2755 => x"ff",
          2756 => x"ff",
          2757 => x"59",
          2758 => x"77",
          2759 => x"81",
          2760 => x"7f",
          2761 => x"f9",
          2762 => x"11",
          2763 => x"38",
          2764 => x"f9",
          2765 => x"7e",
          2766 => x"e1",
          2767 => x"7a",
          2768 => x"bc",
          2769 => x"ff",
          2770 => x"29",
          2771 => x"f9",
          2772 => x"05",
          2773 => x"92",
          2774 => x"60",
          2775 => x"ff",
          2776 => x"80",
          2777 => x"ff",
          2778 => x"38",
          2779 => x"23",
          2780 => x"41",
          2781 => x"84",
          2782 => x"8d",
          2783 => x"f9",
          2784 => x"f9",
          2785 => x"76",
          2786 => x"05",
          2787 => x"5c",
          2788 => x"80",
          2789 => x"ff",
          2790 => x"29",
          2791 => x"27",
          2792 => x"57",
          2793 => x"88",
          2794 => x"34",
          2795 => x"70",
          2796 => x"b8",
          2797 => x"71",
          2798 => x"60",
          2799 => x"33",
          2800 => x"70",
          2801 => x"05",
          2802 => x"34",
          2803 => x"b7",
          2804 => x"40",
          2805 => x"38",
          2806 => x"56",
          2807 => x"52",
          2808 => x"3f",
          2809 => x"80",
          2810 => x"5d",
          2811 => x"38",
          2812 => x"2e",
          2813 => x"f9",
          2814 => x"83",
          2815 => x"76",
          2816 => x"ff",
          2817 => x"38",
          2818 => x"26",
          2819 => x"7d",
          2820 => x"7a",
          2821 => x"05",
          2822 => x"5d",
          2823 => x"83",
          2824 => x"38",
          2825 => x"38",
          2826 => x"71",
          2827 => x"71",
          2828 => x"77",
          2829 => x"84",
          2830 => x"05",
          2831 => x"84",
          2832 => x"41",
          2833 => x"ff",
          2834 => x"29",
          2835 => x"77",
          2836 => x"70",
          2837 => x"76",
          2838 => x"e0",
          2839 => x"de",
          2840 => x"19",
          2841 => x"34",
          2842 => x"c0",
          2843 => x"79",
          2844 => x"17",
          2845 => x"a8",
          2846 => x"5d",
          2847 => x"33",
          2848 => x"80",
          2849 => x"5d",
          2850 => x"06",
          2851 => x"b8",
          2852 => x"59",
          2853 => x"17",
          2854 => x"7c",
          2855 => x"80",
          2856 => x"ff",
          2857 => x"39",
          2858 => x"75",
          2859 => x"81",
          2860 => x"83",
          2861 => x"07",
          2862 => x"39",
          2863 => x"83",
          2864 => x"d4",
          2865 => x"06",
          2866 => x"34",
          2867 => x"9f",
          2868 => x"b8",
          2869 => x"83",
          2870 => x"ff",
          2871 => x"f9",
          2872 => x"83",
          2873 => x"f9",
          2874 => x"56",
          2875 => x"39",
          2876 => x"80",
          2877 => x"34",
          2878 => x"81",
          2879 => x"83",
          2880 => x"f9",
          2881 => x"56",
          2882 => x"39",
          2883 => x"86",
          2884 => x"fe",
          2885 => x"fc",
          2886 => x"b8",
          2887 => x"33",
          2888 => x"83",
          2889 => x"f9",
          2890 => x"83",
          2891 => x"f9",
          2892 => x"83",
          2893 => x"f9",
          2894 => x"83",
          2895 => x"f9",
          2896 => x"07",
          2897 => x"cc",
          2898 => x"06",
          2899 => x"34",
          2900 => x"bd",
          2901 => x"3f",
          2902 => x"83",
          2903 => x"83",
          2904 => x"59",
          2905 => x"84",
          2906 => x"0b",
          2907 => x"ba",
          2908 => x"83",
          2909 => x"70",
          2910 => x"e7",
          2911 => x"3d",
          2912 => x"f9",
          2913 => x"38",
          2914 => x"0c",
          2915 => x"0b",
          2916 => x"04",
          2917 => x"39",
          2918 => x"5c",
          2919 => x"83",
          2920 => x"22",
          2921 => x"84",
          2922 => x"83",
          2923 => x"d1",
          2924 => x"81",
          2925 => x"d8",
          2926 => x"80",
          2927 => x"98",
          2928 => x"ef",
          2929 => x"05",
          2930 => x"58",
          2931 => x"81",
          2932 => x"40",
          2933 => x"83",
          2934 => x"f9",
          2935 => x"9f",
          2936 => x"e2",
          2937 => x"84",
          2938 => x"56",
          2939 => x"57",
          2940 => x"70",
          2941 => x"26",
          2942 => x"84",
          2943 => x"83",
          2944 => x"87",
          2945 => x"22",
          2946 => x"83",
          2947 => x"5d",
          2948 => x"2e",
          2949 => x"06",
          2950 => x"84",
          2951 => x"76",
          2952 => x"56",
          2953 => x"ff",
          2954 => x"24",
          2955 => x"56",
          2956 => x"16",
          2957 => x"81",
          2958 => x"57",
          2959 => x"75",
          2960 => x"06",
          2961 => x"58",
          2962 => x"b0",
          2963 => x"ff",
          2964 => x"42",
          2965 => x"84",
          2966 => x"33",
          2967 => x"70",
          2968 => x"05",
          2969 => x"34",
          2970 => x"b7",
          2971 => x"41",
          2972 => x"38",
          2973 => x"88",
          2974 => x"34",
          2975 => x"70",
          2976 => x"b8",
          2977 => x"71",
          2978 => x"78",
          2979 => x"83",
          2980 => x"88",
          2981 => x"33",
          2982 => x"22",
          2983 => x"5d",
          2984 => x"84",
          2985 => x"ff",
          2986 => x"83",
          2987 => x"23",
          2988 => x"5a",
          2989 => x"76",
          2990 => x"33",
          2991 => x"59",
          2992 => x"80",
          2993 => x"88",
          2994 => x"84",
          2995 => x"56",
          2996 => x"57",
          2997 => x"81",
          2998 => x"33",
          2999 => x"33",
          3000 => x"2e",
          3001 => x"a1",
          3002 => x"bc",
          3003 => x"75",
          3004 => x"7c",
          3005 => x"34",
          3006 => x"77",
          3007 => x"70",
          3008 => x"33",
          3009 => x"7a",
          3010 => x"81",
          3011 => x"77",
          3012 => x"27",
          3013 => x"31",
          3014 => x"a8",
          3015 => x"fc",
          3016 => x"fc",
          3017 => x"23",
          3018 => x"bc",
          3019 => x"18",
          3020 => x"77",
          3021 => x"e9",
          3022 => x"05",
          3023 => x"72",
          3024 => x"9c",
          3025 => x"85",
          3026 => x"d7",
          3027 => x"0c",
          3028 => x"02",
          3029 => x"f8",
          3030 => x"f7",
          3031 => x"74",
          3032 => x"56",
          3033 => x"78",
          3034 => x"04",
          3035 => x"73",
          3036 => x"70",
          3037 => x"2a",
          3038 => x"ec",
          3039 => x"2e",
          3040 => x"7b",
          3041 => x"76",
          3042 => x"85",
          3043 => x"f9",
          3044 => x"71",
          3045 => x"83",
          3046 => x"79",
          3047 => x"83",
          3048 => x"74",
          3049 => x"54",
          3050 => x"0b",
          3051 => x"98",
          3052 => x"38",
          3053 => x"83",
          3054 => x"81",
          3055 => x"27",
          3056 => x"14",
          3057 => x"b6",
          3058 => x"2e",
          3059 => x"86",
          3060 => x"34",
          3061 => x"ff",
          3062 => x"ca",
          3063 => x"83",
          3064 => x"81",
          3065 => x"ff",
          3066 => x"98",
          3067 => x"75",
          3068 => x"06",
          3069 => x"06",
          3070 => x"e7",
          3071 => x"73",
          3072 => x"85",
          3073 => x"34",
          3074 => x"f7",
          3075 => x"83",
          3076 => x"5d",
          3077 => x"f7",
          3078 => x"2e",
          3079 => x"54",
          3080 => x"f7",
          3081 => x"2e",
          3082 => x"54",
          3083 => x"06",
          3084 => x"83",
          3085 => x"2e",
          3086 => x"53",
          3087 => x"83",
          3088 => x"27",
          3089 => x"87",
          3090 => x"54",
          3091 => x"81",
          3092 => x"f7",
          3093 => x"ff",
          3094 => x"f6",
          3095 => x"83",
          3096 => x"72",
          3097 => x"10",
          3098 => x"04",
          3099 => x"2e",
          3100 => x"98",
          3101 => x"fc",
          3102 => x"33",
          3103 => x"74",
          3104 => x"c0",
          3105 => x"73",
          3106 => x"94",
          3107 => x"84",
          3108 => x"f0",
          3109 => x"08",
          3110 => x"72",
          3111 => x"76",
          3112 => x"80",
          3113 => x"57",
          3114 => x"79",
          3115 => x"38",
          3116 => x"81",
          3117 => x"06",
          3118 => x"54",
          3119 => x"80",
          3120 => x"ff",
          3121 => x"72",
          3122 => x"58",
          3123 => x"10",
          3124 => x"83",
          3125 => x"70",
          3126 => x"98",
          3127 => x"fd",
          3128 => x"ff",
          3129 => x"ff",
          3130 => x"78",
          3131 => x"84",
          3132 => x"2e",
          3133 => x"30",
          3134 => x"56",
          3135 => x"81",
          3136 => x"f9",
          3137 => x"10",
          3138 => x"54",
          3139 => x"13",
          3140 => x"73",
          3141 => x"53",
          3142 => x"b8",
          3143 => x"78",
          3144 => x"d4",
          3145 => x"3d",
          3146 => x"54",
          3147 => x"92",
          3148 => x"05",
          3149 => x"fa",
          3150 => x"15",
          3151 => x"34",
          3152 => x"fa",
          3153 => x"72",
          3154 => x"f7",
          3155 => x"fc",
          3156 => x"73",
          3157 => x"38",
          3158 => x"87",
          3159 => x"73",
          3160 => x"9c",
          3161 => x"ff",
          3162 => x"83",
          3163 => x"72",
          3164 => x"06",
          3165 => x"f7",
          3166 => x"33",
          3167 => x"33",
          3168 => x"e7",
          3169 => x"56",
          3170 => x"81",
          3171 => x"81",
          3172 => x"09",
          3173 => x"39",
          3174 => x"98",
          3175 => x"57",
          3176 => x"84",
          3177 => x"39",
          3178 => x"54",
          3179 => x"b8",
          3180 => x"81",
          3181 => x"f7",
          3182 => x"0c",
          3183 => x"70",
          3184 => x"54",
          3185 => x"74",
          3186 => x"06",
          3187 => x"83",
          3188 => x"34",
          3189 => x"06",
          3190 => x"83",
          3191 => x"34",
          3192 => x"83",
          3193 => x"f6",
          3194 => x"84",
          3195 => x"fe",
          3196 => x"90",
          3197 => x"bb",
          3198 => x"ac",
          3199 => x"0d",
          3200 => x"58",
          3201 => x"83",
          3202 => x"34",
          3203 => x"57",
          3204 => x"86",
          3205 => x"9c",
          3206 => x"ce",
          3207 => x"08",
          3208 => x"71",
          3209 => x"87",
          3210 => x"74",
          3211 => x"db",
          3212 => x"ff",
          3213 => x"72",
          3214 => x"87",
          3215 => x"05",
          3216 => x"87",
          3217 => x"2e",
          3218 => x"98",
          3219 => x"87",
          3220 => x"87",
          3221 => x"71",
          3222 => x"ff",
          3223 => x"38",
          3224 => x"d8",
          3225 => x"84",
          3226 => x"ff",
          3227 => x"76",
          3228 => x"52",
          3229 => x"ba",
          3230 => x"3d",
          3231 => x"33",
          3232 => x"08",
          3233 => x"06",
          3234 => x"56",
          3235 => x"2a",
          3236 => x"2a",
          3237 => x"16",
          3238 => x"82",
          3239 => x"80",
          3240 => x"98",
          3241 => x"34",
          3242 => x"87",
          3243 => x"08",
          3244 => x"c0",
          3245 => x"9c",
          3246 => x"81",
          3247 => x"57",
          3248 => x"81",
          3249 => x"a4",
          3250 => x"80",
          3251 => x"80",
          3252 => x"80",
          3253 => x"9c",
          3254 => x"56",
          3255 => x"33",
          3256 => x"71",
          3257 => x"2e",
          3258 => x"52",
          3259 => x"38",
          3260 => x"38",
          3261 => x"81",
          3262 => x"75",
          3263 => x"aa",
          3264 => x"11",
          3265 => x"38",
          3266 => x"70",
          3267 => x"f0",
          3268 => x"3d",
          3269 => x"52",
          3270 => x"ba",
          3271 => x"17",
          3272 => x"ff",
          3273 => x"f9",
          3274 => x"05",
          3275 => x"98",
          3276 => x"80",
          3277 => x"56",
          3278 => x"90",
          3279 => x"90",
          3280 => x"86",
          3281 => x"80",
          3282 => x"56",
          3283 => x"70",
          3284 => x"05",
          3285 => x"83",
          3286 => x"34",
          3287 => x"76",
          3288 => x"56",
          3289 => x"0b",
          3290 => x"98",
          3291 => x"80",
          3292 => x"9c",
          3293 => x"52",
          3294 => x"33",
          3295 => x"75",
          3296 => x"2e",
          3297 => x"52",
          3298 => x"38",
          3299 => x"38",
          3300 => x"90",
          3301 => x"53",
          3302 => x"73",
          3303 => x"c0",
          3304 => x"27",
          3305 => x"38",
          3306 => x"56",
          3307 => x"72",
          3308 => x"a8",
          3309 => x"fe",
          3310 => x"56",
          3311 => x"8c",
          3312 => x"70",
          3313 => x"38",
          3314 => x"74",
          3315 => x"e4",
          3316 => x"77",
          3317 => x"04",
          3318 => x"51",
          3319 => x"f4",
          3320 => x"16",
          3321 => x"34",
          3322 => x"98",
          3323 => x"87",
          3324 => x"98",
          3325 => x"38",
          3326 => x"08",
          3327 => x"71",
          3328 => x"98",
          3329 => x"27",
          3330 => x"2e",
          3331 => x"08",
          3332 => x"98",
          3333 => x"08",
          3334 => x"15",
          3335 => x"52",
          3336 => x"ff",
          3337 => x"08",
          3338 => x"38",
          3339 => x"75",
          3340 => x"06",
          3341 => x"ff",
          3342 => x"e7",
          3343 => x"51",
          3344 => x"04",
          3345 => x"7a",
          3346 => x"ff",
          3347 => x"33",
          3348 => x"83",
          3349 => x"12",
          3350 => x"07",
          3351 => x"59",
          3352 => x"81",
          3353 => x"83",
          3354 => x"2b",
          3355 => x"33",
          3356 => x"57",
          3357 => x"71",
          3358 => x"85",
          3359 => x"2b",
          3360 => x"54",
          3361 => x"81",
          3362 => x"84",
          3363 => x"33",
          3364 => x"70",
          3365 => x"77",
          3366 => x"84",
          3367 => x"86",
          3368 => x"84",
          3369 => x"34",
          3370 => x"08",
          3371 => x"88",
          3372 => x"88",
          3373 => x"34",
          3374 => x"04",
          3375 => x"8b",
          3376 => x"84",
          3377 => x"2b",
          3378 => x"51",
          3379 => x"72",
          3380 => x"70",
          3381 => x"71",
          3382 => x"5a",
          3383 => x"87",
          3384 => x"88",
          3385 => x"13",
          3386 => x"fc",
          3387 => x"71",
          3388 => x"70",
          3389 => x"72",
          3390 => x"fc",
          3391 => x"33",
          3392 => x"74",
          3393 => x"88",
          3394 => x"f8",
          3395 => x"52",
          3396 => x"77",
          3397 => x"84",
          3398 => x"81",
          3399 => x"2b",
          3400 => x"33",
          3401 => x"06",
          3402 => x"5a",
          3403 => x"81",
          3404 => x"17",
          3405 => x"8b",
          3406 => x"70",
          3407 => x"71",
          3408 => x"5a",
          3409 => x"e4",
          3410 => x"88",
          3411 => x"88",
          3412 => x"77",
          3413 => x"70",
          3414 => x"8b",
          3415 => x"82",
          3416 => x"2b",
          3417 => x"52",
          3418 => x"34",
          3419 => x"04",
          3420 => x"08",
          3421 => x"77",
          3422 => x"90",
          3423 => x"f4",
          3424 => x"0b",
          3425 => x"53",
          3426 => x"d2",
          3427 => x"76",
          3428 => x"84",
          3429 => x"34",
          3430 => x"fc",
          3431 => x"0b",
          3432 => x"84",
          3433 => x"80",
          3434 => x"88",
          3435 => x"17",
          3436 => x"f8",
          3437 => x"fc",
          3438 => x"82",
          3439 => x"fe",
          3440 => x"80",
          3441 => x"38",
          3442 => x"83",
          3443 => x"ff",
          3444 => x"11",
          3445 => x"07",
          3446 => x"ff",
          3447 => x"38",
          3448 => x"81",
          3449 => x"81",
          3450 => x"ff",
          3451 => x"5c",
          3452 => x"38",
          3453 => x"55",
          3454 => x"71",
          3455 => x"38",
          3456 => x"77",
          3457 => x"78",
          3458 => x"88",
          3459 => x"56",
          3460 => x"2e",
          3461 => x"73",
          3462 => x"80",
          3463 => x"82",
          3464 => x"78",
          3465 => x"88",
          3466 => x"74",
          3467 => x"fc",
          3468 => x"71",
          3469 => x"84",
          3470 => x"81",
          3471 => x"83",
          3472 => x"7e",
          3473 => x"5c",
          3474 => x"82",
          3475 => x"72",
          3476 => x"18",
          3477 => x"34",
          3478 => x"11",
          3479 => x"71",
          3480 => x"5c",
          3481 => x"85",
          3482 => x"16",
          3483 => x"12",
          3484 => x"2a",
          3485 => x"34",
          3486 => x"08",
          3487 => x"33",
          3488 => x"74",
          3489 => x"86",
          3490 => x"b9",
          3491 => x"84",
          3492 => x"2b",
          3493 => x"59",
          3494 => x"34",
          3495 => x"51",
          3496 => x"0d",
          3497 => x"71",
          3498 => x"05",
          3499 => x"88",
          3500 => x"59",
          3501 => x"76",
          3502 => x"70",
          3503 => x"71",
          3504 => x"05",
          3505 => x"88",
          3506 => x"5f",
          3507 => x"1a",
          3508 => x"fc",
          3509 => x"71",
          3510 => x"70",
          3511 => x"77",
          3512 => x"fc",
          3513 => x"39",
          3514 => x"08",
          3515 => x"77",
          3516 => x"8c",
          3517 => x"fb",
          3518 => x"ba",
          3519 => x"ff",
          3520 => x"80",
          3521 => x"80",
          3522 => x"fe",
          3523 => x"55",
          3524 => x"34",
          3525 => x"15",
          3526 => x"b9",
          3527 => x"81",
          3528 => x"08",
          3529 => x"80",
          3530 => x"70",
          3531 => x"88",
          3532 => x"b9",
          3533 => x"b9",
          3534 => x"76",
          3535 => x"34",
          3536 => x"38",
          3537 => x"67",
          3538 => x"08",
          3539 => x"aa",
          3540 => x"7f",
          3541 => x"84",
          3542 => x"83",
          3543 => x"06",
          3544 => x"7f",
          3545 => x"ff",
          3546 => x"33",
          3547 => x"70",
          3548 => x"70",
          3549 => x"2b",
          3550 => x"71",
          3551 => x"90",
          3552 => x"54",
          3553 => x"5f",
          3554 => x"82",
          3555 => x"2b",
          3556 => x"33",
          3557 => x"90",
          3558 => x"56",
          3559 => x"62",
          3560 => x"77",
          3561 => x"2e",
          3562 => x"62",
          3563 => x"61",
          3564 => x"70",
          3565 => x"71",
          3566 => x"81",
          3567 => x"2b",
          3568 => x"5b",
          3569 => x"76",
          3570 => x"71",
          3571 => x"11",
          3572 => x"8b",
          3573 => x"84",
          3574 => x"2b",
          3575 => x"52",
          3576 => x"77",
          3577 => x"84",
          3578 => x"33",
          3579 => x"83",
          3580 => x"87",
          3581 => x"88",
          3582 => x"41",
          3583 => x"16",
          3584 => x"33",
          3585 => x"81",
          3586 => x"5c",
          3587 => x"1a",
          3588 => x"82",
          3589 => x"2b",
          3590 => x"33",
          3591 => x"70",
          3592 => x"5a",
          3593 => x"1a",
          3594 => x"70",
          3595 => x"71",
          3596 => x"33",
          3597 => x"70",
          3598 => x"5a",
          3599 => x"83",
          3600 => x"1f",
          3601 => x"88",
          3602 => x"83",
          3603 => x"84",
          3604 => x"b9",
          3605 => x"05",
          3606 => x"44",
          3607 => x"7e",
          3608 => x"3d",
          3609 => x"b9",
          3610 => x"f8",
          3611 => x"84",
          3612 => x"84",
          3613 => x"81",
          3614 => x"08",
          3615 => x"85",
          3616 => x"60",
          3617 => x"34",
          3618 => x"22",
          3619 => x"83",
          3620 => x"5a",
          3621 => x"89",
          3622 => x"10",
          3623 => x"f8",
          3624 => x"81",
          3625 => x"08",
          3626 => x"2e",
          3627 => x"2e",
          3628 => x"3f",
          3629 => x"0c",
          3630 => x"b9",
          3631 => x"5e",
          3632 => x"33",
          3633 => x"06",
          3634 => x"40",
          3635 => x"61",
          3636 => x"2a",
          3637 => x"83",
          3638 => x"1f",
          3639 => x"2b",
          3640 => x"06",
          3641 => x"70",
          3642 => x"5b",
          3643 => x"81",
          3644 => x"34",
          3645 => x"7b",
          3646 => x"b9",
          3647 => x"88",
          3648 => x"75",
          3649 => x"54",
          3650 => x"06",
          3651 => x"82",
          3652 => x"2b",
          3653 => x"33",
          3654 => x"90",
          3655 => x"58",
          3656 => x"38",
          3657 => x"83",
          3658 => x"77",
          3659 => x"27",
          3660 => x"ff",
          3661 => x"80",
          3662 => x"80",
          3663 => x"fe",
          3664 => x"5a",
          3665 => x"34",
          3666 => x"1a",
          3667 => x"b9",
          3668 => x"81",
          3669 => x"08",
          3670 => x"80",
          3671 => x"70",
          3672 => x"64",
          3673 => x"34",
          3674 => x"10",
          3675 => x"42",
          3676 => x"61",
          3677 => x"7a",
          3678 => x"ff",
          3679 => x"38",
          3680 => x"bd",
          3681 => x"54",
          3682 => x"0d",
          3683 => x"12",
          3684 => x"07",
          3685 => x"33",
          3686 => x"7e",
          3687 => x"71",
          3688 => x"44",
          3689 => x"45",
          3690 => x"64",
          3691 => x"70",
          3692 => x"71",
          3693 => x"05",
          3694 => x"88",
          3695 => x"42",
          3696 => x"86",
          3697 => x"84",
          3698 => x"12",
          3699 => x"ff",
          3700 => x"5d",
          3701 => x"84",
          3702 => x"33",
          3703 => x"83",
          3704 => x"15",
          3705 => x"2a",
          3706 => x"54",
          3707 => x"84",
          3708 => x"81",
          3709 => x"2b",
          3710 => x"15",
          3711 => x"2a",
          3712 => x"55",
          3713 => x"34",
          3714 => x"11",
          3715 => x"07",
          3716 => x"42",
          3717 => x"51",
          3718 => x"08",
          3719 => x"06",
          3720 => x"f4",
          3721 => x"0b",
          3722 => x"53",
          3723 => x"c0",
          3724 => x"7f",
          3725 => x"84",
          3726 => x"34",
          3727 => x"fc",
          3728 => x"0b",
          3729 => x"84",
          3730 => x"80",
          3731 => x"88",
          3732 => x"1f",
          3733 => x"f8",
          3734 => x"fc",
          3735 => x"82",
          3736 => x"7e",
          3737 => x"c0",
          3738 => x"71",
          3739 => x"05",
          3740 => x"88",
          3741 => x"5e",
          3742 => x"34",
          3743 => x"fc",
          3744 => x"12",
          3745 => x"07",
          3746 => x"33",
          3747 => x"41",
          3748 => x"79",
          3749 => x"05",
          3750 => x"33",
          3751 => x"81",
          3752 => x"42",
          3753 => x"19",
          3754 => x"70",
          3755 => x"71",
          3756 => x"81",
          3757 => x"83",
          3758 => x"63",
          3759 => x"40",
          3760 => x"7b",
          3761 => x"70",
          3762 => x"8b",
          3763 => x"70",
          3764 => x"07",
          3765 => x"48",
          3766 => x"60",
          3767 => x"61",
          3768 => x"39",
          3769 => x"8b",
          3770 => x"84",
          3771 => x"2b",
          3772 => x"52",
          3773 => x"85",
          3774 => x"19",
          3775 => x"8b",
          3776 => x"86",
          3777 => x"2b",
          3778 => x"52",
          3779 => x"05",
          3780 => x"b9",
          3781 => x"33",
          3782 => x"06",
          3783 => x"77",
          3784 => x"b9",
          3785 => x"12",
          3786 => x"07",
          3787 => x"71",
          3788 => x"ff",
          3789 => x"56",
          3790 => x"55",
          3791 => x"34",
          3792 => x"33",
          3793 => x"83",
          3794 => x"12",
          3795 => x"ff",
          3796 => x"58",
          3797 => x"76",
          3798 => x"70",
          3799 => x"71",
          3800 => x"11",
          3801 => x"8b",
          3802 => x"84",
          3803 => x"2b",
          3804 => x"52",
          3805 => x"57",
          3806 => x"34",
          3807 => x"11",
          3808 => x"71",
          3809 => x"33",
          3810 => x"70",
          3811 => x"57",
          3812 => x"87",
          3813 => x"70",
          3814 => x"07",
          3815 => x"5a",
          3816 => x"81",
          3817 => x"1f",
          3818 => x"8b",
          3819 => x"73",
          3820 => x"07",
          3821 => x"5f",
          3822 => x"81",
          3823 => x"1f",
          3824 => x"2b",
          3825 => x"14",
          3826 => x"07",
          3827 => x"5f",
          3828 => x"75",
          3829 => x"70",
          3830 => x"71",
          3831 => x"70",
          3832 => x"05",
          3833 => x"84",
          3834 => x"65",
          3835 => x"5d",
          3836 => x"33",
          3837 => x"83",
          3838 => x"85",
          3839 => x"88",
          3840 => x"7a",
          3841 => x"05",
          3842 => x"84",
          3843 => x"2b",
          3844 => x"14",
          3845 => x"07",
          3846 => x"5c",
          3847 => x"34",
          3848 => x"fc",
          3849 => x"71",
          3850 => x"70",
          3851 => x"75",
          3852 => x"fc",
          3853 => x"33",
          3854 => x"74",
          3855 => x"88",
          3856 => x"f8",
          3857 => x"44",
          3858 => x"74",
          3859 => x"84",
          3860 => x"81",
          3861 => x"2b",
          3862 => x"33",
          3863 => x"06",
          3864 => x"46",
          3865 => x"81",
          3866 => x"5b",
          3867 => x"e5",
          3868 => x"84",
          3869 => x"62",
          3870 => x"51",
          3871 => x"88",
          3872 => x"b7",
          3873 => x"7a",
          3874 => x"58",
          3875 => x"77",
          3876 => x"89",
          3877 => x"3f",
          3878 => x"8c",
          3879 => x"80",
          3880 => x"b6",
          3881 => x"89",
          3882 => x"84",
          3883 => x"b9",
          3884 => x"52",
          3885 => x"3f",
          3886 => x"34",
          3887 => x"fc",
          3888 => x"0b",
          3889 => x"56",
          3890 => x"17",
          3891 => x"f8",
          3892 => x"70",
          3893 => x"58",
          3894 => x"73",
          3895 => x"70",
          3896 => x"05",
          3897 => x"34",
          3898 => x"77",
          3899 => x"39",
          3900 => x"51",
          3901 => x"84",
          3902 => x"ba",
          3903 => x"3d",
          3904 => x"53",
          3905 => x"d3",
          3906 => x"ff",
          3907 => x"ba",
          3908 => x"33",
          3909 => x"3d",
          3910 => x"60",
          3911 => x"5c",
          3912 => x"87",
          3913 => x"73",
          3914 => x"38",
          3915 => x"8c",
          3916 => x"d5",
          3917 => x"ff",
          3918 => x"87",
          3919 => x"38",
          3920 => x"80",
          3921 => x"38",
          3922 => x"8c",
          3923 => x"16",
          3924 => x"55",
          3925 => x"d5",
          3926 => x"02",
          3927 => x"57",
          3928 => x"38",
          3929 => x"81",
          3930 => x"73",
          3931 => x"0c",
          3932 => x"e7",
          3933 => x"06",
          3934 => x"c0",
          3935 => x"79",
          3936 => x"80",
          3937 => x"81",
          3938 => x"0c",
          3939 => x"81",
          3940 => x"56",
          3941 => x"39",
          3942 => x"9b",
          3943 => x"33",
          3944 => x"26",
          3945 => x"53",
          3946 => x"9b",
          3947 => x"0c",
          3948 => x"72",
          3949 => x"9a",
          3950 => x"0c",
          3951 => x"75",
          3952 => x"3d",
          3953 => x"0b",
          3954 => x"04",
          3955 => x"11",
          3956 => x"70",
          3957 => x"80",
          3958 => x"08",
          3959 => x"8c",
          3960 => x"0c",
          3961 => x"08",
          3962 => x"9b",
          3963 => x"ee",
          3964 => x"7c",
          3965 => x"5b",
          3966 => x"06",
          3967 => x"2e",
          3968 => x"81",
          3969 => x"ba",
          3970 => x"59",
          3971 => x"0d",
          3972 => x"b8",
          3973 => x"5a",
          3974 => x"8c",
          3975 => x"38",
          3976 => x"b4",
          3977 => x"a0",
          3978 => x"58",
          3979 => x"38",
          3980 => x"09",
          3981 => x"75",
          3982 => x"51",
          3983 => x"59",
          3984 => x"fb",
          3985 => x"2e",
          3986 => x"18",
          3987 => x"75",
          3988 => x"57",
          3989 => x"b6",
          3990 => x"19",
          3991 => x"0b",
          3992 => x"19",
          3993 => x"80",
          3994 => x"f2",
          3995 => x"0b",
          3996 => x"84",
          3997 => x"74",
          3998 => x"5b",
          3999 => x"2a",
          4000 => x"98",
          4001 => x"90",
          4002 => x"34",
          4003 => x"19",
          4004 => x"a6",
          4005 => x"84",
          4006 => x"05",
          4007 => x"7a",
          4008 => x"fa",
          4009 => x"53",
          4010 => x"d8",
          4011 => x"fd",
          4012 => x"0d",
          4013 => x"81",
          4014 => x"76",
          4015 => x"ba",
          4016 => x"77",
          4017 => x"cc",
          4018 => x"74",
          4019 => x"75",
          4020 => x"19",
          4021 => x"17",
          4022 => x"33",
          4023 => x"83",
          4024 => x"17",
          4025 => x"3f",
          4026 => x"38",
          4027 => x"0c",
          4028 => x"06",
          4029 => x"89",
          4030 => x"5d",
          4031 => x"38",
          4032 => x"56",
          4033 => x"84",
          4034 => x"17",
          4035 => x"3f",
          4036 => x"38",
          4037 => x"0c",
          4038 => x"06",
          4039 => x"7e",
          4040 => x"53",
          4041 => x"38",
          4042 => x"0c",
          4043 => x"a8",
          4044 => x"79",
          4045 => x"33",
          4046 => x"09",
          4047 => x"78",
          4048 => x"51",
          4049 => x"80",
          4050 => x"78",
          4051 => x"75",
          4052 => x"05",
          4053 => x"2b",
          4054 => x"8f",
          4055 => x"81",
          4056 => x"a8",
          4057 => x"79",
          4058 => x"33",
          4059 => x"09",
          4060 => x"78",
          4061 => x"51",
          4062 => x"80",
          4063 => x"78",
          4064 => x"75",
          4065 => x"b8",
          4066 => x"71",
          4067 => x"14",
          4068 => x"33",
          4069 => x"07",
          4070 => x"59",
          4071 => x"54",
          4072 => x"53",
          4073 => x"3f",
          4074 => x"2e",
          4075 => x"ba",
          4076 => x"08",
          4077 => x"08",
          4078 => x"fe",
          4079 => x"82",
          4080 => x"81",
          4081 => x"05",
          4082 => x"f6",
          4083 => x"81",
          4084 => x"70",
          4085 => x"81",
          4086 => x"09",
          4087 => x"8c",
          4088 => x"a8",
          4089 => x"08",
          4090 => x"7d",
          4091 => x"8c",
          4092 => x"b4",
          4093 => x"81",
          4094 => x"81",
          4095 => x"09",
          4096 => x"8c",
          4097 => x"a8",
          4098 => x"5b",
          4099 => x"c5",
          4100 => x"2e",
          4101 => x"54",
          4102 => x"53",
          4103 => x"f1",
          4104 => x"54",
          4105 => x"53",
          4106 => x"3f",
          4107 => x"2e",
          4108 => x"ba",
          4109 => x"08",
          4110 => x"08",
          4111 => x"fb",
          4112 => x"82",
          4113 => x"81",
          4114 => x"05",
          4115 => x"f4",
          4116 => x"81",
          4117 => x"05",
          4118 => x"f3",
          4119 => x"7a",
          4120 => x"3d",
          4121 => x"82",
          4122 => x"9c",
          4123 => x"55",
          4124 => x"24",
          4125 => x"8a",
          4126 => x"3d",
          4127 => x"08",
          4128 => x"58",
          4129 => x"83",
          4130 => x"2e",
          4131 => x"54",
          4132 => x"33",
          4133 => x"08",
          4134 => x"5a",
          4135 => x"ff",
          4136 => x"79",
          4137 => x"5e",
          4138 => x"5a",
          4139 => x"1a",
          4140 => x"3d",
          4141 => x"06",
          4142 => x"1a",
          4143 => x"08",
          4144 => x"38",
          4145 => x"7c",
          4146 => x"81",
          4147 => x"19",
          4148 => x"8c",
          4149 => x"81",
          4150 => x"79",
          4151 => x"fc",
          4152 => x"33",
          4153 => x"f0",
          4154 => x"7d",
          4155 => x"b9",
          4156 => x"ba",
          4157 => x"bb",
          4158 => x"fe",
          4159 => x"89",
          4160 => x"08",
          4161 => x"38",
          4162 => x"56",
          4163 => x"82",
          4164 => x"19",
          4165 => x"3f",
          4166 => x"38",
          4167 => x"0c",
          4168 => x"83",
          4169 => x"77",
          4170 => x"7c",
          4171 => x"9f",
          4172 => x"07",
          4173 => x"83",
          4174 => x"08",
          4175 => x"56",
          4176 => x"81",
          4177 => x"81",
          4178 => x"81",
          4179 => x"09",
          4180 => x"8c",
          4181 => x"70",
          4182 => x"84",
          4183 => x"74",
          4184 => x"55",
          4185 => x"54",
          4186 => x"51",
          4187 => x"80",
          4188 => x"75",
          4189 => x"7d",
          4190 => x"84",
          4191 => x"88",
          4192 => x"8f",
          4193 => x"81",
          4194 => x"81",
          4195 => x"81",
          4196 => x"81",
          4197 => x"09",
          4198 => x"8c",
          4199 => x"70",
          4200 => x"84",
          4201 => x"7e",
          4202 => x"33",
          4203 => x"fb",
          4204 => x"7c",
          4205 => x"3f",
          4206 => x"76",
          4207 => x"33",
          4208 => x"84",
          4209 => x"06",
          4210 => x"83",
          4211 => x"1b",
          4212 => x"8c",
          4213 => x"27",
          4214 => x"74",
          4215 => x"38",
          4216 => x"81",
          4217 => x"5c",
          4218 => x"b8",
          4219 => x"57",
          4220 => x"8c",
          4221 => x"c5",
          4222 => x"34",
          4223 => x"31",
          4224 => x"5d",
          4225 => x"87",
          4226 => x"2e",
          4227 => x"54",
          4228 => x"33",
          4229 => x"e7",
          4230 => x"52",
          4231 => x"7e",
          4232 => x"83",
          4233 => x"ff",
          4234 => x"34",
          4235 => x"34",
          4236 => x"39",
          4237 => x"7a",
          4238 => x"98",
          4239 => x"06",
          4240 => x"7d",
          4241 => x"1d",
          4242 => x"1d",
          4243 => x"1d",
          4244 => x"7c",
          4245 => x"81",
          4246 => x"80",
          4247 => x"08",
          4248 => x"70",
          4249 => x"38",
          4250 => x"56",
          4251 => x"26",
          4252 => x"82",
          4253 => x"f5",
          4254 => x"81",
          4255 => x"08",
          4256 => x"08",
          4257 => x"25",
          4258 => x"73",
          4259 => x"81",
          4260 => x"84",
          4261 => x"81",
          4262 => x"08",
          4263 => x"f0",
          4264 => x"8c",
          4265 => x"08",
          4266 => x"ce",
          4267 => x"08",
          4268 => x"39",
          4269 => x"26",
          4270 => x"51",
          4271 => x"8c",
          4272 => x"ba",
          4273 => x"07",
          4274 => x"8c",
          4275 => x"ff",
          4276 => x"2e",
          4277 => x"74",
          4278 => x"08",
          4279 => x"57",
          4280 => x"8e",
          4281 => x"f5",
          4282 => x"ba",
          4283 => x"08",
          4284 => x"80",
          4285 => x"90",
          4286 => x"94",
          4287 => x"86",
          4288 => x"19",
          4289 => x"34",
          4290 => x"8c",
          4291 => x"8c",
          4292 => x"8c",
          4293 => x"2e",
          4294 => x"78",
          4295 => x"08",
          4296 => x"08",
          4297 => x"04",
          4298 => x"38",
          4299 => x"0d",
          4300 => x"73",
          4301 => x"73",
          4302 => x"73",
          4303 => x"74",
          4304 => x"82",
          4305 => x"53",
          4306 => x"72",
          4307 => x"98",
          4308 => x"18",
          4309 => x"94",
          4310 => x"0c",
          4311 => x"9c",
          4312 => x"8c",
          4313 => x"84",
          4314 => x"ac",
          4315 => x"ac",
          4316 => x"57",
          4317 => x"17",
          4318 => x"56",
          4319 => x"8a",
          4320 => x"08",
          4321 => x"ff",
          4322 => x"cd",
          4323 => x"ba",
          4324 => x"0b",
          4325 => x"38",
          4326 => x"08",
          4327 => x"31",
          4328 => x"aa",
          4329 => x"8a",
          4330 => x"70",
          4331 => x"5a",
          4332 => x"38",
          4333 => x"08",
          4334 => x"38",
          4335 => x"38",
          4336 => x"75",
          4337 => x"22",
          4338 => x"38",
          4339 => x"0c",
          4340 => x"80",
          4341 => x"3d",
          4342 => x"19",
          4343 => x"5c",
          4344 => x"eb",
          4345 => x"82",
          4346 => x"27",
          4347 => x"08",
          4348 => x"84",
          4349 => x"60",
          4350 => x"08",
          4351 => x"ba",
          4352 => x"8c",
          4353 => x"56",
          4354 => x"91",
          4355 => x"ff",
          4356 => x"08",
          4357 => x"ea",
          4358 => x"05",
          4359 => x"8d",
          4360 => x"b0",
          4361 => x"1a",
          4362 => x"57",
          4363 => x"34",
          4364 => x"56",
          4365 => x"81",
          4366 => x"77",
          4367 => x"3f",
          4368 => x"81",
          4369 => x"0c",
          4370 => x"3d",
          4371 => x"53",
          4372 => x"52",
          4373 => x"08",
          4374 => x"83",
          4375 => x"08",
          4376 => x"fe",
          4377 => x"82",
          4378 => x"81",
          4379 => x"05",
          4380 => x"e3",
          4381 => x"22",
          4382 => x"74",
          4383 => x"7c",
          4384 => x"08",
          4385 => x"7d",
          4386 => x"76",
          4387 => x"19",
          4388 => x"84",
          4389 => x"ee",
          4390 => x"7c",
          4391 => x"1e",
          4392 => x"82",
          4393 => x"80",
          4394 => x"d1",
          4395 => x"74",
          4396 => x"38",
          4397 => x"81",
          4398 => x"ba",
          4399 => x"5a",
          4400 => x"5b",
          4401 => x"70",
          4402 => x"81",
          4403 => x"81",
          4404 => x"34",
          4405 => x"ae",
          4406 => x"80",
          4407 => x"74",
          4408 => x"56",
          4409 => x"60",
          4410 => x"80",
          4411 => x"ba",
          4412 => x"81",
          4413 => x"fe",
          4414 => x"94",
          4415 => x"08",
          4416 => x"e1",
          4417 => x"08",
          4418 => x"38",
          4419 => x"b4",
          4420 => x"ba",
          4421 => x"08",
          4422 => x"41",
          4423 => x"a8",
          4424 => x"1a",
          4425 => x"33",
          4426 => x"90",
          4427 => x"81",
          4428 => x"5b",
          4429 => x"33",
          4430 => x"08",
          4431 => x"76",
          4432 => x"74",
          4433 => x"60",
          4434 => x"c1",
          4435 => x"0c",
          4436 => x"0d",
          4437 => x"18",
          4438 => x"06",
          4439 => x"33",
          4440 => x"58",
          4441 => x"33",
          4442 => x"05",
          4443 => x"e6",
          4444 => x"33",
          4445 => x"44",
          4446 => x"79",
          4447 => x"10",
          4448 => x"23",
          4449 => x"77",
          4450 => x"2a",
          4451 => x"90",
          4452 => x"38",
          4453 => x"23",
          4454 => x"41",
          4455 => x"2e",
          4456 => x"39",
          4457 => x"74",
          4458 => x"78",
          4459 => x"05",
          4460 => x"56",
          4461 => x"fd",
          4462 => x"7a",
          4463 => x"04",
          4464 => x"5c",
          4465 => x"84",
          4466 => x"08",
          4467 => x"5d",
          4468 => x"5e",
          4469 => x"1b",
          4470 => x"1b",
          4471 => x"09",
          4472 => x"75",
          4473 => x"51",
          4474 => x"80",
          4475 => x"75",
          4476 => x"b2",
          4477 => x"59",
          4478 => x"19",
          4479 => x"57",
          4480 => x"e5",
          4481 => x"81",
          4482 => x"38",
          4483 => x"81",
          4484 => x"56",
          4485 => x"81",
          4486 => x"5a",
          4487 => x"06",
          4488 => x"38",
          4489 => x"1c",
          4490 => x"8b",
          4491 => x"81",
          4492 => x"5a",
          4493 => x"58",
          4494 => x"38",
          4495 => x"5d",
          4496 => x"7b",
          4497 => x"08",
          4498 => x"fe",
          4499 => x"93",
          4500 => x"08",
          4501 => x"dc",
          4502 => x"08",
          4503 => x"38",
          4504 => x"b4",
          4505 => x"ba",
          4506 => x"08",
          4507 => x"5a",
          4508 => x"dd",
          4509 => x"1c",
          4510 => x"33",
          4511 => x"c5",
          4512 => x"1c",
          4513 => x"55",
          4514 => x"81",
          4515 => x"8d",
          4516 => x"90",
          4517 => x"5e",
          4518 => x"ff",
          4519 => x"f4",
          4520 => x"84",
          4521 => x"38",
          4522 => x"c2",
          4523 => x"1d",
          4524 => x"57",
          4525 => x"38",
          4526 => x"1b",
          4527 => x"40",
          4528 => x"bf",
          4529 => x"81",
          4530 => x"33",
          4531 => x"71",
          4532 => x"80",
          4533 => x"26",
          4534 => x"8a",
          4535 => x"61",
          4536 => x"5b",
          4537 => x"ba",
          4538 => x"de",
          4539 => x"78",
          4540 => x"86",
          4541 => x"2e",
          4542 => x"79",
          4543 => x"7f",
          4544 => x"ff",
          4545 => x"0b",
          4546 => x"04",
          4547 => x"38",
          4548 => x"3d",
          4549 => x"33",
          4550 => x"86",
          4551 => x"1d",
          4552 => x"80",
          4553 => x"17",
          4554 => x"38",
          4555 => x"60",
          4556 => x"05",
          4557 => x"34",
          4558 => x"80",
          4559 => x"56",
          4560 => x"c0",
          4561 => x"3d",
          4562 => x"59",
          4563 => x"70",
          4564 => x"05",
          4565 => x"38",
          4566 => x"79",
          4567 => x"38",
          4568 => x"75",
          4569 => x"2a",
          4570 => x"2a",
          4571 => x"80",
          4572 => x"32",
          4573 => x"d7",
          4574 => x"87",
          4575 => x"58",
          4576 => x"75",
          4577 => x"76",
          4578 => x"2a",
          4579 => x"1f",
          4580 => x"58",
          4581 => x"33",
          4582 => x"16",
          4583 => x"75",
          4584 => x"2e",
          4585 => x"56",
          4586 => x"98",
          4587 => x"71",
          4588 => x"87",
          4589 => x"f8",
          4590 => x"38",
          4591 => x"fe",
          4592 => x"2e",
          4593 => x"56",
          4594 => x"81",
          4595 => x"05",
          4596 => x"84",
          4597 => x"75",
          4598 => x"7e",
          4599 => x"1d",
          4600 => x"8c",
          4601 => x"ed",
          4602 => x"84",
          4603 => x"ba",
          4604 => x"1e",
          4605 => x"76",
          4606 => x"40",
          4607 => x"a3",
          4608 => x"52",
          4609 => x"84",
          4610 => x"ff",
          4611 => x"76",
          4612 => x"70",
          4613 => x"81",
          4614 => x"78",
          4615 => x"c9",
          4616 => x"86",
          4617 => x"83",
          4618 => x"ba",
          4619 => x"87",
          4620 => x"75",
          4621 => x"40",
          4622 => x"57",
          4623 => x"83",
          4624 => x"82",
          4625 => x"52",
          4626 => x"84",
          4627 => x"ff",
          4628 => x"75",
          4629 => x"9c",
          4630 => x"81",
          4631 => x"f4",
          4632 => x"58",
          4633 => x"33",
          4634 => x"15",
          4635 => x"ab",
          4636 => x"8c",
          4637 => x"77",
          4638 => x"3d",
          4639 => x"25",
          4640 => x"b9",
          4641 => x"ec",
          4642 => x"84",
          4643 => x"38",
          4644 => x"08",
          4645 => x"d3",
          4646 => x"2e",
          4647 => x"ba",
          4648 => x"08",
          4649 => x"19",
          4650 => x"41",
          4651 => x"ba",
          4652 => x"85",
          4653 => x"58",
          4654 => x"8c",
          4655 => x"ef",
          4656 => x"58",
          4657 => x"80",
          4658 => x"33",
          4659 => x"ff",
          4660 => x"74",
          4661 => x"98",
          4662 => x"08",
          4663 => x"5b",
          4664 => x"c9",
          4665 => x"52",
          4666 => x"84",
          4667 => x"ff",
          4668 => x"75",
          4669 => x"08",
          4670 => x"5f",
          4671 => x"0b",
          4672 => x"75",
          4673 => x"7c",
          4674 => x"58",
          4675 => x"38",
          4676 => x"5b",
          4677 => x"7b",
          4678 => x"57",
          4679 => x"34",
          4680 => x"81",
          4681 => x"76",
          4682 => x"78",
          4683 => x"80",
          4684 => x"81",
          4685 => x"51",
          4686 => x"58",
          4687 => x"7f",
          4688 => x"fb",
          4689 => x"53",
          4690 => x"52",
          4691 => x"ba",
          4692 => x"8c",
          4693 => x"a8",
          4694 => x"57",
          4695 => x"c9",
          4696 => x"2e",
          4697 => x"54",
          4698 => x"53",
          4699 => x"d1",
          4700 => x"9c",
          4701 => x"74",
          4702 => x"ba",
          4703 => x"57",
          4704 => x"d7",
          4705 => x"d4",
          4706 => x"61",
          4707 => x"3f",
          4708 => x"81",
          4709 => x"83",
          4710 => x"08",
          4711 => x"8a",
          4712 => x"2e",
          4713 => x"fc",
          4714 => x"7f",
          4715 => x"39",
          4716 => x"70",
          4717 => x"38",
          4718 => x"08",
          4719 => x"81",
          4720 => x"c1",
          4721 => x"19",
          4722 => x"33",
          4723 => x"f3",
          4724 => x"5e",
          4725 => x"1c",
          4726 => x"1c",
          4727 => x"70",
          4728 => x"57",
          4729 => x"bc",
          4730 => x"81",
          4731 => x"38",
          4732 => x"ff",
          4733 => x"82",
          4734 => x"70",
          4735 => x"38",
          4736 => x"7a",
          4737 => x"05",
          4738 => x"70",
          4739 => x"08",
          4740 => x"53",
          4741 => x"2e",
          4742 => x"30",
          4743 => x"54",
          4744 => x"2e",
          4745 => x"59",
          4746 => x"81",
          4747 => x"76",
          4748 => x"05",
          4749 => x"1d",
          4750 => x"f3",
          4751 => x"57",
          4752 => x"82",
          4753 => x"33",
          4754 => x"1e",
          4755 => x"33",
          4756 => x"11",
          4757 => x"90",
          4758 => x"33",
          4759 => x"71",
          4760 => x"96",
          4761 => x"41",
          4762 => x"86",
          4763 => x"33",
          4764 => x"84",
          4765 => x"e5",
          4766 => x"11",
          4767 => x"83",
          4768 => x"51",
          4769 => x"08",
          4770 => x"75",
          4771 => x"b3",
          4772 => x"34",
          4773 => x"58",
          4774 => x"78",
          4775 => x"54",
          4776 => x"74",
          4777 => x"25",
          4778 => x"75",
          4779 => x"78",
          4780 => x"56",
          4781 => x"33",
          4782 => x"88",
          4783 => x"54",
          4784 => x"54",
          4785 => x"08",
          4786 => x"27",
          4787 => x"81",
          4788 => x"a0",
          4789 => x"53",
          4790 => x"81",
          4791 => x"13",
          4792 => x"ff",
          4793 => x"2a",
          4794 => x"80",
          4795 => x"5f",
          4796 => x"63",
          4797 => x"65",
          4798 => x"2e",
          4799 => x"2e",
          4800 => x"d9",
          4801 => x"73",
          4802 => x"55",
          4803 => x"42",
          4804 => x"70",
          4805 => x"73",
          4806 => x"ff",
          4807 => x"74",
          4808 => x"80",
          4809 => x"ff",
          4810 => x"9f",
          4811 => x"5b",
          4812 => x"80",
          4813 => x"ff",
          4814 => x"83",
          4815 => x"56",
          4816 => x"38",
          4817 => x"70",
          4818 => x"56",
          4819 => x"5b",
          4820 => x"26",
          4821 => x"74",
          4822 => x"81",
          4823 => x"80",
          4824 => x"81",
          4825 => x"80",
          4826 => x"72",
          4827 => x"46",
          4828 => x"af",
          4829 => x"70",
          4830 => x"54",
          4831 => x"0c",
          4832 => x"42",
          4833 => x"b4",
          4834 => x"8d",
          4835 => x"ff",
          4836 => x"86",
          4837 => x"3d",
          4838 => x"81",
          4839 => x"fe",
          4840 => x"ab",
          4841 => x"8d",
          4842 => x"8c",
          4843 => x"80",
          4844 => x"73",
          4845 => x"2e",
          4846 => x"70",
          4847 => x"dd",
          4848 => x"70",
          4849 => x"7d",
          4850 => x"27",
          4851 => x"f8",
          4852 => x"76",
          4853 => x"76",
          4854 => x"70",
          4855 => x"52",
          4856 => x"2e",
          4857 => x"57",
          4858 => x"56",
          4859 => x"c7",
          4860 => x"ff",
          4861 => x"a0",
          4862 => x"ff",
          4863 => x"38",
          4864 => x"fe",
          4865 => x"2e",
          4866 => x"54",
          4867 => x"38",
          4868 => x"ae",
          4869 => x"0b",
          4870 => x"81",
          4871 => x"f4",
          4872 => x"16",
          4873 => x"5d",
          4874 => x"a0",
          4875 => x"70",
          4876 => x"75",
          4877 => x"bb",
          4878 => x"38",
          4879 => x"70",
          4880 => x"51",
          4881 => x"e0",
          4882 => x"75",
          4883 => x"5a",
          4884 => x"88",
          4885 => x"06",
          4886 => x"70",
          4887 => x"ff",
          4888 => x"81",
          4889 => x"2e",
          4890 => x"77",
          4891 => x"06",
          4892 => x"79",
          4893 => x"38",
          4894 => x"85",
          4895 => x"2a",
          4896 => x"38",
          4897 => x"34",
          4898 => x"8c",
          4899 => x"ba",
          4900 => x"84",
          4901 => x"06",
          4902 => x"06",
          4903 => x"74",
          4904 => x"98",
          4905 => x"42",
          4906 => x"ce",
          4907 => x"70",
          4908 => x"2e",
          4909 => x"38",
          4910 => x"82",
          4911 => x"81",
          4912 => x"73",
          4913 => x"38",
          4914 => x"80",
          4915 => x"76",
          4916 => x"75",
          4917 => x"53",
          4918 => x"07",
          4919 => x"e3",
          4920 => x"1d",
          4921 => x"fe",
          4922 => x"58",
          4923 => x"70",
          4924 => x"80",
          4925 => x"83",
          4926 => x"33",
          4927 => x"07",
          4928 => x"83",
          4929 => x"0c",
          4930 => x"39",
          4931 => x"f0",
          4932 => x"38",
          4933 => x"17",
          4934 => x"2b",
          4935 => x"5e",
          4936 => x"95",
          4937 => x"39",
          4938 => x"2e",
          4939 => x"39",
          4940 => x"0b",
          4941 => x"04",
          4942 => x"ff",
          4943 => x"59",
          4944 => x"83",
          4945 => x"fc",
          4946 => x"b5",
          4947 => x"84",
          4948 => x"70",
          4949 => x"80",
          4950 => x"83",
          4951 => x"81",
          4952 => x"2e",
          4953 => x"83",
          4954 => x"56",
          4955 => x"38",
          4956 => x"70",
          4957 => x"59",
          4958 => x"59",
          4959 => x"54",
          4960 => x"07",
          4961 => x"9f",
          4962 => x"7d",
          4963 => x"17",
          4964 => x"5f",
          4965 => x"79",
          4966 => x"fa",
          4967 => x"83",
          4968 => x"5a",
          4969 => x"80",
          4970 => x"05",
          4971 => x"1b",
          4972 => x"80",
          4973 => x"90",
          4974 => x"5a",
          4975 => x"05",
          4976 => x"34",
          4977 => x"5b",
          4978 => x"9c",
          4979 => x"58",
          4980 => x"06",
          4981 => x"82",
          4982 => x"38",
          4983 => x"3d",
          4984 => x"02",
          4985 => x"42",
          4986 => x"70",
          4987 => x"d7",
          4988 => x"70",
          4989 => x"85",
          4990 => x"2e",
          4991 => x"56",
          4992 => x"10",
          4993 => x"58",
          4994 => x"96",
          4995 => x"06",
          4996 => x"9b",
          4997 => x"b0",
          4998 => x"06",
          4999 => x"2e",
          5000 => x"16",
          5001 => x"18",
          5002 => x"ff",
          5003 => x"81",
          5004 => x"83",
          5005 => x"2e",
          5006 => x"41",
          5007 => x"5b",
          5008 => x"18",
          5009 => x"7a",
          5010 => x"33",
          5011 => x"ba",
          5012 => x"55",
          5013 => x"56",
          5014 => x"84",
          5015 => x"56",
          5016 => x"2e",
          5017 => x"38",
          5018 => x"85",
          5019 => x"83",
          5020 => x"83",
          5021 => x"c3",
          5022 => x"59",
          5023 => x"83",
          5024 => x"ce",
          5025 => x"5a",
          5026 => x"11",
          5027 => x"71",
          5028 => x"72",
          5029 => x"56",
          5030 => x"a0",
          5031 => x"18",
          5032 => x"70",
          5033 => x"58",
          5034 => x"81",
          5035 => x"19",
          5036 => x"23",
          5037 => x"38",
          5038 => x"bb",
          5039 => x"18",
          5040 => x"74",
          5041 => x"5e",
          5042 => x"80",
          5043 => x"71",
          5044 => x"38",
          5045 => x"12",
          5046 => x"07",
          5047 => x"2b",
          5048 => x"58",
          5049 => x"80",
          5050 => x"5d",
          5051 => x"ce",
          5052 => x"5a",
          5053 => x"52",
          5054 => x"3f",
          5055 => x"8c",
          5056 => x"ba",
          5057 => x"26",
          5058 => x"f5",
          5059 => x"f5",
          5060 => x"16",
          5061 => x"0c",
          5062 => x"1d",
          5063 => x"2e",
          5064 => x"8d",
          5065 => x"7d",
          5066 => x"7c",
          5067 => x"70",
          5068 => x"5a",
          5069 => x"58",
          5070 => x"ff",
          5071 => x"18",
          5072 => x"7c",
          5073 => x"34",
          5074 => x"7c",
          5075 => x"23",
          5076 => x"80",
          5077 => x"84",
          5078 => x"8b",
          5079 => x"0d",
          5080 => x"ff",
          5081 => x"91",
          5082 => x"d0",
          5083 => x"fe",
          5084 => x"5f",
          5085 => x"7a",
          5086 => x"81",
          5087 => x"58",
          5088 => x"16",
          5089 => x"9f",
          5090 => x"e0",
          5091 => x"75",
          5092 => x"77",
          5093 => x"ff",
          5094 => x"70",
          5095 => x"58",
          5096 => x"81",
          5097 => x"25",
          5098 => x"39",
          5099 => x"82",
          5100 => x"fe",
          5101 => x"7a",
          5102 => x"2e",
          5103 => x"75",
          5104 => x"25",
          5105 => x"ad",
          5106 => x"38",
          5107 => x"83",
          5108 => x"80",
          5109 => x"84",
          5110 => x"88",
          5111 => x"72",
          5112 => x"71",
          5113 => x"77",
          5114 => x"19",
          5115 => x"ff",
          5116 => x"70",
          5117 => x"9b",
          5118 => x"84",
          5119 => x"42",
          5120 => x"2e",
          5121 => x"34",
          5122 => x"80",
          5123 => x"54",
          5124 => x"33",
          5125 => x"8c",
          5126 => x"81",
          5127 => x"75",
          5128 => x"71",
          5129 => x"7b",
          5130 => x"a8",
          5131 => x"58",
          5132 => x"75",
          5133 => x"25",
          5134 => x"38",
          5135 => x"58",
          5136 => x"84",
          5137 => x"78",
          5138 => x"58",
          5139 => x"80",
          5140 => x"1a",
          5141 => x"38",
          5142 => x"18",
          5143 => x"70",
          5144 => x"05",
          5145 => x"5b",
          5146 => x"c5",
          5147 => x"0b",
          5148 => x"5d",
          5149 => x"7e",
          5150 => x"31",
          5151 => x"80",
          5152 => x"e1",
          5153 => x"58",
          5154 => x"8c",
          5155 => x"75",
          5156 => x"81",
          5157 => x"58",
          5158 => x"8c",
          5159 => x"80",
          5160 => x"58",
          5161 => x"70",
          5162 => x"ff",
          5163 => x"2e",
          5164 => x"38",
          5165 => x"c0",
          5166 => x"5a",
          5167 => x"71",
          5168 => x"40",
          5169 => x"80",
          5170 => x"5a",
          5171 => x"fd",
          5172 => x"e8",
          5173 => x"55",
          5174 => x"d5",
          5175 => x"17",
          5176 => x"33",
          5177 => x"82",
          5178 => x"17",
          5179 => x"d2",
          5180 => x"85",
          5181 => x"18",
          5182 => x"18",
          5183 => x"18",
          5184 => x"75",
          5185 => x"f8",
          5186 => x"82",
          5187 => x"2b",
          5188 => x"88",
          5189 => x"59",
          5190 => x"85",
          5191 => x"cd",
          5192 => x"82",
          5193 => x"2b",
          5194 => x"88",
          5195 => x"40",
          5196 => x"85",
          5197 => x"9d",
          5198 => x"82",
          5199 => x"2b",
          5200 => x"88",
          5201 => x"0c",
          5202 => x"82",
          5203 => x"2b",
          5204 => x"88",
          5205 => x"05",
          5206 => x"40",
          5207 => x"84",
          5208 => x"84",
          5209 => x"84",
          5210 => x"0b",
          5211 => x"83",
          5212 => x"0c",
          5213 => x"17",
          5214 => x"18",
          5215 => x"84",
          5216 => x"06",
          5217 => x"83",
          5218 => x"08",
          5219 => x"8b",
          5220 => x"2e",
          5221 => x"5a",
          5222 => x"2e",
          5223 => x"18",
          5224 => x"ab",
          5225 => x"18",
          5226 => x"8d",
          5227 => x"22",
          5228 => x"17",
          5229 => x"90",
          5230 => x"33",
          5231 => x"71",
          5232 => x"2b",
          5233 => x"d8",
          5234 => x"e8",
          5235 => x"80",
          5236 => x"57",
          5237 => x"5a",
          5238 => x"75",
          5239 => x"05",
          5240 => x"ff",
          5241 => x"3d",
          5242 => x"70",
          5243 => x"76",
          5244 => x"38",
          5245 => x"9f",
          5246 => x"e2",
          5247 => x"80",
          5248 => x"80",
          5249 => x"10",
          5250 => x"55",
          5251 => x"34",
          5252 => x"80",
          5253 => x"7c",
          5254 => x"53",
          5255 => x"ef",
          5256 => x"73",
          5257 => x"04",
          5258 => x"3d",
          5259 => x"81",
          5260 => x"26",
          5261 => x"06",
          5262 => x"80",
          5263 => x"fc",
          5264 => x"5a",
          5265 => x"70",
          5266 => x"59",
          5267 => x"e0",
          5268 => x"ff",
          5269 => x"38",
          5270 => x"54",
          5271 => x"74",
          5272 => x"76",
          5273 => x"30",
          5274 => x"5c",
          5275 => x"81",
          5276 => x"25",
          5277 => x"39",
          5278 => x"60",
          5279 => x"0d",
          5280 => x"33",
          5281 => x"a6",
          5282 => x"3d",
          5283 => x"52",
          5284 => x"08",
          5285 => x"8f",
          5286 => x"84",
          5287 => x"7e",
          5288 => x"5a",
          5289 => x"57",
          5290 => x"ba",
          5291 => x"2e",
          5292 => x"c1",
          5293 => x"77",
          5294 => x"77",
          5295 => x"2e",
          5296 => x"9a",
          5297 => x"70",
          5298 => x"83",
          5299 => x"17",
          5300 => x"0b",
          5301 => x"17",
          5302 => x"34",
          5303 => x"17",
          5304 => x"33",
          5305 => x"66",
          5306 => x"0b",
          5307 => x"34",
          5308 => x"81",
          5309 => x"80",
          5310 => x"7c",
          5311 => x"27",
          5312 => x"83",
          5313 => x"fe",
          5314 => x"70",
          5315 => x"fe",
          5316 => x"57",
          5317 => x"38",
          5318 => x"2a",
          5319 => x"38",
          5320 => x"80",
          5321 => x"79",
          5322 => x"06",
          5323 => x"80",
          5324 => x"a0",
          5325 => x"9b",
          5326 => x"2b",
          5327 => x"5a",
          5328 => x"88",
          5329 => x"82",
          5330 => x"2b",
          5331 => x"88",
          5332 => x"8c",
          5333 => x"41",
          5334 => x"84",
          5335 => x"0b",
          5336 => x"0c",
          5337 => x"80",
          5338 => x"84",
          5339 => x"1a",
          5340 => x"58",
          5341 => x"56",
          5342 => x"81",
          5343 => x"2e",
          5344 => x"ff",
          5345 => x"58",
          5346 => x"38",
          5347 => x"2e",
          5348 => x"c0",
          5349 => x"06",
          5350 => x"81",
          5351 => x"38",
          5352 => x"39",
          5353 => x"39",
          5354 => x"39",
          5355 => x"8c",
          5356 => x"fb",
          5357 => x"7b",
          5358 => x"16",
          5359 => x"71",
          5360 => x"5c",
          5361 => x"27",
          5362 => x"ff",
          5363 => x"5d",
          5364 => x"a7",
          5365 => x"fc",
          5366 => x"2e",
          5367 => x"76",
          5368 => x"8c",
          5369 => x"fe",
          5370 => x"75",
          5371 => x"94",
          5372 => x"55",
          5373 => x"7d",
          5374 => x"80",
          5375 => x"17",
          5376 => x"94",
          5377 => x"2b",
          5378 => x"0b",
          5379 => x"34",
          5380 => x"0b",
          5381 => x"8b",
          5382 => x"0b",
          5383 => x"34",
          5384 => x"81",
          5385 => x"80",
          5386 => x"b4",
          5387 => x"16",
          5388 => x"06",
          5389 => x"16",
          5390 => x"ba",
          5391 => x"85",
          5392 => x"17",
          5393 => x"18",
          5394 => x"38",
          5395 => x"54",
          5396 => x"53",
          5397 => x"81",
          5398 => x"09",
          5399 => x"8c",
          5400 => x"a8",
          5401 => x"5c",
          5402 => x"92",
          5403 => x"2e",
          5404 => x"54",
          5405 => x"53",
          5406 => x"a3",
          5407 => x"74",
          5408 => x"39",
          5409 => x"38",
          5410 => x"2e",
          5411 => x"12",
          5412 => x"7d",
          5413 => x"78",
          5414 => x"5c",
          5415 => x"89",
          5416 => x"f7",
          5417 => x"56",
          5418 => x"0c",
          5419 => x"57",
          5420 => x"7f",
          5421 => x"0d",
          5422 => x"5a",
          5423 => x"2e",
          5424 => x"2e",
          5425 => x"2e",
          5426 => x"22",
          5427 => x"38",
          5428 => x"82",
          5429 => x"82",
          5430 => x"57",
          5431 => x"38",
          5432 => x"31",
          5433 => x"38",
          5434 => x"59",
          5435 => x"e3",
          5436 => x"89",
          5437 => x"83",
          5438 => x"75",
          5439 => x"83",
          5440 => x"59",
          5441 => x"08",
          5442 => x"83",
          5443 => x"29",
          5444 => x"80",
          5445 => x"89",
          5446 => x"81",
          5447 => x"85",
          5448 => x"76",
          5449 => x"ff",
          5450 => x"83",
          5451 => x"59",
          5452 => x"08",
          5453 => x"38",
          5454 => x"1b",
          5455 => x"57",
          5456 => x"ff",
          5457 => x"2b",
          5458 => x"7f",
          5459 => x"70",
          5460 => x"fe",
          5461 => x"8c",
          5462 => x"ba",
          5463 => x"5c",
          5464 => x"75",
          5465 => x"59",
          5466 => x"58",
          5467 => x"b6",
          5468 => x"5d",
          5469 => x"06",
          5470 => x"b8",
          5471 => x"9e",
          5472 => x"2e",
          5473 => x"b4",
          5474 => x"94",
          5475 => x"7f",
          5476 => x"80",
          5477 => x"05",
          5478 => x"34",
          5479 => x"d1",
          5480 => x"77",
          5481 => x"56",
          5482 => x"54",
          5483 => x"53",
          5484 => x"c9",
          5485 => x"7f",
          5486 => x"84",
          5487 => x"19",
          5488 => x"8c",
          5489 => x"27",
          5490 => x"74",
          5491 => x"38",
          5492 => x"08",
          5493 => x"51",
          5494 => x"bb",
          5495 => x"08",
          5496 => x"52",
          5497 => x"ba",
          5498 => x"16",
          5499 => x"ba",
          5500 => x"b8",
          5501 => x"b2",
          5502 => x"0b",
          5503 => x"04",
          5504 => x"84",
          5505 => x"f0",
          5506 => x"40",
          5507 => x"79",
          5508 => x"75",
          5509 => x"74",
          5510 => x"84",
          5511 => x"85",
          5512 => x"55",
          5513 => x"55",
          5514 => x"70",
          5515 => x"56",
          5516 => x"1a",
          5517 => x"27",
          5518 => x"2e",
          5519 => x"5f",
          5520 => x"22",
          5521 => x"56",
          5522 => x"88",
          5523 => x"b1",
          5524 => x"74",
          5525 => x"1b",
          5526 => x"88",
          5527 => x"9c",
          5528 => x"1a",
          5529 => x"05",
          5530 => x"38",
          5531 => x"18",
          5532 => x"85",
          5533 => x"59",
          5534 => x"77",
          5535 => x"76",
          5536 => x"7c",
          5537 => x"a1",
          5538 => x"38",
          5539 => x"57",
          5540 => x"0b",
          5541 => x"58",
          5542 => x"77",
          5543 => x"56",
          5544 => x"1a",
          5545 => x"31",
          5546 => x"94",
          5547 => x"0c",
          5548 => x"5b",
          5549 => x"75",
          5550 => x"90",
          5551 => x"5b",
          5552 => x"84",
          5553 => x"74",
          5554 => x"04",
          5555 => x"38",
          5556 => x"1b",
          5557 => x"84",
          5558 => x"27",
          5559 => x"16",
          5560 => x"83",
          5561 => x"7f",
          5562 => x"81",
          5563 => x"16",
          5564 => x"ba",
          5565 => x"57",
          5566 => x"83",
          5567 => x"ff",
          5568 => x"59",
          5569 => x"76",
          5570 => x"81",
          5571 => x"ef",
          5572 => x"34",
          5573 => x"08",
          5574 => x"33",
          5575 => x"5c",
          5576 => x"81",
          5577 => x"08",
          5578 => x"17",
          5579 => x"55",
          5580 => x"38",
          5581 => x"09",
          5582 => x"b4",
          5583 => x"7f",
          5584 => x"a9",
          5585 => x"1a",
          5586 => x"93",
          5587 => x"b9",
          5588 => x"1b",
          5589 => x"0c",
          5590 => x"52",
          5591 => x"ba",
          5592 => x"fb",
          5593 => x"ab",
          5594 => x"cc",
          5595 => x"ba",
          5596 => x"81",
          5597 => x"70",
          5598 => x"97",
          5599 => x"b8",
          5600 => x"34",
          5601 => x"58",
          5602 => x"38",
          5603 => x"09",
          5604 => x"b4",
          5605 => x"76",
          5606 => x"f9",
          5607 => x"16",
          5608 => x"ba",
          5609 => x"f2",
          5610 => x"ec",
          5611 => x"b8",
          5612 => x"57",
          5613 => x"08",
          5614 => x"83",
          5615 => x"08",
          5616 => x"fe",
          5617 => x"82",
          5618 => x"81",
          5619 => x"05",
          5620 => x"ff",
          5621 => x"0c",
          5622 => x"39",
          5623 => x"84",
          5624 => x"82",
          5625 => x"ba",
          5626 => x"3d",
          5627 => x"2e",
          5628 => x"2e",
          5629 => x"2e",
          5630 => x"22",
          5631 => x"38",
          5632 => x"81",
          5633 => x"2a",
          5634 => x"81",
          5635 => x"57",
          5636 => x"83",
          5637 => x"81",
          5638 => x"17",
          5639 => x"ba",
          5640 => x"59",
          5641 => x"81",
          5642 => x"33",
          5643 => x"34",
          5644 => x"ff",
          5645 => x"18",
          5646 => x"18",
          5647 => x"5c",
          5648 => x"38",
          5649 => x"74",
          5650 => x"74",
          5651 => x"74",
          5652 => x"80",
          5653 => x"a1",
          5654 => x"99",
          5655 => x"80",
          5656 => x"0b",
          5657 => x"94",
          5658 => x"33",
          5659 => x"19",
          5660 => x"3d",
          5661 => x"53",
          5662 => x"52",
          5663 => x"84",
          5664 => x"ba",
          5665 => x"08",
          5666 => x"08",
          5667 => x"fe",
          5668 => x"82",
          5669 => x"81",
          5670 => x"05",
          5671 => x"ff",
          5672 => x"39",
          5673 => x"34",
          5674 => x"34",
          5675 => x"74",
          5676 => x"74",
          5677 => x"74",
          5678 => x"80",
          5679 => x"a1",
          5680 => x"99",
          5681 => x"80",
          5682 => x"0b",
          5683 => x"c4",
          5684 => x"33",
          5685 => x"19",
          5686 => x"51",
          5687 => x"08",
          5688 => x"74",
          5689 => x"f9",
          5690 => x"fe",
          5691 => x"ba",
          5692 => x"80",
          5693 => x"80",
          5694 => x"80",
          5695 => x"16",
          5696 => x"38",
          5697 => x"84",
          5698 => x"8c",
          5699 => x"33",
          5700 => x"8c",
          5701 => x"73",
          5702 => x"3d",
          5703 => x"75",
          5704 => x"05",
          5705 => x"71",
          5706 => x"71",
          5707 => x"33",
          5708 => x"84",
          5709 => x"8c",
          5710 => x"84",
          5711 => x"78",
          5712 => x"53",
          5713 => x"82",
          5714 => x"59",
          5715 => x"80",
          5716 => x"08",
          5717 => x"58",
          5718 => x"ff",
          5719 => x"26",
          5720 => x"06",
          5721 => x"99",
          5722 => x"ff",
          5723 => x"2a",
          5724 => x"06",
          5725 => x"76",
          5726 => x"2a",
          5727 => x"2e",
          5728 => x"58",
          5729 => x"51",
          5730 => x"38",
          5731 => x"ea",
          5732 => x"05",
          5733 => x"84",
          5734 => x"08",
          5735 => x"8c",
          5736 => x"68",
          5737 => x"94",
          5738 => x"ba",
          5739 => x"d7",
          5740 => x"80",
          5741 => x"05",
          5742 => x"59",
          5743 => x"9b",
          5744 => x"2b",
          5745 => x"58",
          5746 => x"19",
          5747 => x"3d",
          5748 => x"2e",
          5749 => x"0b",
          5750 => x"04",
          5751 => x"98",
          5752 => x"98",
          5753 => x"7e",
          5754 => x"8c",
          5755 => x"3d",
          5756 => x"3d",
          5757 => x"53",
          5758 => x"80",
          5759 => x"ba",
          5760 => x"83",
          5761 => x"7f",
          5762 => x"0c",
          5763 => x"79",
          5764 => x"3d",
          5765 => x"51",
          5766 => x"08",
          5767 => x"38",
          5768 => x"b4",
          5769 => x"ba",
          5770 => x"7d",
          5771 => x"b8",
          5772 => x"8b",
          5773 => x"2e",
          5774 => x"b4",
          5775 => x"df",
          5776 => x"33",
          5777 => x"5d",
          5778 => x"82",
          5779 => x"80",
          5780 => x"84",
          5781 => x"08",
          5782 => x"ff",
          5783 => x"59",
          5784 => x"df",
          5785 => x"33",
          5786 => x"42",
          5787 => x"81",
          5788 => x"84",
          5789 => x"a4",
          5790 => x"84",
          5791 => x"38",
          5792 => x"81",
          5793 => x"05",
          5794 => x"78",
          5795 => x"80",
          5796 => x"17",
          5797 => x"7c",
          5798 => x"26",
          5799 => x"38",
          5800 => x"80",
          5801 => x"19",
          5802 => x"34",
          5803 => x"3d",
          5804 => x"80",
          5805 => x"38",
          5806 => x"0b",
          5807 => x"83",
          5808 => x"43",
          5809 => x"8d",
          5810 => x"57",
          5811 => x"5b",
          5812 => x"76",
          5813 => x"7e",
          5814 => x"81",
          5815 => x"ba",
          5816 => x"ff",
          5817 => x"91",
          5818 => x"8c",
          5819 => x"16",
          5820 => x"71",
          5821 => x"5e",
          5822 => x"17",
          5823 => x"07",
          5824 => x"5d",
          5825 => x"3f",
          5826 => x"8c",
          5827 => x"b1",
          5828 => x"b8",
          5829 => x"5e",
          5830 => x"ba",
          5831 => x"8c",
          5832 => x"a8",
          5833 => x"5a",
          5834 => x"83",
          5835 => x"2e",
          5836 => x"54",
          5837 => x"53",
          5838 => x"88",
          5839 => x"ff",
          5840 => x"58",
          5841 => x"e8",
          5842 => x"05",
          5843 => x"5e",
          5844 => x"fd",
          5845 => x"3d",
          5846 => x"33",
          5847 => x"60",
          5848 => x"08",
          5849 => x"7c",
          5850 => x"26",
          5851 => x"80",
          5852 => x"80",
          5853 => x"7b",
          5854 => x"2e",
          5855 => x"2e",
          5856 => x"2e",
          5857 => x"22",
          5858 => x"38",
          5859 => x"81",
          5860 => x"81",
          5861 => x"76",
          5862 => x"54",
          5863 => x"38",
          5864 => x"52",
          5865 => x"38",
          5866 => x"d3",
          5867 => x"77",
          5868 => x"c3",
          5869 => x"81",
          5870 => x"94",
          5871 => x"08",
          5872 => x"98",
          5873 => x"76",
          5874 => x"17",
          5875 => x"81",
          5876 => x"81",
          5877 => x"99",
          5878 => x"84",
          5879 => x"38",
          5880 => x"27",
          5881 => x"14",
          5882 => x"16",
          5883 => x"16",
          5884 => x"0c",
          5885 => x"70",
          5886 => x"fe",
          5887 => x"57",
          5888 => x"06",
          5889 => x"94",
          5890 => x"38",
          5891 => x"80",
          5892 => x"73",
          5893 => x"8c",
          5894 => x"38",
          5895 => x"ba",
          5896 => x"0b",
          5897 => x"73",
          5898 => x"16",
          5899 => x"fe",
          5900 => x"94",
          5901 => x"83",
          5902 => x"38",
          5903 => x"05",
          5904 => x"f6",
          5905 => x"b0",
          5906 => x"5a",
          5907 => x"38",
          5908 => x"73",
          5909 => x"84",
          5910 => x"81",
          5911 => x"84",
          5912 => x"fc",
          5913 => x"fc",
          5914 => x"97",
          5915 => x"84",
          5916 => x"84",
          5917 => x"38",
          5918 => x"73",
          5919 => x"0b",
          5920 => x"8c",
          5921 => x"0d",
          5922 => x"a2",
          5923 => x"52",
          5924 => x"3f",
          5925 => x"8c",
          5926 => x"0c",
          5927 => x"8c",
          5928 => x"52",
          5929 => x"ba",
          5930 => x"80",
          5931 => x"2b",
          5932 => x"86",
          5933 => x"5b",
          5934 => x"9c",
          5935 => x"33",
          5936 => x"5d",
          5937 => x"b3",
          5938 => x"86",
          5939 => x"75",
          5940 => x"8c",
          5941 => x"74",
          5942 => x"0c",
          5943 => x"0c",
          5944 => x"18",
          5945 => x"07",
          5946 => x"ff",
          5947 => x"89",
          5948 => x"08",
          5949 => x"33",
          5950 => x"13",
          5951 => x"76",
          5952 => x"73",
          5953 => x"ba",
          5954 => x"13",
          5955 => x"ba",
          5956 => x"38",
          5957 => x"f8",
          5958 => x"56",
          5959 => x"54",
          5960 => x"53",
          5961 => x"22",
          5962 => x"2e",
          5963 => x"75",
          5964 => x"2e",
          5965 => x"ff",
          5966 => x"53",
          5967 => x"38",
          5968 => x"52",
          5969 => x"52",
          5970 => x"ba",
          5971 => x"72",
          5972 => x"06",
          5973 => x"0c",
          5974 => x"75",
          5975 => x"52",
          5976 => x"ba",
          5977 => x"72",
          5978 => x"06",
          5979 => x"74",
          5980 => x"8c",
          5981 => x"0d",
          5982 => x"e8",
          5983 => x"53",
          5984 => x"54",
          5985 => x"66",
          5986 => x"97",
          5987 => x"ba",
          5988 => x"80",
          5989 => x"0c",
          5990 => x"51",
          5991 => x"08",
          5992 => x"02",
          5993 => x"55",
          5994 => x"80",
          5995 => x"ff",
          5996 => x"0c",
          5997 => x"ba",
          5998 => x"3d",
          5999 => x"95",
          6000 => x"c0",
          6001 => x"84",
          6002 => x"0c",
          6003 => x"94",
          6004 => x"75",
          6005 => x"84",
          6006 => x"84",
          6007 => x"78",
          6008 => x"18",
          6009 => x"59",
          6010 => x"71",
          6011 => x"2e",
          6012 => x"5f",
          6013 => x"75",
          6014 => x"51",
          6015 => x"08",
          6016 => x"5e",
          6017 => x"57",
          6018 => x"7d",
          6019 => x"b8",
          6020 => x"71",
          6021 => x"14",
          6022 => x"33",
          6023 => x"07",
          6024 => x"60",
          6025 => x"05",
          6026 => x"58",
          6027 => x"7a",
          6028 => x"17",
          6029 => x"34",
          6030 => x"0d",
          6031 => x"b8",
          6032 => x"5d",
          6033 => x"ba",
          6034 => x"8c",
          6035 => x"a8",
          6036 => x"5f",
          6037 => x"bd",
          6038 => x"2e",
          6039 => x"54",
          6040 => x"53",
          6041 => x"fb",
          6042 => x"82",
          6043 => x"52",
          6044 => x"ba",
          6045 => x"84",
          6046 => x"38",
          6047 => x"ba",
          6048 => x"81",
          6049 => x"17",
          6050 => x"0c",
          6051 => x"81",
          6052 => x"c8",
          6053 => x"33",
          6054 => x"30",
          6055 => x"ff",
          6056 => x"5f",
          6057 => x"8f",
          6058 => x"60",
          6059 => x"18",
          6060 => x"77",
          6061 => x"60",
          6062 => x"7b",
          6063 => x"38",
          6064 => x"38",
          6065 => x"38",
          6066 => x"59",
          6067 => x"54",
          6068 => x"17",
          6069 => x"17",
          6070 => x"58",
          6071 => x"38",
          6072 => x"08",
          6073 => x"88",
          6074 => x"74",
          6075 => x"26",
          6076 => x"18",
          6077 => x"77",
          6078 => x"34",
          6079 => x"18",
          6080 => x"0c",
          6081 => x"78",
          6082 => x"51",
          6083 => x"08",
          6084 => x"80",
          6085 => x"2e",
          6086 => x"ff",
          6087 => x"52",
          6088 => x"ba",
          6089 => x"08",
          6090 => x"58",
          6091 => x"15",
          6092 => x"07",
          6093 => x"77",
          6094 => x"81",
          6095 => x"84",
          6096 => x"fe",
          6097 => x"fe",
          6098 => x"59",
          6099 => x"0c",
          6100 => x"76",
          6101 => x"8c",
          6102 => x"ba",
          6103 => x"75",
          6104 => x"8c",
          6105 => x"38",
          6106 => x"78",
          6107 => x"ba",
          6108 => x"ba",
          6109 => x"96",
          6110 => x"53",
          6111 => x"3f",
          6112 => x"8c",
          6113 => x"51",
          6114 => x"08",
          6115 => x"80",
          6116 => x"2e",
          6117 => x"ff",
          6118 => x"52",
          6119 => x"ba",
          6120 => x"08",
          6121 => x"58",
          6122 => x"94",
          6123 => x"54",
          6124 => x"79",
          6125 => x"56",
          6126 => x"81",
          6127 => x"18",
          6128 => x"56",
          6129 => x"59",
          6130 => x"08",
          6131 => x"39",
          6132 => x"fd",
          6133 => x"c0",
          6134 => x"3d",
          6135 => x"05",
          6136 => x"3f",
          6137 => x"8c",
          6138 => x"ba",
          6139 => x"4b",
          6140 => x"52",
          6141 => x"8c",
          6142 => x"38",
          6143 => x"2a",
          6144 => x"cd",
          6145 => x"24",
          6146 => x"70",
          6147 => x"ff",
          6148 => x"11",
          6149 => x"07",
          6150 => x"7c",
          6151 => x"2a",
          6152 => x"ed",
          6153 => x"2e",
          6154 => x"84",
          6155 => x"52",
          6156 => x"8c",
          6157 => x"e5",
          6158 => x"51",
          6159 => x"08",
          6160 => x"87",
          6161 => x"0d",
          6162 => x"71",
          6163 => x"07",
          6164 => x"ba",
          6165 => x"ba",
          6166 => x"6f",
          6167 => x"ff",
          6168 => x"51",
          6169 => x"08",
          6170 => x"be",
          6171 => x"25",
          6172 => x"74",
          6173 => x"58",
          6174 => x"17",
          6175 => x"56",
          6176 => x"f5",
          6177 => x"ba",
          6178 => x"17",
          6179 => x"b4",
          6180 => x"83",
          6181 => x"2e",
          6182 => x"54",
          6183 => x"33",
          6184 => x"8c",
          6185 => x"81",
          6186 => x"77",
          6187 => x"78",
          6188 => x"19",
          6189 => x"52",
          6190 => x"ba",
          6191 => x"80",
          6192 => x"09",
          6193 => x"fe",
          6194 => x"53",
          6195 => x"f2",
          6196 => x"08",
          6197 => x"38",
          6198 => x"b4",
          6199 => x"ba",
          6200 => x"08",
          6201 => x"55",
          6202 => x"de",
          6203 => x"18",
          6204 => x"33",
          6205 => x"fe",
          6206 => x"80",
          6207 => x"f6",
          6208 => x"84",
          6209 => x"38",
          6210 => x"e6",
          6211 => x"80",
          6212 => x"51",
          6213 => x"08",
          6214 => x"94",
          6215 => x"27",
          6216 => x"0c",
          6217 => x"84",
          6218 => x"ff",
          6219 => x"79",
          6220 => x"08",
          6221 => x"90",
          6222 => x"3d",
          6223 => x"ff",
          6224 => x"56",
          6225 => x"38",
          6226 => x"0d",
          6227 => x"70",
          6228 => x"ba",
          6229 => x"8b",
          6230 => x"9f",
          6231 => x"84",
          6232 => x"80",
          6233 => x"06",
          6234 => x"38",
          6235 => x"52",
          6236 => x"8c",
          6237 => x"08",
          6238 => x"08",
          6239 => x"8c",
          6240 => x"81",
          6241 => x"83",
          6242 => x"e2",
          6243 => x"05",
          6244 => x"8d",
          6245 => x"b0",
          6246 => x"18",
          6247 => x"57",
          6248 => x"34",
          6249 => x"58",
          6250 => x"81",
          6251 => x"78",
          6252 => x"c9",
          6253 => x"38",
          6254 => x"ff",
          6255 => x"53",
          6256 => x"52",
          6257 => x"84",
          6258 => x"8c",
          6259 => x"a8",
          6260 => x"08",
          6261 => x"5b",
          6262 => x"e1",
          6263 => x"18",
          6264 => x"33",
          6265 => x"39",
          6266 => x"81",
          6267 => x"18",
          6268 => x"7c",
          6269 => x"8c",
          6270 => x"2e",
          6271 => x"81",
          6272 => x"08",
          6273 => x"74",
          6274 => x"84",
          6275 => x"17",
          6276 => x"5c",
          6277 => x"18",
          6278 => x"07",
          6279 => x"78",
          6280 => x"ba",
          6281 => x"17",
          6282 => x"57",
          6283 => x"06",
          6284 => x"56",
          6285 => x"34",
          6286 => x"57",
          6287 => x"90",
          6288 => x"75",
          6289 => x"1a",
          6290 => x"80",
          6291 => x"7c",
          6292 => x"80",
          6293 => x"7a",
          6294 => x"74",
          6295 => x"a0",
          6296 => x"58",
          6297 => x"77",
          6298 => x"56",
          6299 => x"80",
          6300 => x"ff",
          6301 => x"f2",
          6302 => x"80",
          6303 => x"83",
          6304 => x"0b",
          6305 => x"96",
          6306 => x"ba",
          6307 => x"84",
          6308 => x"ba",
          6309 => x"98",
          6310 => x"34",
          6311 => x"34",
          6312 => x"34",
          6313 => x"d9",
          6314 => x"34",
          6315 => x"7d",
          6316 => x"8c",
          6317 => x"9f",
          6318 => x"74",
          6319 => x"57",
          6320 => x"39",
          6321 => x"17",
          6322 => x"cd",
          6323 => x"d8",
          6324 => x"a1",
          6325 => x"18",
          6326 => x"18",
          6327 => x"34",
          6328 => x"7d",
          6329 => x"8c",
          6330 => x"0d",
          6331 => x"5b",
          6332 => x"70",
          6333 => x"56",
          6334 => x"74",
          6335 => x"38",
          6336 => x"52",
          6337 => x"84",
          6338 => x"08",
          6339 => x"8c",
          6340 => x"3d",
          6341 => x"70",
          6342 => x"ba",
          6343 => x"dc",
          6344 => x"a0",
          6345 => x"a0",
          6346 => x"58",
          6347 => x"77",
          6348 => x"55",
          6349 => x"78",
          6350 => x"05",
          6351 => x"34",
          6352 => x"3d",
          6353 => x"3f",
          6354 => x"8c",
          6355 => x"08",
          6356 => x"ba",
          6357 => x"33",
          6358 => x"57",
          6359 => x"17",
          6360 => x"59",
          6361 => x"7f",
          6362 => x"5d",
          6363 => x"05",
          6364 => x"33",
          6365 => x"99",
          6366 => x"ff",
          6367 => x"77",
          6368 => x"81",
          6369 => x"9f",
          6370 => x"81",
          6371 => x"78",
          6372 => x"9f",
          6373 => x"80",
          6374 => x"5e",
          6375 => x"7c",
          6376 => x"7b",
          6377 => x"0c",
          6378 => x"52",
          6379 => x"84",
          6380 => x"08",
          6381 => x"aa",
          6382 => x"ac",
          6383 => x"84",
          6384 => x"08",
          6385 => x"8d",
          6386 => x"58",
          6387 => x"33",
          6388 => x"1a",
          6389 => x"05",
          6390 => x"70",
          6391 => x"89",
          6392 => x"19",
          6393 => x"34",
          6394 => x"06",
          6395 => x"38",
          6396 => x"38",
          6397 => x"71",
          6398 => x"5c",
          6399 => x"fe",
          6400 => x"56",
          6401 => x"17",
          6402 => x"05",
          6403 => x"38",
          6404 => x"76",
          6405 => x"7e",
          6406 => x"b8",
          6407 => x"e3",
          6408 => x"2e",
          6409 => x"b4",
          6410 => x"18",
          6411 => x"15",
          6412 => x"06",
          6413 => x"06",
          6414 => x"7b",
          6415 => x"34",
          6416 => x"81",
          6417 => x"7d",
          6418 => x"56",
          6419 => x"81",
          6420 => x"3d",
          6421 => x"74",
          6422 => x"51",
          6423 => x"08",
          6424 => x"38",
          6425 => x"80",
          6426 => x"38",
          6427 => x"7a",
          6428 => x"81",
          6429 => x"16",
          6430 => x"ba",
          6431 => x"57",
          6432 => x"55",
          6433 => x"e5",
          6434 => x"90",
          6435 => x"52",
          6436 => x"ba",
          6437 => x"80",
          6438 => x"84",
          6439 => x"f9",
          6440 => x"3f",
          6441 => x"0c",
          6442 => x"ba",
          6443 => x"18",
          6444 => x"71",
          6445 => x"5c",
          6446 => x"84",
          6447 => x"08",
          6448 => x"ba",
          6449 => x"54",
          6450 => x"16",
          6451 => x"58",
          6452 => x"81",
          6453 => x"08",
          6454 => x"17",
          6455 => x"55",
          6456 => x"38",
          6457 => x"09",
          6458 => x"b4",
          6459 => x"7b",
          6460 => x"c9",
          6461 => x"54",
          6462 => x"53",
          6463 => x"b1",
          6464 => x"fc",
          6465 => x"18",
          6466 => x"31",
          6467 => x"a0",
          6468 => x"17",
          6469 => x"06",
          6470 => x"08",
          6471 => x"81",
          6472 => x"79",
          6473 => x"02",
          6474 => x"80",
          6475 => x"96",
          6476 => x"ff",
          6477 => x"56",
          6478 => x"38",
          6479 => x"0d",
          6480 => x"d0",
          6481 => x"ba",
          6482 => x"e0",
          6483 => x"a0",
          6484 => x"74",
          6485 => x"33",
          6486 => x"56",
          6487 => x"55",
          6488 => x"fe",
          6489 => x"84",
          6490 => x"ec",
          6491 => x"3d",
          6492 => x"a1",
          6493 => x"84",
          6494 => x"74",
          6495 => x"04",
          6496 => x"05",
          6497 => x"8c",
          6498 => x"38",
          6499 => x"06",
          6500 => x"84",
          6501 => x"2b",
          6502 => x"34",
          6503 => x"34",
          6504 => x"34",
          6505 => x"34",
          6506 => x"78",
          6507 => x"8c",
          6508 => x"0d",
          6509 => x"5b",
          6510 => x"9b",
          6511 => x"ba",
          6512 => x"70",
          6513 => x"51",
          6514 => x"81",
          6515 => x"a4",
          6516 => x"25",
          6517 => x"38",
          6518 => x"80",
          6519 => x"08",
          6520 => x"77",
          6521 => x"7a",
          6522 => x"06",
          6523 => x"b8",
          6524 => x"dc",
          6525 => x"2e",
          6526 => x"b4",
          6527 => x"7c",
          6528 => x"74",
          6529 => x"74",
          6530 => x"18",
          6531 => x"33",
          6532 => x"81",
          6533 => x"75",
          6534 => x"5e",
          6535 => x"0c",
          6536 => x"40",
          6537 => x"fe",
          6538 => x"57",
          6539 => x"8d",
          6540 => x"fe",
          6541 => x"fe",
          6542 => x"53",
          6543 => x"52",
          6544 => x"84",
          6545 => x"06",
          6546 => x"83",
          6547 => x"08",
          6548 => x"74",
          6549 => x"82",
          6550 => x"81",
          6551 => x"16",
          6552 => x"52",
          6553 => x"3f",
          6554 => x"16",
          6555 => x"d2",
          6556 => x"fe",
          6557 => x"74",
          6558 => x"8c",
          6559 => x"e1",
          6560 => x"8c",
          6561 => x"81",
          6562 => x"33",
          6563 => x"27",
          6564 => x"80",
          6565 => x"38",
          6566 => x"57",
          6567 => x"e1",
          6568 => x"3d",
          6569 => x"05",
          6570 => x"3f",
          6571 => x"8c",
          6572 => x"8b",
          6573 => x"05",
          6574 => x"38",
          6575 => x"81",
          6576 => x"78",
          6577 => x"3d",
          6578 => x"18",
          6579 => x"7c",
          6580 => x"ff",
          6581 => x"b5",
          6582 => x"dc",
          6583 => x"ff",
          6584 => x"38",
          6585 => x"33",
          6586 => x"78",
          6587 => x"78",
          6588 => x"33",
          6589 => x"74",
          6590 => x"09",
          6591 => x"06",
          6592 => x"77",
          6593 => x"81",
          6594 => x"38",
          6595 => x"81",
          6596 => x"7b",
          6597 => x"a3",
          6598 => x"06",
          6599 => x"fe",
          6600 => x"56",
          6601 => x"80",
          6602 => x"79",
          6603 => x"2e",
          6604 => x"5a",
          6605 => x"80",
          6606 => x"ef",
          6607 => x"84",
          6608 => x"74",
          6609 => x"3d",
          6610 => x"9e",
          6611 => x"ff",
          6612 => x"86",
          6613 => x"3d",
          6614 => x"fe",
          6615 => x"f4",
          6616 => x"84",
          6617 => x"80",
          6618 => x"59",
          6619 => x"33",
          6620 => x"15",
          6621 => x"0b",
          6622 => x"ec",
          6623 => x"56",
          6624 => x"8a",
          6625 => x"ba",
          6626 => x"fe",
          6627 => x"fe",
          6628 => x"52",
          6629 => x"8c",
          6630 => x"2e",
          6631 => x"ba",
          6632 => x"16",
          6633 => x"77",
          6634 => x"74",
          6635 => x"38",
          6636 => x"81",
          6637 => x"84",
          6638 => x"ff",
          6639 => x"78",
          6640 => x"08",
          6641 => x"e5",
          6642 => x"80",
          6643 => x"2e",
          6644 => x"81",
          6645 => x"fe",
          6646 => x"57",
          6647 => x"86",
          6648 => x"bf",
          6649 => x"a0",
          6650 => x"05",
          6651 => x"38",
          6652 => x"8b",
          6653 => x"81",
          6654 => x"58",
          6655 => x"fd",
          6656 => x"33",
          6657 => x"15",
          6658 => x"6b",
          6659 => x"0b",
          6660 => x"bc",
          6661 => x"ce",
          6662 => x"54",
          6663 => x"18",
          6664 => x"ba",
          6665 => x"80",
          6666 => x"19",
          6667 => x"31",
          6668 => x"38",
          6669 => x"b1",
          6670 => x"e8",
          6671 => x"fe",
          6672 => x"57",
          6673 => x"b6",
          6674 => x"59",
          6675 => x"a1",
          6676 => x"19",
          6677 => x"33",
          6678 => x"39",
          6679 => x"05",
          6680 => x"89",
          6681 => x"08",
          6682 => x"33",
          6683 => x"15",
          6684 => x"78",
          6685 => x"5f",
          6686 => x"56",
          6687 => x"81",
          6688 => x"38",
          6689 => x"06",
          6690 => x"38",
          6691 => x"70",
          6692 => x"87",
          6693 => x"30",
          6694 => x"8c",
          6695 => x"53",
          6696 => x"38",
          6697 => x"82",
          6698 => x"74",
          6699 => x"81",
          6700 => x"75",
          6701 => x"8c",
          6702 => x"ba",
          6703 => x"84",
          6704 => x"19",
          6705 => x"78",
          6706 => x"56",
          6707 => x"90",
          6708 => x"8c",
          6709 => x"33",
          6710 => x"8c",
          6711 => x"38",
          6712 => x"39",
          6713 => x"7d",
          6714 => x"81",
          6715 => x"38",
          6716 => x"dd",
          6717 => x"84",
          6718 => x"81",
          6719 => x"d7",
          6720 => x"7b",
          6721 => x"18",
          6722 => x"33",
          6723 => x"34",
          6724 => x"08",
          6725 => x"38",
          6726 => x"15",
          6727 => x"34",
          6728 => x"ff",
          6729 => x"be",
          6730 => x"54",
          6731 => x"a1",
          6732 => x"0d",
          6733 => x"88",
          6734 => x"5f",
          6735 => x"5b",
          6736 => x"79",
          6737 => x"26",
          6738 => x"38",
          6739 => x"92",
          6740 => x"76",
          6741 => x"84",
          6742 => x"74",
          6743 => x"75",
          6744 => x"ba",
          6745 => x"52",
          6746 => x"ba",
          6747 => x"06",
          6748 => x"38",
          6749 => x"57",
          6750 => x"05",
          6751 => x"b0",
          6752 => x"38",
          6753 => x"38",
          6754 => x"38",
          6755 => x"ff",
          6756 => x"80",
          6757 => x"80",
          6758 => x"7f",
          6759 => x"89",
          6760 => x"89",
          6761 => x"80",
          6762 => x"80",
          6763 => x"74",
          6764 => x"df",
          6765 => x"79",
          6766 => x"84",
          6767 => x"83",
          6768 => x"33",
          6769 => x"57",
          6770 => x"06",
          6771 => x"05",
          6772 => x"80",
          6773 => x"83",
          6774 => x"2b",
          6775 => x"70",
          6776 => x"07",
          6777 => x"12",
          6778 => x"07",
          6779 => x"2b",
          6780 => x"0c",
          6781 => x"44",
          6782 => x"4b",
          6783 => x"27",
          6784 => x"80",
          6785 => x"70",
          6786 => x"83",
          6787 => x"82",
          6788 => x"66",
          6789 => x"4a",
          6790 => x"8a",
          6791 => x"2a",
          6792 => x"56",
          6793 => x"77",
          6794 => x"77",
          6795 => x"58",
          6796 => x"27",
          6797 => x"80",
          6798 => x"84",
          6799 => x"f5",
          6800 => x"8c",
          6801 => x"71",
          6802 => x"43",
          6803 => x"5c",
          6804 => x"05",
          6805 => x"72",
          6806 => x"2e",
          6807 => x"90",
          6808 => x"74",
          6809 => x"31",
          6810 => x"52",
          6811 => x"8c",
          6812 => x"38",
          6813 => x"dd",
          6814 => x"8c",
          6815 => x"f9",
          6816 => x"26",
          6817 => x"39",
          6818 => x"9f",
          6819 => x"81",
          6820 => x"ba",
          6821 => x"98",
          6822 => x"81",
          6823 => x"26",
          6824 => x"06",
          6825 => x"81",
          6826 => x"5f",
          6827 => x"70",
          6828 => x"05",
          6829 => x"57",
          6830 => x"70",
          6831 => x"18",
          6832 => x"18",
          6833 => x"30",
          6834 => x"2e",
          6835 => x"be",
          6836 => x"72",
          6837 => x"4a",
          6838 => x"1c",
          6839 => x"ff",
          6840 => x"9f",
          6841 => x"51",
          6842 => x"ba",
          6843 => x"2a",
          6844 => x"56",
          6845 => x"8e",
          6846 => x"74",
          6847 => x"56",
          6848 => x"ba",
          6849 => x"f9",
          6850 => x"57",
          6851 => x"6e",
          6852 => x"39",
          6853 => x"9d",
          6854 => x"81",
          6855 => x"57",
          6856 => x"0d",
          6857 => x"62",
          6858 => x"60",
          6859 => x"8e",
          6860 => x"61",
          6861 => x"58",
          6862 => x"8b",
          6863 => x"76",
          6864 => x"81",
          6865 => x"ef",
          6866 => x"34",
          6867 => x"8d",
          6868 => x"4b",
          6869 => x"2a",
          6870 => x"61",
          6871 => x"30",
          6872 => x"78",
          6873 => x"92",
          6874 => x"ff",
          6875 => x"ff",
          6876 => x"74",
          6877 => x"34",
          6878 => x"98",
          6879 => x"ff",
          6880 => x"05",
          6881 => x"88",
          6882 => x"7e",
          6883 => x"34",
          6884 => x"84",
          6885 => x"62",
          6886 => x"a7",
          6887 => x"a1",
          6888 => x"aa",
          6889 => x"55",
          6890 => x"2a",
          6891 => x"80",
          6892 => x"05",
          6893 => x"d4",
          6894 => x"58",
          6895 => x"ff",
          6896 => x"fe",
          6897 => x"83",
          6898 => x"81",
          6899 => x"fe",
          6900 => x"8c",
          6901 => x"62",
          6902 => x"57",
          6903 => x"34",
          6904 => x"75",
          6905 => x"38",
          6906 => x"2e",
          6907 => x"76",
          6908 => x"70",
          6909 => x"59",
          6910 => x"76",
          6911 => x"57",
          6912 => x"76",
          6913 => x"79",
          6914 => x"8c",
          6915 => x"57",
          6916 => x"34",
          6917 => x"1b",
          6918 => x"38",
          6919 => x"ff",
          6920 => x"83",
          6921 => x"26",
          6922 => x"53",
          6923 => x"3f",
          6924 => x"74",
          6925 => x"db",
          6926 => x"38",
          6927 => x"8a",
          6928 => x"38",
          6929 => x"83",
          6930 => x"38",
          6931 => x"70",
          6932 => x"78",
          6933 => x"aa",
          6934 => x"78",
          6935 => x"81",
          6936 => x"05",
          6937 => x"43",
          6938 => x"fc",
          6939 => x"34",
          6940 => x"07",
          6941 => x"ba",
          6942 => x"61",
          6943 => x"c7",
          6944 => x"34",
          6945 => x"05",
          6946 => x"62",
          6947 => x"05",
          6948 => x"83",
          6949 => x"7e",
          6950 => x"78",
          6951 => x"f1",
          6952 => x"f7",
          6953 => x"51",
          6954 => x"ba",
          6955 => x"8c",
          6956 => x"0d",
          6957 => x"f9",
          6958 => x"5c",
          6959 => x"91",
          6960 => x"22",
          6961 => x"74",
          6962 => x"56",
          6963 => x"57",
          6964 => x"75",
          6965 => x"fc",
          6966 => x"10",
          6967 => x"5e",
          6968 => x"8c",
          6969 => x"fd",
          6970 => x"38",
          6971 => x"8c",
          6972 => x"38",
          6973 => x"5b",
          6974 => x"c8",
          6975 => x"2e",
          6976 => x"39",
          6977 => x"2a",
          6978 => x"90",
          6979 => x"75",
          6980 => x"34",
          6981 => x"05",
          6982 => x"a1",
          6983 => x"61",
          6984 => x"05",
          6985 => x"a5",
          6986 => x"61",
          6987 => x"75",
          6988 => x"05",
          6989 => x"61",
          6990 => x"34",
          6991 => x"b1",
          6992 => x"80",
          6993 => x"80",
          6994 => x"05",
          6995 => x"e5",
          6996 => x"05",
          6997 => x"34",
          6998 => x"cd",
          6999 => x"76",
          7000 => x"55",
          7001 => x"54",
          7002 => x"be",
          7003 => x"08",
          7004 => x"05",
          7005 => x"76",
          7006 => x"52",
          7007 => x"c3",
          7008 => x"9f",
          7009 => x"f8",
          7010 => x"81",
          7011 => x"05",
          7012 => x"84",
          7013 => x"ff",
          7014 => x"05",
          7015 => x"61",
          7016 => x"34",
          7017 => x"39",
          7018 => x"79",
          7019 => x"61",
          7020 => x"57",
          7021 => x"60",
          7022 => x"5e",
          7023 => x"81",
          7024 => x"81",
          7025 => x"80",
          7026 => x"f2",
          7027 => x"61",
          7028 => x"83",
          7029 => x"7a",
          7030 => x"2a",
          7031 => x"7a",
          7032 => x"05",
          7033 => x"83",
          7034 => x"05",
          7035 => x"76",
          7036 => x"83",
          7037 => x"ff",
          7038 => x"53",
          7039 => x"3f",
          7040 => x"79",
          7041 => x"57",
          7042 => x"7e",
          7043 => x"05",
          7044 => x"38",
          7045 => x"54",
          7046 => x"9a",
          7047 => x"06",
          7048 => x"8d",
          7049 => x"05",
          7050 => x"2e",
          7051 => x"80",
          7052 => x"76",
          7053 => x"3d",
          7054 => x"84",
          7055 => x"8a",
          7056 => x"56",
          7057 => x"08",
          7058 => x"75",
          7059 => x"8e",
          7060 => x"88",
          7061 => x"3d",
          7062 => x"52",
          7063 => x"74",
          7064 => x"9f",
          7065 => x"1c",
          7066 => x"39",
          7067 => x"ff",
          7068 => x"ff",
          7069 => x"cc",
          7070 => x"05",
          7071 => x"38",
          7072 => x"2e",
          7073 => x"24",
          7074 => x"05",
          7075 => x"55",
          7076 => x"18",
          7077 => x"55",
          7078 => x"ff",
          7079 => x"52",
          7080 => x"84",
          7081 => x"2e",
          7082 => x"0c",
          7083 => x"b0",
          7084 => x"76",
          7085 => x"7b",
          7086 => x"2a",
          7087 => x"a5",
          7088 => x"3f",
          7089 => x"0c",
          7090 => x"75",
          7091 => x"53",
          7092 => x"38",
          7093 => x"84",
          7094 => x"83",
          7095 => x"b5",
          7096 => x"80",
          7097 => x"51",
          7098 => x"70",
          7099 => x"80",
          7100 => x"e7",
          7101 => x"39",
          7102 => x"84",
          7103 => x"04",
          7104 => x"02",
          7105 => x"80",
          7106 => x"70",
          7107 => x"3d",
          7108 => x"81",
          7109 => x"e9",
          7110 => x"70",
          7111 => x"3d",
          7112 => x"70",
          7113 => x"70",
          7114 => x"56",
          7115 => x"38",
          7116 => x"71",
          7117 => x"07",
          7118 => x"71",
          7119 => x"88",
          7120 => x"14",
          7121 => x"71",
          7122 => x"82",
          7123 => x"80",
          7124 => x"52",
          7125 => x"70",
          7126 => x"04",
          7127 => x"71",
          7128 => x"83",
          7129 => x"c7",
          7130 => x"57",
          7131 => x"16",
          7132 => x"f1",
          7133 => x"06",
          7134 => x"83",
          7135 => x"d0",
          7136 => x"51",
          7137 => x"ff",
          7138 => x"70",
          7139 => x"b9",
          7140 => x"71",
          7141 => x"52",
          7142 => x"10",
          7143 => x"ef",
          7144 => x"00",
          7145 => x"ff",
          7146 => x"00",
          7147 => x"00",
          7148 => x"00",
          7149 => x"00",
          7150 => x"00",
          7151 => x"00",
          7152 => x"00",
          7153 => x"00",
          7154 => x"00",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"00",
          7372 => x"00",
          7373 => x"00",
          7374 => x"00",
          7375 => x"00",
          7376 => x"00",
          7377 => x"00",
          7378 => x"00",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"69",
          7383 => x"69",
          7384 => x"69",
          7385 => x"6c",
          7386 => x"65",
          7387 => x"63",
          7388 => x"63",
          7389 => x"64",
          7390 => x"64",
          7391 => x"65",
          7392 => x"65",
          7393 => x"69",
          7394 => x"66",
          7395 => x"00",
          7396 => x"65",
          7397 => x"65",
          7398 => x"6e",
          7399 => x"65",
          7400 => x"6c",
          7401 => x"62",
          7402 => x"62",
          7403 => x"69",
          7404 => x"64",
          7405 => x"77",
          7406 => x"2e",
          7407 => x"65",
          7408 => x"63",
          7409 => x"00",
          7410 => x"61",
          7411 => x"20",
          7412 => x"00",
          7413 => x"66",
          7414 => x"6d",
          7415 => x"00",
          7416 => x"69",
          7417 => x"64",
          7418 => x"75",
          7419 => x"61",
          7420 => x"6e",
          7421 => x"00",
          7422 => x"74",
          7423 => x"64",
          7424 => x"6d",
          7425 => x"20",
          7426 => x"74",
          7427 => x"64",
          7428 => x"6b",
          7429 => x"6e",
          7430 => x"6c",
          7431 => x"72",
          7432 => x"62",
          7433 => x"6e",
          7434 => x"00",
          7435 => x"20",
          7436 => x"72",
          7437 => x"2e",
          7438 => x"68",
          7439 => x"6e",
          7440 => x"00",
          7441 => x"61",
          7442 => x"65",
          7443 => x"00",
          7444 => x"73",
          7445 => x"2e",
          7446 => x"69",
          7447 => x"61",
          7448 => x"6f",
          7449 => x"6f",
          7450 => x"6f",
          7451 => x"6f",
          7452 => x"69",
          7453 => x"72",
          7454 => x"6e",
          7455 => x"65",
          7456 => x"69",
          7457 => x"72",
          7458 => x"73",
          7459 => x"25",
          7460 => x"73",
          7461 => x"25",
          7462 => x"73",
          7463 => x"00",
          7464 => x"00",
          7465 => x"00",
          7466 => x"30",
          7467 => x"7c",
          7468 => x"20",
          7469 => x"00",
          7470 => x"20",
          7471 => x"4f",
          7472 => x"20",
          7473 => x"2f",
          7474 => x"31",
          7475 => x"5a",
          7476 => x"20",
          7477 => x"73",
          7478 => x"0a",
          7479 => x"6e",
          7480 => x"20",
          7481 => x"00",
          7482 => x"20",
          7483 => x"72",
          7484 => x"41",
          7485 => x"69",
          7486 => x"74",
          7487 => x"20",
          7488 => x"72",
          7489 => x"41",
          7490 => x"69",
          7491 => x"74",
          7492 => x"20",
          7493 => x"72",
          7494 => x"4f",
          7495 => x"69",
          7496 => x"74",
          7497 => x"6e",
          7498 => x"00",
          7499 => x"20",
          7500 => x"70",
          7501 => x"6e",
          7502 => x"6d",
          7503 => x"6e",
          7504 => x"74",
          7505 => x"00",
          7506 => x"78",
          7507 => x"00",
          7508 => x"70",
          7509 => x"61",
          7510 => x"20",
          7511 => x"69",
          7512 => x"61",
          7513 => x"6c",
          7514 => x"69",
          7515 => x"6c",
          7516 => x"20",
          7517 => x"73",
          7518 => x"69",
          7519 => x"73",
          7520 => x"3a",
          7521 => x"6f",
          7522 => x"00",
          7523 => x"69",
          7524 => x"73",
          7525 => x"00",
          7526 => x"72",
          7527 => x"67",
          7528 => x"65",
          7529 => x"67",
          7530 => x"61",
          7531 => x"00",
          7532 => x"6e",
          7533 => x"40",
          7534 => x"2e",
          7535 => x"61",
          7536 => x"72",
          7537 => x"65",
          7538 => x"00",
          7539 => x"74",
          7540 => x"65",
          7541 => x"78",
          7542 => x"30",
          7543 => x"6c",
          7544 => x"30",
          7545 => x"58",
          7546 => x"72",
          7547 => x"00",
          7548 => x"28",
          7549 => x"25",
          7550 => x"38",
          7551 => x"6f",
          7552 => x"2e",
          7553 => x"20",
          7554 => x"6c",
          7555 => x"2e",
          7556 => x"75",
          7557 => x"72",
          7558 => x"6c",
          7559 => x"64",
          7560 => x"00",
          7561 => x"79",
          7562 => x"74",
          7563 => x"6e",
          7564 => x"65",
          7565 => x"61",
          7566 => x"3f",
          7567 => x"2f",
          7568 => x"64",
          7569 => x"64",
          7570 => x"6f",
          7571 => x"74",
          7572 => x"0a",
          7573 => x"20",
          7574 => x"6e",
          7575 => x"64",
          7576 => x"3a",
          7577 => x"50",
          7578 => x"20",
          7579 => x"41",
          7580 => x"3d",
          7581 => x"00",
          7582 => x"50",
          7583 => x"79",
          7584 => x"41",
          7585 => x"3d",
          7586 => x"00",
          7587 => x"74",
          7588 => x"72",
          7589 => x"73",
          7590 => x"3d",
          7591 => x"00",
          7592 => x"00",
          7593 => x"50",
          7594 => x"20",
          7595 => x"20",
          7596 => x"3d",
          7597 => x"00",
          7598 => x"79",
          7599 => x"6f",
          7600 => x"20",
          7601 => x"3d",
          7602 => x"64",
          7603 => x"20",
          7604 => x"6f",
          7605 => x"4d",
          7606 => x"46",
          7607 => x"2e",
          7608 => x"0a",
          7609 => x"44",
          7610 => x"63",
          7611 => x"20",
          7612 => x"3d",
          7613 => x"64",
          7614 => x"20",
          7615 => x"20",
          7616 => x"20",
          7617 => x"00",
          7618 => x"42",
          7619 => x"20",
          7620 => x"4f",
          7621 => x"00",
          7622 => x"4e",
          7623 => x"20",
          7624 => x"6c",
          7625 => x"2e",
          7626 => x"49",
          7627 => x"20",
          7628 => x"20",
          7629 => x"2e",
          7630 => x"44",
          7631 => x"20",
          7632 => x"73",
          7633 => x"2e",
          7634 => x"41",
          7635 => x"20",
          7636 => x"30",
          7637 => x"20",
          7638 => x"20",
          7639 => x"38",
          7640 => x"2e",
          7641 => x"4e",
          7642 => x"20",
          7643 => x"30",
          7644 => x"20",
          7645 => x"20",
          7646 => x"38",
          7647 => x"2e",
          7648 => x"42",
          7649 => x"20",
          7650 => x"30",
          7651 => x"28",
          7652 => x"43",
          7653 => x"29",
          7654 => x"77",
          7655 => x"00",
          7656 => x"00",
          7657 => x"6d",
          7658 => x"00",
          7659 => x"00",
          7660 => x"00",
          7661 => x"00",
          7662 => x"00",
          7663 => x"00",
          7664 => x"00",
          7665 => x"00",
          7666 => x"00",
          7667 => x"00",
          7668 => x"00",
          7669 => x"00",
          7670 => x"00",
          7671 => x"00",
          7672 => x"00",
          7673 => x"00",
          7674 => x"00",
          7675 => x"00",
          7676 => x"00",
          7677 => x"00",
          7678 => x"00",
          7679 => x"00",
          7680 => x"00",
          7681 => x"00",
          7682 => x"00",
          7683 => x"00",
          7684 => x"00",
          7685 => x"00",
          7686 => x"00",
          7687 => x"00",
          7688 => x"00",
          7689 => x"00",
          7690 => x"00",
          7691 => x"00",
          7692 => x"5b",
          7693 => x"5b",
          7694 => x"5b",
          7695 => x"5b",
          7696 => x"5b",
          7697 => x"5b",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"00",
          7703 => x"61",
          7704 => x"65",
          7705 => x"65",
          7706 => x"79",
          7707 => x"64",
          7708 => x"67",
          7709 => x"72",
          7710 => x"00",
          7711 => x"30",
          7712 => x"0a",
          7713 => x"64",
          7714 => x"65",
          7715 => x"69",
          7716 => x"69",
          7717 => x"4f",
          7718 => x"25",
          7719 => x"5b",
          7720 => x"5b",
          7721 => x"5b",
          7722 => x"5b",
          7723 => x"5b",
          7724 => x"5b",
          7725 => x"5b",
          7726 => x"5b",
          7727 => x"5b",
          7728 => x"5b",
          7729 => x"5b",
          7730 => x"5b",
          7731 => x"5b",
          7732 => x"5b",
          7733 => x"5b",
          7734 => x"5b",
          7735 => x"00",
          7736 => x"00",
          7737 => x"25",
          7738 => x"2c",
          7739 => x"30",
          7740 => x"3a",
          7741 => x"64",
          7742 => x"25",
          7743 => x"64",
          7744 => x"00",
          7745 => x"00",
          7746 => x"3b",
          7747 => x"65",
          7748 => x"72",
          7749 => x"70",
          7750 => x"30",
          7751 => x"77",
          7752 => x"30",
          7753 => x"64",
          7754 => x"00",
          7755 => x"78",
          7756 => x"49",
          7757 => x"61",
          7758 => x"20",
          7759 => x"00",
          7760 => x"78",
          7761 => x"57",
          7762 => x"6f",
          7763 => x"65",
          7764 => x"00",
          7765 => x"2a",
          7766 => x"00",
          7767 => x"5d",
          7768 => x"41",
          7769 => x"fe",
          7770 => x"2e",
          7771 => x"4d",
          7772 => x"54",
          7773 => x"4f",
          7774 => x"20",
          7775 => x"20",
          7776 => x"00",
          7777 => x"00",
          7778 => x"0e",
          7779 => x"00",
          7780 => x"41",
          7781 => x"49",
          7782 => x"4f",
          7783 => x"9d",
          7784 => x"a5",
          7785 => x"ad",
          7786 => x"b5",
          7787 => x"bd",
          7788 => x"c5",
          7789 => x"cd",
          7790 => x"d5",
          7791 => x"dd",
          7792 => x"e5",
          7793 => x"ed",
          7794 => x"f5",
          7795 => x"fd",
          7796 => x"5b",
          7797 => x"3e",
          7798 => x"01",
          7799 => x"00",
          7800 => x"01",
          7801 => x"10",
          7802 => x"c7",
          7803 => x"e4",
          7804 => x"ea",
          7805 => x"ee",
          7806 => x"c9",
          7807 => x"f6",
          7808 => x"ff",
          7809 => x"a3",
          7810 => x"e1",
          7811 => x"f1",
          7812 => x"bf",
          7813 => x"bc",
          7814 => x"91",
          7815 => x"24",
          7816 => x"55",
          7817 => x"5d",
          7818 => x"14",
          7819 => x"00",
          7820 => x"5a",
          7821 => x"60",
          7822 => x"68",
          7823 => x"58",
          7824 => x"6a",
          7825 => x"84",
          7826 => x"b1",
          7827 => x"a3",
          7828 => x"a6",
          7829 => x"1e",
          7830 => x"61",
          7831 => x"20",
          7832 => x"b0",
          7833 => x"7f",
          7834 => x"61",
          7835 => x"f8",
          7836 => x"78",
          7837 => x"06",
          7838 => x"2e",
          7839 => x"4d",
          7840 => x"82",
          7841 => x"87",
          7842 => x"8b",
          7843 => x"8f",
          7844 => x"93",
          7845 => x"97",
          7846 => x"9b",
          7847 => x"9f",
          7848 => x"a2",
          7849 => x"a7",
          7850 => x"ab",
          7851 => x"af",
          7852 => x"b3",
          7853 => x"b7",
          7854 => x"bb",
          7855 => x"f7",
          7856 => x"c3",
          7857 => x"c7",
          7858 => x"cb",
          7859 => x"dd",
          7860 => x"12",
          7861 => x"f4",
          7862 => x"22",
          7863 => x"65",
          7864 => x"66",
          7865 => x"41",
          7866 => x"40",
          7867 => x"89",
          7868 => x"5a",
          7869 => x"5e",
          7870 => x"62",
          7871 => x"66",
          7872 => x"6a",
          7873 => x"6e",
          7874 => x"9d",
          7875 => x"76",
          7876 => x"7a",
          7877 => x"7e",
          7878 => x"82",
          7879 => x"86",
          7880 => x"b1",
          7881 => x"8e",
          7882 => x"b7",
          7883 => x"fe",
          7884 => x"86",
          7885 => x"b1",
          7886 => x"a3",
          7887 => x"cc",
          7888 => x"8f",
          7889 => x"0a",
          7890 => x"f5",
          7891 => x"f9",
          7892 => x"20",
          7893 => x"22",
          7894 => x"0e",
          7895 => x"d0",
          7896 => x"00",
          7897 => x"63",
          7898 => x"5a",
          7899 => x"06",
          7900 => x"08",
          7901 => x"07",
          7902 => x"54",
          7903 => x"60",
          7904 => x"ba",
          7905 => x"ca",
          7906 => x"f8",
          7907 => x"fa",
          7908 => x"90",
          7909 => x"b0",
          7910 => x"b2",
          7911 => x"c3",
          7912 => x"02",
          7913 => x"f3",
          7914 => x"01",
          7915 => x"84",
          7916 => x"1a",
          7917 => x"02",
          7918 => x"02",
          7919 => x"26",
          7920 => x"00",
          7921 => x"02",
          7922 => x"00",
          7923 => x"04",
          7924 => x"00",
          7925 => x"14",
          7926 => x"00",
          7927 => x"2b",
          7928 => x"00",
          7929 => x"30",
          7930 => x"00",
          7931 => x"3c",
          7932 => x"00",
          7933 => x"3d",
          7934 => x"00",
          7935 => x"3f",
          7936 => x"00",
          7937 => x"40",
          7938 => x"00",
          7939 => x"41",
          7940 => x"00",
          7941 => x"42",
          7942 => x"00",
          7943 => x"43",
          7944 => x"00",
          7945 => x"50",
          7946 => x"00",
          7947 => x"51",
          7948 => x"00",
          7949 => x"54",
          7950 => x"00",
          7951 => x"55",
          7952 => x"00",
          7953 => x"79",
          7954 => x"00",
          7955 => x"78",
          7956 => x"00",
          7957 => x"82",
          7958 => x"00",
          7959 => x"83",
          7960 => x"00",
          7961 => x"85",
          7962 => x"00",
          7963 => x"87",
          7964 => x"00",
          7965 => x"88",
          7966 => x"00",
          7967 => x"89",
          7968 => x"00",
          7969 => x"8c",
          7970 => x"00",
          7971 => x"8d",
          7972 => x"00",
          7973 => x"8e",
          7974 => x"00",
          7975 => x"8f",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"01",
          7980 => x"01",
          7981 => x"00",
          7982 => x"00",
          7983 => x"00",
          7984 => x"f5",
          7985 => x"f5",
          7986 => x"01",
          7987 => x"01",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"00",
          7996 => x"00",
          7997 => x"00",
          7998 => x"00",
          7999 => x"00",
          8000 => x"00",
          8001 => x"00",
          8002 => x"00",
          8003 => x"01",
          8004 => x"3b",
          8005 => x"f0",
          8006 => x"76",
          8007 => x"6e",
          8008 => x"66",
          8009 => x"36",
          8010 => x"39",
          8011 => x"f2",
          8012 => x"f0",
          8013 => x"f0",
          8014 => x"3a",
          8015 => x"f0",
          8016 => x"56",
          8017 => x"4e",
          8018 => x"46",
          8019 => x"36",
          8020 => x"39",
          8021 => x"f2",
          8022 => x"f0",
          8023 => x"f0",
          8024 => x"2b",
          8025 => x"f0",
          8026 => x"56",
          8027 => x"4e",
          8028 => x"46",
          8029 => x"26",
          8030 => x"29",
          8031 => x"f8",
          8032 => x"f0",
          8033 => x"f0",
          8034 => x"f0",
          8035 => x"f0",
          8036 => x"16",
          8037 => x"0e",
          8038 => x"06",
          8039 => x"f0",
          8040 => x"1f",
          8041 => x"f0",
          8042 => x"f0",
          8043 => x"f0",
          8044 => x"b5",
          8045 => x"f0",
          8046 => x"a6",
          8047 => x"33",
          8048 => x"43",
          8049 => x"1e",
          8050 => x"a3",
          8051 => x"c4",
          8052 => x"f0",
          8053 => x"f0",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"01",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"e0",
          9090 => x"f9",
          9091 => x"c1",
          9092 => x"e4",
          9093 => x"61",
          9094 => x"69",
          9095 => x"21",
          9096 => x"29",
          9097 => x"01",
          9098 => x"09",
          9099 => x"11",
          9100 => x"19",
          9101 => x"81",
          9102 => x"89",
          9103 => x"91",
          9104 => x"99",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"00",
          9113 => x"00",
          9114 => x"00",
          9115 => x"00",
          9116 => x"00",
          9117 => x"00",
          9118 => x"00",
          9119 => x"00",
          9120 => x"02",
          9121 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"00",
             3 => x"00",
             4 => x"88",
             5 => x"08",
             6 => x"04",
             7 => x"00",
             8 => x"71",
             9 => x"81",
            10 => x"ff",
            11 => x"00",
            12 => x"71",
            13 => x"83",
            14 => x"2b",
            15 => x"0b",
            16 => x"72",
            17 => x"09",
            18 => x"07",
            19 => x"00",
            20 => x"72",
            21 => x"51",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"09",
            26 => x"0a",
            27 => x"51",
            28 => x"72",
            29 => x"51",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"72",
            45 => x"0b",
            46 => x"00",
            47 => x"00",
            48 => x"72",
            49 => x"09",
            50 => x"06",
            51 => x"00",
            52 => x"71",
            53 => x"06",
            54 => x"0b",
            55 => x"51",
            56 => x"72",
            57 => x"81",
            58 => x"51",
            59 => x"00",
            60 => x"72",
            61 => x"81",
            62 => x"53",
            63 => x"00",
            64 => x"71",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"72",
            69 => x"04",
            70 => x"00",
            71 => x"00",
            72 => x"72",
            73 => x"07",
            74 => x"00",
            75 => x"00",
            76 => x"71",
            77 => x"81",
            78 => x"81",
            79 => x"00",
            80 => x"71",
            81 => x"bc",
            82 => x"06",
            83 => x"00",
            84 => x"88",
            85 => x"0b",
            86 => x"88",
            87 => x"0c",
            88 => x"88",
            89 => x"0b",
            90 => x"88",
            91 => x"0c",
            92 => x"72",
            93 => x"81",
            94 => x"73",
            95 => x"07",
            96 => x"72",
            97 => x"09",
            98 => x"06",
            99 => x"06",
           100 => x"05",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"04",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"71",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"04",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"02",
           117 => x"04",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"02",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"0b",
           134 => x"96",
           135 => x"0b",
           136 => x"0b",
           137 => x"d6",
           138 => x"0b",
           139 => x"0b",
           140 => x"96",
           141 => x"0b",
           142 => x"0b",
           143 => x"d7",
           144 => x"0b",
           145 => x"0b",
           146 => x"9b",
           147 => x"0b",
           148 => x"0b",
           149 => x"df",
           150 => x"0b",
           151 => x"0b",
           152 => x"a3",
           153 => x"0b",
           154 => x"0b",
           155 => x"e7",
           156 => x"0b",
           157 => x"0b",
           158 => x"ab",
           159 => x"0b",
           160 => x"0b",
           161 => x"ef",
           162 => x"0b",
           163 => x"0b",
           164 => x"b3",
           165 => x"0b",
           166 => x"0b",
           167 => x"f7",
           168 => x"0b",
           169 => x"0b",
           170 => x"bb",
           171 => x"0b",
           172 => x"0b",
           173 => x"fe",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"04",
           193 => x"0c",
           194 => x"08",
           195 => x"98",
           196 => x"08",
           197 => x"98",
           198 => x"08",
           199 => x"98",
           200 => x"08",
           201 => x"98",
           202 => x"08",
           203 => x"98",
           204 => x"08",
           205 => x"98",
           206 => x"08",
           207 => x"98",
           208 => x"08",
           209 => x"98",
           210 => x"08",
           211 => x"98",
           212 => x"08",
           213 => x"98",
           214 => x"08",
           215 => x"98",
           216 => x"08",
           217 => x"98",
           218 => x"98",
           219 => x"ba",
           220 => x"ba",
           221 => x"84",
           222 => x"84",
           223 => x"04",
           224 => x"2d",
           225 => x"90",
           226 => x"f7",
           227 => x"80",
           228 => x"e3",
           229 => x"c0",
           230 => x"82",
           231 => x"80",
           232 => x"0c",
           233 => x"08",
           234 => x"98",
           235 => x"98",
           236 => x"ba",
           237 => x"ba",
           238 => x"84",
           239 => x"84",
           240 => x"04",
           241 => x"2d",
           242 => x"90",
           243 => x"d4",
           244 => x"80",
           245 => x"f4",
           246 => x"c0",
           247 => x"83",
           248 => x"80",
           249 => x"0c",
           250 => x"08",
           251 => x"98",
           252 => x"98",
           253 => x"ba",
           254 => x"ba",
           255 => x"84",
           256 => x"84",
           257 => x"04",
           258 => x"2d",
           259 => x"90",
           260 => x"99",
           261 => x"80",
           262 => x"e4",
           263 => x"c0",
           264 => x"82",
           265 => x"80",
           266 => x"0c",
           267 => x"08",
           268 => x"98",
           269 => x"98",
           270 => x"ba",
           271 => x"ba",
           272 => x"84",
           273 => x"84",
           274 => x"04",
           275 => x"2d",
           276 => x"90",
           277 => x"db",
           278 => x"80",
           279 => x"b9",
           280 => x"c0",
           281 => x"83",
           282 => x"80",
           283 => x"0c",
           284 => x"08",
           285 => x"98",
           286 => x"98",
           287 => x"ba",
           288 => x"ba",
           289 => x"84",
           290 => x"84",
           291 => x"04",
           292 => x"2d",
           293 => x"90",
           294 => x"94",
           295 => x"80",
           296 => x"9a",
           297 => x"80",
           298 => x"db",
           299 => x"c0",
           300 => x"81",
           301 => x"80",
           302 => x"0c",
           303 => x"08",
           304 => x"98",
           305 => x"98",
           306 => x"04",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"53",
           311 => x"06",
           312 => x"05",
           313 => x"06",
           314 => x"72",
           315 => x"05",
           316 => x"53",
           317 => x"04",
           318 => x"27",
           319 => x"53",
           320 => x"8c",
           321 => x"fc",
           322 => x"05",
           323 => x"d5",
           324 => x"3d",
           325 => x"7c",
           326 => x"80",
           327 => x"80",
           328 => x"80",
           329 => x"32",
           330 => x"51",
           331 => x"b7",
           332 => x"51",
           333 => x"53",
           334 => x"38",
           335 => x"05",
           336 => x"70",
           337 => x"54",
           338 => x"80",
           339 => x"8c",
           340 => x"84",
           341 => x"f5",
           342 => x"05",
           343 => x"58",
           344 => x"8d",
           345 => x"19",
           346 => x"04",
           347 => x"53",
           348 => x"3d",
           349 => x"65",
           350 => x"0c",
           351 => x"32",
           352 => x"72",
           353 => x"38",
           354 => x"c5",
           355 => x"5c",
           356 => x"17",
           357 => x"76",
           358 => x"51",
           359 => x"2e",
           360 => x"32",
           361 => x"9e",
           362 => x"33",
           363 => x"08",
           364 => x"3d",
           365 => x"10",
           366 => x"2b",
           367 => x"0a",
           368 => x"52",
           369 => x"81",
           370 => x"ff",
           371 => x"76",
           372 => x"a5",
           373 => x"73",
           374 => x"58",
           375 => x"39",
           376 => x"7b",
           377 => x"8d",
           378 => x"54",
           379 => x"06",
           380 => x"53",
           381 => x"10",
           382 => x"08",
           383 => x"d8",
           384 => x"51",
           385 => x"5b",
           386 => x"80",
           387 => x"7f",
           388 => x"ff",
           389 => x"ba",
           390 => x"9a",
           391 => x"06",
           392 => x"56",
           393 => x"ba",
           394 => x"70",
           395 => x"51",
           396 => x"56",
           397 => x"84",
           398 => x"06",
           399 => x"77",
           400 => x"05",
           401 => x"2a",
           402 => x"2e",
           403 => x"f8",
           404 => x"8b",
           405 => x"80",
           406 => x"7a",
           407 => x"72",
           408 => x"70",
           409 => x"24",
           410 => x"06",
           411 => x"56",
           412 => x"2e",
           413 => x"2b",
           414 => x"56",
           415 => x"38",
           416 => x"85",
           417 => x"54",
           418 => x"81",
           419 => x"81",
           420 => x"88",
           421 => x"b2",
           422 => x"fc",
           423 => x"40",
           424 => x"52",
           425 => x"84",
           426 => x"70",
           427 => x"24",
           428 => x"80",
           429 => x"0a",
           430 => x"2c",
           431 => x"38",
           432 => x"78",
           433 => x"0a",
           434 => x"74",
           435 => x"70",
           436 => x"81",
           437 => x"d8",
           438 => x"38",
           439 => x"7d",
           440 => x"52",
           441 => x"a5",
           442 => x"81",
           443 => x"7a",
           444 => x"84",
           445 => x"70",
           446 => x"25",
           447 => x"86",
           448 => x"5b",
           449 => x"76",
           450 => x"80",
           451 => x"60",
           452 => x"ff",
           453 => x"fb",
           454 => x"fe",
           455 => x"98",
           456 => x"29",
           457 => x"5e",
           458 => x"87",
           459 => x"fe",
           460 => x"29",
           461 => x"5a",
           462 => x"38",
           463 => x"e2",
           464 => x"06",
           465 => x"fe",
           466 => x"05",
           467 => x"39",
           468 => x"5b",
           469 => x"ab",
           470 => x"57",
           471 => x"75",
           472 => x"78",
           473 => x"05",
           474 => x"e3",
           475 => x"56",
           476 => x"39",
           477 => x"53",
           478 => x"df",
           479 => x"84",
           480 => x"84",
           481 => x"89",
           482 => x"5b",
           483 => x"f9",
           484 => x"05",
           485 => x"41",
           486 => x"87",
           487 => x"ff",
           488 => x"54",
           489 => x"39",
           490 => x"5b",
           491 => x"7f",
           492 => x"06",
           493 => x"38",
           494 => x"8c",
           495 => x"31",
           496 => x"81",
           497 => x"f7",
           498 => x"84",
           499 => x"70",
           500 => x"25",
           501 => x"83",
           502 => x"51",
           503 => x"81",
           504 => x"51",
           505 => x"06",
           506 => x"fa",
           507 => x"31",
           508 => x"80",
           509 => x"90",
           510 => x"51",
           511 => x"73",
           512 => x"39",
           513 => x"e5",
           514 => x"2e",
           515 => x"74",
           516 => x"53",
           517 => x"82",
           518 => x"51",
           519 => x"52",
           520 => x"8c",
           521 => x"31",
           522 => x"7a",
           523 => x"bf",
           524 => x"fe",
           525 => x"75",
           526 => x"3d",
           527 => x"80",
           528 => x"33",
           529 => x"06",
           530 => x"72",
           531 => x"38",
           532 => x"72",
           533 => x"08",
           534 => x"72",
           535 => x"83",
           536 => x"56",
           537 => x"84",
           538 => x"d5",
           539 => x"52",
           540 => x"2d",
           541 => x"38",
           542 => x"8c",
           543 => x"0d",
           544 => x"16",
           545 => x"81",
           546 => x"72",
           547 => x"73",
           548 => x"77",
           549 => x"56",
           550 => x"0d",
           551 => x"53",
           552 => x"72",
           553 => x"84",
           554 => x"ff",
           555 => x"57",
           556 => x"0d",
           557 => x"85",
           558 => x"0d",
           559 => x"2a",
           560 => x"57",
           561 => x"2a",
           562 => x"38",
           563 => x"08",
           564 => x"76",
           565 => x"8c",
           566 => x"0c",
           567 => x"88",
           568 => x"ff",
           569 => x"2d",
           570 => x"38",
           571 => x"0c",
           572 => x"77",
           573 => x"70",
           574 => x"56",
           575 => x"2a",
           576 => x"82",
           577 => x"80",
           578 => x"53",
           579 => x"13",
           580 => x"8c",
           581 => x"73",
           582 => x"04",
           583 => x"17",
           584 => x"17",
           585 => x"0c",
           586 => x"16",
           587 => x"08",
           588 => x"ff",
           589 => x"07",
           590 => x"2e",
           591 => x"85",
           592 => x"8c",
           593 => x"07",
           594 => x"ec",
           595 => x"54",
           596 => x"33",
           597 => x"72",
           598 => x"72",
           599 => x"38",
           600 => x"0d",
           601 => x"7a",
           602 => x"9d",
           603 => x"80",
           604 => x"53",
           605 => x"ff",
           606 => x"ba",
           607 => x"12",
           608 => x"14",
           609 => x"53",
           610 => x"51",
           611 => x"ff",
           612 => x"ff",
           613 => x"fe",
           614 => x"70",
           615 => x"38",
           616 => x"8c",
           617 => x"3d",
           618 => x"72",
           619 => x"72",
           620 => x"38",
           621 => x"0d",
           622 => x"79",
           623 => x"93",
           624 => x"73",
           625 => x"51",
           626 => x"0c",
           627 => x"76",
           628 => x"2e",
           629 => x"05",
           630 => x"09",
           631 => x"71",
           632 => x"72",
           633 => x"8c",
           634 => x"2e",
           635 => x"72",
           636 => x"52",
           637 => x"72",
           638 => x"3d",
           639 => x"86",
           640 => x"79",
           641 => x"84",
           642 => x"81",
           643 => x"84",
           644 => x"08",
           645 => x"08",
           646 => x"75",
           647 => x"b1",
           648 => x"84",
           649 => x"fd",
           650 => x"55",
           651 => x"72",
           652 => x"80",
           653 => x"ff",
           654 => x"13",
           655 => x"ba",
           656 => x"3d",
           657 => x"54",
           658 => x"72",
           659 => x"51",
           660 => x"0c",
           661 => x"78",
           662 => x"2e",
           663 => x"84",
           664 => x"73",
           665 => x"e3",
           666 => x"53",
           667 => x"38",
           668 => x"38",
           669 => x"31",
           670 => x"80",
           671 => x"10",
           672 => x"07",
           673 => x"70",
           674 => x"31",
           675 => x"58",
           676 => x"76",
           677 => x"88",
           678 => x"70",
           679 => x"72",
           680 => x"71",
           681 => x"80",
           682 => x"2b",
           683 => x"81",
           684 => x"82",
           685 => x"55",
           686 => x"70",
           687 => x"31",
           688 => x"32",
           689 => x"31",
           690 => x"0c",
           691 => x"5a",
           692 => x"56",
           693 => x"3d",
           694 => x"70",
           695 => x"3f",
           696 => x"71",
           697 => x"3d",
           698 => x"58",
           699 => x"38",
           700 => x"8c",
           701 => x"2e",
           702 => x"72",
           703 => x"53",
           704 => x"53",
           705 => x"74",
           706 => x"2b",
           707 => x"76",
           708 => x"2a",
           709 => x"31",
           710 => x"7b",
           711 => x"5c",
           712 => x"74",
           713 => x"88",
           714 => x"9f",
           715 => x"7b",
           716 => x"73",
           717 => x"31",
           718 => x"b4",
           719 => x"75",
           720 => x"0d",
           721 => x"57",
           722 => x"33",
           723 => x"81",
           724 => x"0c",
           725 => x"f3",
           726 => x"73",
           727 => x"58",
           728 => x"38",
           729 => x"80",
           730 => x"38",
           731 => x"53",
           732 => x"53",
           733 => x"70",
           734 => x"27",
           735 => x"83",
           736 => x"70",
           737 => x"73",
           738 => x"2e",
           739 => x"0c",
           740 => x"8b",
           741 => x"79",
           742 => x"b0",
           743 => x"81",
           744 => x"55",
           745 => x"58",
           746 => x"56",
           747 => x"53",
           748 => x"fe",
           749 => x"8b",
           750 => x"70",
           751 => x"56",
           752 => x"8c",
           753 => x"0d",
           754 => x"0c",
           755 => x"73",
           756 => x"81",
           757 => x"55",
           758 => x"2e",
           759 => x"83",
           760 => x"89",
           761 => x"56",
           762 => x"e0",
           763 => x"81",
           764 => x"81",
           765 => x"8f",
           766 => x"54",
           767 => x"72",
           768 => x"29",
           769 => x"33",
           770 => x"be",
           771 => x"30",
           772 => x"84",
           773 => x"81",
           774 => x"56",
           775 => x"06",
           776 => x"0c",
           777 => x"2e",
           778 => x"2e",
           779 => x"c6",
           780 => x"58",
           781 => x"84",
           782 => x"82",
           783 => x"33",
           784 => x"80",
           785 => x"0d",
           786 => x"8c",
           787 => x"0c",
           788 => x"93",
           789 => x"be",
           790 => x"ce",
           791 => x"0d",
           792 => x"3f",
           793 => x"51",
           794 => x"83",
           795 => x"3d",
           796 => x"92",
           797 => x"cc",
           798 => x"04",
           799 => x"83",
           800 => x"ee",
           801 => x"d0",
           802 => x"0d",
           803 => x"3f",
           804 => x"51",
           805 => x"83",
           806 => x"3d",
           807 => x"ba",
           808 => x"9c",
           809 => x"04",
           810 => x"83",
           811 => x"ee",
           812 => x"d1",
           813 => x"0d",
           814 => x"3f",
           815 => x"51",
           816 => x"83",
           817 => x"3d",
           818 => x"e2",
           819 => x"0d",
           820 => x"33",
           821 => x"7b",
           822 => x"78",
           823 => x"81",
           824 => x"06",
           825 => x"38",
           826 => x"52",
           827 => x"8c",
           828 => x"2e",
           829 => x"e0",
           830 => x"25",
           831 => x"53",
           832 => x"38",
           833 => x"87",
           834 => x"78",
           835 => x"84",
           836 => x"53",
           837 => x"df",
           838 => x"3d",
           839 => x"c0",
           840 => x"59",
           841 => x"53",
           842 => x"3f",
           843 => x"8c",
           844 => x"80",
           845 => x"17",
           846 => x"74",
           847 => x"08",
           848 => x"ba",
           849 => x"78",
           850 => x"3f",
           851 => x"02",
           852 => x"ff",
           853 => x"fd",
           854 => x"38",
           855 => x"2e",
           856 => x"8a",
           857 => x"ec",
           858 => x"8c",
           859 => x"84",
           860 => x"8a",
           861 => x"61",
           862 => x"33",
           863 => x"5c",
           864 => x"82",
           865 => x"dd",
           866 => x"f7",
           867 => x"38",
           868 => x"a0",
           869 => x"72",
           870 => x"52",
           871 => x"81",
           872 => x"a0",
           873 => x"dc",
           874 => x"3f",
           875 => x"38",
           876 => x"55",
           877 => x"80",
           878 => x"53",
           879 => x"56",
           880 => x"fe",
           881 => x"f0",
           882 => x"81",
           883 => x"83",
           884 => x"18",
           885 => x"b2",
           886 => x"70",
           887 => x"81",
           888 => x"38",
           889 => x"b9",
           890 => x"8f",
           891 => x"dc",
           892 => x"08",
           893 => x"78",
           894 => x"39",
           895 => x"82",
           896 => x"a0",
           897 => x"fe",
           898 => x"27",
           899 => x"e4",
           900 => x"d5",
           901 => x"c5",
           902 => x"99",
           903 => x"3f",
           904 => x"54",
           905 => x"27",
           906 => x"7a",
           907 => x"d2",
           908 => x"84",
           909 => x"ea",
           910 => x"fd",
           911 => x"73",
           912 => x"fe",
           913 => x"ba",
           914 => x"59",
           915 => x"59",
           916 => x"fc",
           917 => x"80",
           918 => x"08",
           919 => x"32",
           920 => x"70",
           921 => x"55",
           922 => x"25",
           923 => x"3f",
           924 => x"98",
           925 => x"9b",
           926 => x"75",
           927 => x"58",
           928 => x"fd",
           929 => x"0c",
           930 => x"87",
           931 => x"3f",
           932 => x"b4",
           933 => x"eb",
           934 => x"51",
           935 => x"2a",
           936 => x"89",
           937 => x"51",
           938 => x"2a",
           939 => x"ad",
           940 => x"51",
           941 => x"2a",
           942 => x"d2",
           943 => x"51",
           944 => x"81",
           945 => x"3f",
           946 => x"83",
           947 => x"3f",
           948 => x"3f",
           949 => x"eb",
           950 => x"3f",
           951 => x"2a",
           952 => x"38",
           953 => x"83",
           954 => x"51",
           955 => x"81",
           956 => x"9c",
           957 => x"3f",
           958 => x"80",
           959 => x"70",
           960 => x"fe",
           961 => x"9b",
           962 => x"9b",
           963 => x"85",
           964 => x"80",
           965 => x"81",
           966 => x"51",
           967 => x"3f",
           968 => x"52",
           969 => x"bd",
           970 => x"d4",
           971 => x"9a",
           972 => x"06",
           973 => x"38",
           974 => x"3f",
           975 => x"80",
           976 => x"70",
           977 => x"fd",
           978 => x"0d",
           979 => x"d1",
           980 => x"81",
           981 => x"81",
           982 => x"61",
           983 => x"51",
           984 => x"d5",
           985 => x"80",
           986 => x"ae",
           987 => x"70",
           988 => x"2e",
           989 => x"88",
           990 => x"82",
           991 => x"5a",
           992 => x"33",
           993 => x"8c",
           994 => x"7b",
           995 => x"9b",
           996 => x"ef",
           997 => x"ff",
           998 => x"8c",
           999 => x"5d",
          1000 => x"8b",
          1001 => x"2e",
          1002 => x"ff",
          1003 => x"38",
          1004 => x"fe",
          1005 => x"e9",
          1006 => x"84",
          1007 => x"38",
          1008 => x"ff",
          1009 => x"ba",
          1010 => x"7a",
          1011 => x"8c",
          1012 => x"8c",
          1013 => x"0b",
          1014 => x"8d",
          1015 => x"38",
          1016 => x"54",
          1017 => x"51",
          1018 => x"84",
          1019 => x"80",
          1020 => x"0a",
          1021 => x"ba",
          1022 => x"70",
          1023 => x"5b",
          1024 => x"83",
          1025 => x"78",
          1026 => x"81",
          1027 => x"38",
          1028 => x"5d",
          1029 => x"81",
          1030 => x"3f",
          1031 => x"7e",
          1032 => x"51",
          1033 => x"80",
          1034 => x"79",
          1035 => x"8c",
          1036 => x"96",
          1037 => x"38",
          1038 => x"34",
          1039 => x"7e",
          1040 => x"8c",
          1041 => x"8c",
          1042 => x"83",
          1043 => x"5f",
          1044 => x"fc",
          1045 => x"51",
          1046 => x"0b",
          1047 => x"53",
          1048 => x"3f",
          1049 => x"38",
          1050 => x"1b",
          1051 => x"80",
          1052 => x"05",
          1053 => x"51",
          1054 => x"53",
          1055 => x"f1",
          1056 => x"b8",
          1057 => x"8c",
          1058 => x"a4",
          1059 => x"41",
          1060 => x"de",
          1061 => x"3f",
          1062 => x"7b",
          1063 => x"83",
          1064 => x"3f",
          1065 => x"fa",
          1066 => x"39",
          1067 => x"fa",
          1068 => x"de",
          1069 => x"3f",
          1070 => x"51",
          1071 => x"c6",
          1072 => x"ff",
          1073 => x"ba",
          1074 => x"68",
          1075 => x"3f",
          1076 => x"08",
          1077 => x"8c",
          1078 => x"d7",
          1079 => x"84",
          1080 => x"c5",
          1081 => x"f9",
          1082 => x"51",
          1083 => x"b8",
          1084 => x"05",
          1085 => x"08",
          1086 => x"fe",
          1087 => x"e9",
          1088 => x"d0",
          1089 => x"52",
          1090 => x"84",
          1091 => x"7e",
          1092 => x"33",
          1093 => x"78",
          1094 => x"05",
          1095 => x"fe",
          1096 => x"e8",
          1097 => x"2e",
          1098 => x"11",
          1099 => x"3f",
          1100 => x"64",
          1101 => x"d7",
          1102 => x"ec",
          1103 => x"cf",
          1104 => x"78",
          1105 => x"26",
          1106 => x"46",
          1107 => x"11",
          1108 => x"3f",
          1109 => x"96",
          1110 => x"ff",
          1111 => x"ba",
          1112 => x"b8",
          1113 => x"05",
          1114 => x"08",
          1115 => x"cc",
          1116 => x"59",
          1117 => x"70",
          1118 => x"7d",
          1119 => x"78",
          1120 => x"51",
          1121 => x"81",
          1122 => x"b8",
          1123 => x"05",
          1124 => x"08",
          1125 => x"fe",
          1126 => x"e8",
          1127 => x"2e",
          1128 => x"11",
          1129 => x"3f",
          1130 => x"ee",
          1131 => x"3f",
          1132 => x"38",
          1133 => x"33",
          1134 => x"39",
          1135 => x"80",
          1136 => x"8c",
          1137 => x"3d",
          1138 => x"51",
          1139 => x"b1",
          1140 => x"d8",
          1141 => x"ec",
          1142 => x"cc",
          1143 => x"78",
          1144 => x"26",
          1145 => x"d1",
          1146 => x"33",
          1147 => x"3d",
          1148 => x"51",
          1149 => x"80",
          1150 => x"80",
          1151 => x"05",
          1152 => x"ff",
          1153 => x"ba",
          1154 => x"39",
          1155 => x"80",
          1156 => x"8c",
          1157 => x"3d",
          1158 => x"51",
          1159 => x"80",
          1160 => x"f8",
          1161 => x"bd",
          1162 => x"84",
          1163 => x"51",
          1164 => x"78",
          1165 => x"79",
          1166 => x"26",
          1167 => x"f4",
          1168 => x"51",
          1169 => x"b9",
          1170 => x"d8",
          1171 => x"52",
          1172 => x"8c",
          1173 => x"ba",
          1174 => x"8e",
          1175 => x"ff",
          1176 => x"ba",
          1177 => x"33",
          1178 => x"83",
          1179 => x"fc",
          1180 => x"a5",
          1181 => x"83",
          1182 => x"83",
          1183 => x"b8",
          1184 => x"05",
          1185 => x"08",
          1186 => x"5c",
          1187 => x"7a",
          1188 => x"9f",
          1189 => x"80",
          1190 => x"38",
          1191 => x"ba",
          1192 => x"66",
          1193 => x"d8",
          1194 => x"39",
          1195 => x"05",
          1196 => x"ff",
          1197 => x"ba",
          1198 => x"64",
          1199 => x"45",
          1200 => x"80",
          1201 => x"8c",
          1202 => x"5e",
          1203 => x"82",
          1204 => x"fe",
          1205 => x"e1",
          1206 => x"2e",
          1207 => x"ce",
          1208 => x"23",
          1209 => x"53",
          1210 => x"84",
          1211 => x"e6",
          1212 => x"ff",
          1213 => x"ba",
          1214 => x"68",
          1215 => x"34",
          1216 => x"b8",
          1217 => x"05",
          1218 => x"08",
          1219 => x"71",
          1220 => x"59",
          1221 => x"81",
          1222 => x"d6",
          1223 => x"52",
          1224 => x"39",
          1225 => x"f3",
          1226 => x"a2",
          1227 => x"f0",
          1228 => x"a1",
          1229 => x"b8",
          1230 => x"22",
          1231 => x"45",
          1232 => x"5c",
          1233 => x"f2",
          1234 => x"f3",
          1235 => x"38",
          1236 => x"39",
          1237 => x"64",
          1238 => x"51",
          1239 => x"39",
          1240 => x"2e",
          1241 => x"fc",
          1242 => x"a2",
          1243 => x"33",
          1244 => x"f2",
          1245 => x"f3",
          1246 => x"38",
          1247 => x"39",
          1248 => x"2e",
          1249 => x"fb",
          1250 => x"7c",
          1251 => x"08",
          1252 => x"33",
          1253 => x"f2",
          1254 => x"f2",
          1255 => x"9c",
          1256 => x"47",
          1257 => x"0b",
          1258 => x"8c",
          1259 => x"52",
          1260 => x"8c",
          1261 => x"87",
          1262 => x"3f",
          1263 => x"0c",
          1264 => x"57",
          1265 => x"9c",
          1266 => x"77",
          1267 => x"75",
          1268 => x"8c",
          1269 => x"0b",
          1270 => x"83",
          1271 => x"bc",
          1272 => x"02",
          1273 => x"84",
          1274 => x"13",
          1275 => x"0c",
          1276 => x"95",
          1277 => x"3f",
          1278 => x"51",
          1279 => x"22",
          1280 => x"84",
          1281 => x"33",
          1282 => x"3f",
          1283 => x"04",
          1284 => x"56",
          1285 => x"81",
          1286 => x"06",
          1287 => x"06",
          1288 => x"81",
          1289 => x"2e",
          1290 => x"73",
          1291 => x"72",
          1292 => x"33",
          1293 => x"70",
          1294 => x"80",
          1295 => x"38",
          1296 => x"81",
          1297 => x"09",
          1298 => x"a2",
          1299 => x"07",
          1300 => x"38",
          1301 => x"71",
          1302 => x"8c",
          1303 => x"2e",
          1304 => x"38",
          1305 => x"81",
          1306 => x"2e",
          1307 => x"15",
          1308 => x"2e",
          1309 => x"39",
          1310 => x"8b",
          1311 => x"86",
          1312 => x"52",
          1313 => x"8c",
          1314 => x"ba",
          1315 => x"3d",
          1316 => x"52",
          1317 => x"98",
          1318 => x"82",
          1319 => x"84",
          1320 => x"26",
          1321 => x"84",
          1322 => x"86",
          1323 => x"26",
          1324 => x"86",
          1325 => x"38",
          1326 => x"87",
          1327 => x"87",
          1328 => x"c0",
          1329 => x"c0",
          1330 => x"c0",
          1331 => x"c0",
          1332 => x"c0",
          1333 => x"c0",
          1334 => x"a4",
          1335 => x"80",
          1336 => x"52",
          1337 => x"0d",
          1338 => x"c0",
          1339 => x"c0",
          1340 => x"87",
          1341 => x"1c",
          1342 => x"79",
          1343 => x"08",
          1344 => x"98",
          1345 => x"87",
          1346 => x"1c",
          1347 => x"7b",
          1348 => x"08",
          1349 => x"0c",
          1350 => x"83",
          1351 => x"57",
          1352 => x"55",
          1353 => x"53",
          1354 => x"d8",
          1355 => x"3d",
          1356 => x"05",
          1357 => x"72",
          1358 => x"8c",
          1359 => x"52",
          1360 => x"38",
          1361 => x"ba",
          1362 => x"51",
          1363 => x"08",
          1364 => x"71",
          1365 => x"72",
          1366 => x"8c",
          1367 => x"52",
          1368 => x"fd",
          1369 => x"88",
          1370 => x"3f",
          1371 => x"98",
          1372 => x"38",
          1373 => x"83",
          1374 => x"8c",
          1375 => x"0d",
          1376 => x"33",
          1377 => x"70",
          1378 => x"94",
          1379 => x"06",
          1380 => x"38",
          1381 => x"51",
          1382 => x"06",
          1383 => x"93",
          1384 => x"73",
          1385 => x"80",
          1386 => x"c0",
          1387 => x"84",
          1388 => x"71",
          1389 => x"70",
          1390 => x"53",
          1391 => x"2a",
          1392 => x"38",
          1393 => x"2a",
          1394 => x"cf",
          1395 => x"8f",
          1396 => x"51",
          1397 => x"83",
          1398 => x"55",
          1399 => x"70",
          1400 => x"83",
          1401 => x"54",
          1402 => x"38",
          1403 => x"2a",
          1404 => x"80",
          1405 => x"81",
          1406 => x"81",
          1407 => x"8a",
          1408 => x"71",
          1409 => x"87",
          1410 => x"86",
          1411 => x"72",
          1412 => x"73",
          1413 => x"0c",
          1414 => x"70",
          1415 => x"72",
          1416 => x"2e",
          1417 => x"52",
          1418 => x"c0",
          1419 => x"81",
          1420 => x"d7",
          1421 => x"80",
          1422 => x"52",
          1423 => x"c0",
          1424 => x"87",
          1425 => x"0c",
          1426 => x"d0",
          1427 => x"f2",
          1428 => x"83",
          1429 => x"08",
          1430 => x"ac",
          1431 => x"9e",
          1432 => x"c0",
          1433 => x"87",
          1434 => x"0c",
          1435 => x"f0",
          1436 => x"f2",
          1437 => x"83",
          1438 => x"08",
          1439 => x"c0",
          1440 => x"87",
          1441 => x"0c",
          1442 => x"88",
          1443 => x"80",
          1444 => x"84",
          1445 => x"82",
          1446 => x"80",
          1447 => x"88",
          1448 => x"80",
          1449 => x"f3",
          1450 => x"90",
          1451 => x"52",
          1452 => x"52",
          1453 => x"87",
          1454 => x"80",
          1455 => x"83",
          1456 => x"34",
          1457 => x"70",
          1458 => x"70",
          1459 => x"83",
          1460 => x"9e",
          1461 => x"51",
          1462 => x"81",
          1463 => x"0b",
          1464 => x"80",
          1465 => x"2e",
          1466 => x"93",
          1467 => x"08",
          1468 => x"52",
          1469 => x"71",
          1470 => x"c0",
          1471 => x"06",
          1472 => x"38",
          1473 => x"80",
          1474 => x"80",
          1475 => x"80",
          1476 => x"f3",
          1477 => x"90",
          1478 => x"52",
          1479 => x"71",
          1480 => x"90",
          1481 => x"53",
          1482 => x"0b",
          1483 => x"80",
          1484 => x"83",
          1485 => x"34",
          1486 => x"06",
          1487 => x"f3",
          1488 => x"90",
          1489 => x"70",
          1490 => x"83",
          1491 => x"08",
          1492 => x"34",
          1493 => x"82",
          1494 => x"51",
          1495 => x"33",
          1496 => x"a0",
          1497 => x"33",
          1498 => x"93",
          1499 => x"f3",
          1500 => x"83",
          1501 => x"38",
          1502 => x"d6",
          1503 => x"84",
          1504 => x"73",
          1505 => x"55",
          1506 => x"33",
          1507 => x"8f",
          1508 => x"f3",
          1509 => x"83",
          1510 => x"38",
          1511 => x"ec",
          1512 => x"3f",
          1513 => x"c4",
          1514 => x"f4",
          1515 => x"b5",
          1516 => x"83",
          1517 => x"83",
          1518 => x"f2",
          1519 => x"ff",
          1520 => x"56",
          1521 => x"9c",
          1522 => x"c0",
          1523 => x"ba",
          1524 => x"ff",
          1525 => x"55",
          1526 => x"33",
          1527 => x"a5",
          1528 => x"88",
          1529 => x"51",
          1530 => x"bd",
          1531 => x"54",
          1532 => x"98",
          1533 => x"c2",
          1534 => x"f3",
          1535 => x"75",
          1536 => x"08",
          1537 => x"54",
          1538 => x"db",
          1539 => x"f3",
          1540 => x"94",
          1541 => x"51",
          1542 => x"c0",
          1543 => x"83",
          1544 => x"83",
          1545 => x"51",
          1546 => x"08",
          1547 => x"af",
          1548 => x"3f",
          1549 => x"c4",
          1550 => x"80",
          1551 => x"51",
          1552 => x"bd",
          1553 => x"54",
          1554 => x"ec",
          1555 => x"93",
          1556 => x"38",
          1557 => x"ff",
          1558 => x"54",
          1559 => x"ec",
          1560 => x"b2",
          1561 => x"80",
          1562 => x"dc",
          1563 => x"f3",
          1564 => x"c7",
          1565 => x"ff",
          1566 => x"54",
          1567 => x"39",
          1568 => x"ac",
          1569 => x"8d",
          1570 => x"38",
          1571 => x"83",
          1572 => x"83",
          1573 => x"fb",
          1574 => x"33",
          1575 => x"cf",
          1576 => x"80",
          1577 => x"f2",
          1578 => x"54",
          1579 => x"af",
          1580 => x"80",
          1581 => x"f2",
          1582 => x"54",
          1583 => x"8f",
          1584 => x"80",
          1585 => x"f2",
          1586 => x"54",
          1587 => x"ef",
          1588 => x"80",
          1589 => x"f2",
          1590 => x"54",
          1591 => x"cf",
          1592 => x"80",
          1593 => x"f2",
          1594 => x"54",
          1595 => x"af",
          1596 => x"80",
          1597 => x"de",
          1598 => x"d9",
          1599 => x"f3",
          1600 => x"cd",
          1601 => x"8e",
          1602 => x"38",
          1603 => x"52",
          1604 => x"ff",
          1605 => x"83",
          1606 => x"83",
          1607 => x"ff",
          1608 => x"83",
          1609 => x"83",
          1610 => x"ff",
          1611 => x"83",
          1612 => x"83",
          1613 => x"04",
          1614 => x"04",
          1615 => x"84",
          1616 => x"08",
          1617 => x"57",
          1618 => x"51",
          1619 => x"08",
          1620 => x"0b",
          1621 => x"f8",
          1622 => x"84",
          1623 => x"76",
          1624 => x"08",
          1625 => x"ba",
          1626 => x"8c",
          1627 => x"80",
          1628 => x"72",
          1629 => x"76",
          1630 => x"83",
          1631 => x"51",
          1632 => x"08",
          1633 => x"77",
          1634 => x"04",
          1635 => x"3f",
          1636 => x"38",
          1637 => x"79",
          1638 => x"08",
          1639 => x"76",
          1640 => x"c7",
          1641 => x"a9",
          1642 => x"3d",
          1643 => x"72",
          1644 => x"2e",
          1645 => x"59",
          1646 => x"80",
          1647 => x"af",
          1648 => x"52",
          1649 => x"ba",
          1650 => x"54",
          1651 => x"82",
          1652 => x"ff",
          1653 => x"38",
          1654 => x"aa",
          1655 => x"3d",
          1656 => x"51",
          1657 => x"80",
          1658 => x"52",
          1659 => x"8c",
          1660 => x"2e",
          1661 => x"06",
          1662 => x"38",
          1663 => x"56",
          1664 => x"15",
          1665 => x"a0",
          1666 => x"75",
          1667 => x"3d",
          1668 => x"ba",
          1669 => x"52",
          1670 => x"8c",
          1671 => x"08",
          1672 => x"cf",
          1673 => x"2e",
          1674 => x"3f",
          1675 => x"84",
          1676 => x"ba",
          1677 => x"55",
          1678 => x"81",
          1679 => x"ab",
          1680 => x"06",
          1681 => x"8c",
          1682 => x"0d",
          1683 => x"3d",
          1684 => x"3d",
          1685 => x"f8",
          1686 => x"83",
          1687 => x"2e",
          1688 => x"8d",
          1689 => x"78",
          1690 => x"fd",
          1691 => x"80",
          1692 => x"08",
          1693 => x"79",
          1694 => x"06",
          1695 => x"70",
          1696 => x"98",
          1697 => x"05",
          1698 => x"70",
          1699 => x"5d",
          1700 => x"57",
          1701 => x"75",
          1702 => x"0a",
          1703 => x"2c",
          1704 => x"38",
          1705 => x"57",
          1706 => x"42",
          1707 => x"de",
          1708 => x"41",
          1709 => x"80",
          1710 => x"34",
          1711 => x"38",
          1712 => x"2c",
          1713 => x"70",
          1714 => x"82",
          1715 => x"53",
          1716 => x"78",
          1717 => x"c8",
          1718 => x"ff",
          1719 => x"81",
          1720 => x"81",
          1721 => x"26",
          1722 => x"82",
          1723 => x"dc",
          1724 => x"ce",
          1725 => x"70",
          1726 => x"bc",
          1727 => x"fe",
          1728 => x"fe",
          1729 => x"fd",
          1730 => x"38",
          1731 => x"d1",
          1732 => x"0c",
          1733 => x"38",
          1734 => x"57",
          1735 => x"08",
          1736 => x"34",
          1737 => x"39",
          1738 => x"2e",
          1739 => x"52",
          1740 => x"d1",
          1741 => x"d1",
          1742 => x"d0",
          1743 => x"cc",
          1744 => x"fc",
          1745 => x"81",
          1746 => x"7b",
          1747 => x"d5",
          1748 => x"8b",
          1749 => x"a8",
          1750 => x"83",
          1751 => x"7c",
          1752 => x"d0",
          1753 => x"38",
          1754 => x"ff",
          1755 => x"52",
          1756 => x"d5",
          1757 => x"85",
          1758 => x"5b",
          1759 => x"ff",
          1760 => x"ff",
          1761 => x"34",
          1762 => x"f3",
          1763 => x"7c",
          1764 => x"11",
          1765 => x"74",
          1766 => x"38",
          1767 => x"ba",
          1768 => x"ba",
          1769 => x"53",
          1770 => x"3f",
          1771 => x"33",
          1772 => x"38",
          1773 => x"ff",
          1774 => x"52",
          1775 => x"d5",
          1776 => x"ed",
          1777 => x"55",
          1778 => x"ff",
          1779 => x"33",
          1780 => x"33",
          1781 => x"af",
          1782 => x"15",
          1783 => x"16",
          1784 => x"3f",
          1785 => x"06",
          1786 => x"75",
          1787 => x"f0",
          1788 => x"d1",
          1789 => x"55",
          1790 => x"33",
          1791 => x"33",
          1792 => x"a9",
          1793 => x"33",
          1794 => x"76",
          1795 => x"7a",
          1796 => x"70",
          1797 => x"57",
          1798 => x"84",
          1799 => x"b2",
          1800 => x"98",
          1801 => x"33",
          1802 => x"f9",
          1803 => x"88",
          1804 => x"80",
          1805 => x"98",
          1806 => x"5a",
          1807 => x"d5",
          1808 => x"ed",
          1809 => x"80",
          1810 => x"cc",
          1811 => x"ff",
          1812 => x"58",
          1813 => x"f0",
          1814 => x"bd",
          1815 => x"80",
          1816 => x"cc",
          1817 => x"fe",
          1818 => x"33",
          1819 => x"77",
          1820 => x"81",
          1821 => x"70",
          1822 => x"57",
          1823 => x"fe",
          1824 => x"74",
          1825 => x"f0",
          1826 => x"3f",
          1827 => x"76",
          1828 => x"06",
          1829 => x"7c",
          1830 => x"f0",
          1831 => x"3f",
          1832 => x"8b",
          1833 => x"06",
          1834 => x"cc",
          1835 => x"38",
          1836 => x"83",
          1837 => x"56",
          1838 => x"87",
          1839 => x"18",
          1840 => x"3f",
          1841 => x"f3",
          1842 => x"a4",
          1843 => x"8b",
          1844 => x"75",
          1845 => x"33",
          1846 => x"80",
          1847 => x"84",
          1848 => x"0c",
          1849 => x"33",
          1850 => x"d5",
          1851 => x"95",
          1852 => x"51",
          1853 => x"08",
          1854 => x"84",
          1855 => x"84",
          1856 => x"55",
          1857 => x"ff",
          1858 => x"d0",
          1859 => x"f5",
          1860 => x"81",
          1861 => x"74",
          1862 => x"08",
          1863 => x"84",
          1864 => x"ae",
          1865 => x"88",
          1866 => x"d0",
          1867 => x"d0",
          1868 => x"cc",
          1869 => x"9f",
          1870 => x"80",
          1871 => x"ba",
          1872 => x"d1",
          1873 => x"56",
          1874 => x"d1",
          1875 => x"d1",
          1876 => x"d1",
          1877 => x"88",
          1878 => x"d0",
          1879 => x"84",
          1880 => x"76",
          1881 => x"f0",
          1882 => x"3f",
          1883 => x"70",
          1884 => x"57",
          1885 => x"38",
          1886 => x"ff",
          1887 => x"29",
          1888 => x"84",
          1889 => x"79",
          1890 => x"08",
          1891 => x"74",
          1892 => x"05",
          1893 => x"5b",
          1894 => x"38",
          1895 => x"17",
          1896 => x"52",
          1897 => x"75",
          1898 => x"05",
          1899 => x"43",
          1900 => x"38",
          1901 => x"34",
          1902 => x"51",
          1903 => x"0a",
          1904 => x"2c",
          1905 => x"60",
          1906 => x"39",
          1907 => x"06",
          1908 => x"38",
          1909 => x"27",
          1910 => x"2c",
          1911 => x"7b",
          1912 => x"75",
          1913 => x"05",
          1914 => x"52",
          1915 => x"81",
          1916 => x"77",
          1917 => x"3d",
          1918 => x"57",
          1919 => x"56",
          1920 => x"84",
          1921 => x"29",
          1922 => x"79",
          1923 => x"60",
          1924 => x"2b",
          1925 => x"5c",
          1926 => x"38",
          1927 => x"ff",
          1928 => x"29",
          1929 => x"84",
          1930 => x"75",
          1931 => x"08",
          1932 => x"75",
          1933 => x"05",
          1934 => x"57",
          1935 => x"38",
          1936 => x"56",
          1937 => x"51",
          1938 => x"08",
          1939 => x"08",
          1940 => x"52",
          1941 => x"d1",
          1942 => x"56",
          1943 => x"d5",
          1944 => x"ad",
          1945 => x"51",
          1946 => x"08",
          1947 => x"84",
          1948 => x"84",
          1949 => x"55",
          1950 => x"3f",
          1951 => x"0c",
          1952 => x"76",
          1953 => x"38",
          1954 => x"52",
          1955 => x"a8",
          1956 => x"81",
          1957 => x"d1",
          1958 => x"24",
          1959 => x"98",
          1960 => x"06",
          1961 => x"ef",
          1962 => x"f8",
          1963 => x"f3",
          1964 => x"74",
          1965 => x"56",
          1966 => x"83",
          1967 => x"55",
          1968 => x"51",
          1969 => x"08",
          1970 => x"83",
          1971 => x"5f",
          1972 => x"da",
          1973 => x"84",
          1974 => x"ac",
          1975 => x"aa",
          1976 => x"d1",
          1977 => x"ff",
          1978 => x"51",
          1979 => x"d1",
          1980 => x"57",
          1981 => x"84",
          1982 => x"a6",
          1983 => x"a0",
          1984 => x"f0",
          1985 => x"3f",
          1986 => x"79",
          1987 => x"06",
          1988 => x"0b",
          1989 => x"d1",
          1990 => x"b4",
          1991 => x"ef",
          1992 => x"cc",
          1993 => x"06",
          1994 => x"ff",
          1995 => x"ff",
          1996 => x"d0",
          1997 => x"2e",
          1998 => x"52",
          1999 => x"d5",
          2000 => x"ed",
          2001 => x"51",
          2002 => x"33",
          2003 => x"34",
          2004 => x"75",
          2005 => x"8c",
          2006 => x"8c",
          2007 => x"75",
          2008 => x"ff",
          2009 => x"cc",
          2010 => x"5e",
          2011 => x"84",
          2012 => x"a5",
          2013 => x"a0",
          2014 => x"f0",
          2015 => x"3f",
          2016 => x"60",
          2017 => x"06",
          2018 => x"c9",
          2019 => x"2b",
          2020 => x"81",
          2021 => x"dd",
          2022 => x"0c",
          2023 => x"83",
          2024 => x"41",
          2025 => x"53",
          2026 => x"3f",
          2027 => x"81",
          2028 => x"82",
          2029 => x"f4",
          2030 => x"54",
          2031 => x"d9",
          2032 => x"8a",
          2033 => x"f8",
          2034 => x"0b",
          2035 => x"d1",
          2036 => x"b4",
          2037 => x"84",
          2038 => x"3f",
          2039 => x"84",
          2040 => x"83",
          2041 => x"7a",
          2042 => x"8c",
          2043 => x"2e",
          2044 => x"ba",
          2045 => x"84",
          2046 => x"ba",
          2047 => x"ba",
          2048 => x"56",
          2049 => x"83",
          2050 => x"f3",
          2051 => x"59",
          2052 => x"87",
          2053 => x"1a",
          2054 => x"3f",
          2055 => x"f3",
          2056 => x"a4",
          2057 => x"a0",
          2058 => x"5e",
          2059 => x"5d",
          2060 => x"df",
          2061 => x"39",
          2062 => x"a5",
          2063 => x"05",
          2064 => x"7a",
          2065 => x"f3",
          2066 => x"80",
          2067 => x"70",
          2068 => x"a4",
          2069 => x"57",
          2070 => x"08",
          2071 => x"10",
          2072 => x"57",
          2073 => x"38",
          2074 => x"34",
          2075 => x"34",
          2076 => x"ff",
          2077 => x"f8",
          2078 => x"c3",
          2079 => x"05",
          2080 => x"8d",
          2081 => x"81",
          2082 => x"2e",
          2083 => x"59",
          2084 => x"80",
          2085 => x"90",
          2086 => x"83",
          2087 => x"23",
          2088 => x"71",
          2089 => x"71",
          2090 => x"78",
          2091 => x"84",
          2092 => x"05",
          2093 => x"75",
          2094 => x"33",
          2095 => x"55",
          2096 => x"34",
          2097 => x"ff",
          2098 => x"0d",
          2099 => x"f9",
          2100 => x"f9",
          2101 => x"05",
          2102 => x"b0",
          2103 => x"81",
          2104 => x"81",
          2105 => x"83",
          2106 => x"59",
          2107 => x"73",
          2108 => x"29",
          2109 => x"ff",
          2110 => x"ff",
          2111 => x"75",
          2112 => x"5c",
          2113 => x"bc",
          2114 => x"29",
          2115 => x"7b",
          2116 => x"55",
          2117 => x"80",
          2118 => x"f9",
          2119 => x"34",
          2120 => x"87",
          2121 => x"33",
          2122 => x"33",
          2123 => x"22",
          2124 => x"5e",
          2125 => x"df",
          2126 => x"ff",
          2127 => x"54",
          2128 => x"0b",
          2129 => x"f9",
          2130 => x"98",
          2131 => x"2b",
          2132 => x"56",
          2133 => x"fd",
          2134 => x"f9",
          2135 => x"10",
          2136 => x"90",
          2137 => x"5e",
          2138 => x"b0",
          2139 => x"70",
          2140 => x"70",
          2141 => x"70",
          2142 => x"60",
          2143 => x"40",
          2144 => x"72",
          2145 => x"57",
          2146 => x"ff",
          2147 => x"ff",
          2148 => x"29",
          2149 => x"78",
          2150 => x"79",
          2151 => x"58",
          2152 => x"5c",
          2153 => x"74",
          2154 => x"39",
          2155 => x"54",
          2156 => x"34",
          2157 => x"34",
          2158 => x"56",
          2159 => x"80",
          2160 => x"ff",
          2161 => x"75",
          2162 => x"51",
          2163 => x"70",
          2164 => x"8c",
          2165 => x"54",
          2166 => x"80",
          2167 => x"72",
          2168 => x"70",
          2169 => x"87",
          2170 => x"f7",
          2171 => x"80",
          2172 => x"0b",
          2173 => x"04",
          2174 => x"0c",
          2175 => x"33",
          2176 => x"b7",
          2177 => x"75",
          2178 => x"80",
          2179 => x"bc",
          2180 => x"a0",
          2181 => x"51",
          2182 => x"83",
          2183 => x"53",
          2184 => x"c4",
          2185 => x"55",
          2186 => x"bc",
          2187 => x"7a",
          2188 => x"7a",
          2189 => x"72",
          2190 => x"22",
          2191 => x"fe",
          2192 => x"82",
          2193 => x"71",
          2194 => x"9f",
          2195 => x"14",
          2196 => x"e0",
          2197 => x"33",
          2198 => x"14",
          2199 => x"38",
          2200 => x"f9",
          2201 => x"55",
          2202 => x"73",
          2203 => x"54",
          2204 => x"b7",
          2205 => x"f9",
          2206 => x"06",
          2207 => x"73",
          2208 => x"31",
          2209 => x"71",
          2210 => x"a3",
          2211 => x"79",
          2212 => x"71",
          2213 => x"75",
          2214 => x"16",
          2215 => x"b8",
          2216 => x"5a",
          2217 => x"77",
          2218 => x"84",
          2219 => x"71",
          2220 => x"72",
          2221 => x"84",
          2222 => x"74",
          2223 => x"22",
          2224 => x"fe",
          2225 => x"fd",
          2226 => x"38",
          2227 => x"f9",
          2228 => x"09",
          2229 => x"31",
          2230 => x"71",
          2231 => x"59",
          2232 => x"83",
          2233 => x"74",
          2234 => x"e0",
          2235 => x"05",
          2236 => x"2e",
          2237 => x"16",
          2238 => x"34",
          2239 => x"f4",
          2240 => x"55",
          2241 => x"15",
          2242 => x"74",
          2243 => x"a9",
          2244 => x"05",
          2245 => x"26",
          2246 => x"b4",
          2247 => x"80",
          2248 => x"71",
          2249 => x"ba",
          2250 => x"0b",
          2251 => x"33",
          2252 => x"80",
          2253 => x"83",
          2254 => x"8c",
          2255 => x"bc",
          2256 => x"9f",
          2257 => x"70",
          2258 => x"f9",
          2259 => x"33",
          2260 => x"25",
          2261 => x"bc",
          2262 => x"86",
          2263 => x"70",
          2264 => x"72",
          2265 => x"f9",
          2266 => x"0c",
          2267 => x"33",
          2268 => x"11",
          2269 => x"38",
          2270 => x"80",
          2271 => x"0d",
          2272 => x"83",
          2273 => x"ff",
          2274 => x"b4",
          2275 => x"bc",
          2276 => x"02",
          2277 => x"b3",
          2278 => x"05",
          2279 => x"33",
          2280 => x"80",
          2281 => x"51",
          2282 => x"09",
          2283 => x"83",
          2284 => x"8c",
          2285 => x"b8",
          2286 => x"70",
          2287 => x"ba",
          2288 => x"f9",
          2289 => x"83",
          2290 => x"b8",
          2291 => x"70",
          2292 => x"f1",
          2293 => x"84",
          2294 => x"83",
          2295 => x"07",
          2296 => x"b4",
          2297 => x"51",
          2298 => x"39",
          2299 => x"85",
          2300 => x"ff",
          2301 => x"fb",
          2302 => x"b8",
          2303 => x"33",
          2304 => x"83",
          2305 => x"f9",
          2306 => x"83",
          2307 => x"f9",
          2308 => x"07",
          2309 => x"cc",
          2310 => x"06",
          2311 => x"34",
          2312 => x"81",
          2313 => x"83",
          2314 => x"f9",
          2315 => x"07",
          2316 => x"94",
          2317 => x"06",
          2318 => x"34",
          2319 => x"81",
          2320 => x"34",
          2321 => x"81",
          2322 => x"f9",
          2323 => x"0d",
          2324 => x"80",
          2325 => x"83",
          2326 => x"84",
          2327 => x"5b",
          2328 => x"78",
          2329 => x"81",
          2330 => x"80",
          2331 => x"f9",
          2332 => x"7c",
          2333 => x"04",
          2334 => x"38",
          2335 => x"0b",
          2336 => x"f9",
          2337 => x"34",
          2338 => x"58",
          2339 => x"ff",
          2340 => x"7b",
          2341 => x"c4",
          2342 => x"b8",
          2343 => x"34",
          2344 => x"f9",
          2345 => x"8f",
          2346 => x"82",
          2347 => x"80",
          2348 => x"83",
          2349 => x"ba",
          2350 => x"b9",
          2351 => x"56",
          2352 => x"52",
          2353 => x"3f",
          2354 => x"5a",
          2355 => x"84",
          2356 => x"83",
          2357 => x"81",
          2358 => x"8d",
          2359 => x"dd",
          2360 => x"c7",
          2361 => x"0b",
          2362 => x"bc",
          2363 => x"83",
          2364 => x"80",
          2365 => x"84",
          2366 => x"bc",
          2367 => x"81",
          2368 => x"f0",
          2369 => x"8c",
          2370 => x"ff",
          2371 => x"51",
          2372 => x"8c",
          2373 => x"f0",
          2374 => x"fe",
          2375 => x"ff",
          2376 => x"0d",
          2377 => x"84",
          2378 => x"83",
          2379 => x"87",
          2380 => x"22",
          2381 => x"05",
          2382 => x"92",
          2383 => x"72",
          2384 => x"2e",
          2385 => x"b9",
          2386 => x"75",
          2387 => x"80",
          2388 => x"bd",
          2389 => x"54",
          2390 => x"a0",
          2391 => x"83",
          2392 => x"72",
          2393 => x"75",
          2394 => x"bc",
          2395 => x"83",
          2396 => x"18",
          2397 => x"ff",
          2398 => x"bd",
          2399 => x"57",
          2400 => x"98",
          2401 => x"ff",
          2402 => x"99",
          2403 => x"81",
          2404 => x"f9",
          2405 => x"72",
          2406 => x"33",
          2407 => x"80",
          2408 => x"0d",
          2409 => x"8d",
          2410 => x"09",
          2411 => x"81",
          2412 => x"f9",
          2413 => x"be",
          2414 => x"33",
          2415 => x"06",
          2416 => x"a0",
          2417 => x"81",
          2418 => x"ff",
          2419 => x"a5",
          2420 => x"54",
          2421 => x"fa",
          2422 => x"f2",
          2423 => x"3f",
          2424 => x"3d",
          2425 => x"81",
          2426 => x"33",
          2427 => x"53",
          2428 => x"f9",
          2429 => x"d5",
          2430 => x"ff",
          2431 => x"a5",
          2432 => x"34",
          2433 => x"bd",
          2434 => x"3f",
          2435 => x"ef",
          2436 => x"0d",
          2437 => x"88",
          2438 => x"b8",
          2439 => x"78",
          2440 => x"24",
          2441 => x"b9",
          2442 => x"84",
          2443 => x"83",
          2444 => x"58",
          2445 => x"87",
          2446 => x"80",
          2447 => x"ba",
          2448 => x"42",
          2449 => x"83",
          2450 => x"05",
          2451 => x"87",
          2452 => x"80",
          2453 => x"ba",
          2454 => x"29",
          2455 => x"f9",
          2456 => x"81",
          2457 => x"76",
          2458 => x"81",
          2459 => x"19",
          2460 => x"0b",
          2461 => x"04",
          2462 => x"79",
          2463 => x"9b",
          2464 => x"cc",
          2465 => x"84",
          2466 => x"83",
          2467 => x"5e",
          2468 => x"87",
          2469 => x"80",
          2470 => x"ba",
          2471 => x"59",
          2472 => x"83",
          2473 => x"5b",
          2474 => x"b0",
          2475 => x"70",
          2476 => x"83",
          2477 => x"44",
          2478 => x"33",
          2479 => x"1f",
          2480 => x"77",
          2481 => x"bd",
          2482 => x"9c",
          2483 => x"b7",
          2484 => x"78",
          2485 => x"38",
          2486 => x"0b",
          2487 => x"04",
          2488 => x"19",
          2489 => x"84",
          2490 => x"77",
          2491 => x"90",
          2492 => x"80",
          2493 => x"0b",
          2494 => x"04",
          2495 => x"0b",
          2496 => x"33",
          2497 => x"33",
          2498 => x"84",
          2499 => x"80",
          2500 => x"f9",
          2501 => x"71",
          2502 => x"83",
          2503 => x"33",
          2504 => x"f9",
          2505 => x"34",
          2506 => x"06",
          2507 => x"33",
          2508 => x"58",
          2509 => x"98",
          2510 => x"89",
          2511 => x"3f",
          2512 => x"ae",
          2513 => x"bd",
          2514 => x"bc",
          2515 => x"a0",
          2516 => x"51",
          2517 => x"ff",
          2518 => x"51",
          2519 => x"a4",
          2520 => x"57",
          2521 => x"75",
          2522 => x"80",
          2523 => x"84",
          2524 => x"8e",
          2525 => x"81",
          2526 => x"84",
          2527 => x"83",
          2528 => x"83",
          2529 => x"83",
          2530 => x"80",
          2531 => x"84",
          2532 => x"78",
          2533 => x"a7",
          2534 => x"80",
          2535 => x"bd",
          2536 => x"29",
          2537 => x"f9",
          2538 => x"05",
          2539 => x"92",
          2540 => x"5c",
          2541 => x"81",
          2542 => x"83",
          2543 => x"34",
          2544 => x"06",
          2545 => x"05",
          2546 => x"87",
          2547 => x"80",
          2548 => x"ba",
          2549 => x"42",
          2550 => x"34",
          2551 => x"62",
          2552 => x"87",
          2553 => x"80",
          2554 => x"ba",
          2555 => x"29",
          2556 => x"f9",
          2557 => x"34",
          2558 => x"58",
          2559 => x"b8",
          2560 => x"ff",
          2561 => x"83",
          2562 => x"58",
          2563 => x"bb",
          2564 => x"83",
          2565 => x"38",
          2566 => x"f9",
          2567 => x"26",
          2568 => x"c6",
          2569 => x"0b",
          2570 => x"51",
          2571 => x"8c",
          2572 => x"bc",
          2573 => x"ff",
          2574 => x"ff",
          2575 => x"a0",
          2576 => x"41",
          2577 => x"ff",
          2578 => x"45",
          2579 => x"82",
          2580 => x"06",
          2581 => x"06",
          2582 => x"84",
          2583 => x"1b",
          2584 => x"bd",
          2585 => x"29",
          2586 => x"83",
          2587 => x"33",
          2588 => x"f9",
          2589 => x"34",
          2590 => x"06",
          2591 => x"33",
          2592 => x"40",
          2593 => x"de",
          2594 => x"ff",
          2595 => x"ac",
          2596 => x"92",
          2597 => x"f9",
          2598 => x"06",
          2599 => x"38",
          2600 => x"33",
          2601 => x"06",
          2602 => x"06",
          2603 => x"5b",
          2604 => x"a3",
          2605 => x"33",
          2606 => x"22",
          2607 => x"56",
          2608 => x"83",
          2609 => x"5a",
          2610 => x"b0",
          2611 => x"70",
          2612 => x"83",
          2613 => x"5b",
          2614 => x"33",
          2615 => x"05",
          2616 => x"7f",
          2617 => x"bd",
          2618 => x"b9",
          2619 => x"0c",
          2620 => x"17",
          2621 => x"7a",
          2622 => x"ff",
          2623 => x"39",
          2624 => x"0b",
          2625 => x"04",
          2626 => x"b8",
          2627 => x"bc",
          2628 => x"bd",
          2629 => x"f4",
          2630 => x"dc",
          2631 => x"cd",
          2632 => x"fb",
          2633 => x"11",
          2634 => x"79",
          2635 => x"ca",
          2636 => x"23",
          2637 => x"33",
          2638 => x"34",
          2639 => x"33",
          2640 => x"f9",
          2641 => x"f9",
          2642 => x"72",
          2643 => x"88",
          2644 => x"05",
          2645 => x"bd",
          2646 => x"29",
          2647 => x"f9",
          2648 => x"76",
          2649 => x"b8",
          2650 => x"34",
          2651 => x"06",
          2652 => x"33",
          2653 => x"42",
          2654 => x"de",
          2655 => x"06",
          2656 => x"38",
          2657 => x"e2",
          2658 => x"bd",
          2659 => x"84",
          2660 => x"f3",
          2661 => x"75",
          2662 => x"ea",
          2663 => x"0c",
          2664 => x"33",
          2665 => x"33",
          2666 => x"33",
          2667 => x"b9",
          2668 => x"f4",
          2669 => x"f5",
          2670 => x"f6",
          2671 => x"33",
          2672 => x"84",
          2673 => x"09",
          2674 => x"bd",
          2675 => x"33",
          2676 => x"8c",
          2677 => x"ed",
          2678 => x"3f",
          2679 => x"83",
          2680 => x"60",
          2681 => x"83",
          2682 => x"fe",
          2683 => x"33",
          2684 => x"77",
          2685 => x"84",
          2686 => x"41",
          2687 => x"10",
          2688 => x"08",
          2689 => x"80",
          2690 => x"33",
          2691 => x"70",
          2692 => x"42",
          2693 => x"34",
          2694 => x"56",
          2695 => x"b9",
          2696 => x"06",
          2697 => x"75",
          2698 => x"f9",
          2699 => x"83",
          2700 => x"70",
          2701 => x"2e",
          2702 => x"83",
          2703 => x"0b",
          2704 => x"33",
          2705 => x"57",
          2706 => x"17",
          2707 => x"f9",
          2708 => x"80",
          2709 => x"33",
          2710 => x"70",
          2711 => x"41",
          2712 => x"34",
          2713 => x"5b",
          2714 => x"b9",
          2715 => x"81",
          2716 => x"33",
          2717 => x"33",
          2718 => x"80",
          2719 => x"5a",
          2720 => x"ff",
          2721 => x"ff",
          2722 => x"7e",
          2723 => x"80",
          2724 => x"39",
          2725 => x"2e",
          2726 => x"58",
          2727 => x"d9",
          2728 => x"fb",
          2729 => x"75",
          2730 => x"e1",
          2731 => x"05",
          2732 => x"5e",
          2733 => x"57",
          2734 => x"39",
          2735 => x"2e",
          2736 => x"83",
          2737 => x"b7",
          2738 => x"75",
          2739 => x"83",
          2740 => x"e4",
          2741 => x"0b",
          2742 => x"76",
          2743 => x"b9",
          2744 => x"e3",
          2745 => x"17",
          2746 => x"33",
          2747 => x"84",
          2748 => x"2e",
          2749 => x"75",
          2750 => x"52",
          2751 => x"3f",
          2752 => x"57",
          2753 => x"b9",
          2754 => x"06",
          2755 => x"81",
          2756 => x"81",
          2757 => x"5b",
          2758 => x"38",
          2759 => x"76",
          2760 => x"77",
          2761 => x"83",
          2762 => x"ff",
          2763 => x"b4",
          2764 => x"34",
          2765 => x"5f",
          2766 => x"b9",
          2767 => x"5b",
          2768 => x"f9",
          2769 => x"81",
          2770 => x"74",
          2771 => x"83",
          2772 => x"29",
          2773 => x"f8",
          2774 => x"5d",
          2775 => x"83",
          2776 => x"57",
          2777 => x"b7",
          2778 => x"d6",
          2779 => x"ba",
          2780 => x"31",
          2781 => x"38",
          2782 => x"27",
          2783 => x"83",
          2784 => x"83",
          2785 => x"76",
          2786 => x"81",
          2787 => x"29",
          2788 => x"a0",
          2789 => x"81",
          2790 => x"71",
          2791 => x"7f",
          2792 => x"1a",
          2793 => x"b8",
          2794 => x"5d",
          2795 => x"7c",
          2796 => x"84",
          2797 => x"71",
          2798 => x"77",
          2799 => x"17",
          2800 => x"7b",
          2801 => x"81",
          2802 => x"5e",
          2803 => x"84",
          2804 => x"43",
          2805 => x"99",
          2806 => x"33",
          2807 => x"80",
          2808 => x"b1",
          2809 => x"b8",
          2810 => x"33",
          2811 => x"94",
          2812 => x"78",
          2813 => x"83",
          2814 => x"06",
          2815 => x"5c",
          2816 => x"b7",
          2817 => x"89",
          2818 => x"76",
          2819 => x"61",
          2820 => x"38",
          2821 => x"62",
          2822 => x"1f",
          2823 => x"79",
          2824 => x"ac",
          2825 => x"a4",
          2826 => x"2b",
          2827 => x"07",
          2828 => x"57",
          2829 => x"70",
          2830 => x"84",
          2831 => x"38",
          2832 => x"33",
          2833 => x"81",
          2834 => x"73",
          2835 => x"77",
          2836 => x"1b",
          2837 => x"75",
          2838 => x"f4",
          2839 => x"98",
          2840 => x"e0",
          2841 => x"5a",
          2842 => x"f4",
          2843 => x"34",
          2844 => x"81",
          2845 => x"f4",
          2846 => x"06",
          2847 => x"b8",
          2848 => x"2b",
          2849 => x"58",
          2850 => x"81",
          2851 => x"f9",
          2852 => x"06",
          2853 => x"be",
          2854 => x"33",
          2855 => x"b8",
          2856 => x"b7",
          2857 => x"ee",
          2858 => x"56",
          2859 => x"70",
          2860 => x"39",
          2861 => x"85",
          2862 => x"e5",
          2863 => x"06",
          2864 => x"34",
          2865 => x"f9",
          2866 => x"b8",
          2867 => x"81",
          2868 => x"f9",
          2869 => x"0b",
          2870 => x"81",
          2871 => x"83",
          2872 => x"75",
          2873 => x"83",
          2874 => x"07",
          2875 => x"fd",
          2876 => x"06",
          2877 => x"b8",
          2878 => x"33",
          2879 => x"75",
          2880 => x"83",
          2881 => x"07",
          2882 => x"c5",
          2883 => x"06",
          2884 => x"34",
          2885 => x"81",
          2886 => x"f9",
          2887 => x"b8",
          2888 => x"75",
          2889 => x"83",
          2890 => x"75",
          2891 => x"83",
          2892 => x"75",
          2893 => x"83",
          2894 => x"75",
          2895 => x"83",
          2896 => x"d0",
          2897 => x"fd",
          2898 => x"bf",
          2899 => x"b8",
          2900 => x"f9",
          2901 => x"c9",
          2902 => x"33",
          2903 => x"33",
          2904 => x"33",
          2905 => x"0b",
          2906 => x"81",
          2907 => x"84",
          2908 => x"77",
          2909 => x"33",
          2910 => x"56",
          2911 => x"9c",
          2912 => x"fe",
          2913 => x"a1",
          2914 => x"88",
          2915 => x"80",
          2916 => x"0d",
          2917 => x"e9",
          2918 => x"5c",
          2919 => x"10",
          2920 => x"05",
          2921 => x"0b",
          2922 => x"0b",
          2923 => x"51",
          2924 => x"70",
          2925 => x"e6",
          2926 => x"34",
          2927 => x"ef",
          2928 => x"3f",
          2929 => x"ff",
          2930 => x"06",
          2931 => x"52",
          2932 => x"33",
          2933 => x"75",
          2934 => x"83",
          2935 => x"70",
          2936 => x"f0",
          2937 => x"05",
          2938 => x"59",
          2939 => x"75",
          2940 => x"33",
          2941 => x"77",
          2942 => x"33",
          2943 => x"06",
          2944 => x"11",
          2945 => x"ba",
          2946 => x"70",
          2947 => x"33",
          2948 => x"81",
          2949 => x"ff",
          2950 => x"24",
          2951 => x"56",
          2952 => x"16",
          2953 => x"81",
          2954 => x"76",
          2955 => x"33",
          2956 => x"ff",
          2957 => x"7b",
          2958 => x"57",
          2959 => x"38",
          2960 => x"ff",
          2961 => x"79",
          2962 => x"a3",
          2963 => x"81",
          2964 => x"42",
          2965 => x"38",
          2966 => x"17",
          2967 => x"7b",
          2968 => x"81",
          2969 => x"5f",
          2970 => x"84",
          2971 => x"59",
          2972 => x"b1",
          2973 => x"b8",
          2974 => x"5d",
          2975 => x"7d",
          2976 => x"84",
          2977 => x"71",
          2978 => x"75",
          2979 => x"39",
          2980 => x"b8",
          2981 => x"bc",
          2982 => x"ba",
          2983 => x"5f",
          2984 => x"38",
          2985 => x"06",
          2986 => x"27",
          2987 => x"ba",
          2988 => x"58",
          2989 => x"57",
          2990 => x"80",
          2991 => x"52",
          2992 => x"38",
          2993 => x"eb",
          2994 => x"05",
          2995 => x"40",
          2996 => x"75",
          2997 => x"09",
          2998 => x"bd",
          2999 => x"bc",
          3000 => x"ff",
          3001 => x"f6",
          3002 => x"f9",
          3003 => x"56",
          3004 => x"39",
          3005 => x"bc",
          3006 => x"56",
          3007 => x"76",
          3008 => x"b8",
          3009 => x"75",
          3010 => x"70",
          3011 => x"33",
          3012 => x"76",
          3013 => x"7b",
          3014 => x"f1",
          3015 => x"34",
          3016 => x"23",
          3017 => x"ba",
          3018 => x"f9",
          3019 => x"be",
          3020 => x"33",
          3021 => x"34",
          3022 => x"97",
          3023 => x"54",
          3024 => x"db",
          3025 => x"0c",
          3026 => x"51",
          3027 => x"8c",
          3028 => x"0d",
          3029 => x"83",
          3030 => x"83",
          3031 => x"59",
          3032 => x"14",
          3033 => x"59",
          3034 => x"0d",
          3035 => x"53",
          3036 => x"32",
          3037 => x"9f",
          3038 => x"f7",
          3039 => x"81",
          3040 => x"54",
          3041 => x"25",
          3042 => x"2e",
          3043 => x"83",
          3044 => x"72",
          3045 => x"05",
          3046 => x"71",
          3047 => x"06",
          3048 => x"58",
          3049 => x"f0",
          3050 => x"80",
          3051 => x"c0",
          3052 => x"f6",
          3053 => x"76",
          3054 => x"70",
          3055 => x"74",
          3056 => x"ac",
          3057 => x"f7",
          3058 => x"76",
          3059 => x"2e",
          3060 => x"15",
          3061 => x"81",
          3062 => x"f7",
          3063 => x"33",
          3064 => x"70",
          3065 => x"27",
          3066 => x"70",
          3067 => x"54",
          3068 => x"ff",
          3069 => x"81",
          3070 => x"85",
          3071 => x"34",
          3072 => x"2e",
          3073 => x"e6",
          3074 => x"83",
          3075 => x"70",
          3076 => x"33",
          3077 => x"83",
          3078 => x"ff",
          3079 => x"33",
          3080 => x"83",
          3081 => x"ff",
          3082 => x"33",
          3083 => x"ff",
          3084 => x"38",
          3085 => x"81",
          3086 => x"06",
          3087 => x"38",
          3088 => x"74",
          3089 => x"08",
          3090 => x"08",
          3091 => x"38",
          3092 => x"83",
          3093 => x"81",
          3094 => x"fe",
          3095 => x"77",
          3096 => x"53",
          3097 => x"10",
          3098 => x"08",
          3099 => x"80",
          3100 => x"c0",
          3101 => x"27",
          3102 => x"92",
          3103 => x"38",
          3104 => x"87",
          3105 => x"0c",
          3106 => x"2e",
          3107 => x"54",
          3108 => x"81",
          3109 => x"ec",
          3110 => x"38",
          3111 => x"c3",
          3112 => x"39",
          3113 => x"56",
          3114 => x"38",
          3115 => x"b4",
          3116 => x"79",
          3117 => x"ff",
          3118 => x"2b",
          3119 => x"73",
          3120 => x"81",
          3121 => x"87",
          3122 => x"57",
          3123 => x"78",
          3124 => x"11",
          3125 => x"05",
          3126 => x"c0",
          3127 => x"57",
          3128 => x"2e",
          3129 => x"59",
          3130 => x"39",
          3131 => x"0b",
          3132 => x"81",
          3133 => x"70",
          3134 => x"59",
          3135 => x"09",
          3136 => x"2e",
          3137 => x"10",
          3138 => x"5d",
          3139 => x"81",
          3140 => x"93",
          3141 => x"33",
          3142 => x"84",
          3143 => x"38",
          3144 => x"cc",
          3145 => x"8f",
          3146 => x"f0",
          3147 => x"2e",
          3148 => x"81",
          3149 => x"34",
          3150 => x"d4",
          3151 => x"15",
          3152 => x"34",
          3153 => x"53",
          3154 => x"83",
          3155 => x"27",
          3156 => x"54",
          3157 => x"fc",
          3158 => x"05",
          3159 => x"74",
          3160 => x"98",
          3161 => x"81",
          3162 => x"0b",
          3163 => x"39",
          3164 => x"81",
          3165 => x"83",
          3166 => x"e5",
          3167 => x"e6",
          3168 => x"f7",
          3169 => x"5e",
          3170 => x"09",
          3171 => x"7a",
          3172 => x"2e",
          3173 => x"93",
          3174 => x"f8",
          3175 => x"33",
          3176 => x"73",
          3177 => x"ac",
          3178 => x"58",
          3179 => x"84",
          3180 => x"39",
          3181 => x"2e",
          3182 => x"ec",
          3183 => x"33",
          3184 => x"5a",
          3185 => x"55",
          3186 => x"ff",
          3187 => x"27",
          3188 => x"bc",
          3189 => x"ff",
          3190 => x"27",
          3191 => x"bd",
          3192 => x"52",
          3193 => x"59",
          3194 => x"39",
          3195 => x"51",
          3196 => x"f8",
          3197 => x"fc",
          3198 => x"f5",
          3199 => x"3d",
          3200 => x"54",
          3201 => x"34",
          3202 => x"72",
          3203 => x"56",
          3204 => x"0b",
          3205 => x"98",
          3206 => x"80",
          3207 => x"9c",
          3208 => x"52",
          3209 => x"33",
          3210 => x"75",
          3211 => x"2e",
          3212 => x"52",
          3213 => x"38",
          3214 => x"38",
          3215 => x"90",
          3216 => x"53",
          3217 => x"73",
          3218 => x"c0",
          3219 => x"27",
          3220 => x"38",
          3221 => x"56",
          3222 => x"72",
          3223 => x"a3",
          3224 => x"fe",
          3225 => x"77",
          3226 => x"04",
          3227 => x"54",
          3228 => x"d4",
          3229 => x"84",
          3230 => x"f9",
          3231 => x"05",
          3232 => x"98",
          3233 => x"80",
          3234 => x"56",
          3235 => x"90",
          3236 => x"90",
          3237 => x"86",
          3238 => x"75",
          3239 => x"52",
          3240 => x"f4",
          3241 => x"16",
          3242 => x"34",
          3243 => x"98",
          3244 => x"87",
          3245 => x"98",
          3246 => x"38",
          3247 => x"08",
          3248 => x"72",
          3249 => x"98",
          3250 => x"27",
          3251 => x"2e",
          3252 => x"08",
          3253 => x"98",
          3254 => x"08",
          3255 => x"15",
          3256 => x"53",
          3257 => x"ff",
          3258 => x"08",
          3259 => x"df",
          3260 => x"d7",
          3261 => x"75",
          3262 => x"38",
          3263 => x"76",
          3264 => x"80",
          3265 => x"92",
          3266 => x"72",
          3267 => x"26",
          3268 => x"89",
          3269 => x"e8",
          3270 => x"84",
          3271 => x"ff",
          3272 => x"76",
          3273 => x"39",
          3274 => x"a7",
          3275 => x"f4",
          3276 => x"80",
          3277 => x"51",
          3278 => x"73",
          3279 => x"76",
          3280 => x"73",
          3281 => x"08",
          3282 => x"55",
          3283 => x"71",
          3284 => x"81",
          3285 => x"38",
          3286 => x"16",
          3287 => x"e2",
          3288 => x"08",
          3289 => x"80",
          3290 => x"c0",
          3291 => x"56",
          3292 => x"98",
          3293 => x"08",
          3294 => x"15",
          3295 => x"53",
          3296 => x"fe",
          3297 => x"08",
          3298 => x"cd",
          3299 => x"c5",
          3300 => x"ce",
          3301 => x"08",
          3302 => x"75",
          3303 => x"87",
          3304 => x"74",
          3305 => x"db",
          3306 => x"ff",
          3307 => x"56",
          3308 => x"2e",
          3309 => x"72",
          3310 => x"06",
          3311 => x"ba",
          3312 => x"17",
          3313 => x"da",
          3314 => x"52",
          3315 => x"83",
          3316 => x"3f",
          3317 => x"0d",
          3318 => x"08",
          3319 => x"83",
          3320 => x"81",
          3321 => x"e8",
          3322 => x"f4",
          3323 => x"54",
          3324 => x"c0",
          3325 => x"f6",
          3326 => x"9c",
          3327 => x"38",
          3328 => x"c0",
          3329 => x"74",
          3330 => x"ff",
          3331 => x"9c",
          3332 => x"c0",
          3333 => x"9c",
          3334 => x"81",
          3335 => x"52",
          3336 => x"81",
          3337 => x"a4",
          3338 => x"98",
          3339 => x"38",
          3340 => x"ff",
          3341 => x"39",
          3342 => x"54",
          3343 => x"90",
          3344 => x"0d",
          3345 => x"08",
          3346 => x"ff",
          3347 => x"70",
          3348 => x"71",
          3349 => x"81",
          3350 => x"2b",
          3351 => x"57",
          3352 => x"24",
          3353 => x"33",
          3354 => x"83",
          3355 => x"12",
          3356 => x"07",
          3357 => x"80",
          3358 => x"33",
          3359 => x"83",
          3360 => x"52",
          3361 => x"73",
          3362 => x"34",
          3363 => x"12",
          3364 => x"07",
          3365 => x"51",
          3366 => x"34",
          3367 => x"0b",
          3368 => x"34",
          3369 => x"14",
          3370 => x"fc",
          3371 => x"71",
          3372 => x"70",
          3373 => x"72",
          3374 => x"0d",
          3375 => x"71",
          3376 => x"11",
          3377 => x"88",
          3378 => x"54",
          3379 => x"34",
          3380 => x"08",
          3381 => x"33",
          3382 => x"56",
          3383 => x"33",
          3384 => x"70",
          3385 => x"86",
          3386 => x"b9",
          3387 => x"33",
          3388 => x"06",
          3389 => x"76",
          3390 => x"b9",
          3391 => x"12",
          3392 => x"07",
          3393 => x"71",
          3394 => x"ff",
          3395 => x"54",
          3396 => x"52",
          3397 => x"34",
          3398 => x"33",
          3399 => x"83",
          3400 => x"12",
          3401 => x"ff",
          3402 => x"55",
          3403 => x"70",
          3404 => x"70",
          3405 => x"71",
          3406 => x"05",
          3407 => x"2b",
          3408 => x"52",
          3409 => x"fc",
          3410 => x"71",
          3411 => x"70",
          3412 => x"34",
          3413 => x"08",
          3414 => x"71",
          3415 => x"05",
          3416 => x"88",
          3417 => x"5c",
          3418 => x"15",
          3419 => x"0d",
          3420 => x"fc",
          3421 => x"38",
          3422 => x"fb",
          3423 => x"ff",
          3424 => x"80",
          3425 => x"80",
          3426 => x"fe",
          3427 => x"55",
          3428 => x"34",
          3429 => x"15",
          3430 => x"b9",
          3431 => x"81",
          3432 => x"08",
          3433 => x"80",
          3434 => x"70",
          3435 => x"88",
          3436 => x"b9",
          3437 => x"b9",
          3438 => x"76",
          3439 => x"34",
          3440 => x"52",
          3441 => x"8e",
          3442 => x"70",
          3443 => x"83",
          3444 => x"84",
          3445 => x"2b",
          3446 => x"81",
          3447 => x"cc",
          3448 => x"33",
          3449 => x"70",
          3450 => x"83",
          3451 => x"53",
          3452 => x"8a",
          3453 => x"73",
          3454 => x"33",
          3455 => x"c1",
          3456 => x"38",
          3457 => x"2b",
          3458 => x"71",
          3459 => x"06",
          3460 => x"79",
          3461 => x"74",
          3462 => x"78",
          3463 => x"2e",
          3464 => x"2b",
          3465 => x"70",
          3466 => x"76",
          3467 => x"b9",
          3468 => x"53",
          3469 => x"34",
          3470 => x"33",
          3471 => x"70",
          3472 => x"05",
          3473 => x"2a",
          3474 => x"75",
          3475 => x"53",
          3476 => x"08",
          3477 => x"15",
          3478 => x"86",
          3479 => x"2b",
          3480 => x"5c",
          3481 => x"72",
          3482 => x"70",
          3483 => x"87",
          3484 => x"88",
          3485 => x"15",
          3486 => x"fc",
          3487 => x"12",
          3488 => x"07",
          3489 => x"75",
          3490 => x"84",
          3491 => x"05",
          3492 => x"88",
          3493 => x"57",
          3494 => x"15",
          3495 => x"05",
          3496 => x"3d",
          3497 => x"33",
          3498 => x"79",
          3499 => x"71",
          3500 => x"5b",
          3501 => x"34",
          3502 => x"08",
          3503 => x"33",
          3504 => x"74",
          3505 => x"71",
          3506 => x"5d",
          3507 => x"86",
          3508 => x"b9",
          3509 => x"33",
          3510 => x"06",
          3511 => x"75",
          3512 => x"b9",
          3513 => x"f1",
          3514 => x"fc",
          3515 => x"38",
          3516 => x"ba",
          3517 => x"51",
          3518 => x"84",
          3519 => x"84",
          3520 => x"a0",
          3521 => x"80",
          3522 => x"51",
          3523 => x"08",
          3524 => x"16",
          3525 => x"84",
          3526 => x"84",
          3527 => x"34",
          3528 => x"fc",
          3529 => x"fe",
          3530 => x"06",
          3531 => x"74",
          3532 => x"84",
          3533 => x"84",
          3534 => x"55",
          3535 => x"15",
          3536 => x"dd",
          3537 => x"65",
          3538 => x"fc",
          3539 => x"84",
          3540 => x"38",
          3541 => x"54",
          3542 => x"05",
          3543 => x"ff",
          3544 => x"06",
          3545 => x"ff",
          3546 => x"70",
          3547 => x"07",
          3548 => x"06",
          3549 => x"83",
          3550 => x"33",
          3551 => x"70",
          3552 => x"53",
          3553 => x"5e",
          3554 => x"38",
          3555 => x"88",
          3556 => x"70",
          3557 => x"71",
          3558 => x"56",
          3559 => x"7a",
          3560 => x"58",
          3561 => x"80",
          3562 => x"77",
          3563 => x"59",
          3564 => x"1e",
          3565 => x"2b",
          3566 => x"33",
          3567 => x"90",
          3568 => x"57",
          3569 => x"38",
          3570 => x"33",
          3571 => x"7a",
          3572 => x"71",
          3573 => x"05",
          3574 => x"88",
          3575 => x"48",
          3576 => x"56",
          3577 => x"34",
          3578 => x"11",
          3579 => x"71",
          3580 => x"33",
          3581 => x"70",
          3582 => x"57",
          3583 => x"87",
          3584 => x"70",
          3585 => x"07",
          3586 => x"5a",
          3587 => x"81",
          3588 => x"1f",
          3589 => x"8b",
          3590 => x"73",
          3591 => x"07",
          3592 => x"5f",
          3593 => x"81",
          3594 => x"1f",
          3595 => x"2b",
          3596 => x"14",
          3597 => x"07",
          3598 => x"5f",
          3599 => x"75",
          3600 => x"70",
          3601 => x"71",
          3602 => x"70",
          3603 => x"05",
          3604 => x"84",
          3605 => x"65",
          3606 => x"5d",
          3607 => x"38",
          3608 => x"95",
          3609 => x"84",
          3610 => x"b9",
          3611 => x"52",
          3612 => x"3f",
          3613 => x"34",
          3614 => x"fc",
          3615 => x"0b",
          3616 => x"5c",
          3617 => x"1d",
          3618 => x"f8",
          3619 => x"70",
          3620 => x"5c",
          3621 => x"77",
          3622 => x"70",
          3623 => x"05",
          3624 => x"34",
          3625 => x"fc",
          3626 => x"80",
          3627 => x"80",
          3628 => x"9b",
          3629 => x"8c",
          3630 => x"84",
          3631 => x"11",
          3632 => x"12",
          3633 => x"ff",
          3634 => x"5e",
          3635 => x"34",
          3636 => x"88",
          3637 => x"7b",
          3638 => x"70",
          3639 => x"88",
          3640 => x"f8",
          3641 => x"06",
          3642 => x"5e",
          3643 => x"76",
          3644 => x"05",
          3645 => x"63",
          3646 => x"84",
          3647 => x"ed",
          3648 => x"7b",
          3649 => x"42",
          3650 => x"ff",
          3651 => x"06",
          3652 => x"88",
          3653 => x"70",
          3654 => x"71",
          3655 => x"58",
          3656 => x"f7",
          3657 => x"fa",
          3658 => x"38",
          3659 => x"7b",
          3660 => x"84",
          3661 => x"a0",
          3662 => x"80",
          3663 => x"51",
          3664 => x"08",
          3665 => x"1b",
          3666 => x"84",
          3667 => x"84",
          3668 => x"34",
          3669 => x"fc",
          3670 => x"fe",
          3671 => x"06",
          3672 => x"74",
          3673 => x"05",
          3674 => x"10",
          3675 => x"05",
          3676 => x"81",
          3677 => x"80",
          3678 => x"ff",
          3679 => x"c0",
          3680 => x"82",
          3681 => x"7f",
          3682 => x"3d",
          3683 => x"83",
          3684 => x"2b",
          3685 => x"12",
          3686 => x"07",
          3687 => x"33",
          3688 => x"43",
          3689 => x"5c",
          3690 => x"7a",
          3691 => x"08",
          3692 => x"33",
          3693 => x"74",
          3694 => x"71",
          3695 => x"41",
          3696 => x"64",
          3697 => x"34",
          3698 => x"81",
          3699 => x"ff",
          3700 => x"5a",
          3701 => x"34",
          3702 => x"11",
          3703 => x"71",
          3704 => x"81",
          3705 => x"88",
          3706 => x"45",
          3707 => x"34",
          3708 => x"33",
          3709 => x"83",
          3710 => x"83",
          3711 => x"88",
          3712 => x"55",
          3713 => x"18",
          3714 => x"82",
          3715 => x"2b",
          3716 => x"2b",
          3717 => x"05",
          3718 => x"fc",
          3719 => x"ff",
          3720 => x"ff",
          3721 => x"80",
          3722 => x"80",
          3723 => x"fe",
          3724 => x"56",
          3725 => x"34",
          3726 => x"16",
          3727 => x"b9",
          3728 => x"81",
          3729 => x"08",
          3730 => x"80",
          3731 => x"70",
          3732 => x"88",
          3733 => x"b9",
          3734 => x"b9",
          3735 => x"7f",
          3736 => x"34",
          3737 => x"fc",
          3738 => x"33",
          3739 => x"79",
          3740 => x"71",
          3741 => x"48",
          3742 => x"05",
          3743 => x"b9",
          3744 => x"85",
          3745 => x"2b",
          3746 => x"15",
          3747 => x"2a",
          3748 => x"40",
          3749 => x"87",
          3750 => x"70",
          3751 => x"07",
          3752 => x"59",
          3753 => x"81",
          3754 => x"1f",
          3755 => x"2b",
          3756 => x"33",
          3757 => x"70",
          3758 => x"05",
          3759 => x"5d",
          3760 => x"34",
          3761 => x"08",
          3762 => x"71",
          3763 => x"05",
          3764 => x"2b",
          3765 => x"2a",
          3766 => x"5b",
          3767 => x"34",
          3768 => x"b3",
          3769 => x"71",
          3770 => x"05",
          3771 => x"88",
          3772 => x"5a",
          3773 => x"79",
          3774 => x"70",
          3775 => x"71",
          3776 => x"05",
          3777 => x"88",
          3778 => x"5e",
          3779 => x"86",
          3780 => x"84",
          3781 => x"12",
          3782 => x"ff",
          3783 => x"55",
          3784 => x"84",
          3785 => x"81",
          3786 => x"2b",
          3787 => x"33",
          3788 => x"8f",
          3789 => x"2a",
          3790 => x"5e",
          3791 => x"17",
          3792 => x"70",
          3793 => x"71",
          3794 => x"81",
          3795 => x"ff",
          3796 => x"5e",
          3797 => x"34",
          3798 => x"08",
          3799 => x"33",
          3800 => x"74",
          3801 => x"71",
          3802 => x"05",
          3803 => x"88",
          3804 => x"49",
          3805 => x"57",
          3806 => x"1d",
          3807 => x"84",
          3808 => x"2b",
          3809 => x"14",
          3810 => x"07",
          3811 => x"40",
          3812 => x"7b",
          3813 => x"16",
          3814 => x"2b",
          3815 => x"2a",
          3816 => x"79",
          3817 => x"70",
          3818 => x"71",
          3819 => x"05",
          3820 => x"2b",
          3821 => x"5d",
          3822 => x"75",
          3823 => x"70",
          3824 => x"8b",
          3825 => x"82",
          3826 => x"2b",
          3827 => x"5d",
          3828 => x"34",
          3829 => x"08",
          3830 => x"33",
          3831 => x"56",
          3832 => x"7e",
          3833 => x"3f",
          3834 => x"61",
          3835 => x"06",
          3836 => x"19",
          3837 => x"71",
          3838 => x"33",
          3839 => x"70",
          3840 => x"55",
          3841 => x"85",
          3842 => x"1e",
          3843 => x"8b",
          3844 => x"86",
          3845 => x"2b",
          3846 => x"48",
          3847 => x"05",
          3848 => x"b9",
          3849 => x"33",
          3850 => x"06",
          3851 => x"78",
          3852 => x"b9",
          3853 => x"12",
          3854 => x"07",
          3855 => x"71",
          3856 => x"ff",
          3857 => x"5d",
          3858 => x"40",
          3859 => x"34",
          3860 => x"33",
          3861 => x"83",
          3862 => x"12",
          3863 => x"ff",
          3864 => x"58",
          3865 => x"78",
          3866 => x"06",
          3867 => x"54",
          3868 => x"5f",
          3869 => x"38",
          3870 => x"08",
          3871 => x"df",
          3872 => x"ef",
          3873 => x"0d",
          3874 => x"58",
          3875 => x"54",
          3876 => x"0c",
          3877 => x"d3",
          3878 => x"ba",
          3879 => x"53",
          3880 => x"fe",
          3881 => x"0c",
          3882 => x"0b",
          3883 => x"84",
          3884 => x"76",
          3885 => x"96",
          3886 => x"75",
          3887 => x"b9",
          3888 => x"81",
          3889 => x"08",
          3890 => x"87",
          3891 => x"b9",
          3892 => x"07",
          3893 => x"2a",
          3894 => x"34",
          3895 => x"22",
          3896 => x"08",
          3897 => x"15",
          3898 => x"54",
          3899 => x"cc",
          3900 => x"33",
          3901 => x"38",
          3902 => x"84",
          3903 => x"fe",
          3904 => x"83",
          3905 => x"51",
          3906 => x"81",
          3907 => x"84",
          3908 => x"12",
          3909 => x"84",
          3910 => x"7e",
          3911 => x"5a",
          3912 => x"26",
          3913 => x"54",
          3914 => x"bd",
          3915 => x"98",
          3916 => x"51",
          3917 => x"81",
          3918 => x"38",
          3919 => x"e2",
          3920 => x"fc",
          3921 => x"83",
          3922 => x"ba",
          3923 => x"80",
          3924 => x"5a",
          3925 => x"38",
          3926 => x"60",
          3927 => x"5c",
          3928 => x"87",
          3929 => x"73",
          3930 => x"38",
          3931 => x"8c",
          3932 => x"d6",
          3933 => x"ff",
          3934 => x"87",
          3935 => x"38",
          3936 => x"80",
          3937 => x"38",
          3938 => x"8c",
          3939 => x"16",
          3940 => x"55",
          3941 => x"d5",
          3942 => x"05",
          3943 => x"05",
          3944 => x"73",
          3945 => x"33",
          3946 => x"73",
          3947 => x"8c",
          3948 => x"38",
          3949 => x"2e",
          3950 => x"8c",
          3951 => x"0a",
          3952 => x"86",
          3953 => x"80",
          3954 => x"0d",
          3955 => x"8c",
          3956 => x"08",
          3957 => x"70",
          3958 => x"8c",
          3959 => x"98",
          3960 => x"72",
          3961 => x"71",
          3962 => x"ff",
          3963 => x"73",
          3964 => x"0d",
          3965 => x"71",
          3966 => x"81",
          3967 => x"83",
          3968 => x"52",
          3969 => x"84",
          3970 => x"81",
          3971 => x"3d",
          3972 => x"53",
          3973 => x"52",
          3974 => x"ba",
          3975 => x"d9",
          3976 => x"34",
          3977 => x"31",
          3978 => x"5c",
          3979 => x"9b",
          3980 => x"2e",
          3981 => x"54",
          3982 => x"33",
          3983 => x"57",
          3984 => x"fe",
          3985 => x"81",
          3986 => x"b8",
          3987 => x"80",
          3988 => x"17",
          3989 => x"84",
          3990 => x"b7",
          3991 => x"d2",
          3992 => x"ba",
          3993 => x"34",
          3994 => x"80",
          3995 => x"c1",
          3996 => x"0b",
          3997 => x"55",
          3998 => x"2a",
          3999 => x"90",
          4000 => x"74",
          4001 => x"34",
          4002 => x"19",
          4003 => x"a5",
          4004 => x"84",
          4005 => x"74",
          4006 => x"81",
          4007 => x"54",
          4008 => x"51",
          4009 => x"80",
          4010 => x"fb",
          4011 => x"2e",
          4012 => x"3d",
          4013 => x"56",
          4014 => x"08",
          4015 => x"84",
          4016 => x"ff",
          4017 => x"81",
          4018 => x"38",
          4019 => x"38",
          4020 => x"a8",
          4021 => x"b4",
          4022 => x"17",
          4023 => x"06",
          4024 => x"b8",
          4025 => x"e3",
          4026 => x"85",
          4027 => x"18",
          4028 => x"ff",
          4029 => x"70",
          4030 => x"5d",
          4031 => x"b5",
          4032 => x"5c",
          4033 => x"06",
          4034 => x"b8",
          4035 => x"93",
          4036 => x"85",
          4037 => x"18",
          4038 => x"ff",
          4039 => x"2b",
          4040 => x"2a",
          4041 => x"ae",
          4042 => x"8c",
          4043 => x"2a",
          4044 => x"08",
          4045 => x"18",
          4046 => x"2e",
          4047 => x"54",
          4048 => x"33",
          4049 => x"08",
          4050 => x"5a",
          4051 => x"38",
          4052 => x"b8",
          4053 => x"88",
          4054 => x"5b",
          4055 => x"09",
          4056 => x"2a",
          4057 => x"08",
          4058 => x"18",
          4059 => x"2e",
          4060 => x"54",
          4061 => x"33",
          4062 => x"08",
          4063 => x"5a",
          4064 => x"38",
          4065 => x"05",
          4066 => x"33",
          4067 => x"81",
          4068 => x"75",
          4069 => x"06",
          4070 => x"5e",
          4071 => x"81",
          4072 => x"70",
          4073 => x"e2",
          4074 => x"7b",
          4075 => x"84",
          4076 => x"17",
          4077 => x"8c",
          4078 => x"27",
          4079 => x"74",
          4080 => x"38",
          4081 => x"08",
          4082 => x"51",
          4083 => x"39",
          4084 => x"17",
          4085 => x"f6",
          4086 => x"2e",
          4087 => x"ba",
          4088 => x"08",
          4089 => x"18",
          4090 => x"5e",
          4091 => x"ba",
          4092 => x"54",
          4093 => x"53",
          4094 => x"3f",
          4095 => x"2e",
          4096 => x"ba",
          4097 => x"08",
          4098 => x"08",
          4099 => x"fd",
          4100 => x"82",
          4101 => x"81",
          4102 => x"05",
          4103 => x"f4",
          4104 => x"81",
          4105 => x"70",
          4106 => x"da",
          4107 => x"7d",
          4108 => x"84",
          4109 => x"17",
          4110 => x"8c",
          4111 => x"27",
          4112 => x"74",
          4113 => x"38",
          4114 => x"08",
          4115 => x"51",
          4116 => x"39",
          4117 => x"08",
          4118 => x"51",
          4119 => x"5b",
          4120 => x"f2",
          4121 => x"59",
          4122 => x"75",
          4123 => x"33",
          4124 => x"78",
          4125 => x"82",
          4126 => x"90",
          4127 => x"1a",
          4128 => x"08",
          4129 => x"38",
          4130 => x"7c",
          4131 => x"81",
          4132 => x"19",
          4133 => x"8c",
          4134 => x"81",
          4135 => x"79",
          4136 => x"06",
          4137 => x"58",
          4138 => x"2a",
          4139 => x"83",
          4140 => x"90",
          4141 => x"81",
          4142 => x"a8",
          4143 => x"1a",
          4144 => x"e1",
          4145 => x"7c",
          4146 => x"38",
          4147 => x"81",
          4148 => x"ba",
          4149 => x"58",
          4150 => x"58",
          4151 => x"83",
          4152 => x"11",
          4153 => x"7e",
          4154 => x"5c",
          4155 => x"75",
          4156 => x"79",
          4157 => x"7a",
          4158 => x"34",
          4159 => x"70",
          4160 => x"1b",
          4161 => x"b7",
          4162 => x"5e",
          4163 => x"06",
          4164 => x"b8",
          4165 => x"83",
          4166 => x"85",
          4167 => x"1a",
          4168 => x"79",
          4169 => x"1b",
          4170 => x"55",
          4171 => x"2b",
          4172 => x"71",
          4173 => x"0b",
          4174 => x"1a",
          4175 => x"08",
          4176 => x"38",
          4177 => x"53",
          4178 => x"3f",
          4179 => x"2e",
          4180 => x"ba",
          4181 => x"08",
          4182 => x"08",
          4183 => x"5c",
          4184 => x"33",
          4185 => x"81",
          4186 => x"33",
          4187 => x"08",
          4188 => x"58",
          4189 => x"38",
          4190 => x"7b",
          4191 => x"7a",
          4192 => x"71",
          4193 => x"34",
          4194 => x"39",
          4195 => x"53",
          4196 => x"3f",
          4197 => x"2e",
          4198 => x"ba",
          4199 => x"08",
          4200 => x"08",
          4201 => x"5e",
          4202 => x"19",
          4203 => x"06",
          4204 => x"53",
          4205 => x"c2",
          4206 => x"54",
          4207 => x"1a",
          4208 => x"5c",
          4209 => x"81",
          4210 => x"08",
          4211 => x"a8",
          4212 => x"ba",
          4213 => x"7e",
          4214 => x"55",
          4215 => x"e3",
          4216 => x"52",
          4217 => x"7c",
          4218 => x"53",
          4219 => x"52",
          4220 => x"ba",
          4221 => x"fb",
          4222 => x"1a",
          4223 => x"08",
          4224 => x"08",
          4225 => x"fb",
          4226 => x"82",
          4227 => x"81",
          4228 => x"19",
          4229 => x"fa",
          4230 => x"76",
          4231 => x"3f",
          4232 => x"10",
          4233 => x"ff",
          4234 => x"1f",
          4235 => x"1f",
          4236 => x"88",
          4237 => x"06",
          4238 => x"70",
          4239 => x"0a",
          4240 => x"7d",
          4241 => x"b9",
          4242 => x"ba",
          4243 => x"bb",
          4244 => x"0d",
          4245 => x"7a",
          4246 => x"76",
          4247 => x"1a",
          4248 => x"08",
          4249 => x"d7",
          4250 => x"76",
          4251 => x"76",
          4252 => x"26",
          4253 => x"f0",
          4254 => x"2e",
          4255 => x"8c",
          4256 => x"8c",
          4257 => x"80",
          4258 => x"55",
          4259 => x"09",
          4260 => x"74",
          4261 => x"04",
          4262 => x"8c",
          4263 => x"51",
          4264 => x"ba",
          4265 => x"8c",
          4266 => x"2e",
          4267 => x"8c",
          4268 => x"dd",
          4269 => x"76",
          4270 => x"79",
          4271 => x"ba",
          4272 => x"84",
          4273 => x"72",
          4274 => x"ba",
          4275 => x"73",
          4276 => x"80",
          4277 => x"81",
          4278 => x"1a",
          4279 => x"57",
          4280 => x"fe",
          4281 => x"51",
          4282 => x"84",
          4283 => x"8c",
          4284 => x"7a",
          4285 => x"75",
          4286 => x"05",
          4287 => x"26",
          4288 => x"84",
          4289 => x"1a",
          4290 => x"0c",
          4291 => x"ba",
          4292 => x"ba",
          4293 => x"80",
          4294 => x"52",
          4295 => x"8c",
          4296 => x"8c",
          4297 => x"0d",
          4298 => x"b9",
          4299 => x"3d",
          4300 => x"58",
          4301 => x"38",
          4302 => x"38",
          4303 => x"55",
          4304 => x"75",
          4305 => x"2a",
          4306 => x"56",
          4307 => x"08",
          4308 => x"98",
          4309 => x"2e",
          4310 => x"19",
          4311 => x"05",
          4312 => x"ba",
          4313 => x"0b",
          4314 => x"04",
          4315 => x"ff",
          4316 => x"2b",
          4317 => x"9c",
          4318 => x"54",
          4319 => x"38",
          4320 => x"19",
          4321 => x"0c",
          4322 => x"ec",
          4323 => x"84",
          4324 => x"81",
          4325 => x"9e",
          4326 => x"8c",
          4327 => x"76",
          4328 => x"ff",
          4329 => x"0c",
          4330 => x"7f",
          4331 => x"5c",
          4332 => x"86",
          4333 => x"17",
          4334 => x"b2",
          4335 => x"9d",
          4336 => x"58",
          4337 => x"1a",
          4338 => x"f5",
          4339 => x"18",
          4340 => x"0c",
          4341 => x"8f",
          4342 => x"8a",
          4343 => x"06",
          4344 => x"51",
          4345 => x"5d",
          4346 => x"08",
          4347 => x"8c",
          4348 => x"08",
          4349 => x"38",
          4350 => x"17",
          4351 => x"84",
          4352 => x"ba",
          4353 => x"82",
          4354 => x"ff",
          4355 => x"08",
          4356 => x"8c",
          4357 => x"80",
          4358 => x"fe",
          4359 => x"27",
          4360 => x"29",
          4361 => x"b4",
          4362 => x"78",
          4363 => x"58",
          4364 => x"74",
          4365 => x"27",
          4366 => x"53",
          4367 => x"b2",
          4368 => x"38",
          4369 => x"18",
          4370 => x"8f",
          4371 => x"08",
          4372 => x"33",
          4373 => x"8c",
          4374 => x"08",
          4375 => x"1a",
          4376 => x"27",
          4377 => x"7b",
          4378 => x"38",
          4379 => x"08",
          4380 => x"51",
          4381 => x"19",
          4382 => x"55",
          4383 => x"38",
          4384 => x"1a",
          4385 => x"75",
          4386 => x"22",
          4387 => x"98",
          4388 => x"0b",
          4389 => x"04",
          4390 => x"84",
          4391 => x"98",
          4392 => x"2e",
          4393 => x"5a",
          4394 => x"82",
          4395 => x"55",
          4396 => x"94",
          4397 => x"52",
          4398 => x"84",
          4399 => x"ff",
          4400 => x"76",
          4401 => x"08",
          4402 => x"82",
          4403 => x"70",
          4404 => x"1d",
          4405 => x"78",
          4406 => x"71",
          4407 => x"55",
          4408 => x"43",
          4409 => x"75",
          4410 => x"5d",
          4411 => x"84",
          4412 => x"08",
          4413 => x"75",
          4414 => x"0c",
          4415 => x"19",
          4416 => x"51",
          4417 => x"8c",
          4418 => x"ef",
          4419 => x"34",
          4420 => x"84",
          4421 => x"1a",
          4422 => x"33",
          4423 => x"fe",
          4424 => x"a0",
          4425 => x"19",
          4426 => x"fe",
          4427 => x"06",
          4428 => x"06",
          4429 => x"18",
          4430 => x"1f",
          4431 => x"5e",
          4432 => x"55",
          4433 => x"75",
          4434 => x"38",
          4435 => x"1d",
          4436 => x"3d",
          4437 => x"8d",
          4438 => x"81",
          4439 => x"19",
          4440 => x"07",
          4441 => x"77",
          4442 => x"f3",
          4443 => x"83",
          4444 => x"11",
          4445 => x"52",
          4446 => x"38",
          4447 => x"79",
          4448 => x"62",
          4449 => x"8c",
          4450 => x"86",
          4451 => x"2e",
          4452 => x"dd",
          4453 => x"63",
          4454 => x"5e",
          4455 => x"ff",
          4456 => x"c0",
          4457 => x"57",
          4458 => x"05",
          4459 => x"7f",
          4460 => x"59",
          4461 => x"2e",
          4462 => x"0c",
          4463 => x"0d",
          4464 => x"5c",
          4465 => x"3f",
          4466 => x"8c",
          4467 => x"40",
          4468 => x"1b",
          4469 => x"b4",
          4470 => x"83",
          4471 => x"2e",
          4472 => x"54",
          4473 => x"33",
          4474 => x"08",
          4475 => x"57",
          4476 => x"81",
          4477 => x"58",
          4478 => x"8b",
          4479 => x"06",
          4480 => x"81",
          4481 => x"2a",
          4482 => x"ef",
          4483 => x"2e",
          4484 => x"7d",
          4485 => x"75",
          4486 => x"05",
          4487 => x"ff",
          4488 => x"e4",
          4489 => x"ab",
          4490 => x"38",
          4491 => x"70",
          4492 => x"05",
          4493 => x"5a",
          4494 => x"dc",
          4495 => x"ff",
          4496 => x"52",
          4497 => x"8c",
          4498 => x"2e",
          4499 => x"0c",
          4500 => x"1b",
          4501 => x"51",
          4502 => x"8c",
          4503 => x"a4",
          4504 => x"34",
          4505 => x"84",
          4506 => x"1c",
          4507 => x"33",
          4508 => x"fd",
          4509 => x"a0",
          4510 => x"1b",
          4511 => x"fd",
          4512 => x"ab",
          4513 => x"42",
          4514 => x"2a",
          4515 => x"38",
          4516 => x"70",
          4517 => x"59",
          4518 => x"81",
          4519 => x"51",
          4520 => x"5a",
          4521 => x"d9",
          4522 => x"fe",
          4523 => x"ac",
          4524 => x"33",
          4525 => x"c7",
          4526 => x"9a",
          4527 => x"42",
          4528 => x"70",
          4529 => x"55",
          4530 => x"18",
          4531 => x"33",
          4532 => x"75",
          4533 => x"fe",
          4534 => x"a1",
          4535 => x"10",
          4536 => x"1b",
          4537 => x"84",
          4538 => x"fe",
          4539 => x"8c",
          4540 => x"70",
          4541 => x"80",
          4542 => x"38",
          4543 => x"41",
          4544 => x"81",
          4545 => x"84",
          4546 => x"0d",
          4547 => x"bc",
          4548 => x"ea",
          4549 => x"13",
          4550 => x"5e",
          4551 => x"8c",
          4552 => x"74",
          4553 => x"10",
          4554 => x"f4",
          4555 => x"8c",
          4556 => x"81",
          4557 => x"59",
          4558 => x"02",
          4559 => x"58",
          4560 => x"80",
          4561 => x"94",
          4562 => x"58",
          4563 => x"77",
          4564 => x"81",
          4565 => x"ef",
          4566 => x"7a",
          4567 => x"b8",
          4568 => x"58",
          4569 => x"81",
          4570 => x"90",
          4571 => x"60",
          4572 => x"a1",
          4573 => x"25",
          4574 => x"38",
          4575 => x"57",
          4576 => x"b9",
          4577 => x"74",
          4578 => x"84",
          4579 => x"77",
          4580 => x"7a",
          4581 => x"79",
          4582 => x"81",
          4583 => x"38",
          4584 => x"a0",
          4585 => x"16",
          4586 => x"38",
          4587 => x"19",
          4588 => x"34",
          4589 => x"51",
          4590 => x"8b",
          4591 => x"27",
          4592 => x"e4",
          4593 => x"08",
          4594 => x"09",
          4595 => x"db",
          4596 => x"02",
          4597 => x"58",
          4598 => x"5b",
          4599 => x"8c",
          4600 => x"ba",
          4601 => x"51",
          4602 => x"56",
          4603 => x"84",
          4604 => x"98",
          4605 => x"08",
          4606 => x"33",
          4607 => x"82",
          4608 => x"18",
          4609 => x"3f",
          4610 => x"38",
          4611 => x"0c",
          4612 => x"08",
          4613 => x"2e",
          4614 => x"25",
          4615 => x"81",
          4616 => x"2e",
          4617 => x"ee",
          4618 => x"84",
          4619 => x"38",
          4620 => x"38",
          4621 => x"1b",
          4622 => x"08",
          4623 => x"38",
          4624 => x"84",
          4625 => x"1c",
          4626 => x"3f",
          4627 => x"38",
          4628 => x"0c",
          4629 => x"0b",
          4630 => x"70",
          4631 => x"74",
          4632 => x"7b",
          4633 => x"57",
          4634 => x"ff",
          4635 => x"08",
          4636 => x"7c",
          4637 => x"34",
          4638 => x"98",
          4639 => x"80",
          4640 => x"fe",
          4641 => x"51",
          4642 => x"56",
          4643 => x"c7",
          4644 => x"18",
          4645 => x"51",
          4646 => x"77",
          4647 => x"84",
          4648 => x"18",
          4649 => x"a0",
          4650 => x"33",
          4651 => x"84",
          4652 => x"7f",
          4653 => x"53",
          4654 => x"ba",
          4655 => x"fe",
          4656 => x"56",
          4657 => x"81",
          4658 => x"5a",
          4659 => x"06",
          4660 => x"38",
          4661 => x"41",
          4662 => x"1c",
          4663 => x"33",
          4664 => x"82",
          4665 => x"1c",
          4666 => x"3f",
          4667 => x"38",
          4668 => x"0c",
          4669 => x"1c",
          4670 => x"06",
          4671 => x"8f",
          4672 => x"34",
          4673 => x"34",
          4674 => x"5a",
          4675 => x"8b",
          4676 => x"1b",
          4677 => x"33",
          4678 => x"05",
          4679 => x"75",
          4680 => x"57",
          4681 => x"38",
          4682 => x"38",
          4683 => x"76",
          4684 => x"34",
          4685 => x"7d",
          4686 => x"08",
          4687 => x"38",
          4688 => x"38",
          4689 => x"08",
          4690 => x"33",
          4691 => x"84",
          4692 => x"ba",
          4693 => x"08",
          4694 => x"08",
          4695 => x"fb",
          4696 => x"82",
          4697 => x"81",
          4698 => x"05",
          4699 => x"cf",
          4700 => x"76",
          4701 => x"56",
          4702 => x"fa",
          4703 => x"57",
          4704 => x"fa",
          4705 => x"fe",
          4706 => x"53",
          4707 => x"92",
          4708 => x"09",
          4709 => x"08",
          4710 => x"1d",
          4711 => x"27",
          4712 => x"82",
          4713 => x"56",
          4714 => x"58",
          4715 => x"87",
          4716 => x"81",
          4717 => x"fe",
          4718 => x"1c",
          4719 => x"52",
          4720 => x"fc",
          4721 => x"a0",
          4722 => x"18",
          4723 => x"39",
          4724 => x"40",
          4725 => x"98",
          4726 => x"ac",
          4727 => x"80",
          4728 => x"22",
          4729 => x"2e",
          4730 => x"22",
          4731 => x"95",
          4732 => x"ff",
          4733 => x"26",
          4734 => x"11",
          4735 => x"d4",
          4736 => x"30",
          4737 => x"94",
          4738 => x"80",
          4739 => x"1c",
          4740 => x"56",
          4741 => x"85",
          4742 => x"70",
          4743 => x"5b",
          4744 => x"80",
          4745 => x"05",
          4746 => x"70",
          4747 => x"8a",
          4748 => x"88",
          4749 => x"96",
          4750 => x"81",
          4751 => x"81",
          4752 => x"0b",
          4753 => x"11",
          4754 => x"89",
          4755 => x"13",
          4756 => x"9c",
          4757 => x"71",
          4758 => x"14",
          4759 => x"33",
          4760 => x"33",
          4761 => x"5f",
          4762 => x"77",
          4763 => x"16",
          4764 => x"7b",
          4765 => x"81",
          4766 => x"96",
          4767 => x"57",
          4768 => x"07",
          4769 => x"8c",
          4770 => x"ff",
          4771 => x"81",
          4772 => x"7a",
          4773 => x"05",
          4774 => x"5b",
          4775 => x"57",
          4776 => x"39",
          4777 => x"80",
          4778 => x"57",
          4779 => x"81",
          4780 => x"08",
          4781 => x"1f",
          4782 => x"fe",
          4783 => x"59",
          4784 => x"5a",
          4785 => x"1c",
          4786 => x"76",
          4787 => x"72",
          4788 => x"38",
          4789 => x"55",
          4790 => x"34",
          4791 => x"89",
          4792 => x"79",
          4793 => x"83",
          4794 => x"70",
          4795 => x"5d",
          4796 => x"0d",
          4797 => x"80",
          4798 => x"af",
          4799 => x"dc",
          4800 => x"81",
          4801 => x"0c",
          4802 => x"42",
          4803 => x"73",
          4804 => x"61",
          4805 => x"53",
          4806 => x"73",
          4807 => x"ff",
          4808 => x"56",
          4809 => x"83",
          4810 => x"30",
          4811 => x"57",
          4812 => x"74",
          4813 => x"80",
          4814 => x"0b",
          4815 => x"06",
          4816 => x"ab",
          4817 => x"16",
          4818 => x"54",
          4819 => x"06",
          4820 => x"fe",
          4821 => x"5d",
          4822 => x"70",
          4823 => x"73",
          4824 => x"39",
          4825 => x"70",
          4826 => x"55",
          4827 => x"70",
          4828 => x"72",
          4829 => x"32",
          4830 => x"51",
          4831 => x"1d",
          4832 => x"41",
          4833 => x"38",
          4834 => x"81",
          4835 => x"83",
          4836 => x"38",
          4837 => x"93",
          4838 => x"70",
          4839 => x"2e",
          4840 => x"0b",
          4841 => x"de",
          4842 => x"ba",
          4843 => x"73",
          4844 => x"25",
          4845 => x"80",
          4846 => x"62",
          4847 => x"2e",
          4848 => x"30",
          4849 => x"59",
          4850 => x"75",
          4851 => x"84",
          4852 => x"38",
          4853 => x"38",
          4854 => x"22",
          4855 => x"2a",
          4856 => x"ae",
          4857 => x"17",
          4858 => x"19",
          4859 => x"fe",
          4860 => x"ff",
          4861 => x"7a",
          4862 => x"ff",
          4863 => x"f1",
          4864 => x"19",
          4865 => x"ae",
          4866 => x"05",
          4867 => x"8f",
          4868 => x"7c",
          4869 => x"8b",
          4870 => x"70",
          4871 => x"72",
          4872 => x"78",
          4873 => x"54",
          4874 => x"74",
          4875 => x"32",
          4876 => x"54",
          4877 => x"83",
          4878 => x"83",
          4879 => x"30",
          4880 => x"07",
          4881 => x"83",
          4882 => x"38",
          4883 => x"07",
          4884 => x"56",
          4885 => x"fc",
          4886 => x"15",
          4887 => x"74",
          4888 => x"76",
          4889 => x"88",
          4890 => x"58",
          4891 => x"83",
          4892 => x"38",
          4893 => x"9d",
          4894 => x"2e",
          4895 => x"82",
          4896 => x"85",
          4897 => x"1d",
          4898 => x"ba",
          4899 => x"84",
          4900 => x"38",
          4901 => x"81",
          4902 => x"81",
          4903 => x"38",
          4904 => x"82",
          4905 => x"73",
          4906 => x"f9",
          4907 => x"11",
          4908 => x"a0",
          4909 => x"85",
          4910 => x"39",
          4911 => x"09",
          4912 => x"54",
          4913 => x"a0",
          4914 => x"23",
          4915 => x"54",
          4916 => x"73",
          4917 => x"13",
          4918 => x"a0",
          4919 => x"51",
          4920 => x"ab",
          4921 => x"08",
          4922 => x"06",
          4923 => x"33",
          4924 => x"74",
          4925 => x"08",
          4926 => x"11",
          4927 => x"2b",
          4928 => x"7d",
          4929 => x"1d",
          4930 => x"b7",
          4931 => x"fe",
          4932 => x"88",
          4933 => x"76",
          4934 => x"82",
          4935 => x"59",
          4936 => x"fd",
          4937 => x"98",
          4938 => x"88",
          4939 => x"d6",
          4940 => x"80",
          4941 => x"0d",
          4942 => x"81",
          4943 => x"1d",
          4944 => x"79",
          4945 => x"5a",
          4946 => x"83",
          4947 => x"3f",
          4948 => x"06",
          4949 => x"78",
          4950 => x"06",
          4951 => x"74",
          4952 => x"80",
          4953 => x"0b",
          4954 => x"06",
          4955 => x"e0",
          4956 => x"19",
          4957 => x"54",
          4958 => x"06",
          4959 => x"15",
          4960 => x"82",
          4961 => x"ff",
          4962 => x"38",
          4963 => x"e0",
          4964 => x"56",
          4965 => x"74",
          4966 => x"55",
          4967 => x"39",
          4968 => x"06",
          4969 => x"38",
          4970 => x"a0",
          4971 => x"81",
          4972 => x"33",
          4973 => x"71",
          4974 => x"0c",
          4975 => x"a0",
          4976 => x"74",
          4977 => x"5a",
          4978 => x"ff",
          4979 => x"33",
          4980 => x"81",
          4981 => x"74",
          4982 => x"f2",
          4983 => x"93",
          4984 => x"69",
          4985 => x"42",
          4986 => x"08",
          4987 => x"85",
          4988 => x"33",
          4989 => x"2e",
          4990 => x"ba",
          4991 => x"33",
          4992 => x"75",
          4993 => x"08",
          4994 => x"85",
          4995 => x"fe",
          4996 => x"2e",
          4997 => x"bb",
          4998 => x"ff",
          4999 => x"80",
          5000 => x"75",
          5001 => x"81",
          5002 => x"51",
          5003 => x"08",
          5004 => x"56",
          5005 => x"80",
          5006 => x"06",
          5007 => x"80",
          5008 => x"b4",
          5009 => x"54",
          5010 => x"18",
          5011 => x"84",
          5012 => x"ff",
          5013 => x"84",
          5014 => x"33",
          5015 => x"07",
          5016 => x"d5",
          5017 => x"8b",
          5018 => x"61",
          5019 => x"2e",
          5020 => x"26",
          5021 => x"80",
          5022 => x"5e",
          5023 => x"06",
          5024 => x"80",
          5025 => x"57",
          5026 => x"83",
          5027 => x"2b",
          5028 => x"70",
          5029 => x"07",
          5030 => x"75",
          5031 => x"82",
          5032 => x"11",
          5033 => x"8d",
          5034 => x"78",
          5035 => x"c5",
          5036 => x"18",
          5037 => x"c4",
          5038 => x"87",
          5039 => x"c9",
          5040 => x"40",
          5041 => x"06",
          5042 => x"38",
          5043 => x"33",
          5044 => x"a4",
          5045 => x"82",
          5046 => x"2b",
          5047 => x"88",
          5048 => x"5a",
          5049 => x"33",
          5050 => x"07",
          5051 => x"81",
          5052 => x"05",
          5053 => x"78",
          5054 => x"b4",
          5055 => x"ba",
          5056 => x"84",
          5057 => x"f5",
          5058 => x"ff",
          5059 => x"9f",
          5060 => x"82",
          5061 => x"19",
          5062 => x"7b",
          5063 => x"83",
          5064 => x"5c",
          5065 => x"38",
          5066 => x"55",
          5067 => x"19",
          5068 => x"56",
          5069 => x"8d",
          5070 => x"38",
          5071 => x"90",
          5072 => x"34",
          5073 => x"77",
          5074 => x"5d",
          5075 => x"18",
          5076 => x"0c",
          5077 => x"77",
          5078 => x"04",
          5079 => x"3d",
          5080 => x"81",
          5081 => x"26",
          5082 => x"06",
          5083 => x"87",
          5084 => x"fc",
          5085 => x"5b",
          5086 => x"70",
          5087 => x"5a",
          5088 => x"e0",
          5089 => x"ff",
          5090 => x"38",
          5091 => x"55",
          5092 => x"75",
          5093 => x"77",
          5094 => x"30",
          5095 => x"5d",
          5096 => x"38",
          5097 => x"7c",
          5098 => x"a9",
          5099 => x"77",
          5100 => x"7d",
          5101 => x"39",
          5102 => x"e9",
          5103 => x"59",
          5104 => x"80",
          5105 => x"83",
          5106 => x"a6",
          5107 => x"59",
          5108 => x"7a",
          5109 => x"33",
          5110 => x"71",
          5111 => x"70",
          5112 => x"33",
          5113 => x"40",
          5114 => x"ff",
          5115 => x"25",
          5116 => x"33",
          5117 => x"31",
          5118 => x"05",
          5119 => x"5b",
          5120 => x"80",
          5121 => x"18",
          5122 => x"55",
          5123 => x"81",
          5124 => x"17",
          5125 => x"ba",
          5126 => x"55",
          5127 => x"58",
          5128 => x"33",
          5129 => x"58",
          5130 => x"06",
          5131 => x"57",
          5132 => x"38",
          5133 => x"80",
          5134 => x"bc",
          5135 => x"82",
          5136 => x"0b",
          5137 => x"7b",
          5138 => x"81",
          5139 => x"77",
          5140 => x"84",
          5141 => x"d1",
          5142 => x"ee",
          5143 => x"7b",
          5144 => x"81",
          5145 => x"1b",
          5146 => x"80",
          5147 => x"85",
          5148 => x"40",
          5149 => x"33",
          5150 => x"71",
          5151 => x"77",
          5152 => x"2e",
          5153 => x"8d",
          5154 => x"ba",
          5155 => x"58",
          5156 => x"0b",
          5157 => x"5d",
          5158 => x"ba",
          5159 => x"0b",
          5160 => x"5a",
          5161 => x"7a",
          5162 => x"31",
          5163 => x"80",
          5164 => x"e1",
          5165 => x"e5",
          5166 => x"05",
          5167 => x"33",
          5168 => x"42",
          5169 => x"75",
          5170 => x"57",
          5171 => x"58",
          5172 => x"80",
          5173 => x"57",
          5174 => x"f9",
          5175 => x"b4",
          5176 => x"17",
          5177 => x"06",
          5178 => x"b8",
          5179 => x"b0",
          5180 => x"2e",
          5181 => x"b4",
          5182 => x"84",
          5183 => x"b6",
          5184 => x"5e",
          5185 => x"06",
          5186 => x"33",
          5187 => x"88",
          5188 => x"07",
          5189 => x"41",
          5190 => x"8b",
          5191 => x"f8",
          5192 => x"33",
          5193 => x"88",
          5194 => x"07",
          5195 => x"44",
          5196 => x"8a",
          5197 => x"f8",
          5198 => x"33",
          5199 => x"88",
          5200 => x"07",
          5201 => x"1e",
          5202 => x"33",
          5203 => x"88",
          5204 => x"07",
          5205 => x"90",
          5206 => x"45",
          5207 => x"34",
          5208 => x"7c",
          5209 => x"23",
          5210 => x"80",
          5211 => x"7b",
          5212 => x"7f",
          5213 => x"b4",
          5214 => x"81",
          5215 => x"3f",
          5216 => x"81",
          5217 => x"08",
          5218 => x"18",
          5219 => x"27",
          5220 => x"82",
          5221 => x"08",
          5222 => x"80",
          5223 => x"8a",
          5224 => x"fc",
          5225 => x"e2",
          5226 => x"5a",
          5227 => x"17",
          5228 => x"e4",
          5229 => x"71",
          5230 => x"14",
          5231 => x"33",
          5232 => x"82",
          5233 => x"f5",
          5234 => x"f9",
          5235 => x"75",
          5236 => x"77",
          5237 => x"75",
          5238 => x"39",
          5239 => x"08",
          5240 => x"51",
          5241 => x"f0",
          5242 => x"64",
          5243 => x"ff",
          5244 => x"e9",
          5245 => x"70",
          5246 => x"80",
          5247 => x"2e",
          5248 => x"54",
          5249 => x"10",
          5250 => x"55",
          5251 => x"74",
          5252 => x"38",
          5253 => x"0c",
          5254 => x"80",
          5255 => x"51",
          5256 => x"54",
          5257 => x"0d",
          5258 => x"92",
          5259 => x"70",
          5260 => x"89",
          5261 => x"ff",
          5262 => x"2e",
          5263 => x"e5",
          5264 => x"59",
          5265 => x"78",
          5266 => x"12",
          5267 => x"38",
          5268 => x"54",
          5269 => x"89",
          5270 => x"57",
          5271 => x"54",
          5272 => x"38",
          5273 => x"70",
          5274 => x"07",
          5275 => x"38",
          5276 => x"7b",
          5277 => x"98",
          5278 => x"79",
          5279 => x"3d",
          5280 => x"05",
          5281 => x"2e",
          5282 => x"9d",
          5283 => x"05",
          5284 => x"8c",
          5285 => x"2e",
          5286 => x"75",
          5287 => x"04",
          5288 => x"52",
          5289 => x"08",
          5290 => x"81",
          5291 => x"80",
          5292 => x"83",
          5293 => x"38",
          5294 => x"38",
          5295 => x"80",
          5296 => x"33",
          5297 => x"61",
          5298 => x"7d",
          5299 => x"8e",
          5300 => x"a1",
          5301 => x"91",
          5302 => x"17",
          5303 => x"9a",
          5304 => x"7d",
          5305 => x"38",
          5306 => x"80",
          5307 => x"1c",
          5308 => x"55",
          5309 => x"2e",
          5310 => x"7d",
          5311 => x"7c",
          5312 => x"26",
          5313 => x"0c",
          5314 => x"33",
          5315 => x"25",
          5316 => x"5e",
          5317 => x"82",
          5318 => x"84",
          5319 => x"91",
          5320 => x"7d",
          5321 => x"5a",
          5322 => x"81",
          5323 => x"77",
          5324 => x"08",
          5325 => x"67",
          5326 => x"88",
          5327 => x"57",
          5328 => x"7a",
          5329 => x"33",
          5330 => x"88",
          5331 => x"07",
          5332 => x"60",
          5333 => x"52",
          5334 => x"22",
          5335 => x"80",
          5336 => x"1a",
          5337 => x"74",
          5338 => x"2e",
          5339 => x"8a",
          5340 => x"5b",
          5341 => x"25",
          5342 => x"38",
          5343 => x"80",
          5344 => x"51",
          5345 => x"08",
          5346 => x"83",
          5347 => x"ff",
          5348 => x"56",
          5349 => x"91",
          5350 => x"2a",
          5351 => x"b8",
          5352 => x"ed",
          5353 => x"e5",
          5354 => x"dd",
          5355 => x"ba",
          5356 => x"76",
          5357 => x"76",
          5358 => x"95",
          5359 => x"2b",
          5360 => x"5e",
          5361 => x"7b",
          5362 => x"51",
          5363 => x"08",
          5364 => x"81",
          5365 => x"2e",
          5366 => x"ff",
          5367 => x"52",
          5368 => x"ba",
          5369 => x"08",
          5370 => x"5b",
          5371 => x"16",
          5372 => x"07",
          5373 => x"7a",
          5374 => x"39",
          5375 => x"95",
          5376 => x"33",
          5377 => x"90",
          5378 => x"80",
          5379 => x"17",
          5380 => x"cc",
          5381 => x"0b",
          5382 => x"80",
          5383 => x"17",
          5384 => x"09",
          5385 => x"39",
          5386 => x"5d",
          5387 => x"83",
          5388 => x"81",
          5389 => x"b8",
          5390 => x"a3",
          5391 => x"2e",
          5392 => x"b4",
          5393 => x"90",
          5394 => x"bc",
          5395 => x"81",
          5396 => x"70",
          5397 => x"a4",
          5398 => x"2e",
          5399 => x"ba",
          5400 => x"08",
          5401 => x"08",
          5402 => x"ff",
          5403 => x"82",
          5404 => x"81",
          5405 => x"05",
          5406 => x"ff",
          5407 => x"39",
          5408 => x"af",
          5409 => x"a2",
          5410 => x"80",
          5411 => x"9c",
          5412 => x"77",
          5413 => x"22",
          5414 => x"56",
          5415 => x"75",
          5416 => x"56",
          5417 => x"76",
          5418 => x"79",
          5419 => x"08",
          5420 => x"81",
          5421 => x"3d",
          5422 => x"5d",
          5423 => x"80",
          5424 => x"80",
          5425 => x"80",
          5426 => x"1b",
          5427 => x"b7",
          5428 => x"76",
          5429 => x"74",
          5430 => x"06",
          5431 => x"ed",
          5432 => x"71",
          5433 => x"ef",
          5434 => x"60",
          5435 => x"81",
          5436 => x"76",
          5437 => x"75",
          5438 => x"81",
          5439 => x"2e",
          5440 => x"60",
          5441 => x"1a",
          5442 => x"27",
          5443 => x"78",
          5444 => x"74",
          5445 => x"7c",
          5446 => x"83",
          5447 => x"27",
          5448 => x"54",
          5449 => x"51",
          5450 => x"08",
          5451 => x"57",
          5452 => x"19",
          5453 => x"9e",
          5454 => x"b8",
          5455 => x"05",
          5456 => x"34",
          5457 => x"89",
          5458 => x"19",
          5459 => x"1a",
          5460 => x"7b",
          5461 => x"ba",
          5462 => x"84",
          5463 => x"74",
          5464 => x"57",
          5465 => x"31",
          5466 => x"7b",
          5467 => x"2e",
          5468 => x"71",
          5469 => x"81",
          5470 => x"53",
          5471 => x"ff",
          5472 => x"80",
          5473 => x"75",
          5474 => x"60",
          5475 => x"79",
          5476 => x"77",
          5477 => x"81",
          5478 => x"59",
          5479 => x"fe",
          5480 => x"33",
          5481 => x"16",
          5482 => x"81",
          5483 => x"70",
          5484 => x"9e",
          5485 => x"08",
          5486 => x"38",
          5487 => x"b4",
          5488 => x"ba",
          5489 => x"08",
          5490 => x"55",
          5491 => x"d4",
          5492 => x"1a",
          5493 => x"33",
          5494 => x"fe",
          5495 => x"1a",
          5496 => x"08",
          5497 => x"84",
          5498 => x"81",
          5499 => x"84",
          5500 => x"fb",
          5501 => x"fb",
          5502 => x"81",
          5503 => x"0d",
          5504 => x"0b",
          5505 => x"04",
          5506 => x"40",
          5507 => x"57",
          5508 => x"56",
          5509 => x"55",
          5510 => x"22",
          5511 => x"2e",
          5512 => x"76",
          5513 => x"33",
          5514 => x"33",
          5515 => x"87",
          5516 => x"94",
          5517 => x"77",
          5518 => x"80",
          5519 => x"06",
          5520 => x"11",
          5521 => x"5a",
          5522 => x"38",
          5523 => x"84",
          5524 => x"38",
          5525 => x"98",
          5526 => x"74",
          5527 => x"08",
          5528 => x"98",
          5529 => x"fe",
          5530 => x"f0",
          5531 => x"b0",
          5532 => x"2e",
          5533 => x"2a",
          5534 => x"38",
          5535 => x"38",
          5536 => x"53",
          5537 => x"9b",
          5538 => x"a1",
          5539 => x"56",
          5540 => x"80",
          5541 => x"57",
          5542 => x"33",
          5543 => x"16",
          5544 => x"83",
          5545 => x"79",
          5546 => x"1e",
          5547 => x"1f",
          5548 => x"5e",
          5549 => x"56",
          5550 => x"38",
          5551 => x"07",
          5552 => x"75",
          5553 => x"04",
          5554 => x"0d",
          5555 => x"c8",
          5556 => x"9c",
          5557 => x"06",
          5558 => x"79",
          5559 => x"b4",
          5560 => x"0b",
          5561 => x"7f",
          5562 => x"38",
          5563 => x"81",
          5564 => x"84",
          5565 => x"ff",
          5566 => x"7b",
          5567 => x"83",
          5568 => x"7e",
          5569 => x"38",
          5570 => x"70",
          5571 => x"75",
          5572 => x"19",
          5573 => x"16",
          5574 => x"17",
          5575 => x"81",
          5576 => x"09",
          5577 => x"8c",
          5578 => x"a8",
          5579 => x"5d",
          5580 => x"f0",
          5581 => x"2e",
          5582 => x"54",
          5583 => x"53",
          5584 => x"98",
          5585 => x"94",
          5586 => x"26",
          5587 => x"81",
          5588 => x"94",
          5589 => x"1c",
          5590 => x"08",
          5591 => x"84",
          5592 => x"08",
          5593 => x"fd",
          5594 => x"ab",
          5595 => x"84",
          5596 => x"39",
          5597 => x"16",
          5598 => x"ff",
          5599 => x"81",
          5600 => x"17",
          5601 => x"31",
          5602 => x"89",
          5603 => x"2e",
          5604 => x"54",
          5605 => x"53",
          5606 => x"96",
          5607 => x"81",
          5608 => x"84",
          5609 => x"f9",
          5610 => x"f9",
          5611 => x"53",
          5612 => x"52",
          5613 => x"8c",
          5614 => x"08",
          5615 => x"17",
          5616 => x"27",
          5617 => x"77",
          5618 => x"38",
          5619 => x"08",
          5620 => x"51",
          5621 => x"12",
          5622 => x"f4",
          5623 => x"0b",
          5624 => x"04",
          5625 => x"84",
          5626 => x"f5",
          5627 => x"80",
          5628 => x"80",
          5629 => x"80",
          5630 => x"19",
          5631 => x"b5",
          5632 => x"79",
          5633 => x"86",
          5634 => x"2e",
          5635 => x"5a",
          5636 => x"38",
          5637 => x"38",
          5638 => x"81",
          5639 => x"84",
          5640 => x"ff",
          5641 => x"75",
          5642 => x"11",
          5643 => x"18",
          5644 => x"83",
          5645 => x"9a",
          5646 => x"9b",
          5647 => x"19",
          5648 => x"c1",
          5649 => x"34",
          5650 => x"34",
          5651 => x"34",
          5652 => x"34",
          5653 => x"34",
          5654 => x"0b",
          5655 => x"34",
          5656 => x"81",
          5657 => x"96",
          5658 => x"19",
          5659 => x"90",
          5660 => x"8d",
          5661 => x"08",
          5662 => x"33",
          5663 => x"56",
          5664 => x"84",
          5665 => x"17",
          5666 => x"8c",
          5667 => x"27",
          5668 => x"74",
          5669 => x"38",
          5670 => x"08",
          5671 => x"51",
          5672 => x"e8",
          5673 => x"18",
          5674 => x"18",
          5675 => x"34",
          5676 => x"34",
          5677 => x"34",
          5678 => x"34",
          5679 => x"34",
          5680 => x"0b",
          5681 => x"34",
          5682 => x"81",
          5683 => x"94",
          5684 => x"19",
          5685 => x"90",
          5686 => x"33",
          5687 => x"8c",
          5688 => x"38",
          5689 => x"39",
          5690 => x"fb",
          5691 => x"84",
          5692 => x"74",
          5693 => x"72",
          5694 => x"71",
          5695 => x"84",
          5696 => x"96",
          5697 => x"75",
          5698 => x"ba",
          5699 => x"13",
          5700 => x"ba",
          5701 => x"38",
          5702 => x"f6",
          5703 => x"5b",
          5704 => x"81",
          5705 => x"52",
          5706 => x"38",
          5707 => x"e8",
          5708 => x"70",
          5709 => x"ba",
          5710 => x"0b",
          5711 => x"04",
          5712 => x"06",
          5713 => x"38",
          5714 => x"05",
          5715 => x"38",
          5716 => x"79",
          5717 => x"05",
          5718 => x"33",
          5719 => x"99",
          5720 => x"ff",
          5721 => x"70",
          5722 => x"81",
          5723 => x"9f",
          5724 => x"81",
          5725 => x"74",
          5726 => x"9f",
          5727 => x"80",
          5728 => x"5b",
          5729 => x"7a",
          5730 => x"f7",
          5731 => x"39",
          5732 => x"cc",
          5733 => x"3f",
          5734 => x"8c",
          5735 => x"ba",
          5736 => x"5c",
          5737 => x"c5",
          5738 => x"84",
          5739 => x"80",
          5740 => x"5a",
          5741 => x"b2",
          5742 => x"57",
          5743 => x"63",
          5744 => x"88",
          5745 => x"57",
          5746 => x"98",
          5747 => x"98",
          5748 => x"84",
          5749 => x"85",
          5750 => x"0d",
          5751 => x"71",
          5752 => x"07",
          5753 => x"7a",
          5754 => x"ba",
          5755 => x"9e",
          5756 => x"e6",
          5757 => x"80",
          5758 => x"52",
          5759 => x"84",
          5760 => x"08",
          5761 => x"0c",
          5762 => x"3d",
          5763 => x"58",
          5764 => x"d8",
          5765 => x"7a",
          5766 => x"8c",
          5767 => x"92",
          5768 => x"56",
          5769 => x"84",
          5770 => x"5d",
          5771 => x"53",
          5772 => x"ff",
          5773 => x"80",
          5774 => x"76",
          5775 => x"80",
          5776 => x"12",
          5777 => x"33",
          5778 => x"2e",
          5779 => x"0c",
          5780 => x"3f",
          5781 => x"8c",
          5782 => x"51",
          5783 => x"08",
          5784 => x"80",
          5785 => x"12",
          5786 => x"33",
          5787 => x"2e",
          5788 => x"38",
          5789 => x"ff",
          5790 => x"59",
          5791 => x"b4",
          5792 => x"78",
          5793 => x"b8",
          5794 => x"3f",
          5795 => x"79",
          5796 => x"81",
          5797 => x"57",
          5798 => x"78",
          5799 => x"9c",
          5800 => x"18",
          5801 => x"ff",
          5802 => x"75",
          5803 => x"e6",
          5804 => x"34",
          5805 => x"bd",
          5806 => x"80",
          5807 => x"10",
          5808 => x"33",
          5809 => x"2e",
          5810 => x"33",
          5811 => x"1a",
          5812 => x"57",
          5813 => x"5f",
          5814 => x"34",
          5815 => x"38",
          5816 => x"76",
          5817 => x"38",
          5818 => x"ba",
          5819 => x"95",
          5820 => x"2b",
          5821 => x"56",
          5822 => x"94",
          5823 => x"2b",
          5824 => x"5a",
          5825 => x"ce",
          5826 => x"ba",
          5827 => x"ff",
          5828 => x"53",
          5829 => x"52",
          5830 => x"84",
          5831 => x"ba",
          5832 => x"08",
          5833 => x"08",
          5834 => x"fc",
          5835 => x"82",
          5836 => x"81",
          5837 => x"05",
          5838 => x"ff",
          5839 => x"39",
          5840 => x"5c",
          5841 => x"d1",
          5842 => x"fc",
          5843 => x"59",
          5844 => x"06",
          5845 => x"e5",
          5846 => x"79",
          5847 => x"77",
          5848 => x"3d",
          5849 => x"33",
          5850 => x"78",
          5851 => x"59",
          5852 => x"0c",
          5853 => x"0d",
          5854 => x"80",
          5855 => x"80",
          5856 => x"80",
          5857 => x"16",
          5858 => x"a0",
          5859 => x"75",
          5860 => x"72",
          5861 => x"76",
          5862 => x"08",
          5863 => x"cc",
          5864 => x"2b",
          5865 => x"f7",
          5866 => x"ba",
          5867 => x"15",
          5868 => x"ba",
          5869 => x"26",
          5870 => x"70",
          5871 => x"17",
          5872 => x"82",
          5873 => x"38",
          5874 => x"94",
          5875 => x"2a",
          5876 => x"2e",
          5877 => x"ff",
          5878 => x"54",
          5879 => x"a3",
          5880 => x"74",
          5881 => x"9c",
          5882 => x"98",
          5883 => x"91",
          5884 => x"8c",
          5885 => x"33",
          5886 => x"73",
          5887 => x"55",
          5888 => x"81",
          5889 => x"0c",
          5890 => x"90",
          5891 => x"33",
          5892 => x"34",
          5893 => x"2e",
          5894 => x"85",
          5895 => x"84",
          5896 => x"80",
          5897 => x"54",
          5898 => x"98",
          5899 => x"38",
          5900 => x"57",
          5901 => x"76",
          5902 => x"a9",
          5903 => x"fe",
          5904 => x"80",
          5905 => x"29",
          5906 => x"11",
          5907 => x"df",
          5908 => x"39",
          5909 => x"3f",
          5910 => x"39",
          5911 => x"3f",
          5912 => x"72",
          5913 => x"56",
          5914 => x"ff",
          5915 => x"54",
          5916 => x"38",
          5917 => x"ed",
          5918 => x"0c",
          5919 => x"82",
          5920 => x"ba",
          5921 => x"3d",
          5922 => x"2e",
          5923 => x"05",
          5924 => x"9b",
          5925 => x"ba",
          5926 => x"76",
          5927 => x"0c",
          5928 => x"7d",
          5929 => x"84",
          5930 => x"08",
          5931 => x"98",
          5932 => x"38",
          5933 => x"06",
          5934 => x"38",
          5935 => x"12",
          5936 => x"33",
          5937 => x"2e",
          5938 => x"58",
          5939 => x"52",
          5940 => x"ba",
          5941 => x"38",
          5942 => x"76",
          5943 => x"76",
          5944 => x"94",
          5945 => x"2b",
          5946 => x"5a",
          5947 => x"55",
          5948 => x"74",
          5949 => x"72",
          5950 => x"86",
          5951 => x"71",
          5952 => x"57",
          5953 => x"84",
          5954 => x"81",
          5955 => x"84",
          5956 => x"dc",
          5957 => x"39",
          5958 => x"89",
          5959 => x"08",
          5960 => x"33",
          5961 => x"14",
          5962 => x"78",
          5963 => x"59",
          5964 => x"80",
          5965 => x"51",
          5966 => x"08",
          5967 => x"b5",
          5968 => x"76",
          5969 => x"72",
          5970 => x"84",
          5971 => x"70",
          5972 => x"08",
          5973 => x"8c",
          5974 => x"53",
          5975 => x"72",
          5976 => x"84",
          5977 => x"70",
          5978 => x"08",
          5979 => x"52",
          5980 => x"ba",
          5981 => x"3d",
          5982 => x"fd",
          5983 => x"06",
          5984 => x"08",
          5985 => x"0d",
          5986 => x"53",
          5987 => x"84",
          5988 => x"08",
          5989 => x"8c",
          5990 => x"75",
          5991 => x"8c",
          5992 => x"38",
          5993 => x"2b",
          5994 => x"76",
          5995 => x"51",
          5996 => x"8c",
          5997 => x"84",
          5998 => x"ed",
          5999 => x"53",
          6000 => x"51",
          6001 => x"5a",
          6002 => x"75",
          6003 => x"11",
          6004 => x"75",
          6005 => x"79",
          6006 => x"04",
          6007 => x"5b",
          6008 => x"a8",
          6009 => x"5d",
          6010 => x"1d",
          6011 => x"76",
          6012 => x"78",
          6013 => x"54",
          6014 => x"33",
          6015 => x"8c",
          6016 => x"81",
          6017 => x"5b",
          6018 => x"5e",
          6019 => x"17",
          6020 => x"33",
          6021 => x"81",
          6022 => x"75",
          6023 => x"06",
          6024 => x"05",
          6025 => x"ff",
          6026 => x"53",
          6027 => x"38",
          6028 => x"84",
          6029 => x"18",
          6030 => x"3d",
          6031 => x"53",
          6032 => x"52",
          6033 => x"84",
          6034 => x"ba",
          6035 => x"08",
          6036 => x"08",
          6037 => x"fe",
          6038 => x"82",
          6039 => x"81",
          6040 => x"05",
          6041 => x"fe",
          6042 => x"39",
          6043 => x"75",
          6044 => x"84",
          6045 => x"38",
          6046 => x"f7",
          6047 => x"84",
          6048 => x"05",
          6049 => x"9c",
          6050 => x"7f",
          6051 => x"33",
          6052 => x"fe",
          6053 => x"11",
          6054 => x"70",
          6055 => x"83",
          6056 => x"59",
          6057 => x"fe",
          6058 => x"81",
          6059 => x"94",
          6060 => x"58",
          6061 => x"82",
          6062 => x"0d",
          6063 => x"9f",
          6064 => x"97",
          6065 => x"8f",
          6066 => x"59",
          6067 => x"80",
          6068 => x"91",
          6069 => x"90",
          6070 => x"55",
          6071 => x"c4",
          6072 => x"18",
          6073 => x"38",
          6074 => x"81",
          6075 => x"74",
          6076 => x"88",
          6077 => x"0c",
          6078 => x"18",
          6079 => x"91",
          6080 => x"8c",
          6081 => x"78",
          6082 => x"76",
          6083 => x"8c",
          6084 => x"2e",
          6085 => x"81",
          6086 => x"08",
          6087 => x"73",
          6088 => x"84",
          6089 => x"16",
          6090 => x"55",
          6091 => x"81",
          6092 => x"81",
          6093 => x"54",
          6094 => x"39",
          6095 => x"3f",
          6096 => x"73",
          6097 => x"56",
          6098 => x"33",
          6099 => x"18",
          6100 => x"52",
          6101 => x"ba",
          6102 => x"84",
          6103 => x"38",
          6104 => x"ba",
          6105 => x"a1",
          6106 => x"08",
          6107 => x"84",
          6108 => x"84",
          6109 => x"81",
          6110 => x"ff",
          6111 => x"c7",
          6112 => x"ba",
          6113 => x"76",
          6114 => x"8c",
          6115 => x"2e",
          6116 => x"81",
          6117 => x"08",
          6118 => x"73",
          6119 => x"84",
          6120 => x"16",
          6121 => x"55",
          6122 => x"15",
          6123 => x"07",
          6124 => x"77",
          6125 => x"74",
          6126 => x"39",
          6127 => x"90",
          6128 => x"82",
          6129 => x"33",
          6130 => x"8c",
          6131 => x"fa",
          6132 => x"54",
          6133 => x"56",
          6134 => x"db",
          6135 => x"9c",
          6136 => x"fb",
          6137 => x"ba",
          6138 => x"84",
          6139 => x"7d",
          6140 => x"70",
          6141 => x"ba",
          6142 => x"de",
          6143 => x"85",
          6144 => x"77",
          6145 => x"7b",
          6146 => x"33",
          6147 => x"7b",
          6148 => x"9b",
          6149 => x"2b",
          6150 => x"58",
          6151 => x"84",
          6152 => x"80",
          6153 => x"7b",
          6154 => x"41",
          6155 => x"70",
          6156 => x"ba",
          6157 => x"fe",
          6158 => x"74",
          6159 => x"8c",
          6160 => x"38",
          6161 => x"3d",
          6162 => x"33",
          6163 => x"7d",
          6164 => x"84",
          6165 => x"84",
          6166 => x"08",
          6167 => x"74",
          6168 => x"78",
          6169 => x"8c",
          6170 => x"2e",
          6171 => x"80",
          6172 => x"38",
          6173 => x"08",
          6174 => x"9c",
          6175 => x"82",
          6176 => x"fe",
          6177 => x"84",
          6178 => x"b8",
          6179 => x"5a",
          6180 => x"38",
          6181 => x"7a",
          6182 => x"81",
          6183 => x"17",
          6184 => x"ba",
          6185 => x"56",
          6186 => x"56",
          6187 => x"e5",
          6188 => x"90",
          6189 => x"80",
          6190 => x"84",
          6191 => x"08",
          6192 => x"2e",
          6193 => x"56",
          6194 => x"08",
          6195 => x"fe",
          6196 => x"8c",
          6197 => x"a6",
          6198 => x"34",
          6199 => x"84",
          6200 => x"18",
          6201 => x"33",
          6202 => x"fe",
          6203 => x"a0",
          6204 => x"17",
          6205 => x"58",
          6206 => x"27",
          6207 => x"fe",
          6208 => x"5a",
          6209 => x"cb",
          6210 => x"fd",
          6211 => x"2e",
          6212 => x"76",
          6213 => x"8c",
          6214 => x"11",
          6215 => x"7b",
          6216 => x"18",
          6217 => x"7b",
          6218 => x"26",
          6219 => x"39",
          6220 => x"8c",
          6221 => x"fd",
          6222 => x"9f",
          6223 => x"51",
          6224 => x"08",
          6225 => x"8a",
          6226 => x"3d",
          6227 => x"3d",
          6228 => x"84",
          6229 => x"08",
          6230 => x"0c",
          6231 => x"08",
          6232 => x"02",
          6233 => x"81",
          6234 => x"b9",
          6235 => x"70",
          6236 => x"ba",
          6237 => x"8c",
          6238 => x"8c",
          6239 => x"ba",
          6240 => x"75",
          6241 => x"08",
          6242 => x"80",
          6243 => x"fe",
          6244 => x"27",
          6245 => x"29",
          6246 => x"b4",
          6247 => x"79",
          6248 => x"58",
          6249 => x"74",
          6250 => x"27",
          6251 => x"53",
          6252 => x"ee",
          6253 => x"df",
          6254 => x"56",
          6255 => x"08",
          6256 => x"33",
          6257 => x"56",
          6258 => x"ba",
          6259 => x"08",
          6260 => x"18",
          6261 => x"33",
          6262 => x"fe",
          6263 => x"a0",
          6264 => x"17",
          6265 => x"ca",
          6266 => x"55",
          6267 => x"9c",
          6268 => x"52",
          6269 => x"ba",
          6270 => x"80",
          6271 => x"08",
          6272 => x"8c",
          6273 => x"53",
          6274 => x"3f",
          6275 => x"9c",
          6276 => x"5a",
          6277 => x"81",
          6278 => x"81",
          6279 => x"55",
          6280 => x"84",
          6281 => x"8a",
          6282 => x"06",
          6283 => x"81",
          6284 => x"1f",
          6285 => x"57",
          6286 => x"7d",
          6287 => x"58",
          6288 => x"59",
          6289 => x"cf",
          6290 => x"34",
          6291 => x"7d",
          6292 => x"77",
          6293 => x"5b",
          6294 => x"55",
          6295 => x"59",
          6296 => x"57",
          6297 => x"33",
          6298 => x"16",
          6299 => x"0b",
          6300 => x"83",
          6301 => x"80",
          6302 => x"7a",
          6303 => x"74",
          6304 => x"81",
          6305 => x"92",
          6306 => x"84",
          6307 => x"56",
          6308 => x"84",
          6309 => x"0b",
          6310 => x"17",
          6311 => x"18",
          6312 => x"18",
          6313 => x"80",
          6314 => x"16",
          6315 => x"34",
          6316 => x"ba",
          6317 => x"0c",
          6318 => x"55",
          6319 => x"2a",
          6320 => x"fd",
          6321 => x"cc",
          6322 => x"80",
          6323 => x"80",
          6324 => x"fe",
          6325 => x"94",
          6326 => x"95",
          6327 => x"16",
          6328 => x"34",
          6329 => x"ba",
          6330 => x"3d",
          6331 => x"59",
          6332 => x"79",
          6333 => x"26",
          6334 => x"38",
          6335 => x"af",
          6336 => x"05",
          6337 => x"3f",
          6338 => x"8c",
          6339 => x"ba",
          6340 => x"a6",
          6341 => x"3d",
          6342 => x"84",
          6343 => x"08",
          6344 => x"81",
          6345 => x"38",
          6346 => x"58",
          6347 => x"33",
          6348 => x"15",
          6349 => x"b0",
          6350 => x"81",
          6351 => x"59",
          6352 => x"b3",
          6353 => x"d5",
          6354 => x"ba",
          6355 => x"3d",
          6356 => x"84",
          6357 => x"76",
          6358 => x"57",
          6359 => x"82",
          6360 => x"5d",
          6361 => x"80",
          6362 => x"72",
          6363 => x"81",
          6364 => x"5b",
          6365 => x"77",
          6366 => x"81",
          6367 => x"58",
          6368 => x"70",
          6369 => x"70",
          6370 => x"09",
          6371 => x"38",
          6372 => x"07",
          6373 => x"7a",
          6374 => x"1e",
          6375 => x"38",
          6376 => x"39",
          6377 => x"7f",
          6378 => x"05",
          6379 => x"3f",
          6380 => x"8c",
          6381 => x"6c",
          6382 => x"fe",
          6383 => x"3f",
          6384 => x"8c",
          6385 => x"0b",
          6386 => x"05",
          6387 => x"57",
          6388 => x"ff",
          6389 => x"cb",
          6390 => x"33",
          6391 => x"7e",
          6392 => x"8b",
          6393 => x"1e",
          6394 => x"81",
          6395 => x"c5",
          6396 => x"bd",
          6397 => x"33",
          6398 => x"58",
          6399 => x"38",
          6400 => x"5e",
          6401 => x"8a",
          6402 => x"08",
          6403 => x"b5",
          6404 => x"08",
          6405 => x"5f",
          6406 => x"53",
          6407 => x"fe",
          6408 => x"80",
          6409 => x"77",
          6410 => x"d8",
          6411 => x"81",
          6412 => x"81",
          6413 => x"ff",
          6414 => x"34",
          6415 => x"18",
          6416 => x"09",
          6417 => x"5e",
          6418 => x"2a",
          6419 => x"57",
          6420 => x"aa",
          6421 => x"56",
          6422 => x"78",
          6423 => x"8c",
          6424 => x"f5",
          6425 => x"57",
          6426 => x"b4",
          6427 => x"7e",
          6428 => x"38",
          6429 => x"81",
          6430 => x"84",
          6431 => x"ff",
          6432 => x"77",
          6433 => x"5a",
          6434 => x"34",
          6435 => x"80",
          6436 => x"84",
          6437 => x"08",
          6438 => x"74",
          6439 => x"74",
          6440 => x"9d",
          6441 => x"8c",
          6442 => x"84",
          6443 => x"95",
          6444 => x"2b",
          6445 => x"56",
          6446 => x"08",
          6447 => x"8c",
          6448 => x"84",
          6449 => x"81",
          6450 => x"81",
          6451 => x"81",
          6452 => x"09",
          6453 => x"8c",
          6454 => x"a8",
          6455 => x"59",
          6456 => x"a0",
          6457 => x"2e",
          6458 => x"54",
          6459 => x"53",
          6460 => x"e1",
          6461 => x"81",
          6462 => x"70",
          6463 => x"e1",
          6464 => x"08",
          6465 => x"83",
          6466 => x"08",
          6467 => x"74",
          6468 => x"82",
          6469 => x"81",
          6470 => x"17",
          6471 => x"52",
          6472 => x"3f",
          6473 => x"0d",
          6474 => x"05",
          6475 => x"53",
          6476 => x"51",
          6477 => x"08",
          6478 => x"8a",
          6479 => x"3d",
          6480 => x"3d",
          6481 => x"84",
          6482 => x"08",
          6483 => x"81",
          6484 => x"38",
          6485 => x"12",
          6486 => x"51",
          6487 => x"78",
          6488 => x"51",
          6489 => x"08",
          6490 => x"04",
          6491 => x"96",
          6492 => x"ff",
          6493 => x"55",
          6494 => x"38",
          6495 => x"0d",
          6496 => x"d0",
          6497 => x"ba",
          6498 => x"e0",
          6499 => x"a0",
          6500 => x"60",
          6501 => x"90",
          6502 => x"17",
          6503 => x"17",
          6504 => x"17",
          6505 => x"17",
          6506 => x"34",
          6507 => x"ba",
          6508 => x"3d",
          6509 => x"5d",
          6510 => x"52",
          6511 => x"84",
          6512 => x"30",
          6513 => x"25",
          6514 => x"38",
          6515 => x"81",
          6516 => x"80",
          6517 => x"8c",
          6518 => x"78",
          6519 => x"11",
          6520 => x"08",
          6521 => x"33",
          6522 => x"81",
          6523 => x"53",
          6524 => x"fe",
          6525 => x"80",
          6526 => x"76",
          6527 => x"38",
          6528 => x"56",
          6529 => x"56",
          6530 => x"75",
          6531 => x"12",
          6532 => x"07",
          6533 => x"2b",
          6534 => x"5d",
          6535 => x"8c",
          6536 => x"80",
          6537 => x"55",
          6538 => x"08",
          6539 => x"81",
          6540 => x"06",
          6541 => x"57",
          6542 => x"08",
          6543 => x"33",
          6544 => x"59",
          6545 => x"81",
          6546 => x"08",
          6547 => x"17",
          6548 => x"55",
          6549 => x"38",
          6550 => x"09",
          6551 => x"b4",
          6552 => x"7a",
          6553 => x"e2",
          6554 => x"b8",
          6555 => x"da",
          6556 => x"2e",
          6557 => x"52",
          6558 => x"ba",
          6559 => x"fe",
          6560 => x"ba",
          6561 => x"18",
          6562 => x"75",
          6563 => x"78",
          6564 => x"58",
          6565 => x"f2",
          6566 => x"5c",
          6567 => x"fc",
          6568 => x"e1",
          6569 => x"b4",
          6570 => x"eb",
          6571 => x"ba",
          6572 => x"5d",
          6573 => x"81",
          6574 => x"f4",
          6575 => x"70",
          6576 => x"9f",
          6577 => x"90",
          6578 => x"81",
          6579 => x"75",
          6580 => x"81",
          6581 => x"83",
          6582 => x"9f",
          6583 => x"ff",
          6584 => x"e0",
          6585 => x"9c",
          6586 => x"58",
          6587 => x"56",
          6588 => x"70",
          6589 => x"58",
          6590 => x"2e",
          6591 => x"ff",
          6592 => x"ff",
          6593 => x"26",
          6594 => x"8f",
          6595 => x"70",
          6596 => x"76",
          6597 => x"1a",
          6598 => x"ff",
          6599 => x"26",
          6600 => x"86",
          6601 => x"79",
          6602 => x"56",
          6603 => x"a0",
          6604 => x"1a",
          6605 => x"47",
          6606 => x"fe",
          6607 => x"55",
          6608 => x"38",
          6609 => x"a1",
          6610 => x"51",
          6611 => x"83",
          6612 => x"38",
          6613 => x"a1",
          6614 => x"56",
          6615 => x"fe",
          6616 => x"55",
          6617 => x"79",
          6618 => x"7e",
          6619 => x"58",
          6620 => x"ff",
          6621 => x"81",
          6622 => x"d9",
          6623 => x"74",
          6624 => x"fe",
          6625 => x"84",
          6626 => x"06",
          6627 => x"2e",
          6628 => x"76",
          6629 => x"ba",
          6630 => x"75",
          6631 => x"84",
          6632 => x"98",
          6633 => x"08",
          6634 => x"55",
          6635 => x"d7",
          6636 => x"52",
          6637 => x"3f",
          6638 => x"38",
          6639 => x"0c",
          6640 => x"17",
          6641 => x"81",
          6642 => x"70",
          6643 => x"80",
          6644 => x"79",
          6645 => x"51",
          6646 => x"08",
          6647 => x"ff",
          6648 => x"fd",
          6649 => x"38",
          6650 => x"81",
          6651 => x"f4",
          6652 => x"34",
          6653 => x"70",
          6654 => x"05",
          6655 => x"2e",
          6656 => x"58",
          6657 => x"ff",
          6658 => x"39",
          6659 => x"81",
          6660 => x"d7",
          6661 => x"fd",
          6662 => x"81",
          6663 => x"81",
          6664 => x"84",
          6665 => x"06",
          6666 => x"83",
          6667 => x"08",
          6668 => x"8a",
          6669 => x"2e",
          6670 => x"fd",
          6671 => x"51",
          6672 => x"08",
          6673 => x"fd",
          6674 => x"58",
          6675 => x"fe",
          6676 => x"a0",
          6677 => x"18",
          6678 => x"a9",
          6679 => x"88",
          6680 => x"57",
          6681 => x"76",
          6682 => x"74",
          6683 => x"86",
          6684 => x"78",
          6685 => x"73",
          6686 => x"33",
          6687 => x"2e",
          6688 => x"9c",
          6689 => x"81",
          6690 => x"8c",
          6691 => x"2b",
          6692 => x"fd",
          6693 => x"70",
          6694 => x"ba",
          6695 => x"42",
          6696 => x"88",
          6697 => x"38",
          6698 => x"59",
          6699 => x"3f",
          6700 => x"08",
          6701 => x"ba",
          6702 => x"84",
          6703 => x"38",
          6704 => x"81",
          6705 => x"74",
          6706 => x"87",
          6707 => x"0c",
          6708 => x"ba",
          6709 => x"15",
          6710 => x"ba",
          6711 => x"ad",
          6712 => x"a7",
          6713 => x"7a",
          6714 => x"38",
          6715 => x"e6",
          6716 => x"fe",
          6717 => x"56",
          6718 => x"77",
          6719 => x"74",
          6720 => x"55",
          6721 => x"88",
          6722 => x"17",
          6723 => x"18",
          6724 => x"16",
          6725 => x"e9",
          6726 => x"84",
          6727 => x"16",
          6728 => x"54",
          6729 => x"fe",
          6730 => x"81",
          6731 => x"ff",
          6732 => x"3d",
          6733 => x"02",
          6734 => x"42",
          6735 => x"5f",
          6736 => x"38",
          6737 => x"9f",
          6738 => x"9b",
          6739 => x"85",
          6740 => x"80",
          6741 => x"10",
          6742 => x"5a",
          6743 => x"34",
          6744 => x"84",
          6745 => x"81",
          6746 => x"84",
          6747 => x"81",
          6748 => x"ab",
          6749 => x"8a",
          6750 => x"fc",
          6751 => x"d0",
          6752 => x"98",
          6753 => x"90",
          6754 => x"88",
          6755 => x"83",
          6756 => x"84",
          6757 => x"81",
          6758 => x"1f",
          6759 => x"7e",
          6760 => x"70",
          6761 => x"60",
          6762 => x"70",
          6763 => x"57",
          6764 => x"84",
          6765 => x"52",
          6766 => x"57",
          6767 => x"60",
          6768 => x"05",
          6769 => x"8e",
          6770 => x"81",
          6771 => x"61",
          6772 => x"62",
          6773 => x"18",
          6774 => x"90",
          6775 => x"33",
          6776 => x"71",
          6777 => x"82",
          6778 => x"2b",
          6779 => x"88",
          6780 => x"3d",
          6781 => x"0c",
          6782 => x"5a",
          6783 => x"79",
          6784 => x"81",
          6785 => x"2a",
          6786 => x"2e",
          6787 => x"64",
          6788 => x"47",
          6789 => x"30",
          6790 => x"2e",
          6791 => x"8c",
          6792 => x"22",
          6793 => x"74",
          6794 => x"56",
          6795 => x"57",
          6796 => x"75",
          6797 => x"fd",
          6798 => x"10",
          6799 => x"9f",
          6800 => x"ba",
          6801 => x"05",
          6802 => x"4c",
          6803 => x"81",
          6804 => x"68",
          6805 => x"06",
          6806 => x"83",
          6807 => x"77",
          6808 => x"57",
          6809 => x"7c",
          6810 => x"31",
          6811 => x"ba",
          6812 => x"f6",
          6813 => x"82",
          6814 => x"ba",
          6815 => x"89",
          6816 => x"c0",
          6817 => x"a3",
          6818 => x"0c",
          6819 => x"04",
          6820 => x"84",
          6821 => x"ba",
          6822 => x"70",
          6823 => x"89",
          6824 => x"ff",
          6825 => x"2e",
          6826 => x"fc",
          6827 => x"7a",
          6828 => x"81",
          6829 => x"59",
          6830 => x"17",
          6831 => x"9f",
          6832 => x"e0",
          6833 => x"76",
          6834 => x"78",
          6835 => x"ff",
          6836 => x"70",
          6837 => x"4a",
          6838 => x"81",
          6839 => x"25",
          6840 => x"39",
          6841 => x"79",
          6842 => x"84",
          6843 => x"83",
          6844 => x"40",
          6845 => x"55",
          6846 => x"38",
          6847 => x"81",
          6848 => x"ff",
          6849 => x"56",
          6850 => x"93",
          6851 => x"82",
          6852 => x"8b",
          6853 => x"26",
          6854 => x"5b",
          6855 => x"8e",
          6856 => x"3d",
          6857 => x"55",
          6858 => x"f5",
          6859 => x"5b",
          6860 => x"80",
          6861 => x"05",
          6862 => x"38",
          6863 => x"55",
          6864 => x"70",
          6865 => x"74",
          6866 => x"65",
          6867 => x"61",
          6868 => x"06",
          6869 => x"88",
          6870 => x"81",
          6871 => x"70",
          6872 => x"34",
          6873 => x"61",
          6874 => x"ff",
          6875 => x"ff",
          6876 => x"34",
          6877 => x"05",
          6878 => x"61",
          6879 => x"34",
          6880 => x"9b",
          6881 => x"7e",
          6882 => x"34",
          6883 => x"05",
          6884 => x"0c",
          6885 => x"34",
          6886 => x"61",
          6887 => x"34",
          6888 => x"61",
          6889 => x"06",
          6890 => x"88",
          6891 => x"ff",
          6892 => x"a6",
          6893 => x"e5",
          6894 => x"05",
          6895 => x"34",
          6896 => x"83",
          6897 => x"60",
          6898 => x"34",
          6899 => x"51",
          6900 => x"ba",
          6901 => x"5c",
          6902 => x"61",
          6903 => x"58",
          6904 => x"63",
          6905 => x"c0",
          6906 => x"81",
          6907 => x"34",
          6908 => x"64",
          6909 => x"2a",
          6910 => x"34",
          6911 => x"7c",
          6912 => x"38",
          6913 => x"52",
          6914 => x"ba",
          6915 => x"61",
          6916 => x"58",
          6917 => x"78",
          6918 => x"c9",
          6919 => x"2e",
          6920 => x"2e",
          6921 => x"66",
          6922 => x"7a",
          6923 => x"d2",
          6924 => x"38",
          6925 => x"75",
          6926 => x"93",
          6927 => x"26",
          6928 => x"83",
          6929 => x"61",
          6930 => x"b3",
          6931 => x"75",
          6932 => x"59",
          6933 => x"ff",
          6934 => x"47",
          6935 => x"34",
          6936 => x"83",
          6937 => x"6c",
          6938 => x"51",
          6939 => x"05",
          6940 => x"bf",
          6941 => x"84",
          6942 => x"7e",
          6943 => x"83",
          6944 => x"05",
          6945 => x"c9",
          6946 => x"34",
          6947 => x"cb",
          6948 => x"61",
          6949 => x"5f",
          6950 => x"54",
          6951 => x"c2",
          6952 => x"08",
          6953 => x"79",
          6954 => x"84",
          6955 => x"ba",
          6956 => x"3d",
          6957 => x"55",
          6958 => x"45",
          6959 => x"78",
          6960 => x"c0",
          6961 => x"38",
          6962 => x"c0",
          6963 => x"57",
          6964 => x"76",
          6965 => x"51",
          6966 => x"08",
          6967 => x"2a",
          6968 => x"ba",
          6969 => x"47",
          6970 => x"cb",
          6971 => x"ba",
          6972 => x"e6",
          6973 => x"2a",
          6974 => x"f8",
          6975 => x"80",
          6976 => x"ab",
          6977 => x"88",
          6978 => x"75",
          6979 => x"34",
          6980 => x"05",
          6981 => x"c3",
          6982 => x"34",
          6983 => x"cc",
          6984 => x"a4",
          6985 => x"61",
          6986 => x"78",
          6987 => x"56",
          6988 => x"ac",
          6989 => x"80",
          6990 => x"05",
          6991 => x"61",
          6992 => x"34",
          6993 => x"61",
          6994 => x"c2",
          6995 => x"83",
          6996 => x"81",
          6997 => x"58",
          6998 => x"f9",
          6999 => x"33",
          7000 => x"15",
          7001 => x"81",
          7002 => x"fe",
          7003 => x"8c",
          7004 => x"61",
          7005 => x"34",
          7006 => x"60",
          7007 => x"fc",
          7008 => x"0c",
          7009 => x"04",
          7010 => x"70",
          7011 => x"81",
          7012 => x"61",
          7013 => x"34",
          7014 => x"87",
          7015 => x"ff",
          7016 => x"05",
          7017 => x"b1",
          7018 => x"52",
          7019 => x"80",
          7020 => x"05",
          7021 => x"38",
          7022 => x"05",
          7023 => x"70",
          7024 => x"70",
          7025 => x"34",
          7026 => x"80",
          7027 => x"c1",
          7028 => x"61",
          7029 => x"5b",
          7030 => x"88",
          7031 => x"34",
          7032 => x"ea",
          7033 => x"61",
          7034 => x"ec",
          7035 => x"34",
          7036 => x"61",
          7037 => x"34",
          7038 => x"1f",
          7039 => x"b2",
          7040 => x"52",
          7041 => x"61",
          7042 => x"0d",
          7043 => x"ff",
          7044 => x"b8",
          7045 => x"05",
          7046 => x"ff",
          7047 => x"81",
          7048 => x"74",
          7049 => x"81",
          7050 => x"8a",
          7051 => x"38",
          7052 => x"38",
          7053 => x"8e",
          7054 => x"02",
          7055 => x"77",
          7056 => x"08",
          7057 => x"17",
          7058 => x"77",
          7059 => x"24",
          7060 => x"19",
          7061 => x"8b",
          7062 => x"17",
          7063 => x"3f",
          7064 => x"07",
          7065 => x"81",
          7066 => x"d3",
          7067 => x"3f",
          7068 => x"80",
          7069 => x"80",
          7070 => x"81",
          7071 => x"f4",
          7072 => x"8a",
          7073 => x"76",
          7074 => x"8c",
          7075 => x"16",
          7076 => x"84",
          7077 => x"7c",
          7078 => x"3d",
          7079 => x"05",
          7080 => x"3f",
          7081 => x"7a",
          7082 => x"8c",
          7083 => x"ff",
          7084 => x"52",
          7085 => x"74",
          7086 => x"9f",
          7087 => x"ff",
          7088 => x"eb",
          7089 => x"8c",
          7090 => x"0d",
          7091 => x"52",
          7092 => x"90",
          7093 => x"71",
          7094 => x"04",
          7095 => x"83",
          7096 => x"73",
          7097 => x"22",
          7098 => x"12",
          7099 => x"71",
          7100 => x"83",
          7101 => x"e1",
          7102 => x"06",
          7103 => x"0d",
          7104 => x"22",
          7105 => x"51",
          7106 => x"38",
          7107 => x"84",
          7108 => x"09",
          7109 => x"26",
          7110 => x"05",
          7111 => x"84",
          7112 => x"51",
          7113 => x"38",
          7114 => x"d0",
          7115 => x"d9",
          7116 => x"75",
          7117 => x"26",
          7118 => x"38",
          7119 => x"71",
          7120 => x"70",
          7121 => x"38",
          7122 => x"70",
          7123 => x"70",
          7124 => x"55",
          7125 => x"51",
          7126 => x"0d",
          7127 => x"39",
          7128 => x"10",
          7129 => x"04",
          7130 => x"06",
          7131 => x"b0",
          7132 => x"51",
          7133 => x"ff",
          7134 => x"70",
          7135 => x"39",
          7136 => x"57",
          7137 => x"ff",
          7138 => x"16",
          7139 => x"ff",
          7140 => x"76",
          7141 => x"58",
          7142 => x"31",
          7143 => x"fe",
          7144 => x"ff",
          7145 => x"ff",
          7146 => x"00",
          7147 => x"00",
          7148 => x"00",
          7149 => x"00",
          7150 => x"00",
          7151 => x"00",
          7152 => x"00",
          7153 => x"00",
          7154 => x"00",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"00",
          7372 => x"00",
          7373 => x"00",
          7374 => x"00",
          7375 => x"00",
          7376 => x"00",
          7377 => x"00",
          7378 => x"00",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"64",
          7383 => x"64",
          7384 => x"66",
          7385 => x"66",
          7386 => x"66",
          7387 => x"6d",
          7388 => x"6d",
          7389 => x"6d",
          7390 => x"6d",
          7391 => x"6d",
          7392 => x"6d",
          7393 => x"68",
          7394 => x"68",
          7395 => x"00",
          7396 => x"72",
          7397 => x"72",
          7398 => x"69",
          7399 => x"74",
          7400 => x"63",
          7401 => x"74",
          7402 => x"6d",
          7403 => x"6b",
          7404 => x"65",
          7405 => x"6f",
          7406 => x"72",
          7407 => x"6d",
          7408 => x"6e",
          7409 => x"2e",
          7410 => x"6d",
          7411 => x"6e",
          7412 => x"00",
          7413 => x"66",
          7414 => x"20",
          7415 => x"00",
          7416 => x"20",
          7417 => x"65",
          7418 => x"6f",
          7419 => x"72",
          7420 => x"61",
          7421 => x"2e",
          7422 => x"61",
          7423 => x"65",
          7424 => x"6f",
          7425 => x"65",
          7426 => x"73",
          7427 => x"6e",
          7428 => x"73",
          7429 => x"20",
          7430 => x"62",
          7431 => x"44",
          7432 => x"6d",
          7433 => x"69",
          7434 => x"00",
          7435 => x"73",
          7436 => x"70",
          7437 => x"64",
          7438 => x"20",
          7439 => x"69",
          7440 => x"00",
          7441 => x"20",
          7442 => x"20",
          7443 => x"00",
          7444 => x"73",
          7445 => x"64",
          7446 => x"6c",
          7447 => x"6e",
          7448 => x"4e",
          7449 => x"66",
          7450 => x"4e",
          7451 => x"66",
          7452 => x"44",
          7453 => x"20",
          7454 => x"49",
          7455 => x"20",
          7456 => x"44",
          7457 => x"6f",
          7458 => x"65",
          7459 => x"0a",
          7460 => x"65",
          7461 => x"20",
          7462 => x"65",
          7463 => x"00",
          7464 => x"00",
          7465 => x"58",
          7466 => x"25",
          7467 => x"20",
          7468 => x"20",
          7469 => x"00",
          7470 => x"20",
          7471 => x"7a",
          7472 => x"73",
          7473 => x"32",
          7474 => x"76",
          7475 => x"20",
          7476 => x"76",
          7477 => x"25",
          7478 => x"0a",
          7479 => x"49",
          7480 => x"74",
          7481 => x"72",
          7482 => x"31",
          7483 => x"65",
          7484 => x"55",
          7485 => x"20",
          7486 => x"70",
          7487 => x"30",
          7488 => x"65",
          7489 => x"55",
          7490 => x"20",
          7491 => x"70",
          7492 => x"4c",
          7493 => x"65",
          7494 => x"49",
          7495 => x"20",
          7496 => x"70",
          7497 => x"69",
          7498 => x"74",
          7499 => x"72",
          7500 => x"75",
          7501 => x"69",
          7502 => x"69",
          7503 => x"45",
          7504 => x"20",
          7505 => x"2e",
          7506 => x"65",
          7507 => x"00",
          7508 => x"7a",
          7509 => x"46",
          7510 => x"6f",
          7511 => x"6c",
          7512 => x"63",
          7513 => x"70",
          7514 => x"6e",
          7515 => x"61",
          7516 => x"2a",
          7517 => x"25",
          7518 => x"20",
          7519 => x"69",
          7520 => x"30",
          7521 => x"63",
          7522 => x"00",
          7523 => x"62",
          7524 => x"25",
          7525 => x"00",
          7526 => x"20",
          7527 => x"6e",
          7528 => x"52",
          7529 => x"6e",
          7530 => x"63",
          7531 => x"2e",
          7532 => x"69",
          7533 => x"20",
          7534 => x"20",
          7535 => x"43",
          7536 => x"75",
          7537 => x"64",
          7538 => x"0a",
          7539 => x"75",
          7540 => x"64",
          7541 => x"6c",
          7542 => x"25",
          7543 => x"38",
          7544 => x"25",
          7545 => x"34",
          7546 => x"61",
          7547 => x"00",
          7548 => x"78",
          7549 => x"3e",
          7550 => x"30",
          7551 => x"43",
          7552 => x"2e",
          7553 => x"58",
          7554 => x"43",
          7555 => x"2e",
          7556 => x"44",
          7557 => x"6f",
          7558 => x"70",
          7559 => x"25",
          7560 => x"73",
          7561 => x"72",
          7562 => x"73",
          7563 => x"6e",
          7564 => x"63",
          7565 => x"6d",
          7566 => x"3f",
          7567 => x"64",
          7568 => x"25",
          7569 => x"25",
          7570 => x"43",
          7571 => x"61",
          7572 => x"3a",
          7573 => x"73",
          7574 => x"65",
          7575 => x"41",
          7576 => x"73",
          7577 => x"43",
          7578 => x"74",
          7579 => x"20",
          7580 => x"20",
          7581 => x"00",
          7582 => x"43",
          7583 => x"72",
          7584 => x"20",
          7585 => x"20",
          7586 => x"00",
          7587 => x"53",
          7588 => x"61",
          7589 => x"65",
          7590 => x"20",
          7591 => x"00",
          7592 => x"3a",
          7593 => x"5a",
          7594 => x"20",
          7595 => x"20",
          7596 => x"20",
          7597 => x"00",
          7598 => x"53",
          7599 => x"6c",
          7600 => x"71",
          7601 => x"20",
          7602 => x"34",
          7603 => x"20",
          7604 => x"62",
          7605 => x"41",
          7606 => x"20",
          7607 => x"64",
          7608 => x"7a",
          7609 => x"53",
          7610 => x"6f",
          7611 => x"20",
          7612 => x"20",
          7613 => x"34",
          7614 => x"20",
          7615 => x"20",
          7616 => x"20",
          7617 => x"4c",
          7618 => x"57",
          7619 => x"20",
          7620 => x"42",
          7621 => x"00",
          7622 => x"49",
          7623 => x"4c",
          7624 => x"65",
          7625 => x"29",
          7626 => x"54",
          7627 => x"20",
          7628 => x"73",
          7629 => x"29",
          7630 => x"53",
          7631 => x"20",
          7632 => x"65",
          7633 => x"29",
          7634 => x"52",
          7635 => x"20",
          7636 => x"25",
          7637 => x"20",
          7638 => x"20",
          7639 => x"30",
          7640 => x"29",
          7641 => x"49",
          7642 => x"4d",
          7643 => x"25",
          7644 => x"20",
          7645 => x"4d",
          7646 => x"30",
          7647 => x"29",
          7648 => x"57",
          7649 => x"20",
          7650 => x"25",
          7651 => x"20",
          7652 => x"6f",
          7653 => x"67",
          7654 => x"6f",
          7655 => x"00",
          7656 => x"6c",
          7657 => x"75",
          7658 => x"00",
          7659 => x"00",
          7660 => x"00",
          7661 => x"01",
          7662 => x"00",
          7663 => x"00",
          7664 => x"01",
          7665 => x"00",
          7666 => x"00",
          7667 => x"01",
          7668 => x"00",
          7669 => x"00",
          7670 => x"01",
          7671 => x"00",
          7672 => x"00",
          7673 => x"01",
          7674 => x"00",
          7675 => x"00",
          7676 => x"04",
          7677 => x"00",
          7678 => x"00",
          7679 => x"04",
          7680 => x"00",
          7681 => x"00",
          7682 => x"04",
          7683 => x"00",
          7684 => x"00",
          7685 => x"04",
          7686 => x"00",
          7687 => x"00",
          7688 => x"03",
          7689 => x"00",
          7690 => x"00",
          7691 => x"03",
          7692 => x"1b",
          7693 => x"1b",
          7694 => x"1b",
          7695 => x"1b",
          7696 => x"1b",
          7697 => x"1b",
          7698 => x"0e",
          7699 => x"0b",
          7700 => x"06",
          7701 => x"04",
          7702 => x"02",
          7703 => x"43",
          7704 => x"70",
          7705 => x"74",
          7706 => x"72",
          7707 => x"20",
          7708 => x"6e",
          7709 => x"6f",
          7710 => x"00",
          7711 => x"25",
          7712 => x"73",
          7713 => x"65",
          7714 => x"73",
          7715 => x"68",
          7716 => x"66",
          7717 => x"45",
          7718 => x"3e",
          7719 => x"1b",
          7720 => x"1b",
          7721 => x"1b",
          7722 => x"1b",
          7723 => x"1b",
          7724 => x"1b",
          7725 => x"1b",
          7726 => x"1b",
          7727 => x"1b",
          7728 => x"1b",
          7729 => x"1b",
          7730 => x"1b",
          7731 => x"1b",
          7732 => x"1b",
          7733 => x"1b",
          7734 => x"1b",
          7735 => x"00",
          7736 => x"00",
          7737 => x"2c",
          7738 => x"64",
          7739 => x"25",
          7740 => x"44",
          7741 => x"25",
          7742 => x"2c",
          7743 => x"25",
          7744 => x"3a",
          7745 => x"2c",
          7746 => x"64",
          7747 => x"52",
          7748 => x"75",
          7749 => x"55",
          7750 => x"25",
          7751 => x"44",
          7752 => x"25",
          7753 => x"48",
          7754 => x"00",
          7755 => x"65",
          7756 => x"20",
          7757 => x"42",
          7758 => x"2c",
          7759 => x"64",
          7760 => x"65",
          7761 => x"20",
          7762 => x"4e",
          7763 => x"64",
          7764 => x"00",
          7765 => x"22",
          7766 => x"00",
          7767 => x"5b",
          7768 => x"46",
          7769 => x"eb",
          7770 => x"35",
          7771 => x"41",
          7772 => x"41",
          7773 => x"4e",
          7774 => x"20",
          7775 => x"20",
          7776 => x"00",
          7777 => x"00",
          7778 => x"09",
          7779 => x"1e",
          7780 => x"8e",
          7781 => x"49",
          7782 => x"99",
          7783 => x"9c",
          7784 => x"a5",
          7785 => x"ac",
          7786 => x"b4",
          7787 => x"bc",
          7788 => x"c4",
          7789 => x"cc",
          7790 => x"d4",
          7791 => x"dc",
          7792 => x"e4",
          7793 => x"ec",
          7794 => x"f4",
          7795 => x"fc",
          7796 => x"3d",
          7797 => x"3c",
          7798 => x"00",
          7799 => x"01",
          7800 => x"00",
          7801 => x"00",
          7802 => x"00",
          7803 => x"00",
          7804 => x"00",
          7805 => x"00",
          7806 => x"00",
          7807 => x"00",
          7808 => x"00",
          7809 => x"00",
          7810 => x"00",
          7811 => x"00",
          7812 => x"00",
          7813 => x"00",
          7814 => x"25",
          7815 => x"25",
          7816 => x"25",
          7817 => x"25",
          7818 => x"25",
          7819 => x"25",
          7820 => x"25",
          7821 => x"25",
          7822 => x"25",
          7823 => x"25",
          7824 => x"25",
          7825 => x"25",
          7826 => x"03",
          7827 => x"03",
          7828 => x"03",
          7829 => x"22",
          7830 => x"22",
          7831 => x"23",
          7832 => x"00",
          7833 => x"20",
          7834 => x"00",
          7835 => x"00",
          7836 => x"01",
          7837 => x"01",
          7838 => x"01",
          7839 => x"00",
          7840 => x"01",
          7841 => x"01",
          7842 => x"01",
          7843 => x"01",
          7844 => x"01",
          7845 => x"01",
          7846 => x"01",
          7847 => x"01",
          7848 => x"01",
          7849 => x"01",
          7850 => x"01",
          7851 => x"01",
          7852 => x"01",
          7853 => x"01",
          7854 => x"01",
          7855 => x"01",
          7856 => x"01",
          7857 => x"01",
          7858 => x"01",
          7859 => x"01",
          7860 => x"01",
          7861 => x"01",
          7862 => x"02",
          7863 => x"2c",
          7864 => x"2c",
          7865 => x"02",
          7866 => x"00",
          7867 => x"01",
          7868 => x"02",
          7869 => x"02",
          7870 => x"02",
          7871 => x"02",
          7872 => x"02",
          7873 => x"02",
          7874 => x"01",
          7875 => x"02",
          7876 => x"02",
          7877 => x"02",
          7878 => x"02",
          7879 => x"02",
          7880 => x"01",
          7881 => x"02",
          7882 => x"01",
          7883 => x"03",
          7884 => x"03",
          7885 => x"03",
          7886 => x"03",
          7887 => x"03",
          7888 => x"03",
          7889 => x"00",
          7890 => x"03",
          7891 => x"03",
          7892 => x"03",
          7893 => x"01",
          7894 => x"01",
          7895 => x"04",
          7896 => x"00",
          7897 => x"2c",
          7898 => x"01",
          7899 => x"06",
          7900 => x"06",
          7901 => x"00",
          7902 => x"1f",
          7903 => x"1f",
          7904 => x"1f",
          7905 => x"1f",
          7906 => x"1f",
          7907 => x"1f",
          7908 => x"1f",
          7909 => x"1f",
          7910 => x"1f",
          7911 => x"1f",
          7912 => x"06",
          7913 => x"1f",
          7914 => x"00",
          7915 => x"21",
          7916 => x"05",
          7917 => x"01",
          7918 => x"01",
          7919 => x"08",
          7920 => x"00",
          7921 => x"01",
          7922 => x"00",
          7923 => x"01",
          7924 => x"00",
          7925 => x"01",
          7926 => x"00",
          7927 => x"01",
          7928 => x"00",
          7929 => x"01",
          7930 => x"00",
          7931 => x"01",
          7932 => x"00",
          7933 => x"01",
          7934 => x"00",
          7935 => x"01",
          7936 => x"00",
          7937 => x"01",
          7938 => x"00",
          7939 => x"01",
          7940 => x"00",
          7941 => x"01",
          7942 => x"00",
          7943 => x"01",
          7944 => x"00",
          7945 => x"01",
          7946 => x"00",
          7947 => x"01",
          7948 => x"00",
          7949 => x"01",
          7950 => x"00",
          7951 => x"01",
          7952 => x"00",
          7953 => x"01",
          7954 => x"00",
          7955 => x"01",
          7956 => x"00",
          7957 => x"01",
          7958 => x"00",
          7959 => x"01",
          7960 => x"00",
          7961 => x"01",
          7962 => x"00",
          7963 => x"01",
          7964 => x"00",
          7965 => x"01",
          7966 => x"00",
          7967 => x"01",
          7968 => x"00",
          7969 => x"01",
          7970 => x"00",
          7971 => x"01",
          7972 => x"00",
          7973 => x"01",
          7974 => x"00",
          7975 => x"01",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"00",
          7980 => x"00",
          7981 => x"01",
          7982 => x"00",
          7983 => x"00",
          7984 => x"05",
          7985 => x"05",
          7986 => x"01",
          7987 => x"01",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"00",
          7996 => x"00",
          7997 => x"00",
          7998 => x"00",
          7999 => x"00",
          8000 => x"00",
          8001 => x"00",
          8002 => x"00",
          8003 => x"00",
          8004 => x"f0",
          8005 => x"5d",
          8006 => x"75",
          8007 => x"6d",
          8008 => x"65",
          8009 => x"35",
          8010 => x"30",
          8011 => x"f1",
          8012 => x"f0",
          8013 => x"84",
          8014 => x"f0",
          8015 => x"5d",
          8016 => x"55",
          8017 => x"4d",
          8018 => x"45",
          8019 => x"35",
          8020 => x"30",
          8021 => x"f1",
          8022 => x"f0",
          8023 => x"84",
          8024 => x"f0",
          8025 => x"7d",
          8026 => x"55",
          8027 => x"4d",
          8028 => x"45",
          8029 => x"25",
          8030 => x"20",
          8031 => x"f9",
          8032 => x"f0",
          8033 => x"89",
          8034 => x"f0",
          8035 => x"1d",
          8036 => x"15",
          8037 => x"0d",
          8038 => x"05",
          8039 => x"f0",
          8040 => x"f0",
          8041 => x"f0",
          8042 => x"f0",
          8043 => x"84",
          8044 => x"f0",
          8045 => x"b7",
          8046 => x"39",
          8047 => x"1d",
          8048 => x"74",
          8049 => x"7a",
          8050 => x"9d",
          8051 => x"c3",
          8052 => x"f0",
          8053 => x"84",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"f8",
          8068 => x"f3",
          8069 => x"f4",
          8070 => x"f1",
          8071 => x"f2",
          8072 => x"80",
          8073 => x"81",
          8074 => x"82",
          8075 => x"83",
          8076 => x"84",
          8077 => x"85",
          8078 => x"86",
          8079 => x"87",
          8080 => x"88",
          8081 => x"89",
          8082 => x"f6",
          8083 => x"7f",
          8084 => x"f9",
          8085 => x"e0",
          8086 => x"e1",
          8087 => x"71",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"50",
          9089 => x"cc",
          9090 => x"f8",
          9091 => x"e1",
          9092 => x"e3",
          9093 => x"00",
          9094 => x"68",
          9095 => x"20",
          9096 => x"28",
          9097 => x"55",
          9098 => x"08",
          9099 => x"10",
          9100 => x"18",
          9101 => x"c7",
          9102 => x"88",
          9103 => x"90",
          9104 => x"98",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"00",
          9113 => x"00",
          9114 => x"00",
          9115 => x"00",
          9116 => x"00",
          9117 => x"00",
          9118 => x"00",
          9119 => x"00",
          9120 => x"00",
          9121 => x"01",
        others => X"00"
    );

    shared variable RAM4 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"80",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"09",
             9 => x"83",
            10 => x"00",
            11 => x"00",
            12 => x"73",
            13 => x"83",
            14 => x"ff",
            15 => x"00",
            16 => x"73",
            17 => x"06",
            18 => x"00",
            19 => x"00",
            20 => x"53",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"72",
            26 => x"06",
            27 => x"00",
            28 => x"53",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"00",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"04",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"0b",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"2a",
            49 => x"05",
            50 => x"00",
            51 => x"00",
            52 => x"83",
            53 => x"2b",
            54 => x"51",
            55 => x"00",
            56 => x"70",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"70",
            61 => x"06",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"51",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"06",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"09",
            77 => x"2a",
            78 => x"00",
            79 => x"00",
            80 => x"be",
            81 => x"08",
            82 => x"00",
            83 => x"00",
            84 => x"75",
            85 => x"50",
            86 => x"88",
            87 => x"00",
            88 => x"75",
            89 => x"50",
            90 => x"88",
            91 => x"00",
            92 => x"0a",
            93 => x"06",
            94 => x"06",
            95 => x"00",
            96 => x"0a",
            97 => x"71",
            98 => x"05",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"52",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"51",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"8c",
           134 => x"04",
           135 => x"0b",
           136 => x"8c",
           137 => x"04",
           138 => x"0b",
           139 => x"8d",
           140 => x"04",
           141 => x"0b",
           142 => x"8d",
           143 => x"04",
           144 => x"0b",
           145 => x"8e",
           146 => x"04",
           147 => x"0b",
           148 => x"8e",
           149 => x"04",
           150 => x"0b",
           151 => x"8f",
           152 => x"04",
           153 => x"0b",
           154 => x"8f",
           155 => x"04",
           156 => x"0b",
           157 => x"90",
           158 => x"04",
           159 => x"0b",
           160 => x"90",
           161 => x"04",
           162 => x"0b",
           163 => x"91",
           164 => x"04",
           165 => x"0b",
           166 => x"91",
           167 => x"04",
           168 => x"0b",
           169 => x"92",
           170 => x"04",
           171 => x"0b",
           172 => x"92",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"98",
           193 => x"98",
           194 => x"ba",
           195 => x"98",
           196 => x"ba",
           197 => x"98",
           198 => x"ba",
           199 => x"98",
           200 => x"ba",
           201 => x"98",
           202 => x"ba",
           203 => x"98",
           204 => x"ba",
           205 => x"98",
           206 => x"ba",
           207 => x"98",
           208 => x"ba",
           209 => x"98",
           210 => x"ba",
           211 => x"98",
           212 => x"ba",
           213 => x"98",
           214 => x"ba",
           215 => x"98",
           216 => x"ba",
           217 => x"ba",
           218 => x"84",
           219 => x"84",
           220 => x"04",
           221 => x"2d",
           222 => x"90",
           223 => x"ca",
           224 => x"80",
           225 => x"c9",
           226 => x"c0",
           227 => x"82",
           228 => x"80",
           229 => x"0c",
           230 => x"08",
           231 => x"98",
           232 => x"98",
           233 => x"ba",
           234 => x"ba",
           235 => x"84",
           236 => x"84",
           237 => x"04",
           238 => x"2d",
           239 => x"90",
           240 => x"87",
           241 => x"80",
           242 => x"f3",
           243 => x"c0",
           244 => x"82",
           245 => x"80",
           246 => x"0c",
           247 => x"08",
           248 => x"98",
           249 => x"98",
           250 => x"ba",
           251 => x"ba",
           252 => x"84",
           253 => x"84",
           254 => x"04",
           255 => x"2d",
           256 => x"90",
           257 => x"d1",
           258 => x"80",
           259 => x"e6",
           260 => x"c0",
           261 => x"82",
           262 => x"80",
           263 => x"0c",
           264 => x"08",
           265 => x"98",
           266 => x"98",
           267 => x"ba",
           268 => x"ba",
           269 => x"84",
           270 => x"84",
           271 => x"04",
           272 => x"2d",
           273 => x"90",
           274 => x"c8",
           275 => x"80",
           276 => x"a4",
           277 => x"c0",
           278 => x"83",
           279 => x"80",
           280 => x"0c",
           281 => x"08",
           282 => x"98",
           283 => x"98",
           284 => x"ba",
           285 => x"ba",
           286 => x"84",
           287 => x"84",
           288 => x"04",
           289 => x"2d",
           290 => x"90",
           291 => x"e9",
           292 => x"80",
           293 => x"d7",
           294 => x"c0",
           295 => x"b1",
           296 => x"c0",
           297 => x"81",
           298 => x"80",
           299 => x"0c",
           300 => x"08",
           301 => x"98",
           302 => x"98",
           303 => x"ba",
           304 => x"ba",
           305 => x"3c",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"ff",
           311 => x"83",
           312 => x"fc",
           313 => x"80",
           314 => x"06",
           315 => x"0a",
           316 => x"51",
           317 => x"f8",
           318 => x"05",
           319 => x"04",
           320 => x"00",
           321 => x"84",
           322 => x"84",
           323 => x"86",
           324 => x"7a",
           325 => x"06",
           326 => x"57",
           327 => x"06",
           328 => x"8a",
           329 => x"2a",
           330 => x"25",
           331 => x"75",
           332 => x"08",
           333 => x"ae",
           334 => x"81",
           335 => x"32",
           336 => x"51",
           337 => x"38",
           338 => x"ba",
           339 => x"0b",
           340 => x"04",
           341 => x"84",
           342 => x"0a",
           343 => x"52",
           344 => x"73",
           345 => x"0d",
           346 => x"05",
           347 => x"85",
           348 => x"63",
           349 => x"1f",
           350 => x"81",
           351 => x"54",
           352 => x"d2",
           353 => x"80",
           354 => x"54",
           355 => x"d0",
           356 => x"38",
           357 => x"25",
           358 => x"80",
           359 => x"81",
           360 => x"2e",
           361 => x"7b",
           362 => x"1d",
           363 => x"91",
           364 => x"78",
           365 => x"98",
           366 => x"80",
           367 => x"2c",
           368 => x"24",
           369 => x"72",
           370 => x"58",
           371 => x"76",
           372 => x"81",
           373 => x"33",
           374 => x"9e",
           375 => x"3f",
           376 => x"ff",
           377 => x"06",
           378 => x"74",
           379 => x"17",
           380 => x"72",
           381 => x"73",
           382 => x"80",
           383 => x"76",
           384 => x"58",
           385 => x"39",
           386 => x"5a",
           387 => x"83",
           388 => x"84",
           389 => x"93",
           390 => x"ff",
           391 => x"05",
           392 => x"84",
           393 => x"7e",
           394 => x"75",
           395 => x"08",
           396 => x"7d",
           397 => x"b2",
           398 => x"38",
           399 => x"80",
           400 => x"86",
           401 => x"80",
           402 => x"29",
           403 => x"2e",
           404 => x"fc",
           405 => x"58",
           406 => x"55",
           407 => x"2c",
           408 => x"73",
           409 => x"f7",
           410 => x"41",
           411 => x"80",
           412 => x"90",
           413 => x"06",
           414 => x"96",
           415 => x"73",
           416 => x"06",
           417 => x"2a",
           418 => x"7e",
           419 => x"7a",
           420 => x"2e",
           421 => x"29",
           422 => x"5a",
           423 => x"7c",
           424 => x"78",
           425 => x"05",
           426 => x"80",
           427 => x"72",
           428 => x"80",
           429 => x"98",
           430 => x"9d",
           431 => x"3f",
           432 => x"ff",
           433 => x"55",
           434 => x"2a",
           435 => x"2e",
           436 => x"84",
           437 => x"ca",
           438 => x"38",
           439 => x"7c",
           440 => x"87",
           441 => x"09",
           442 => x"5b",
           443 => x"78",
           444 => x"05",
           445 => x"75",
           446 => x"51",
           447 => x"07",
           448 => x"5b",
           449 => x"7a",
           450 => x"90",
           451 => x"83",
           452 => x"5a",
           453 => x"77",
           454 => x"70",
           455 => x"80",
           456 => x"2c",
           457 => x"7a",
           458 => x"7a",
           459 => x"80",
           460 => x"2c",
           461 => x"b3",
           462 => x"3f",
           463 => x"ff",
           464 => x"2e",
           465 => x"81",
           466 => x"e2",
           467 => x"06",
           468 => x"fe",
           469 => x"05",
           470 => x"39",
           471 => x"07",
           472 => x"80",
           473 => x"80",
           474 => x"5d",
           475 => x"fb",
           476 => x"70",
           477 => x"82",
           478 => x"5b",
           479 => x"7a",
           480 => x"f8",
           481 => x"07",
           482 => x"f7",
           483 => x"84",
           484 => x"58",
           485 => x"51",
           486 => x"83",
           487 => x"2b",
           488 => x"87",
           489 => x"58",
           490 => x"39",
           491 => x"81",
           492 => x"cf",
           493 => x"ba",
           494 => x"71",
           495 => x"7a",
           496 => x"76",
           497 => x"78",
           498 => x"05",
           499 => x"74",
           500 => x"51",
           501 => x"b0",
           502 => x"09",
           503 => x"76",
           504 => x"81",
           505 => x"38",
           506 => x"71",
           507 => x"83",
           508 => x"fa",
           509 => x"ad",
           510 => x"54",
           511 => x"ad",
           512 => x"82",
           513 => x"80",
           514 => x"78",
           515 => x"5a",
           516 => x"51",
           517 => x"a0",
           518 => x"78",
           519 => x"ba",
           520 => x"71",
           521 => x"39",
           522 => x"ff",
           523 => x"39",
           524 => x"53",
           525 => x"84",
           526 => x"55",
           527 => x"11",
           528 => x"81",
           529 => x"56",
           530 => x"d5",
           531 => x"53",
           532 => x"f0",
           533 => x"53",
           534 => x"2e",
           535 => x"05",
           536 => x"38",
           537 => x"84",
           538 => x"08",
           539 => x"74",
           540 => x"83",
           541 => x"ba",
           542 => x"3d",
           543 => x"85",
           544 => x"70",
           545 => x"56",
           546 => x"38",
           547 => x"72",
           548 => x"76",
           549 => x"3d",
           550 => x"33",
           551 => x"52",
           552 => x"2d",
           553 => x"38",
           554 => x"54",
           555 => x"3d",
           556 => x"51",
           557 => x"3d",
           558 => x"81",
           559 => x"56",
           560 => x"82",
           561 => x"ac",
           562 => x"16",
           563 => x"76",
           564 => x"0c",
           565 => x"16",
           566 => x"0c",
           567 => x"81",
           568 => x"73",
           569 => x"e3",
           570 => x"16",
           571 => x"0d",
           572 => x"06",
           573 => x"56",
           574 => x"86",
           575 => x"72",
           576 => x"2e",
           577 => x"53",
           578 => x"81",
           579 => x"05",
           580 => x"54",
           581 => x"0d",
           582 => x"85",
           583 => x"8c",
           584 => x"8c",
           585 => x"94",
           586 => x"8c",
           587 => x"25",
           588 => x"90",
           589 => x"ff",
           590 => x"72",
           591 => x"ba",
           592 => x"a0",
           593 => x"54",
           594 => x"71",
           595 => x"53",
           596 => x"52",
           597 => x"70",
           598 => x"f0",
           599 => x"3d",
           600 => x"71",
           601 => x"2e",
           602 => x"70",
           603 => x"05",
           604 => x"34",
           605 => x"84",
           606 => x"70",
           607 => x"70",
           608 => x"13",
           609 => x"11",
           610 => x"13",
           611 => x"34",
           612 => x"39",
           613 => x"71",
           614 => x"f7",
           615 => x"ba",
           616 => x"fd",
           617 => x"54",
           618 => x"70",
           619 => x"f0",
           620 => x"3d",
           621 => x"71",
           622 => x"2e",
           623 => x"33",
           624 => x"11",
           625 => x"8c",
           626 => x"0d",
           627 => x"80",
           628 => x"81",
           629 => x"2e",
           630 => x"54",
           631 => x"53",
           632 => x"ba",
           633 => x"80",
           634 => x"51",
           635 => x"33",
           636 => x"38",
           637 => x"86",
           638 => x"0c",
           639 => x"77",
           640 => x"3f",
           641 => x"08",
           642 => x"3f",
           643 => x"8c",
           644 => x"8c",
           645 => x"53",
           646 => x"fe",
           647 => x"73",
           648 => x"04",
           649 => x"54",
           650 => x"38",
           651 => x"70",
           652 => x"71",
           653 => x"ff",
           654 => x"84",
           655 => x"fd",
           656 => x"53",
           657 => x"72",
           658 => x"11",
           659 => x"8c",
           660 => x"0d",
           661 => x"80",
           662 => x"3f",
           663 => x"53",
           664 => x"80",
           665 => x"31",
           666 => x"cb",
           667 => x"c3",
           668 => x"72",
           669 => x"55",
           670 => x"72",
           671 => x"77",
           672 => x"2c",
           673 => x"71",
           674 => x"55",
           675 => x"10",
           676 => x"0c",
           677 => x"76",
           678 => x"70",
           679 => x"90",
           680 => x"fe",
           681 => x"83",
           682 => x"70",
           683 => x"25",
           684 => x"2a",
           685 => x"06",
           686 => x"71",
           687 => x"81",
           688 => x"74",
           689 => x"8c",
           690 => x"56",
           691 => x"56",
           692 => x"86",
           693 => x"77",
           694 => x"94",
           695 => x"74",
           696 => x"85",
           697 => x"7a",
           698 => x"8b",
           699 => x"ba",
           700 => x"80",
           701 => x"3f",
           702 => x"73",
           703 => x"80",
           704 => x"12",
           705 => x"71",
           706 => x"74",
           707 => x"9f",
           708 => x"72",
           709 => x"06",
           710 => x"1c",
           711 => x"53",
           712 => x"0c",
           713 => x"78",
           714 => x"2c",
           715 => x"73",
           716 => x"75",
           717 => x"fc",
           718 => x"32",
           719 => x"3d",
           720 => x"5b",
           721 => x"70",
           722 => x"09",
           723 => x"78",
           724 => x"2e",
           725 => x"38",
           726 => x"14",
           727 => x"db",
           728 => x"27",
           729 => x"89",
           730 => x"55",
           731 => x"51",
           732 => x"13",
           733 => x"73",
           734 => x"81",
           735 => x"16",
           736 => x"56",
           737 => x"80",
           738 => x"7a",
           739 => x"0c",
           740 => x"70",
           741 => x"73",
           742 => x"38",
           743 => x"55",
           744 => x"90",
           745 => x"81",
           746 => x"14",
           747 => x"27",
           748 => x"0c",
           749 => x"15",
           750 => x"80",
           751 => x"ba",
           752 => x"3d",
           753 => x"7b",
           754 => x"59",
           755 => x"38",
           756 => x"55",
           757 => x"ad",
           758 => x"81",
           759 => x"77",
           760 => x"80",
           761 => x"80",
           762 => x"70",
           763 => x"70",
           764 => x"27",
           765 => x"06",
           766 => x"38",
           767 => x"76",
           768 => x"70",
           769 => x"ff",
           770 => x"75",
           771 => x"75",
           772 => x"04",
           773 => x"33",
           774 => x"81",
           775 => x"78",
           776 => x"e2",
           777 => x"f8",
           778 => x"27",
           779 => x"88",
           780 => x"75",
           781 => x"04",
           782 => x"70",
           783 => x"39",
           784 => x"3d",
           785 => x"ba",
           786 => x"8c",
           787 => x"71",
           788 => x"83",
           789 => x"83",
           790 => x"3d",
           791 => x"b3",
           792 => x"8c",
           793 => x"04",
           794 => x"83",
           795 => x"ef",
           796 => x"cf",
           797 => x"0d",
           798 => x"3f",
           799 => x"51",
           800 => x"83",
           801 => x"3d",
           802 => x"db",
           803 => x"d4",
           804 => x"04",
           805 => x"83",
           806 => x"ee",
           807 => x"d1",
           808 => x"0d",
           809 => x"3f",
           810 => x"51",
           811 => x"83",
           812 => x"3d",
           813 => x"83",
           814 => x"f0",
           815 => x"04",
           816 => x"83",
           817 => x"ed",
           818 => x"3d",
           819 => x"05",
           820 => x"70",
           821 => x"59",
           822 => x"38",
           823 => x"ff",
           824 => x"e2",
           825 => x"70",
           826 => x"ba",
           827 => x"80",
           828 => x"af",
           829 => x"80",
           830 => x"06",
           831 => x"aa",
           832 => x"74",
           833 => x"52",
           834 => x"3f",
           835 => x"bc",
           836 => x"df",
           837 => x"96",
           838 => x"87",
           839 => x"08",
           840 => x"80",
           841 => x"97",
           842 => x"ba",
           843 => x"74",
           844 => x"75",
           845 => x"52",
           846 => x"8c",
           847 => x"84",
           848 => x"53",
           849 => x"f8",
           850 => x"7c",
           851 => x"59",
           852 => x"51",
           853 => x"8b",
           854 => x"81",
           855 => x"0c",
           856 => x"d5",
           857 => x"ba",
           858 => x"2d",
           859 => x"0c",
           860 => x"7f",
           861 => x"05",
           862 => x"5c",
           863 => x"83",
           864 => x"51",
           865 => x"dd",
           866 => x"b2",
           867 => x"7c",
           868 => x"53",
           869 => x"33",
           870 => x"3f",
           871 => x"54",
           872 => x"26",
           873 => x"b8",
           874 => x"c0",
           875 => x"80",
           876 => x"55",
           877 => x"81",
           878 => x"06",
           879 => x"80",
           880 => x"d5",
           881 => x"3f",
           882 => x"38",
           883 => x"78",
           884 => x"9d",
           885 => x"2b",
           886 => x"2e",
           887 => x"c3",
           888 => x"fe",
           889 => x"0c",
           890 => x"51",
           891 => x"f0",
           892 => x"3f",
           893 => x"da",
           894 => x"3f",
           895 => x"54",
           896 => x"27",
           897 => x"7a",
           898 => x"d2",
           899 => x"84",
           900 => x"ea",
           901 => x"fe",
           902 => x"d0",
           903 => x"53",
           904 => x"79",
           905 => x"72",
           906 => x"83",
           907 => x"14",
           908 => x"51",
           909 => x"38",
           910 => x"52",
           911 => x"56",
           912 => x"84",
           913 => x"88",
           914 => x"a0",
           915 => x"06",
           916 => x"39",
           917 => x"8c",
           918 => x"a0",
           919 => x"30",
           920 => x"51",
           921 => x"80",
           922 => x"83",
           923 => x"70",
           924 => x"72",
           925 => x"73",
           926 => x"57",
           927 => x"38",
           928 => x"8c",
           929 => x"0d",
           930 => x"d1",
           931 => x"d3",
           932 => x"9c",
           933 => x"06",
           934 => x"82",
           935 => x"82",
           936 => x"06",
           937 => x"84",
           938 => x"81",
           939 => x"06",
           940 => x"86",
           941 => x"80",
           942 => x"06",
           943 => x"2a",
           944 => x"e9",
           945 => x"9c",
           946 => x"94",
           947 => x"d1",
           948 => x"9b",
           949 => x"fc",
           950 => x"88",
           951 => x"c6",
           952 => x"3f",
           953 => x"80",
           954 => x"70",
           955 => x"ff",
           956 => x"ac",
           957 => x"3f",
           958 => x"2a",
           959 => x"2e",
           960 => x"51",
           961 => x"9b",
           962 => x"72",
           963 => x"71",
           964 => x"39",
           965 => x"b0",
           966 => x"dc",
           967 => x"51",
           968 => x"ff",
           969 => x"83",
           970 => x"51",
           971 => x"81",
           972 => x"e6",
           973 => x"a4",
           974 => x"3f",
           975 => x"2a",
           976 => x"2e",
           977 => x"3d",
           978 => x"84",
           979 => x"51",
           980 => x"08",
           981 => x"78",
           982 => x"a8",
           983 => x"83",
           984 => x"48",
           985 => x"eb",
           986 => x"33",
           987 => x"80",
           988 => x"83",
           989 => x"7d",
           990 => x"5a",
           991 => x"79",
           992 => x"06",
           993 => x"5a",
           994 => x"7b",
           995 => x"83",
           996 => x"e7",
           997 => x"ba",
           998 => x"52",
           999 => x"08",
          1000 => x"81",
          1001 => x"81",
          1002 => x"c4",
          1003 => x"2e",
          1004 => x"51",
          1005 => x"5e",
          1006 => x"d3",
          1007 => x"3d",
          1008 => x"84",
          1009 => x"5c",
          1010 => x"ba",
          1011 => x"ba",
          1012 => x"81",
          1013 => x"2e",
          1014 => x"ec",
          1015 => x"7b",
          1016 => x"7c",
          1017 => x"58",
          1018 => x"55",
          1019 => x"80",
          1020 => x"84",
          1021 => x"09",
          1022 => x"51",
          1023 => x"26",
          1024 => x"59",
          1025 => x"70",
          1026 => x"95",
          1027 => x"07",
          1028 => x"2e",
          1029 => x"aa",
          1030 => x"3f",
          1031 => x"7e",
          1032 => x"ef",
          1033 => x"59",
          1034 => x"d5",
          1035 => x"89",
          1036 => x"c5",
          1037 => x"80",
          1038 => x"52",
          1039 => x"ba",
          1040 => x"ba",
          1041 => x"0b",
          1042 => x"06",
          1043 => x"06",
          1044 => x"9c",
          1045 => x"0b",
          1046 => x"9c",
          1047 => x"ce",
          1048 => x"b7",
          1049 => x"85",
          1050 => x"fd",
          1051 => x"9c",
          1052 => x"ec",
          1053 => x"83",
          1054 => x"e4",
          1055 => x"bb",
          1056 => x"ba",
          1057 => x"fb",
          1058 => x"41",
          1059 => x"51",
          1060 => x"b2",
          1061 => x"56",
          1062 => x"53",
          1063 => x"e8",
          1064 => x"3f",
          1065 => x"ef",
          1066 => x"3f",
          1067 => x"fa",
          1068 => x"8b",
          1069 => x"c0",
          1070 => x"fa",
          1071 => x"53",
          1072 => x"84",
          1073 => x"38",
          1074 => x"f0",
          1075 => x"8c",
          1076 => x"ba",
          1077 => x"d0",
          1078 => x"ff",
          1079 => x"eb",
          1080 => x"2e",
          1081 => x"94",
          1082 => x"04",
          1083 => x"80",
          1084 => x"8c",
          1085 => x"3d",
          1086 => x"51",
          1087 => x"86",
          1088 => x"78",
          1089 => x"3f",
          1090 => x"52",
          1091 => x"7e",
          1092 => x"38",
          1093 => x"84",
          1094 => x"3d",
          1095 => x"51",
          1096 => x"80",
          1097 => x"f0",
          1098 => x"aa",
          1099 => x"38",
          1100 => x"83",
          1101 => x"d5",
          1102 => x"51",
          1103 => x"59",
          1104 => x"9f",
          1105 => x"70",
          1106 => x"84",
          1107 => x"e6",
          1108 => x"f8",
          1109 => x"53",
          1110 => x"84",
          1111 => x"38",
          1112 => x"80",
          1113 => x"8c",
          1114 => x"d7",
          1115 => x"5d",
          1116 => x"65",
          1117 => x"7a",
          1118 => x"54",
          1119 => x"dc",
          1120 => x"5c",
          1121 => x"39",
          1122 => x"80",
          1123 => x"8c",
          1124 => x"3d",
          1125 => x"51",
          1126 => x"80",
          1127 => x"f8",
          1128 => x"be",
          1129 => x"f6",
          1130 => x"b0",
          1131 => x"93",
          1132 => x"5b",
          1133 => x"eb",
          1134 => x"ff",
          1135 => x"ba",
          1136 => x"b8",
          1137 => x"05",
          1138 => x"08",
          1139 => x"83",
          1140 => x"d5",
          1141 => x"51",
          1142 => x"59",
          1143 => x"9f",
          1144 => x"49",
          1145 => x"05",
          1146 => x"b8",
          1147 => x"05",
          1148 => x"08",
          1149 => x"02",
          1150 => x"81",
          1151 => x"53",
          1152 => x"84",
          1153 => x"af",
          1154 => x"ff",
          1155 => x"ba",
          1156 => x"b8",
          1157 => x"05",
          1158 => x"08",
          1159 => x"fe",
          1160 => x"e6",
          1161 => x"38",
          1162 => x"90",
          1163 => x"59",
          1164 => x"7a",
          1165 => x"79",
          1166 => x"3f",
          1167 => x"05",
          1168 => x"08",
          1169 => x"88",
          1170 => x"08",
          1171 => x"ba",
          1172 => x"84",
          1173 => x"f4",
          1174 => x"53",
          1175 => x"84",
          1176 => x"90",
          1177 => x"38",
          1178 => x"fe",
          1179 => x"e5",
          1180 => x"38",
          1181 => x"2e",
          1182 => x"47",
          1183 => x"80",
          1184 => x"8c",
          1185 => x"5c",
          1186 => x"5c",
          1187 => x"07",
          1188 => x"79",
          1189 => x"83",
          1190 => x"d6",
          1191 => x"53",
          1192 => x"83",
          1193 => x"ef",
          1194 => x"84",
          1195 => x"53",
          1196 => x"84",
          1197 => x"38",
          1198 => x"05",
          1199 => x"ff",
          1200 => x"ba",
          1201 => x"64",
          1202 => x"70",
          1203 => x"3d",
          1204 => x"51",
          1205 => x"80",
          1206 => x"80",
          1207 => x"40",
          1208 => x"11",
          1209 => x"3f",
          1210 => x"f1",
          1211 => x"53",
          1212 => x"84",
          1213 => x"38",
          1214 => x"7c",
          1215 => x"39",
          1216 => x"80",
          1217 => x"8c",
          1218 => x"64",
          1219 => x"46",
          1220 => x"09",
          1221 => x"83",
          1222 => x"b8",
          1223 => x"8c",
          1224 => x"3f",
          1225 => x"d4",
          1226 => x"fe",
          1227 => x"e0",
          1228 => x"2e",
          1229 => x"05",
          1230 => x"78",
          1231 => x"33",
          1232 => x"83",
          1233 => x"83",
          1234 => x"a1",
          1235 => x"b5",
          1236 => x"3f",
          1237 => x"f0",
          1238 => x"cc",
          1239 => x"80",
          1240 => x"49",
          1241 => x"d3",
          1242 => x"92",
          1243 => x"83",
          1244 => x"83",
          1245 => x"9b",
          1246 => x"dd",
          1247 => x"80",
          1248 => x"47",
          1249 => x"5d",
          1250 => x"e8",
          1251 => x"8e",
          1252 => x"83",
          1253 => x"83",
          1254 => x"fb",
          1255 => x"05",
          1256 => x"80",
          1257 => x"94",
          1258 => x"80",
          1259 => x"ba",
          1260 => x"55",
          1261 => x"b5",
          1262 => x"77",
          1263 => x"56",
          1264 => x"da",
          1265 => x"2b",
          1266 => x"52",
          1267 => x"ba",
          1268 => x"83",
          1269 => x"80",
          1270 => x"81",
          1271 => x"83",
          1272 => x"5e",
          1273 => x"88",
          1274 => x"f0",
          1275 => x"3f",
          1276 => x"fc",
          1277 => x"fc",
          1278 => x"70",
          1279 => x"d3",
          1280 => x"15",
          1281 => x"f8",
          1282 => x"80",
          1283 => x"56",
          1284 => x"2e",
          1285 => x"ff",
          1286 => x"81",
          1287 => x"70",
          1288 => x"a0",
          1289 => x"54",
          1290 => x"52",
          1291 => x"72",
          1292 => x"54",
          1293 => x"70",
          1294 => x"86",
          1295 => x"73",
          1296 => x"2e",
          1297 => x"70",
          1298 => x"76",
          1299 => x"88",
          1300 => x"34",
          1301 => x"ba",
          1302 => x"80",
          1303 => x"be",
          1304 => x"70",
          1305 => x"a2",
          1306 => x"81",
          1307 => x"81",
          1308 => x"dc",
          1309 => x"08",
          1310 => x"0c",
          1311 => x"05",
          1312 => x"ba",
          1313 => x"84",
          1314 => x"fc",
          1315 => x"05",
          1316 => x"81",
          1317 => x"54",
          1318 => x"38",
          1319 => x"97",
          1320 => x"54",
          1321 => x"38",
          1322 => x"bb",
          1323 => x"55",
          1324 => x"d9",
          1325 => x"73",
          1326 => x"0b",
          1327 => x"87",
          1328 => x"87",
          1329 => x"87",
          1330 => x"87",
          1331 => x"87",
          1332 => x"87",
          1333 => x"98",
          1334 => x"0c",
          1335 => x"80",
          1336 => x"3d",
          1337 => x"87",
          1338 => x"87",
          1339 => x"23",
          1340 => x"82",
          1341 => x"5a",
          1342 => x"b0",
          1343 => x"c0",
          1344 => x"34",
          1345 => x"86",
          1346 => x"5c",
          1347 => x"a0",
          1348 => x"7d",
          1349 => x"7b",
          1350 => x"33",
          1351 => x"33",
          1352 => x"33",
          1353 => x"83",
          1354 => x"8f",
          1355 => x"93",
          1356 => x"38",
          1357 => x"ba",
          1358 => x"51",
          1359 => x"86",
          1360 => x"84",
          1361 => x"72",
          1362 => x"8c",
          1363 => x"52",
          1364 => x"38",
          1365 => x"ba",
          1366 => x"51",
          1367 => x"39",
          1368 => x"71",
          1369 => x"ce",
          1370 => x"70",
          1371 => x"eb",
          1372 => x"52",
          1373 => x"ba",
          1374 => x"3d",
          1375 => x"c4",
          1376 => x"55",
          1377 => x"c0",
          1378 => x"81",
          1379 => x"8c",
          1380 => x"51",
          1381 => x"81",
          1382 => x"71",
          1383 => x"38",
          1384 => x"94",
          1385 => x"87",
          1386 => x"74",
          1387 => x"04",
          1388 => x"51",
          1389 => x"06",
          1390 => x"93",
          1391 => x"c0",
          1392 => x"96",
          1393 => x"70",
          1394 => x"02",
          1395 => x"2a",
          1396 => x"34",
          1397 => x"78",
          1398 => x"57",
          1399 => x"15",
          1400 => x"06",
          1401 => x"ff",
          1402 => x"96",
          1403 => x"70",
          1404 => x"70",
          1405 => x"72",
          1406 => x"2e",
          1407 => x"52",
          1408 => x"51",
          1409 => x"2e",
          1410 => x"73",
          1411 => x"57",
          1412 => x"8c",
          1413 => x"2a",
          1414 => x"38",
          1415 => x"80",
          1416 => x"06",
          1417 => x"87",
          1418 => x"70",
          1419 => x"38",
          1420 => x"9e",
          1421 => x"52",
          1422 => x"87",
          1423 => x"0c",
          1424 => x"cc",
          1425 => x"f2",
          1426 => x"83",
          1427 => x"08",
          1428 => x"a0",
          1429 => x"9e",
          1430 => x"c0",
          1431 => x"87",
          1432 => x"0c",
          1433 => x"ec",
          1434 => x"f2",
          1435 => x"83",
          1436 => x"08",
          1437 => x"80",
          1438 => x"87",
          1439 => x"0c",
          1440 => x"84",
          1441 => x"f3",
          1442 => x"34",
          1443 => x"70",
          1444 => x"70",
          1445 => x"34",
          1446 => x"70",
          1447 => x"70",
          1448 => x"83",
          1449 => x"9e",
          1450 => x"51",
          1451 => x"81",
          1452 => x"0b",
          1453 => x"80",
          1454 => x"2e",
          1455 => x"90",
          1456 => x"08",
          1457 => x"52",
          1458 => x"71",
          1459 => x"c0",
          1460 => x"06",
          1461 => x"38",
          1462 => x"80",
          1463 => x"84",
          1464 => x"80",
          1465 => x"f3",
          1466 => x"90",
          1467 => x"52",
          1468 => x"52",
          1469 => x"87",
          1470 => x"80",
          1471 => x"83",
          1472 => x"34",
          1473 => x"70",
          1474 => x"70",
          1475 => x"83",
          1476 => x"9e",
          1477 => x"52",
          1478 => x"52",
          1479 => x"9e",
          1480 => x"2a",
          1481 => x"80",
          1482 => x"84",
          1483 => x"2e",
          1484 => x"99",
          1485 => x"f0",
          1486 => x"83",
          1487 => x"9e",
          1488 => x"52",
          1489 => x"71",
          1490 => x"90",
          1491 => x"9c",
          1492 => x"fd",
          1493 => x"8c",
          1494 => x"8c",
          1495 => x"d9",
          1496 => x"8e",
          1497 => x"f3",
          1498 => x"83",
          1499 => x"38",
          1500 => x"ff",
          1501 => x"84",
          1502 => x"75",
          1503 => x"54",
          1504 => x"33",
          1505 => x"8d",
          1506 => x"f3",
          1507 => x"83",
          1508 => x"38",
          1509 => x"f4",
          1510 => x"81",
          1511 => x"b3",
          1512 => x"d9",
          1513 => x"f2",
          1514 => x"ff",
          1515 => x"52",
          1516 => x"3f",
          1517 => x"83",
          1518 => x"51",
          1519 => x"08",
          1520 => x"ca",
          1521 => x"84",
          1522 => x"84",
          1523 => x"51",
          1524 => x"33",
          1525 => x"8e",
          1526 => x"c3",
          1527 => x"f3",
          1528 => x"75",
          1529 => x"08",
          1530 => x"54",
          1531 => x"db",
          1532 => x"51",
          1533 => x"83",
          1534 => x"52",
          1535 => x"8c",
          1536 => x"31",
          1537 => x"83",
          1538 => x"83",
          1539 => x"ff",
          1540 => x"f0",
          1541 => x"51",
          1542 => x"52",
          1543 => x"3f",
          1544 => x"ec",
          1545 => x"f8",
          1546 => x"b3",
          1547 => x"93",
          1548 => x"da",
          1549 => x"f3",
          1550 => x"75",
          1551 => x"08",
          1552 => x"54",
          1553 => x"da",
          1554 => x"f3",
          1555 => x"8d",
          1556 => x"51",
          1557 => x"33",
          1558 => x"fe",
          1559 => x"bf",
          1560 => x"75",
          1561 => x"83",
          1562 => x"83",
          1563 => x"fc",
          1564 => x"51",
          1565 => x"33",
          1566 => x"d7",
          1567 => x"dc",
          1568 => x"f3",
          1569 => x"86",
          1570 => x"52",
          1571 => x"3f",
          1572 => x"2e",
          1573 => x"98",
          1574 => x"b1",
          1575 => x"73",
          1576 => x"83",
          1577 => x"11",
          1578 => x"b1",
          1579 => x"75",
          1580 => x"83",
          1581 => x"11",
          1582 => x"b1",
          1583 => x"73",
          1584 => x"83",
          1585 => x"11",
          1586 => x"b0",
          1587 => x"74",
          1588 => x"83",
          1589 => x"11",
          1590 => x"b0",
          1591 => x"75",
          1592 => x"83",
          1593 => x"11",
          1594 => x"b0",
          1595 => x"73",
          1596 => x"83",
          1597 => x"83",
          1598 => x"83",
          1599 => x"f9",
          1600 => x"02",
          1601 => x"8c",
          1602 => x"05",
          1603 => x"51",
          1604 => x"04",
          1605 => x"3f",
          1606 => x"51",
          1607 => x"04",
          1608 => x"3f",
          1609 => x"51",
          1610 => x"04",
          1611 => x"3f",
          1612 => x"0c",
          1613 => x"0c",
          1614 => x"96",
          1615 => x"3d",
          1616 => x"70",
          1617 => x"08",
          1618 => x"8c",
          1619 => x"ff",
          1620 => x"80",
          1621 => x"3f",
          1622 => x"38",
          1623 => x"8c",
          1624 => x"84",
          1625 => x"ba",
          1626 => x"55",
          1627 => x"70",
          1628 => x"78",
          1629 => x"38",
          1630 => x"53",
          1631 => x"8c",
          1632 => x"38",
          1633 => x"0d",
          1634 => x"f0",
          1635 => x"e8",
          1636 => x"3f",
          1637 => x"3d",
          1638 => x"34",
          1639 => x"ad",
          1640 => x"0c",
          1641 => x"ab",
          1642 => x"5d",
          1643 => x"a0",
          1644 => x"3d",
          1645 => x"f4",
          1646 => x"bf",
          1647 => x"79",
          1648 => x"84",
          1649 => x"33",
          1650 => x"73",
          1651 => x"81",
          1652 => x"c2",
          1653 => x"0c",
          1654 => x"aa",
          1655 => x"05",
          1656 => x"08",
          1657 => x"78",
          1658 => x"ba",
          1659 => x"80",
          1660 => x"ff",
          1661 => x"fa",
          1662 => x"05",
          1663 => x"81",
          1664 => x"73",
          1665 => x"38",
          1666 => x"8d",
          1667 => x"84",
          1668 => x"08",
          1669 => x"ba",
          1670 => x"f8",
          1671 => x"82",
          1672 => x"80",
          1673 => x"d8",
          1674 => x"0b",
          1675 => x"84",
          1676 => x"58",
          1677 => x"52",
          1678 => x"ff",
          1679 => x"81",
          1680 => x"ba",
          1681 => x"3d",
          1682 => x"b9",
          1683 => x"b4",
          1684 => x"f3",
          1685 => x"74",
          1686 => x"80",
          1687 => x"91",
          1688 => x"57",
          1689 => x"90",
          1690 => x"5f",
          1691 => x"8c",
          1692 => x"56",
          1693 => x"ff",
          1694 => x"2b",
          1695 => x"70",
          1696 => x"2c",
          1697 => x"05",
          1698 => x"5c",
          1699 => x"81",
          1700 => x"78",
          1701 => x"80",
          1702 => x"98",
          1703 => x"cb",
          1704 => x"56",
          1705 => x"33",
          1706 => x"83",
          1707 => x"56",
          1708 => x"76",
          1709 => x"c4",
          1710 => x"99",
          1711 => x"98",
          1712 => x"2b",
          1713 => x"70",
          1714 => x"5f",
          1715 => x"7a",
          1716 => x"d1",
          1717 => x"76",
          1718 => x"29",
          1719 => x"70",
          1720 => x"95",
          1721 => x"70",
          1722 => x"de",
          1723 => x"25",
          1724 => x"18",
          1725 => x"ff",
          1726 => x"38",
          1727 => x"2e",
          1728 => x"56",
          1729 => x"e9",
          1730 => x"84",
          1731 => x"7f",
          1732 => x"b0",
          1733 => x"05",
          1734 => x"15",
          1735 => x"c8",
          1736 => x"d9",
          1737 => x"80",
          1738 => x"08",
          1739 => x"84",
          1740 => x"84",
          1741 => x"d1",
          1742 => x"d1",
          1743 => x"27",
          1744 => x"52",
          1745 => x"34",
          1746 => x"b5",
          1747 => x"2e",
          1748 => x"f3",
          1749 => x"8f",
          1750 => x"75",
          1751 => x"d1",
          1752 => x"b6",
          1753 => x"51",
          1754 => x"08",
          1755 => x"84",
          1756 => x"b5",
          1757 => x"05",
          1758 => x"81",
          1759 => x"51",
          1760 => x"d0",
          1761 => x"83",
          1762 => x"38",
          1763 => x"fc",
          1764 => x"38",
          1765 => x"a8",
          1766 => x"84",
          1767 => x"84",
          1768 => x"05",
          1769 => x"9a",
          1770 => x"d0",
          1771 => x"9e",
          1772 => x"51",
          1773 => x"08",
          1774 => x"84",
          1775 => x"b3",
          1776 => x"05",
          1777 => x"81",
          1778 => x"d0",
          1779 => x"cc",
          1780 => x"fa",
          1781 => x"81",
          1782 => x"7b",
          1783 => x"ae",
          1784 => x"ff",
          1785 => x"55",
          1786 => x"d5",
          1787 => x"84",
          1788 => x"52",
          1789 => x"d0",
          1790 => x"cc",
          1791 => x"ff",
          1792 => x"d0",
          1793 => x"74",
          1794 => x"5b",
          1795 => x"2b",
          1796 => x"43",
          1797 => x"38",
          1798 => x"ff",
          1799 => x"70",
          1800 => x"cc",
          1801 => x"24",
          1802 => x"52",
          1803 => x"81",
          1804 => x"70",
          1805 => x"56",
          1806 => x"84",
          1807 => x"b1",
          1808 => x"81",
          1809 => x"d1",
          1810 => x"25",
          1811 => x"16",
          1812 => x"d5",
          1813 => x"b1",
          1814 => x"81",
          1815 => x"d1",
          1816 => x"25",
          1817 => x"18",
          1818 => x"52",
          1819 => x"75",
          1820 => x"05",
          1821 => x"5b",
          1822 => x"38",
          1823 => x"55",
          1824 => x"d5",
          1825 => x"de",
          1826 => x"57",
          1827 => x"ff",
          1828 => x"33",
          1829 => x"d5",
          1830 => x"b6",
          1831 => x"f4",
          1832 => x"ff",
          1833 => x"d1",
          1834 => x"d8",
          1835 => x"10",
          1836 => x"5e",
          1837 => x"2b",
          1838 => x"81",
          1839 => x"ca",
          1840 => x"83",
          1841 => x"f3",
          1842 => x"74",
          1843 => x"56",
          1844 => x"f4",
          1845 => x"38",
          1846 => x"0b",
          1847 => x"8c",
          1848 => x"d0",
          1849 => x"84",
          1850 => x"af",
          1851 => x"a0",
          1852 => x"f0",
          1853 => x"3f",
          1854 => x"75",
          1855 => x"06",
          1856 => x"51",
          1857 => x"d1",
          1858 => x"34",
          1859 => x"0b",
          1860 => x"55",
          1861 => x"f0",
          1862 => x"3f",
          1863 => x"ff",
          1864 => x"52",
          1865 => x"d1",
          1866 => x"d1",
          1867 => x"74",
          1868 => x"9f",
          1869 => x"34",
          1870 => x"84",
          1871 => x"84",
          1872 => x"5c",
          1873 => x"84",
          1874 => x"84",
          1875 => x"84",
          1876 => x"52",
          1877 => x"d1",
          1878 => x"2c",
          1879 => x"56",
          1880 => x"d5",
          1881 => x"9e",
          1882 => x"2b",
          1883 => x"5d",
          1884 => x"f0",
          1885 => x"51",
          1886 => x"0a",
          1887 => x"2c",
          1888 => x"74",
          1889 => x"f0",
          1890 => x"3f",
          1891 => x"0a",
          1892 => x"33",
          1893 => x"b9",
          1894 => x"81",
          1895 => x"08",
          1896 => x"3f",
          1897 => x"0a",
          1898 => x"33",
          1899 => x"e6",
          1900 => x"77",
          1901 => x"33",
          1902 => x"80",
          1903 => x"98",
          1904 => x"5b",
          1905 => x"b6",
          1906 => x"ff",
          1907 => x"b8",
          1908 => x"75",
          1909 => x"98",
          1910 => x"38",
          1911 => x"34",
          1912 => x"0a",
          1913 => x"33",
          1914 => x"38",
          1915 => x"34",
          1916 => x"b3",
          1917 => x"33",
          1918 => x"17",
          1919 => x"57",
          1920 => x"0a",
          1921 => x"2c",
          1922 => x"58",
          1923 => x"98",
          1924 => x"06",
          1925 => x"a8",
          1926 => x"51",
          1927 => x"0a",
          1928 => x"2c",
          1929 => x"75",
          1930 => x"f0",
          1931 => x"3f",
          1932 => x"0a",
          1933 => x"33",
          1934 => x"b9",
          1935 => x"08",
          1936 => x"75",
          1937 => x"8c",
          1938 => x"8c",
          1939 => x"75",
          1940 => x"84",
          1941 => x"56",
          1942 => x"84",
          1943 => x"a9",
          1944 => x"a0",
          1945 => x"f0",
          1946 => x"3f",
          1947 => x"7a",
          1948 => x"06",
          1949 => x"da",
          1950 => x"f8",
          1951 => x"38",
          1952 => x"ca",
          1953 => x"08",
          1954 => x"ff",
          1955 => x"29",
          1956 => x"84",
          1957 => x"76",
          1958 => x"70",
          1959 => x"ff",
          1960 => x"25",
          1961 => x"f3",
          1962 => x"83",
          1963 => x"55",
          1964 => x"58",
          1965 => x"0b",
          1966 => x"08",
          1967 => x"74",
          1968 => x"f8",
          1969 => x"0b",
          1970 => x"3d",
          1971 => x"80",
          1972 => x"16",
          1973 => x"ff",
          1974 => x"ff",
          1975 => x"84",
          1976 => x"81",
          1977 => x"7b",
          1978 => x"84",
          1979 => x"57",
          1980 => x"38",
          1981 => x"ff",
          1982 => x"52",
          1983 => x"d5",
          1984 => x"e6",
          1985 => x"5a",
          1986 => x"ff",
          1987 => x"80",
          1988 => x"84",
          1989 => x"0c",
          1990 => x"a9",
          1991 => x"d1",
          1992 => x"ff",
          1993 => x"51",
          1994 => x"81",
          1995 => x"d1",
          1996 => x"80",
          1997 => x"08",
          1998 => x"84",
          1999 => x"a5",
          2000 => x"88",
          2001 => x"d0",
          2002 => x"d0",
          2003 => x"39",
          2004 => x"ba",
          2005 => x"ba",
          2006 => x"53",
          2007 => x"3f",
          2008 => x"d1",
          2009 => x"58",
          2010 => x"38",
          2011 => x"ff",
          2012 => x"52",
          2013 => x"d5",
          2014 => x"f6",
          2015 => x"41",
          2016 => x"ff",
          2017 => x"d7",
          2018 => x"82",
          2019 => x"05",
          2020 => x"80",
          2021 => x"7b",
          2022 => x"10",
          2023 => x"41",
          2024 => x"75",
          2025 => x"9a",
          2026 => x"70",
          2027 => x"27",
          2028 => x"34",
          2029 => x"05",
          2030 => x"81",
          2031 => x"52",
          2032 => x"f3",
          2033 => x"80",
          2034 => x"84",
          2035 => x"0c",
          2036 => x"52",
          2037 => x"c7",
          2038 => x"38",
          2039 => x"5d",
          2040 => x"52",
          2041 => x"ba",
          2042 => x"7b",
          2043 => x"84",
          2044 => x"3f",
          2045 => x"84",
          2046 => x"84",
          2047 => x"58",
          2048 => x"06",
          2049 => x"83",
          2050 => x"58",
          2051 => x"2b",
          2052 => x"81",
          2053 => x"9a",
          2054 => x"83",
          2055 => x"f3",
          2056 => x"74",
          2057 => x"06",
          2058 => x"80",
          2059 => x"fe",
          2060 => x"e6",
          2061 => x"ff",
          2062 => x"81",
          2063 => x"93",
          2064 => x"83",
          2065 => x"51",
          2066 => x"33",
          2067 => x"f3",
          2068 => x"56",
          2069 => x"8c",
          2070 => x"70",
          2071 => x"08",
          2072 => x"82",
          2073 => x"fc",
          2074 => x"fc",
          2075 => x"51",
          2076 => x"38",
          2077 => x"80",
          2078 => x"c7",
          2079 => x"81",
          2080 => x"38",
          2081 => x"82",
          2082 => x"80",
          2083 => x"57",
          2084 => x"2e",
          2085 => x"75",
          2086 => x"ba",
          2087 => x"2b",
          2088 => x"07",
          2089 => x"5b",
          2090 => x"70",
          2091 => x"84",
          2092 => x"38",
          2093 => x"b8",
          2094 => x"31",
          2095 => x"15",
          2096 => x"34",
          2097 => x"3d",
          2098 => x"83",
          2099 => x"83",
          2100 => x"74",
          2101 => x"a3",
          2102 => x"70",
          2103 => x"70",
          2104 => x"70",
          2105 => x"5d",
          2106 => x"73",
          2107 => x"75",
          2108 => x"81",
          2109 => x"83",
          2110 => x"70",
          2111 => x"5b",
          2112 => x"f9",
          2113 => x"7d",
          2114 => x"5c",
          2115 => x"7d",
          2116 => x"38",
          2117 => x"83",
          2118 => x"56",
          2119 => x"59",
          2120 => x"80",
          2121 => x"ff",
          2122 => x"ba",
          2123 => x"57",
          2124 => x"81",
          2125 => x"81",
          2126 => x"54",
          2127 => x"80",
          2128 => x"83",
          2129 => x"70",
          2130 => x"88",
          2131 => x"56",
          2132 => x"38",
          2133 => x"83",
          2134 => x"70",
          2135 => x"71",
          2136 => x"11",
          2137 => x"a3",
          2138 => x"33",
          2139 => x"33",
          2140 => x"22",
          2141 => x"29",
          2142 => x"5f",
          2143 => x"38",
          2144 => x"19",
          2145 => x"81",
          2146 => x"ff",
          2147 => x"75",
          2148 => x"7b",
          2149 => x"53",
          2150 => x"5b",
          2151 => x"06",
          2152 => x"39",
          2153 => x"9a",
          2154 => x"9c",
          2155 => x"74",
          2156 => x"73",
          2157 => x"94",
          2158 => x"ff",
          2159 => x"55",
          2160 => x"85",
          2161 => x"83",
          2162 => x"e0",
          2163 => x"87",
          2164 => x"07",
          2165 => x"70",
          2166 => x"53",
          2167 => x"08",
          2168 => x"72",
          2169 => x"81",
          2170 => x"34",
          2171 => x"80",
          2172 => x"0d",
          2173 => x"8c",
          2174 => x"05",
          2175 => x"84",
          2176 => x"53",
          2177 => x"b8",
          2178 => x"f9",
          2179 => x"a3",
          2180 => x"5f",
          2181 => x"70",
          2182 => x"33",
          2183 => x"83",
          2184 => x"05",
          2185 => x"f9",
          2186 => x"06",
          2187 => x"72",
          2188 => x"53",
          2189 => x"ba",
          2190 => x"b7",
          2191 => x"26",
          2192 => x"76",
          2193 => x"9f",
          2194 => x"70",
          2195 => x"e0",
          2196 => x"54",
          2197 => x"81",
          2198 => x"e3",
          2199 => x"83",
          2200 => x"54",
          2201 => x"74",
          2202 => x"14",
          2203 => x"84",
          2204 => x"83",
          2205 => x"ff",
          2206 => x"54",
          2207 => x"74",
          2208 => x"71",
          2209 => x"87",
          2210 => x"80",
          2211 => x"06",
          2212 => x"57",
          2213 => x"de",
          2214 => x"84",
          2215 => x"05",
          2216 => x"33",
          2217 => x"15",
          2218 => x"33",
          2219 => x"55",
          2220 => x"72",
          2221 => x"04",
          2222 => x"ba",
          2223 => x"b7",
          2224 => x"27",
          2225 => x"dd",
          2226 => x"83",
          2227 => x"2e",
          2228 => x"76",
          2229 => x"71",
          2230 => x"52",
          2231 => x"38",
          2232 => x"15",
          2233 => x"0b",
          2234 => x"81",
          2235 => x"80",
          2236 => x"e0",
          2237 => x"57",
          2238 => x"fd",
          2239 => x"33",
          2240 => x"be",
          2241 => x"33",
          2242 => x"fc",
          2243 => x"84",
          2244 => x"86",
          2245 => x"c4",
          2246 => x"b8",
          2247 => x"38",
          2248 => x"84",
          2249 => x"80",
          2250 => x"bc",
          2251 => x"72",
          2252 => x"70",
          2253 => x"ba",
          2254 => x"f9",
          2255 => x"70",
          2256 => x"54",
          2257 => x"83",
          2258 => x"ff",
          2259 => x"75",
          2260 => x"f9",
          2261 => x"0c",
          2262 => x"33",
          2263 => x"2c",
          2264 => x"83",
          2265 => x"8c",
          2266 => x"bd",
          2267 => x"ff",
          2268 => x"83",
          2269 => x"34",
          2270 => x"3d",
          2271 => x"34",
          2272 => x"33",
          2273 => x"fe",
          2274 => x"f9",
          2275 => x"0d",
          2276 => x"26",
          2277 => x"d0",
          2278 => x"b8",
          2279 => x"2b",
          2280 => x"07",
          2281 => x"2e",
          2282 => x"0b",
          2283 => x"ba",
          2284 => x"f9",
          2285 => x"51",
          2286 => x"84",
          2287 => x"83",
          2288 => x"70",
          2289 => x"f9",
          2290 => x"51",
          2291 => x"80",
          2292 => x"0b",
          2293 => x"04",
          2294 => x"84",
          2295 => x"ff",
          2296 => x"07",
          2297 => x"a5",
          2298 => x"06",
          2299 => x"34",
          2300 => x"81",
          2301 => x"f9",
          2302 => x"b8",
          2303 => x"70",
          2304 => x"83",
          2305 => x"70",
          2306 => x"83",
          2307 => x"d0",
          2308 => x"fe",
          2309 => x"bf",
          2310 => x"b8",
          2311 => x"33",
          2312 => x"70",
          2313 => x"83",
          2314 => x"c0",
          2315 => x"fe",
          2316 => x"af",
          2317 => x"b8",
          2318 => x"33",
          2319 => x"b8",
          2320 => x"33",
          2321 => x"83",
          2322 => x"3d",
          2323 => x"05",
          2324 => x"33",
          2325 => x"33",
          2326 => x"5d",
          2327 => x"38",
          2328 => x"2e",
          2329 => x"34",
          2330 => x"83",
          2331 => x"23",
          2332 => x"0d",
          2333 => x"db",
          2334 => x"81",
          2335 => x"83",
          2336 => x"bd",
          2337 => x"79",
          2338 => x"b7",
          2339 => x"55",
          2340 => x"e3",
          2341 => x"84",
          2342 => x"84",
          2343 => x"83",
          2344 => x"34",
          2345 => x"b8",
          2346 => x"34",
          2347 => x"0b",
          2348 => x"f9",
          2349 => x"84",
          2350 => x"33",
          2351 => x"7a",
          2352 => x"80",
          2353 => x"5a",
          2354 => x"10",
          2355 => x"59",
          2356 => x"3f",
          2357 => x"b9",
          2358 => x"26",
          2359 => x"80",
          2360 => x"80",
          2361 => x"f9",
          2362 => x"7c",
          2363 => x"04",
          2364 => x"0b",
          2365 => x"f9",
          2366 => x"34",
          2367 => x"f7",
          2368 => x"ba",
          2369 => x"fe",
          2370 => x"f0",
          2371 => x"ba",
          2372 => x"f7",
          2373 => x"51",
          2374 => x"81",
          2375 => x"3d",
          2376 => x"33",
          2377 => x"33",
          2378 => x"12",
          2379 => x"ba",
          2380 => x"29",
          2381 => x"f8",
          2382 => x"57",
          2383 => x"89",
          2384 => x"81",
          2385 => x"38",
          2386 => x"b8",
          2387 => x"f9",
          2388 => x"56",
          2389 => x"a3",
          2390 => x"33",
          2391 => x"22",
          2392 => x"53",
          2393 => x"f9",
          2394 => x"54",
          2395 => x"80",
          2396 => x"81",
          2397 => x"f9",
          2398 => x"5b",
          2399 => x"84",
          2400 => x"81",
          2401 => x"81",
          2402 => x"77",
          2403 => x"83",
          2404 => x"53",
          2405 => x"84",
          2406 => x"38",
          2407 => x"3d",
          2408 => x"75",
          2409 => x"2e",
          2410 => x"52",
          2411 => x"83",
          2412 => x"f9",
          2413 => x"13",
          2414 => x"81",
          2415 => x"52",
          2416 => x"70",
          2417 => x"26",
          2418 => x"fd",
          2419 => x"06",
          2420 => x"fe",
          2421 => x"fe",
          2422 => x"de",
          2423 => x"89",
          2424 => x"09",
          2425 => x"bd",
          2426 => x"05",
          2427 => x"83",
          2428 => x"fc",
          2429 => x"81",
          2430 => x"fe",
          2431 => x"bd",
          2432 => x"f9",
          2433 => x"e2",
          2434 => x"51",
          2435 => x"3d",
          2436 => x"b9",
          2437 => x"81",
          2438 => x"38",
          2439 => x"8a",
          2440 => x"84",
          2441 => x"38",
          2442 => x"33",
          2443 => x"05",
          2444 => x"33",
          2445 => x"b8",
          2446 => x"f9",
          2447 => x"5a",
          2448 => x"34",
          2449 => x"62",
          2450 => x"7f",
          2451 => x"b8",
          2452 => x"f9",
          2453 => x"72",
          2454 => x"83",
          2455 => x"34",
          2456 => x"58",
          2457 => x"b8",
          2458 => x"ff",
          2459 => x"80",
          2460 => x"0d",
          2461 => x"b7",
          2462 => x"2e",
          2463 => x"89",
          2464 => x"0c",
          2465 => x"33",
          2466 => x"05",
          2467 => x"33",
          2468 => x"b8",
          2469 => x"f9",
          2470 => x"5f",
          2471 => x"34",
          2472 => x"19",
          2473 => x"a3",
          2474 => x"33",
          2475 => x"22",
          2476 => x"11",
          2477 => x"b8",
          2478 => x"81",
          2479 => x"60",
          2480 => x"f9",
          2481 => x"0c",
          2482 => x"82",
          2483 => x"38",
          2484 => x"a8",
          2485 => x"80",
          2486 => x"0d",
          2487 => x"d0",
          2488 => x"38",
          2489 => x"57",
          2490 => x"b9",
          2491 => x"59",
          2492 => x"80",
          2493 => x"0d",
          2494 => x"80",
          2495 => x"80",
          2496 => x"bd",
          2497 => x"40",
          2498 => x"a0",
          2499 => x"83",
          2500 => x"72",
          2501 => x"78",
          2502 => x"bc",
          2503 => x"83",
          2504 => x"1b",
          2505 => x"ff",
          2506 => x"bd",
          2507 => x"43",
          2508 => x"84",
          2509 => x"fe",
          2510 => x"fa",
          2511 => x"fe",
          2512 => x"f9",
          2513 => x"f9",
          2514 => x"a3",
          2515 => x"40",
          2516 => x"83",
          2517 => x"5a",
          2518 => x"86",
          2519 => x"1a",
          2520 => x"56",
          2521 => x"39",
          2522 => x"0b",
          2523 => x"b9",
          2524 => x"34",
          2525 => x"0b",
          2526 => x"04",
          2527 => x"34",
          2528 => x"34",
          2529 => x"34",
          2530 => x"0b",
          2531 => x"04",
          2532 => x"fa",
          2533 => x"b8",
          2534 => x"f9",
          2535 => x"75",
          2536 => x"83",
          2537 => x"29",
          2538 => x"f8",
          2539 => x"5b",
          2540 => x"78",
          2541 => x"75",
          2542 => x"bd",
          2543 => x"ff",
          2544 => x"29",
          2545 => x"33",
          2546 => x"b8",
          2547 => x"f9",
          2548 => x"5e",
          2549 => x"18",
          2550 => x"29",
          2551 => x"33",
          2552 => x"b8",
          2553 => x"f9",
          2554 => x"72",
          2555 => x"83",
          2556 => x"05",
          2557 => x"5c",
          2558 => x"84",
          2559 => x"38",
          2560 => x"34",
          2561 => x"06",
          2562 => x"78",
          2563 => x"2e",
          2564 => x"a8",
          2565 => x"83",
          2566 => x"b4",
          2567 => x"83",
          2568 => x"80",
          2569 => x"81",
          2570 => x"ba",
          2571 => x"f9",
          2572 => x"81",
          2573 => x"81",
          2574 => x"a3",
          2575 => x"5c",
          2576 => x"ff",
          2577 => x"53",
          2578 => x"2e",
          2579 => x"ff",
          2580 => x"ff",
          2581 => x"40",
          2582 => x"80",
          2583 => x"f9",
          2584 => x"71",
          2585 => x"0b",
          2586 => x"bc",
          2587 => x"83",
          2588 => x"1a",
          2589 => x"ff",
          2590 => x"bd",
          2591 => x"5a",
          2592 => x"98",
          2593 => x"81",
          2594 => x"81",
          2595 => x"77",
          2596 => x"83",
          2597 => x"ff",
          2598 => x"a7",
          2599 => x"80",
          2600 => x"ff",
          2601 => x"ff",
          2602 => x"43",
          2603 => x"87",
          2604 => x"80",
          2605 => x"ba",
          2606 => x"5e",
          2607 => x"34",
          2608 => x"1e",
          2609 => x"a3",
          2610 => x"33",
          2611 => x"22",
          2612 => x"11",
          2613 => x"b8",
          2614 => x"81",
          2615 => x"79",
          2616 => x"f9",
          2617 => x"84",
          2618 => x"8c",
          2619 => x"be",
          2620 => x"33",
          2621 => x"81",
          2622 => x"ca",
          2623 => x"80",
          2624 => x"0d",
          2625 => x"84",
          2626 => x"f9",
          2627 => x"f9",
          2628 => x"fc",
          2629 => x"3d",
          2630 => x"8a",
          2631 => x"2e",
          2632 => x"81",
          2633 => x"34",
          2634 => x"80",
          2635 => x"05",
          2636 => x"17",
          2637 => x"7b",
          2638 => x"80",
          2639 => x"5c",
          2640 => x"83",
          2641 => x"72",
          2642 => x"b8",
          2643 => x"80",
          2644 => x"f9",
          2645 => x"71",
          2646 => x"83",
          2647 => x"33",
          2648 => x"f9",
          2649 => x"05",
          2650 => x"ff",
          2651 => x"bd",
          2652 => x"5a",
          2653 => x"98",
          2654 => x"ff",
          2655 => x"a2",
          2656 => x"90",
          2657 => x"f9",
          2658 => x"0c",
          2659 => x"2e",
          2660 => x"56",
          2661 => x"51",
          2662 => x"8c",
          2663 => x"f4",
          2664 => x"f5",
          2665 => x"f6",
          2666 => x"ff",
          2667 => x"b9",
          2668 => x"b9",
          2669 => x"b9",
          2670 => x"8d",
          2671 => x"38",
          2672 => x"2e",
          2673 => x"f9",
          2674 => x"bc",
          2675 => x"e4",
          2676 => x"fe",
          2677 => x"f8",
          2678 => x"06",
          2679 => x"41",
          2680 => x"52",
          2681 => x"3f",
          2682 => x"8d",
          2683 => x"5b",
          2684 => x"10",
          2685 => x"57",
          2686 => x"75",
          2687 => x"7e",
          2688 => x"7d",
          2689 => x"bc",
          2690 => x"31",
          2691 => x"5a",
          2692 => x"bc",
          2693 => x"33",
          2694 => x"84",
          2695 => x"ff",
          2696 => x"5f",
          2697 => x"83",
          2698 => x"0b",
          2699 => x"33",
          2700 => x"80",
          2701 => x"75",
          2702 => x"80",
          2703 => x"bc",
          2704 => x"57",
          2705 => x"81",
          2706 => x"fc",
          2707 => x"7f",
          2708 => x"bd",
          2709 => x"31",
          2710 => x"5a",
          2711 => x"bd",
          2712 => x"33",
          2713 => x"84",
          2714 => x"09",
          2715 => x"80",
          2716 => x"bc",
          2717 => x"a0",
          2718 => x"51",
          2719 => x"83",
          2720 => x"87",
          2721 => x"5d",
          2722 => x"38",
          2723 => x"f2",
          2724 => x"80",
          2725 => x"22",
          2726 => x"fb",
          2727 => x"34",
          2728 => x"56",
          2729 => x"b9",
          2730 => x"7c",
          2731 => x"59",
          2732 => x"75",
          2733 => x"a2",
          2734 => x"80",
          2735 => x"33",
          2736 => x"84",
          2737 => x"56",
          2738 => x"76",
          2739 => x"83",
          2740 => x"80",
          2741 => x"76",
          2742 => x"84",
          2743 => x"83",
          2744 => x"81",
          2745 => x"8d",
          2746 => x"0b",
          2747 => x"80",
          2748 => x"56",
          2749 => x"81",
          2750 => x"f3",
          2751 => x"33",
          2752 => x"84",
          2753 => x"ff",
          2754 => x"70",
          2755 => x"70",
          2756 => x"52",
          2757 => x"83",
          2758 => x"23",
          2759 => x"5f",
          2760 => x"76",
          2761 => x"33",
          2762 => x"f9",
          2763 => x"bd",
          2764 => x"33",
          2765 => x"84",
          2766 => x"40",
          2767 => x"83",
          2768 => x"70",
          2769 => x"71",
          2770 => x"05",
          2771 => x"7e",
          2772 => x"83",
          2773 => x"5f",
          2774 => x"79",
          2775 => x"5d",
          2776 => x"84",
          2777 => x"8e",
          2778 => x"f9",
          2779 => x"7c",
          2780 => x"e5",
          2781 => x"76",
          2782 => x"75",
          2783 => x"06",
          2784 => x"5a",
          2785 => x"31",
          2786 => x"71",
          2787 => x"a3",
          2788 => x"7f",
          2789 => x"71",
          2790 => x"79",
          2791 => x"de",
          2792 => x"84",
          2793 => x"05",
          2794 => x"33",
          2795 => x"18",
          2796 => x"33",
          2797 => x"58",
          2798 => x"e0",
          2799 => x"33",
          2800 => x"70",
          2801 => x"05",
          2802 => x"33",
          2803 => x"1d",
          2804 => x"ff",
          2805 => x"8d",
          2806 => x"38",
          2807 => x"d8",
          2808 => x"84",
          2809 => x"8d",
          2810 => x"2e",
          2811 => x"75",
          2812 => x"38",
          2813 => x"ff",
          2814 => x"5c",
          2815 => x"84",
          2816 => x"f6",
          2817 => x"60",
          2818 => x"26",
          2819 => x"f2",
          2820 => x"29",
          2821 => x"70",
          2822 => x"05",
          2823 => x"8b",
          2824 => x"8b",
          2825 => x"98",
          2826 => x"2b",
          2827 => x"5f",
          2828 => x"77",
          2829 => x"70",
          2830 => x"ee",
          2831 => x"ff",
          2832 => x"60",
          2833 => x"7d",
          2834 => x"5a",
          2835 => x"31",
          2836 => x"40",
          2837 => x"26",
          2838 => x"84",
          2839 => x"e0",
          2840 => x"05",
          2841 => x"26",
          2842 => x"19",
          2843 => x"34",
          2844 => x"38",
          2845 => x"ff",
          2846 => x"f9",
          2847 => x"84",
          2848 => x"07",
          2849 => x"09",
          2850 => x"83",
          2851 => x"ff",
          2852 => x"f9",
          2853 => x"1e",
          2854 => x"84",
          2855 => x"84",
          2856 => x"fa",
          2857 => x"07",
          2858 => x"18",
          2859 => x"fb",
          2860 => x"06",
          2861 => x"34",
          2862 => x"fb",
          2863 => x"b8",
          2864 => x"81",
          2865 => x"f9",
          2866 => x"33",
          2867 => x"83",
          2868 => x"f1",
          2869 => x"70",
          2870 => x"39",
          2871 => x"56",
          2872 => x"39",
          2873 => x"90",
          2874 => x"fe",
          2875 => x"ef",
          2876 => x"f9",
          2877 => x"b8",
          2878 => x"56",
          2879 => x"39",
          2880 => x"a0",
          2881 => x"fe",
          2882 => x"fe",
          2883 => x"b8",
          2884 => x"33",
          2885 => x"83",
          2886 => x"f9",
          2887 => x"56",
          2888 => x"39",
          2889 => x"56",
          2890 => x"39",
          2891 => x"56",
          2892 => x"39",
          2893 => x"56",
          2894 => x"39",
          2895 => x"80",
          2896 => x"34",
          2897 => x"81",
          2898 => x"f9",
          2899 => x"83",
          2900 => x"d2",
          2901 => x"f4",
          2902 => x"f5",
          2903 => x"f6",
          2904 => x"80",
          2905 => x"39",
          2906 => x"0b",
          2907 => x"04",
          2908 => x"bd",
          2909 => x"05",
          2910 => x"42",
          2911 => x"51",
          2912 => x"08",
          2913 => x"b9",
          2914 => x"34",
          2915 => x"3d",
          2916 => x"ef",
          2917 => x"11",
          2918 => x"7b",
          2919 => x"ca",
          2920 => x"80",
          2921 => x"80",
          2922 => x"81",
          2923 => x"33",
          2924 => x"56",
          2925 => x"bd",
          2926 => x"3f",
          2927 => x"de",
          2928 => x"33",
          2929 => x"72",
          2930 => x"75",
          2931 => x"80",
          2932 => x"38",
          2933 => x"39",
          2934 => x"09",
          2935 => x"57",
          2936 => x"81",
          2937 => x"59",
          2938 => x"38",
          2939 => x"ff",
          2940 => x"81",
          2941 => x"bc",
          2942 => x"ff",
          2943 => x"29",
          2944 => x"f9",
          2945 => x"05",
          2946 => x"92",
          2947 => x"77",
          2948 => x"ff",
          2949 => x"7b",
          2950 => x"33",
          2951 => x"ff",
          2952 => x"7c",
          2953 => x"80",
          2954 => x"ff",
          2955 => x"38",
          2956 => x"34",
          2957 => x"22",
          2958 => x"90",
          2959 => x"81",
          2960 => x"5f",
          2961 => x"87",
          2962 => x"7f",
          2963 => x"41",
          2964 => x"ea",
          2965 => x"e0",
          2966 => x"33",
          2967 => x"70",
          2968 => x"05",
          2969 => x"33",
          2970 => x"1d",
          2971 => x"ec",
          2972 => x"84",
          2973 => x"05",
          2974 => x"33",
          2975 => x"18",
          2976 => x"33",
          2977 => x"58",
          2978 => x"fa",
          2979 => x"84",
          2980 => x"f9",
          2981 => x"f9",
          2982 => x"5c",
          2983 => x"d2",
          2984 => x"ff",
          2985 => x"61",
          2986 => x"f9",
          2987 => x"19",
          2988 => x"80",
          2989 => x"b8",
          2990 => x"12",
          2991 => x"8d",
          2992 => x"34",
          2993 => x"81",
          2994 => x"59",
          2995 => x"38",
          2996 => x"2e",
          2997 => x"f9",
          2998 => x"f9",
          2999 => x"76",
          3000 => x"38",
          3001 => x"83",
          3002 => x"1a",
          3003 => x"e7",
          3004 => x"f9",
          3005 => x"58",
          3006 => x"80",
          3007 => x"f9",
          3008 => x"34",
          3009 => x"76",
          3010 => x"b8",
          3011 => x"79",
          3012 => x"79",
          3013 => x"23",
          3014 => x"bc",
          3015 => x"ba",
          3016 => x"f9",
          3017 => x"83",
          3018 => x"f9",
          3019 => x"1a",
          3020 => x"91",
          3021 => x"02",
          3022 => x"54",
          3023 => x"51",
          3024 => x"8c",
          3025 => x"73",
          3026 => x"ba",
          3027 => x"3d",
          3028 => x"0b",
          3029 => x"06",
          3030 => x"55",
          3031 => x"81",
          3032 => x"74",
          3033 => x"3d",
          3034 => x"82",
          3035 => x"73",
          3036 => x"70",
          3037 => x"83",
          3038 => x"7b",
          3039 => x"7b",
          3040 => x"80",
          3041 => x"80",
          3042 => x"33",
          3043 => x"33",
          3044 => x"80",
          3045 => x"5d",
          3046 => x"ff",
          3047 => x"55",
          3048 => x"81",
          3049 => x"34",
          3050 => x"87",
          3051 => x"2e",
          3052 => x"57",
          3053 => x"14",
          3054 => x"f9",
          3055 => x"f7",
          3056 => x"83",
          3057 => x"72",
          3058 => x"ff",
          3059 => x"c0",
          3060 => x"79",
          3061 => x"83",
          3062 => x"14",
          3063 => x"14",
          3064 => x"74",
          3065 => x"33",
          3066 => x"56",
          3067 => x"81",
          3068 => x"70",
          3069 => x"2e",
          3070 => x"e5",
          3071 => x"80",
          3072 => x"f7",
          3073 => x"33",
          3074 => x"33",
          3075 => x"e7",
          3076 => x"56",
          3077 => x"81",
          3078 => x"16",
          3079 => x"38",
          3080 => x"81",
          3081 => x"16",
          3082 => x"81",
          3083 => x"8d",
          3084 => x"72",
          3085 => x"ff",
          3086 => x"8c",
          3087 => x"81",
          3088 => x"e0",
          3089 => x"9c",
          3090 => x"ec",
          3091 => x"08",
          3092 => x"70",
          3093 => x"27",
          3094 => x"34",
          3095 => x"19",
          3096 => x"72",
          3097 => x"79",
          3098 => x"73",
          3099 => x"87",
          3100 => x"7d",
          3101 => x"f8",
          3102 => x"83",
          3103 => x"34",
          3104 => x"94",
          3105 => x"81",
          3106 => x"33",
          3107 => x"34",
          3108 => x"f7",
          3109 => x"9c",
          3110 => x"80",
          3111 => x"8a",
          3112 => x"74",
          3113 => x"9b",
          3114 => x"83",
          3115 => x"38",
          3116 => x"81",
          3117 => x"98",
          3118 => x"38",
          3119 => x"70",
          3120 => x"06",
          3121 => x"53",
          3122 => x"38",
          3123 => x"76",
          3124 => x"9c",
          3125 => x"87",
          3126 => x"0c",
          3127 => x"81",
          3128 => x"06",
          3129 => x"9b",
          3130 => x"80",
          3131 => x"72",
          3132 => x"32",
          3133 => x"40",
          3134 => x"2e",
          3135 => x"ff",
          3136 => x"10",
          3137 => x"33",
          3138 => x"38",
          3139 => x"57",
          3140 => x"83",
          3141 => x"38",
          3142 => x"91",
          3143 => x"51",
          3144 => x"0c",
          3145 => x"81",
          3146 => x"ff",
          3147 => x"33",
          3148 => x"15",
          3149 => x"f7",
          3150 => x"c0",
          3151 => x"15",
          3152 => x"06",
          3153 => x"38",
          3154 => x"75",
          3155 => x"06",
          3156 => x"fb",
          3157 => x"fa",
          3158 => x"55",
          3159 => x"c0",
          3160 => x"76",
          3161 => x"ff",
          3162 => x"ca",
          3163 => x"09",
          3164 => x"72",
          3165 => x"f7",
          3166 => x"f7",
          3167 => x"83",
          3168 => x"5c",
          3169 => x"2e",
          3170 => x"59",
          3171 => x"81",
          3172 => x"fd",
          3173 => x"54",
          3174 => x"83",
          3175 => x"54",
          3176 => x"f7",
          3177 => x"33",
          3178 => x"73",
          3179 => x"95",
          3180 => x"84",
          3181 => x"f7",
          3182 => x"ff",
          3183 => x"57",
          3184 => x"80",
          3185 => x"81",
          3186 => x"73",
          3187 => x"f9",
          3188 => x"81",
          3189 => x"75",
          3190 => x"f9",
          3191 => x"81",
          3192 => x"ff",
          3193 => x"95",
          3194 => x"f0",
          3195 => x"83",
          3196 => x"59",
          3197 => x"51",
          3198 => x"f9",
          3199 => x"08",
          3200 => x"14",
          3201 => x"e0",
          3202 => x"08",
          3203 => x"80",
          3204 => x"c0",
          3205 => x"56",
          3206 => x"98",
          3207 => x"08",
          3208 => x"15",
          3209 => x"53",
          3210 => x"fe",
          3211 => x"08",
          3212 => x"cd",
          3213 => x"c5",
          3214 => x"ce",
          3215 => x"08",
          3216 => x"75",
          3217 => x"87",
          3218 => x"74",
          3219 => x"db",
          3220 => x"ff",
          3221 => x"56",
          3222 => x"2e",
          3223 => x"72",
          3224 => x"38",
          3225 => x"0d",
          3226 => x"58",
          3227 => x"e4",
          3228 => x"77",
          3229 => x"04",
          3230 => x"a7",
          3231 => x"f4",
          3232 => x"80",
          3233 => x"51",
          3234 => x"73",
          3235 => x"72",
          3236 => x"73",
          3237 => x"53",
          3238 => x"08",
          3239 => x"83",
          3240 => x"81",
          3241 => x"e8",
          3242 => x"f4",
          3243 => x"54",
          3244 => x"c0",
          3245 => x"f6",
          3246 => x"9c",
          3247 => x"38",
          3248 => x"c0",
          3249 => x"74",
          3250 => x"ff",
          3251 => x"9c",
          3252 => x"c0",
          3253 => x"9c",
          3254 => x"81",
          3255 => x"53",
          3256 => x"81",
          3257 => x"a4",
          3258 => x"80",
          3259 => x"80",
          3260 => x"38",
          3261 => x"d5",
          3262 => x"57",
          3263 => x"84",
          3264 => x"27",
          3265 => x"33",
          3266 => x"72",
          3267 => x"0c",
          3268 => x"e4",
          3269 => x"77",
          3270 => x"04",
          3271 => x"54",
          3272 => x"ab",
          3273 => x"05",
          3274 => x"83",
          3275 => x"fc",
          3276 => x"07",
          3277 => x"34",
          3278 => x"34",
          3279 => x"34",
          3280 => x"98",
          3281 => x"57",
          3282 => x"38",
          3283 => x"70",
          3284 => x"f0",
          3285 => x"82",
          3286 => x"80",
          3287 => x"98",
          3288 => x"34",
          3289 => x"87",
          3290 => x"08",
          3291 => x"c0",
          3292 => x"9c",
          3293 => x"81",
          3294 => x"57",
          3295 => x"81",
          3296 => x"a4",
          3297 => x"80",
          3298 => x"80",
          3299 => x"80",
          3300 => x"9c",
          3301 => x"56",
          3302 => x"33",
          3303 => x"71",
          3304 => x"2e",
          3305 => x"52",
          3306 => x"72",
          3307 => x"80",
          3308 => x"53",
          3309 => x"ff",
          3310 => x"84",
          3311 => x"ff",
          3312 => x"76",
          3313 => x"56",
          3314 => x"0b",
          3315 => x"d3",
          3316 => x"3d",
          3317 => x"98",
          3318 => x"0b",
          3319 => x"0b",
          3320 => x"80",
          3321 => x"83",
          3322 => x"05",
          3323 => x"87",
          3324 => x"2e",
          3325 => x"98",
          3326 => x"87",
          3327 => x"87",
          3328 => x"70",
          3329 => x"71",
          3330 => x"98",
          3331 => x"87",
          3332 => x"98",
          3333 => x"38",
          3334 => x"08",
          3335 => x"71",
          3336 => x"98",
          3337 => x"27",
          3338 => x"91",
          3339 => x"81",
          3340 => x"ff",
          3341 => x"57",
          3342 => x"e5",
          3343 => x"3d",
          3344 => x"fc",
          3345 => x"83",
          3346 => x"11",
          3347 => x"2b",
          3348 => x"33",
          3349 => x"90",
          3350 => x"5d",
          3351 => x"71",
          3352 => x"11",
          3353 => x"71",
          3354 => x"81",
          3355 => x"2b",
          3356 => x"52",
          3357 => x"13",
          3358 => x"71",
          3359 => x"2a",
          3360 => x"34",
          3361 => x"13",
          3362 => x"84",
          3363 => x"2b",
          3364 => x"54",
          3365 => x"14",
          3366 => x"80",
          3367 => x"13",
          3368 => x"84",
          3369 => x"b9",
          3370 => x"33",
          3371 => x"07",
          3372 => x"74",
          3373 => x"3d",
          3374 => x"33",
          3375 => x"75",
          3376 => x"71",
          3377 => x"58",
          3378 => x"12",
          3379 => x"fc",
          3380 => x"12",
          3381 => x"07",
          3382 => x"12",
          3383 => x"07",
          3384 => x"77",
          3385 => x"84",
          3386 => x"12",
          3387 => x"ff",
          3388 => x"52",
          3389 => x"84",
          3390 => x"81",
          3391 => x"2b",
          3392 => x"33",
          3393 => x"8f",
          3394 => x"2a",
          3395 => x"54",
          3396 => x"14",
          3397 => x"70",
          3398 => x"71",
          3399 => x"81",
          3400 => x"ff",
          3401 => x"53",
          3402 => x"34",
          3403 => x"08",
          3404 => x"33",
          3405 => x"74",
          3406 => x"98",
          3407 => x"5d",
          3408 => x"25",
          3409 => x"33",
          3410 => x"07",
          3411 => x"75",
          3412 => x"fc",
          3413 => x"33",
          3414 => x"74",
          3415 => x"71",
          3416 => x"5c",
          3417 => x"82",
          3418 => x"3d",
          3419 => x"b9",
          3420 => x"8f",
          3421 => x"51",
          3422 => x"84",
          3423 => x"a0",
          3424 => x"80",
          3425 => x"51",
          3426 => x"08",
          3427 => x"16",
          3428 => x"84",
          3429 => x"84",
          3430 => x"34",
          3431 => x"fc",
          3432 => x"fe",
          3433 => x"06",
          3434 => x"74",
          3435 => x"84",
          3436 => x"84",
          3437 => x"55",
          3438 => x"15",
          3439 => x"7b",
          3440 => x"27",
          3441 => x"05",
          3442 => x"70",
          3443 => x"08",
          3444 => x"88",
          3445 => x"55",
          3446 => x"80",
          3447 => x"70",
          3448 => x"07",
          3449 => x"70",
          3450 => x"56",
          3451 => x"27",
          3452 => x"75",
          3453 => x"13",
          3454 => x"75",
          3455 => x"85",
          3456 => x"83",
          3457 => x"33",
          3458 => x"ff",
          3459 => x"70",
          3460 => x"51",
          3461 => x"51",
          3462 => x"75",
          3463 => x"83",
          3464 => x"07",
          3465 => x"5a",
          3466 => x"84",
          3467 => x"53",
          3468 => x"14",
          3469 => x"70",
          3470 => x"07",
          3471 => x"74",
          3472 => x"88",
          3473 => x"52",
          3474 => x"06",
          3475 => x"fc",
          3476 => x"81",
          3477 => x"19",
          3478 => x"8b",
          3479 => x"58",
          3480 => x"34",
          3481 => x"08",
          3482 => x"33",
          3483 => x"70",
          3484 => x"86",
          3485 => x"b9",
          3486 => x"85",
          3487 => x"2b",
          3488 => x"52",
          3489 => x"34",
          3490 => x"78",
          3491 => x"71",
          3492 => x"5c",
          3493 => x"85",
          3494 => x"84",
          3495 => x"8b",
          3496 => x"15",
          3497 => x"07",
          3498 => x"33",
          3499 => x"5a",
          3500 => x"12",
          3501 => x"fc",
          3502 => x"12",
          3503 => x"07",
          3504 => x"33",
          3505 => x"58",
          3506 => x"70",
          3507 => x"84",
          3508 => x"12",
          3509 => x"ff",
          3510 => x"57",
          3511 => x"84",
          3512 => x"fe",
          3513 => x"b9",
          3514 => x"a0",
          3515 => x"84",
          3516 => x"77",
          3517 => x"08",
          3518 => x"04",
          3519 => x"0c",
          3520 => x"82",
          3521 => x"f4",
          3522 => x"fc",
          3523 => x"81",
          3524 => x"76",
          3525 => x"34",
          3526 => x"17",
          3527 => x"b9",
          3528 => x"05",
          3529 => x"ff",
          3530 => x"56",
          3531 => x"34",
          3532 => x"10",
          3533 => x"55",
          3534 => x"83",
          3535 => x"fe",
          3536 => x"0d",
          3537 => x"b9",
          3538 => x"2e",
          3539 => x"af",
          3540 => x"81",
          3541 => x"fb",
          3542 => x"ff",
          3543 => x"ff",
          3544 => x"83",
          3545 => x"11",
          3546 => x"2b",
          3547 => x"ff",
          3548 => x"73",
          3549 => x"12",
          3550 => x"2b",
          3551 => x"44",
          3552 => x"52",
          3553 => x"fd",
          3554 => x"71",
          3555 => x"19",
          3556 => x"2b",
          3557 => x"56",
          3558 => x"38",
          3559 => x"1b",
          3560 => x"60",
          3561 => x"58",
          3562 => x"18",
          3563 => x"76",
          3564 => x"8b",
          3565 => x"70",
          3566 => x"71",
          3567 => x"53",
          3568 => x"ba",
          3569 => x"12",
          3570 => x"07",
          3571 => x"33",
          3572 => x"7e",
          3573 => x"71",
          3574 => x"57",
          3575 => x"59",
          3576 => x"1d",
          3577 => x"84",
          3578 => x"2b",
          3579 => x"14",
          3580 => x"07",
          3581 => x"40",
          3582 => x"7b",
          3583 => x"16",
          3584 => x"2b",
          3585 => x"2a",
          3586 => x"79",
          3587 => x"70",
          3588 => x"71",
          3589 => x"05",
          3590 => x"2b",
          3591 => x"5d",
          3592 => x"75",
          3593 => x"70",
          3594 => x"8b",
          3595 => x"82",
          3596 => x"2b",
          3597 => x"5d",
          3598 => x"34",
          3599 => x"08",
          3600 => x"33",
          3601 => x"56",
          3602 => x"7e",
          3603 => x"3f",
          3604 => x"61",
          3605 => x"06",
          3606 => x"b6",
          3607 => x"0c",
          3608 => x"0b",
          3609 => x"84",
          3610 => x"60",
          3611 => x"9f",
          3612 => x"7e",
          3613 => x"b9",
          3614 => x"81",
          3615 => x"08",
          3616 => x"87",
          3617 => x"b9",
          3618 => x"07",
          3619 => x"2a",
          3620 => x"34",
          3621 => x"22",
          3622 => x"08",
          3623 => x"15",
          3624 => x"b9",
          3625 => x"76",
          3626 => x"7f",
          3627 => x"f4",
          3628 => x"ba",
          3629 => x"1c",
          3630 => x"71",
          3631 => x"81",
          3632 => x"ff",
          3633 => x"5b",
          3634 => x"1c",
          3635 => x"7c",
          3636 => x"34",
          3637 => x"08",
          3638 => x"71",
          3639 => x"ff",
          3640 => x"ff",
          3641 => x"57",
          3642 => x"34",
          3643 => x"83",
          3644 => x"5b",
          3645 => x"61",
          3646 => x"51",
          3647 => x"39",
          3648 => x"06",
          3649 => x"ff",
          3650 => x"ff",
          3651 => x"71",
          3652 => x"1b",
          3653 => x"2b",
          3654 => x"54",
          3655 => x"f9",
          3656 => x"24",
          3657 => x"8f",
          3658 => x"61",
          3659 => x"39",
          3660 => x"0c",
          3661 => x"82",
          3662 => x"f4",
          3663 => x"fc",
          3664 => x"81",
          3665 => x"7e",
          3666 => x"34",
          3667 => x"19",
          3668 => x"b9",
          3669 => x"05",
          3670 => x"ff",
          3671 => x"44",
          3672 => x"89",
          3673 => x"10",
          3674 => x"f8",
          3675 => x"34",
          3676 => x"39",
          3677 => x"83",
          3678 => x"fb",
          3679 => x"2e",
          3680 => x"3f",
          3681 => x"95",
          3682 => x"33",
          3683 => x"83",
          3684 => x"87",
          3685 => x"2b",
          3686 => x"15",
          3687 => x"2a",
          3688 => x"53",
          3689 => x"34",
          3690 => x"fc",
          3691 => x"12",
          3692 => x"07",
          3693 => x"33",
          3694 => x"5b",
          3695 => x"73",
          3696 => x"05",
          3697 => x"33",
          3698 => x"81",
          3699 => x"5c",
          3700 => x"1e",
          3701 => x"82",
          3702 => x"2b",
          3703 => x"33",
          3704 => x"70",
          3705 => x"57",
          3706 => x"1d",
          3707 => x"70",
          3708 => x"71",
          3709 => x"33",
          3710 => x"70",
          3711 => x"5c",
          3712 => x"83",
          3713 => x"1f",
          3714 => x"88",
          3715 => x"83",
          3716 => x"84",
          3717 => x"b9",
          3718 => x"ff",
          3719 => x"84",
          3720 => x"a0",
          3721 => x"80",
          3722 => x"51",
          3723 => x"08",
          3724 => x"17",
          3725 => x"84",
          3726 => x"84",
          3727 => x"34",
          3728 => x"fc",
          3729 => x"fe",
          3730 => x"06",
          3731 => x"61",
          3732 => x"84",
          3733 => x"84",
          3734 => x"5d",
          3735 => x"1c",
          3736 => x"54",
          3737 => x"1a",
          3738 => x"07",
          3739 => x"33",
          3740 => x"5c",
          3741 => x"84",
          3742 => x"84",
          3743 => x"33",
          3744 => x"83",
          3745 => x"87",
          3746 => x"88",
          3747 => x"59",
          3748 => x"64",
          3749 => x"1d",
          3750 => x"2b",
          3751 => x"2a",
          3752 => x"7f",
          3753 => x"70",
          3754 => x"8b",
          3755 => x"70",
          3756 => x"07",
          3757 => x"77",
          3758 => x"5a",
          3759 => x"17",
          3760 => x"fc",
          3761 => x"33",
          3762 => x"74",
          3763 => x"88",
          3764 => x"88",
          3765 => x"41",
          3766 => x"05",
          3767 => x"fa",
          3768 => x"33",
          3769 => x"79",
          3770 => x"71",
          3771 => x"5e",
          3772 => x"34",
          3773 => x"08",
          3774 => x"33",
          3775 => x"74",
          3776 => x"71",
          3777 => x"56",
          3778 => x"60",
          3779 => x"34",
          3780 => x"81",
          3781 => x"ff",
          3782 => x"58",
          3783 => x"34",
          3784 => x"33",
          3785 => x"83",
          3786 => x"12",
          3787 => x"2b",
          3788 => x"88",
          3789 => x"42",
          3790 => x"83",
          3791 => x"1f",
          3792 => x"2b",
          3793 => x"33",
          3794 => x"81",
          3795 => x"54",
          3796 => x"7c",
          3797 => x"fc",
          3798 => x"12",
          3799 => x"07",
          3800 => x"33",
          3801 => x"78",
          3802 => x"71",
          3803 => x"57",
          3804 => x"5a",
          3805 => x"85",
          3806 => x"17",
          3807 => x"8b",
          3808 => x"86",
          3809 => x"2b",
          3810 => x"52",
          3811 => x"34",
          3812 => x"08",
          3813 => x"88",
          3814 => x"88",
          3815 => x"34",
          3816 => x"08",
          3817 => x"33",
          3818 => x"74",
          3819 => x"88",
          3820 => x"45",
          3821 => x"34",
          3822 => x"08",
          3823 => x"71",
          3824 => x"05",
          3825 => x"88",
          3826 => x"45",
          3827 => x"1a",
          3828 => x"fc",
          3829 => x"12",
          3830 => x"62",
          3831 => x"5d",
          3832 => x"fa",
          3833 => x"05",
          3834 => x"ff",
          3835 => x"86",
          3836 => x"2b",
          3837 => x"1c",
          3838 => x"07",
          3839 => x"41",
          3840 => x"61",
          3841 => x"70",
          3842 => x"71",
          3843 => x"05",
          3844 => x"88",
          3845 => x"5f",
          3846 => x"86",
          3847 => x"84",
          3848 => x"12",
          3849 => x"ff",
          3850 => x"55",
          3851 => x"84",
          3852 => x"81",
          3853 => x"2b",
          3854 => x"33",
          3855 => x"8f",
          3856 => x"2a",
          3857 => x"58",
          3858 => x"1e",
          3859 => x"70",
          3860 => x"71",
          3861 => x"81",
          3862 => x"ff",
          3863 => x"49",
          3864 => x"34",
          3865 => x"ff",
          3866 => x"52",
          3867 => x"08",
          3868 => x"93",
          3869 => x"8c",
          3870 => x"51",
          3871 => x"27",
          3872 => x"3d",
          3873 => x"08",
          3874 => x"77",
          3875 => x"8c",
          3876 => x"e4",
          3877 => x"84",
          3878 => x"77",
          3879 => x"51",
          3880 => x"8c",
          3881 => x"f4",
          3882 => x"0b",
          3883 => x"53",
          3884 => x"b6",
          3885 => x"76",
          3886 => x"84",
          3887 => x"34",
          3888 => x"fc",
          3889 => x"0b",
          3890 => x"84",
          3891 => x"80",
          3892 => x"88",
          3893 => x"17",
          3894 => x"f8",
          3895 => x"fc",
          3896 => x"82",
          3897 => x"77",
          3898 => x"fe",
          3899 => x"05",
          3900 => x"87",
          3901 => x"71",
          3902 => x"04",
          3903 => x"52",
          3904 => x"71",
          3905 => x"08",
          3906 => x"72",
          3907 => x"88",
          3908 => x"0c",
          3909 => x"7c",
          3910 => x"33",
          3911 => x"74",
          3912 => x"33",
          3913 => x"73",
          3914 => x"c0",
          3915 => x"76",
          3916 => x"08",
          3917 => x"a7",
          3918 => x"73",
          3919 => x"74",
          3920 => x"2e",
          3921 => x"84",
          3922 => x"84",
          3923 => x"06",
          3924 => x"ac",
          3925 => x"7e",
          3926 => x"5a",
          3927 => x"26",
          3928 => x"54",
          3929 => x"bd",
          3930 => x"98",
          3931 => x"51",
          3932 => x"81",
          3933 => x"38",
          3934 => x"e2",
          3935 => x"fc",
          3936 => x"83",
          3937 => x"ba",
          3938 => x"80",
          3939 => x"5a",
          3940 => x"38",
          3941 => x"84",
          3942 => x"9f",
          3943 => x"71",
          3944 => x"12",
          3945 => x"53",
          3946 => x"98",
          3947 => x"96",
          3948 => x"83",
          3949 => x"ba",
          3950 => x"80",
          3951 => x"0c",
          3952 => x"0c",
          3953 => x"3d",
          3954 => x"92",
          3955 => x"71",
          3956 => x"51",
          3957 => x"98",
          3958 => x"c0",
          3959 => x"81",
          3960 => x"52",
          3961 => x"2e",
          3962 => x"54",
          3963 => x"3d",
          3964 => x"33",
          3965 => x"09",
          3966 => x"75",
          3967 => x"80",
          3968 => x"3f",
          3969 => x"38",
          3970 => x"8c",
          3971 => x"08",
          3972 => x"33",
          3973 => x"84",
          3974 => x"06",
          3975 => x"19",
          3976 => x"08",
          3977 => x"08",
          3978 => x"ff",
          3979 => x"82",
          3980 => x"81",
          3981 => x"18",
          3982 => x"33",
          3983 => x"06",
          3984 => x"76",
          3985 => x"38",
          3986 => x"57",
          3987 => x"ff",
          3988 => x"0b",
          3989 => x"84",
          3990 => x"80",
          3991 => x"0b",
          3992 => x"19",
          3993 => x"34",
          3994 => x"80",
          3995 => x"e1",
          3996 => x"08",
          3997 => x"88",
          3998 => x"74",
          3999 => x"34",
          4000 => x"19",
          4001 => x"a4",
          4002 => x"84",
          4003 => x"75",
          4004 => x"55",
          4005 => x"08",
          4006 => x"81",
          4007 => x"33",
          4008 => x"34",
          4009 => x"51",
          4010 => x"80",
          4011 => x"f3",
          4012 => x"56",
          4013 => x"17",
          4014 => x"77",
          4015 => x"04",
          4016 => x"2e",
          4017 => x"a5",
          4018 => x"dd",
          4019 => x"2a",
          4020 => x"5b",
          4021 => x"83",
          4022 => x"81",
          4023 => x"53",
          4024 => x"f8",
          4025 => x"2e",
          4026 => x"b4",
          4027 => x"83",
          4028 => x"1c",
          4029 => x"53",
          4030 => x"2e",
          4031 => x"71",
          4032 => x"81",
          4033 => x"53",
          4034 => x"f8",
          4035 => x"2e",
          4036 => x"b4",
          4037 => x"83",
          4038 => x"88",
          4039 => x"84",
          4040 => x"fe",
          4041 => x"ba",
          4042 => x"88",
          4043 => x"17",
          4044 => x"83",
          4045 => x"7b",
          4046 => x"81",
          4047 => x"17",
          4048 => x"8c",
          4049 => x"81",
          4050 => x"df",
          4051 => x"05",
          4052 => x"71",
          4053 => x"57",
          4054 => x"2e",
          4055 => x"87",
          4056 => x"17",
          4057 => x"83",
          4058 => x"7b",
          4059 => x"81",
          4060 => x"17",
          4061 => x"8c",
          4062 => x"81",
          4063 => x"f7",
          4064 => x"77",
          4065 => x"12",
          4066 => x"07",
          4067 => x"2b",
          4068 => x"80",
          4069 => x"5c",
          4070 => x"04",
          4071 => x"17",
          4072 => x"f6",
          4073 => x"08",
          4074 => x"38",
          4075 => x"b4",
          4076 => x"ba",
          4077 => x"08",
          4078 => x"55",
          4079 => x"f7",
          4080 => x"18",
          4081 => x"33",
          4082 => x"df",
          4083 => x"b8",
          4084 => x"5c",
          4085 => x"7b",
          4086 => x"84",
          4087 => x"17",
          4088 => x"a0",
          4089 => x"33",
          4090 => x"84",
          4091 => x"81",
          4092 => x"70",
          4093 => x"bb",
          4094 => x"7b",
          4095 => x"84",
          4096 => x"17",
          4097 => x"8c",
          4098 => x"27",
          4099 => x"74",
          4100 => x"38",
          4101 => x"08",
          4102 => x"51",
          4103 => x"39",
          4104 => x"17",
          4105 => x"f4",
          4106 => x"08",
          4107 => x"38",
          4108 => x"b4",
          4109 => x"ba",
          4110 => x"08",
          4111 => x"55",
          4112 => x"84",
          4113 => x"18",
          4114 => x"33",
          4115 => x"ec",
          4116 => x"18",
          4117 => x"33",
          4118 => x"81",
          4119 => x"39",
          4120 => x"57",
          4121 => x"38",
          4122 => x"78",
          4123 => x"74",
          4124 => x"2e",
          4125 => x"0c",
          4126 => x"a8",
          4127 => x"1a",
          4128 => x"b6",
          4129 => x"7c",
          4130 => x"38",
          4131 => x"81",
          4132 => x"ba",
          4133 => x"58",
          4134 => x"58",
          4135 => x"fe",
          4136 => x"06",
          4137 => x"88",
          4138 => x"0b",
          4139 => x"0c",
          4140 => x"09",
          4141 => x"2a",
          4142 => x"b4",
          4143 => x"85",
          4144 => x"5d",
          4145 => x"bd",
          4146 => x"52",
          4147 => x"84",
          4148 => x"ff",
          4149 => x"79",
          4150 => x"2b",
          4151 => x"83",
          4152 => x"06",
          4153 => x"5e",
          4154 => x"56",
          4155 => x"5a",
          4156 => x"5b",
          4157 => x"1a",
          4158 => x"16",
          4159 => x"b4",
          4160 => x"2e",
          4161 => x"71",
          4162 => x"81",
          4163 => x"53",
          4164 => x"f0",
          4165 => x"2e",
          4166 => x"b4",
          4167 => x"38",
          4168 => x"81",
          4169 => x"7a",
          4170 => x"84",
          4171 => x"06",
          4172 => x"81",
          4173 => x"a8",
          4174 => x"1a",
          4175 => x"dd",
          4176 => x"70",
          4177 => x"9b",
          4178 => x"7f",
          4179 => x"84",
          4180 => x"19",
          4181 => x"1b",
          4182 => x"56",
          4183 => x"19",
          4184 => x"38",
          4185 => x"19",
          4186 => x"8c",
          4187 => x"81",
          4188 => x"83",
          4189 => x"05",
          4190 => x"38",
          4191 => x"06",
          4192 => x"76",
          4193 => x"cb",
          4194 => x"70",
          4195 => x"8b",
          4196 => x"7c",
          4197 => x"84",
          4198 => x"19",
          4199 => x"1b",
          4200 => x"40",
          4201 => x"82",
          4202 => x"81",
          4203 => x"1e",
          4204 => x"ee",
          4205 => x"81",
          4206 => x"81",
          4207 => x"81",
          4208 => x"09",
          4209 => x"8c",
          4210 => x"70",
          4211 => x"84",
          4212 => x"74",
          4213 => x"33",
          4214 => x"fc",
          4215 => x"76",
          4216 => x"3f",
          4217 => x"76",
          4218 => x"33",
          4219 => x"84",
          4220 => x"06",
          4221 => x"83",
          4222 => x"1b",
          4223 => x"8c",
          4224 => x"27",
          4225 => x"74",
          4226 => x"38",
          4227 => x"81",
          4228 => x"5a",
          4229 => x"53",
          4230 => x"f3",
          4231 => x"76",
          4232 => x"83",
          4233 => x"b8",
          4234 => x"b9",
          4235 => x"fd",
          4236 => x"fc",
          4237 => x"33",
          4238 => x"f0",
          4239 => x"58",
          4240 => x"75",
          4241 => x"79",
          4242 => x"7a",
          4243 => x"3d",
          4244 => x"5a",
          4245 => x"57",
          4246 => x"9c",
          4247 => x"19",
          4248 => x"80",
          4249 => x"38",
          4250 => x"08",
          4251 => x"77",
          4252 => x"51",
          4253 => x"80",
          4254 => x"ba",
          4255 => x"ba",
          4256 => x"07",
          4257 => x"55",
          4258 => x"2e",
          4259 => x"55",
          4260 => x"0d",
          4261 => x"ba",
          4262 => x"79",
          4263 => x"84",
          4264 => x"ba",
          4265 => x"ff",
          4266 => x"ba",
          4267 => x"fe",
          4268 => x"08",
          4269 => x"52",
          4270 => x"84",
          4271 => x"38",
          4272 => x"70",
          4273 => x"84",
          4274 => x"55",
          4275 => x"08",
          4276 => x"54",
          4277 => x"9c",
          4278 => x"70",
          4279 => x"2e",
          4280 => x"78",
          4281 => x"08",
          4282 => x"ba",
          4283 => x"55",
          4284 => x"38",
          4285 => x"fe",
          4286 => x"78",
          4287 => x"0c",
          4288 => x"84",
          4289 => x"8c",
          4290 => x"84",
          4291 => x"84",
          4292 => x"73",
          4293 => x"7a",
          4294 => x"ba",
          4295 => x"ba",
          4296 => x"3d",
          4297 => x"ff",
          4298 => x"f8",
          4299 => x"55",
          4300 => x"df",
          4301 => x"d7",
          4302 => x"08",
          4303 => x"56",
          4304 => x"85",
          4305 => x"5a",
          4306 => x"17",
          4307 => x"0c",
          4308 => x"80",
          4309 => x"98",
          4310 => x"b8",
          4311 => x"84",
          4312 => x"82",
          4313 => x"0d",
          4314 => x"2e",
          4315 => x"89",
          4316 => x"38",
          4317 => x"14",
          4318 => x"8d",
          4319 => x"b0",
          4320 => x"19",
          4321 => x"51",
          4322 => x"55",
          4323 => x"38",
          4324 => x"ff",
          4325 => x"ba",
          4326 => x"73",
          4327 => x"38",
          4328 => x"8c",
          4329 => x"0d",
          4330 => x"05",
          4331 => x"27",
          4332 => x"98",
          4333 => x"2e",
          4334 => x"7a",
          4335 => x"57",
          4336 => x"88",
          4337 => x"81",
          4338 => x"90",
          4339 => x"18",
          4340 => x"0c",
          4341 => x"0c",
          4342 => x"2a",
          4343 => x"76",
          4344 => x"08",
          4345 => x"8c",
          4346 => x"ba",
          4347 => x"19",
          4348 => x"91",
          4349 => x"94",
          4350 => x"3f",
          4351 => x"84",
          4352 => x"38",
          4353 => x"2e",
          4354 => x"8c",
          4355 => x"ba",
          4356 => x"7d",
          4357 => x"08",
          4358 => x"78",
          4359 => x"71",
          4360 => x"7b",
          4361 => x"80",
          4362 => x"05",
          4363 => x"38",
          4364 => x"75",
          4365 => x"1c",
          4366 => x"e4",
          4367 => x"e7",
          4368 => x"98",
          4369 => x"0c",
          4370 => x"19",
          4371 => x"1a",
          4372 => x"ba",
          4373 => x"8c",
          4374 => x"a8",
          4375 => x"08",
          4376 => x"5c",
          4377 => x"db",
          4378 => x"1a",
          4379 => x"33",
          4380 => x"8a",
          4381 => x"06",
          4382 => x"a7",
          4383 => x"9c",
          4384 => x"58",
          4385 => x"19",
          4386 => x"05",
          4387 => x"81",
          4388 => x"0d",
          4389 => x"5c",
          4390 => x"70",
          4391 => x"80",
          4392 => x"75",
          4393 => x"2e",
          4394 => x"58",
          4395 => x"81",
          4396 => x"19",
          4397 => x"3f",
          4398 => x"38",
          4399 => x"0c",
          4400 => x"1c",
          4401 => x"2e",
          4402 => x"06",
          4403 => x"86",
          4404 => x"30",
          4405 => x"25",
          4406 => x"57",
          4407 => x"06",
          4408 => x"38",
          4409 => x"ff",
          4410 => x"3f",
          4411 => x"8c",
          4412 => x"56",
          4413 => x"8c",
          4414 => x"b4",
          4415 => x"33",
          4416 => x"ba",
          4417 => x"fe",
          4418 => x"1a",
          4419 => x"31",
          4420 => x"a0",
          4421 => x"19",
          4422 => x"06",
          4423 => x"08",
          4424 => x"81",
          4425 => x"57",
          4426 => x"81",
          4427 => x"81",
          4428 => x"8d",
          4429 => x"90",
          4430 => x"5e",
          4431 => x"ff",
          4432 => x"56",
          4433 => x"be",
          4434 => x"98",
          4435 => x"94",
          4436 => x"39",
          4437 => x"09",
          4438 => x"9b",
          4439 => x"2b",
          4440 => x"38",
          4441 => x"29",
          4442 => x"5b",
          4443 => x"81",
          4444 => x"07",
          4445 => x"c5",
          4446 => x"38",
          4447 => x"75",
          4448 => x"57",
          4449 => x"70",
          4450 => x"80",
          4451 => x"fe",
          4452 => x"80",
          4453 => x"06",
          4454 => x"ff",
          4455 => x"fe",
          4456 => x"8b",
          4457 => x"29",
          4458 => x"40",
          4459 => x"19",
          4460 => x"7e",
          4461 => x"1d",
          4462 => x"3d",
          4463 => x"08",
          4464 => x"cf",
          4465 => x"ba",
          4466 => x"70",
          4467 => x"b8",
          4468 => x"58",
          4469 => x"38",
          4470 => x"78",
          4471 => x"81",
          4472 => x"1b",
          4473 => x"8c",
          4474 => x"81",
          4475 => x"76",
          4476 => x"33",
          4477 => x"38",
          4478 => x"ff",
          4479 => x"76",
          4480 => x"83",
          4481 => x"81",
          4482 => x"8f",
          4483 => x"78",
          4484 => x"2a",
          4485 => x"81",
          4486 => x"81",
          4487 => x"76",
          4488 => x"38",
          4489 => x"a7",
          4490 => x"78",
          4491 => x"81",
          4492 => x"1a",
          4493 => x"81",
          4494 => x"81",
          4495 => x"80",
          4496 => x"ba",
          4497 => x"80",
          4498 => x"8c",
          4499 => x"b4",
          4500 => x"33",
          4501 => x"ba",
          4502 => x"fe",
          4503 => x"1c",
          4504 => x"31",
          4505 => x"a0",
          4506 => x"1b",
          4507 => x"06",
          4508 => x"08",
          4509 => x"81",
          4510 => x"57",
          4511 => x"39",
          4512 => x"06",
          4513 => x"86",
          4514 => x"93",
          4515 => x"06",
          4516 => x"0c",
          4517 => x"38",
          4518 => x"7b",
          4519 => x"08",
          4520 => x"fc",
          4521 => x"2e",
          4522 => x"0b",
          4523 => x"19",
          4524 => x"06",
          4525 => x"33",
          4526 => x"59",
          4527 => x"33",
          4528 => x"5b",
          4529 => x"8c",
          4530 => x"71",
          4531 => x"57",
          4532 => x"81",
          4533 => x"81",
          4534 => x"7a",
          4535 => x"81",
          4536 => x"75",
          4537 => x"06",
          4538 => x"58",
          4539 => x"33",
          4540 => x"75",
          4541 => x"8d",
          4542 => x"41",
          4543 => x"70",
          4544 => x"39",
          4545 => x"3d",
          4546 => x"ff",
          4547 => x"39",
          4548 => x"ab",
          4549 => x"5d",
          4550 => x"74",
          4551 => x"5d",
          4552 => x"70",
          4553 => x"74",
          4554 => x"40",
          4555 => x"70",
          4556 => x"05",
          4557 => x"38",
          4558 => x"06",
          4559 => x"38",
          4560 => x"0b",
          4561 => x"7b",
          4562 => x"55",
          4563 => x"70",
          4564 => x"74",
          4565 => x"38",
          4566 => x"2e",
          4567 => x"8f",
          4568 => x"76",
          4569 => x"72",
          4570 => x"57",
          4571 => x"a0",
          4572 => x"80",
          4573 => x"ca",
          4574 => x"05",
          4575 => x"55",
          4576 => x"55",
          4577 => x"78",
          4578 => x"38",
          4579 => x"76",
          4580 => x"38",
          4581 => x"38",
          4582 => x"a2",
          4583 => x"74",
          4584 => x"81",
          4585 => x"8e",
          4586 => x"81",
          4587 => x"77",
          4588 => x"7d",
          4589 => x"08",
          4590 => x"7b",
          4591 => x"80",
          4592 => x"8c",
          4593 => x"2e",
          4594 => x"80",
          4595 => x"08",
          4596 => x"57",
          4597 => x"81",
          4598 => x"52",
          4599 => x"84",
          4600 => x"7d",
          4601 => x"08",
          4602 => x"38",
          4603 => x"59",
          4604 => x"18",
          4605 => x"18",
          4606 => x"06",
          4607 => x"b8",
          4608 => x"a4",
          4609 => x"85",
          4610 => x"19",
          4611 => x"1e",
          4612 => x"e5",
          4613 => x"80",
          4614 => x"2e",
          4615 => x"7b",
          4616 => x"51",
          4617 => x"56",
          4618 => x"88",
          4619 => x"89",
          4620 => x"ff",
          4621 => x"1e",
          4622 => x"af",
          4623 => x"7f",
          4624 => x"b8",
          4625 => x"9c",
          4626 => x"85",
          4627 => x"1d",
          4628 => x"a0",
          4629 => x"76",
          4630 => x"55",
          4631 => x"08",
          4632 => x"05",
          4633 => x"34",
          4634 => x"1e",
          4635 => x"5a",
          4636 => x"1d",
          4637 => x"0c",
          4638 => x"70",
          4639 => x"74",
          4640 => x"7d",
          4641 => x"08",
          4642 => x"fd",
          4643 => x"b4",
          4644 => x"33",
          4645 => x"08",
          4646 => x"38",
          4647 => x"b4",
          4648 => x"74",
          4649 => x"18",
          4650 => x"38",
          4651 => x"39",
          4652 => x"31",
          4653 => x"84",
          4654 => x"08",
          4655 => x"08",
          4656 => x"75",
          4657 => x"05",
          4658 => x"ff",
          4659 => x"e4",
          4660 => x"43",
          4661 => x"b4",
          4662 => x"1c",
          4663 => x"06",
          4664 => x"b8",
          4665 => x"dc",
          4666 => x"85",
          4667 => x"1d",
          4668 => x"8c",
          4669 => x"ff",
          4670 => x"34",
          4671 => x"1c",
          4672 => x"1c",
          4673 => x"77",
          4674 => x"2e",
          4675 => x"81",
          4676 => x"18",
          4677 => x"81",
          4678 => x"75",
          4679 => x"ff",
          4680 => x"cb",
          4681 => x"b3",
          4682 => x"58",
          4683 => x"7b",
          4684 => x"52",
          4685 => x"8c",
          4686 => x"f1",
          4687 => x"a9",
          4688 => x"1c",
          4689 => x"1d",
          4690 => x"56",
          4691 => x"84",
          4692 => x"1c",
          4693 => x"8c",
          4694 => x"27",
          4695 => x"61",
          4696 => x"38",
          4697 => x"08",
          4698 => x"51",
          4699 => x"39",
          4700 => x"43",
          4701 => x"06",
          4702 => x"70",
          4703 => x"38",
          4704 => x"5d",
          4705 => x"08",
          4706 => x"cf",
          4707 => x"2e",
          4708 => x"8c",
          4709 => x"a8",
          4710 => x"08",
          4711 => x"7e",
          4712 => x"08",
          4713 => x"41",
          4714 => x"fc",
          4715 => x"39",
          4716 => x"fc",
          4717 => x"b4",
          4718 => x"61",
          4719 => x"3f",
          4720 => x"08",
          4721 => x"81",
          4722 => x"e3",
          4723 => x"08",
          4724 => x"34",
          4725 => x"38",
          4726 => x"38",
          4727 => x"70",
          4728 => x"78",
          4729 => x"70",
          4730 => x"82",
          4731 => x"83",
          4732 => x"ff",
          4733 => x"76",
          4734 => x"79",
          4735 => x"70",
          4736 => x"18",
          4737 => x"34",
          4738 => x"9c",
          4739 => x"58",
          4740 => x"74",
          4741 => x"32",
          4742 => x"55",
          4743 => x"72",
          4744 => x"81",
          4745 => x"77",
          4746 => x"58",
          4747 => x"18",
          4748 => x"34",
          4749 => x"77",
          4750 => x"34",
          4751 => x"80",
          4752 => x"8c",
          4753 => x"73",
          4754 => x"8b",
          4755 => x"08",
          4756 => x"33",
          4757 => x"81",
          4758 => x"75",
          4759 => x"16",
          4760 => x"07",
          4761 => x"55",
          4762 => x"98",
          4763 => x"54",
          4764 => x"04",
          4765 => x"1d",
          4766 => x"5b",
          4767 => x"74",
          4768 => x"ba",
          4769 => x"81",
          4770 => x"27",
          4771 => x"73",
          4772 => x"78",
          4773 => x"56",
          4774 => x"5c",
          4775 => x"ba",
          4776 => x"07",
          4777 => x"55",
          4778 => x"34",
          4779 => x"1f",
          4780 => x"89",
          4781 => x"2e",
          4782 => x"57",
          4783 => x"11",
          4784 => x"9c",
          4785 => x"88",
          4786 => x"53",
          4787 => x"8a",
          4788 => x"06",
          4789 => x"5a",
          4790 => x"71",
          4791 => x"56",
          4792 => x"72",
          4793 => x"30",
          4794 => x"53",
          4795 => x"3d",
          4796 => x"5c",
          4797 => x"74",
          4798 => x"80",
          4799 => x"2e",
          4800 => x"1d",
          4801 => x"41",
          4802 => x"38",
          4803 => x"57",
          4804 => x"55",
          4805 => x"0c",
          4806 => x"ff",
          4807 => x"18",
          4808 => x"73",
          4809 => x"70",
          4810 => x"07",
          4811 => x"38",
          4812 => x"74",
          4813 => x"a8",
          4814 => x"ff",
          4815 => x"81",
          4816 => x"81",
          4817 => x"56",
          4818 => x"ff",
          4819 => x"81",
          4820 => x"18",
          4821 => x"70",
          4822 => x"57",
          4823 => x"cb",
          4824 => x"30",
          4825 => x"58",
          4826 => x"14",
          4827 => x"55",
          4828 => x"dc",
          4829 => x"07",
          4830 => x"88",
          4831 => x"3d",
          4832 => x"90",
          4833 => x"51",
          4834 => x"08",
          4835 => x"8d",
          4836 => x"0c",
          4837 => x"33",
          4838 => x"80",
          4839 => x"80",
          4840 => x"51",
          4841 => x"84",
          4842 => x"81",
          4843 => x"80",
          4844 => x"7d",
          4845 => x"80",
          4846 => x"af",
          4847 => x"70",
          4848 => x"54",
          4849 => x"9f",
          4850 => x"2e",
          4851 => x"d1",
          4852 => x"a7",
          4853 => x"70",
          4854 => x"9f",
          4855 => x"7c",
          4856 => x"ff",
          4857 => x"77",
          4858 => x"2e",
          4859 => x"83",
          4860 => x"56",
          4861 => x"83",
          4862 => x"82",
          4863 => x"77",
          4864 => x"78",
          4865 => x"fe",
          4866 => x"2e",
          4867 => x"54",
          4868 => x"38",
          4869 => x"74",
          4870 => x"53",
          4871 => x"88",
          4872 => x"57",
          4873 => x"38",
          4874 => x"ae",
          4875 => x"5a",
          4876 => x"72",
          4877 => x"26",
          4878 => x"70",
          4879 => x"7c",
          4880 => x"2e",
          4881 => x"83",
          4882 => x"83",
          4883 => x"76",
          4884 => x"81",
          4885 => x"77",
          4886 => x"53",
          4887 => x"57",
          4888 => x"7c",
          4889 => x"06",
          4890 => x"7d",
          4891 => x"e3",
          4892 => x"75",
          4893 => x"80",
          4894 => x"7d",
          4895 => x"2e",
          4896 => x"ab",
          4897 => x"84",
          4898 => x"54",
          4899 => x"ac",
          4900 => x"09",
          4901 => x"2a",
          4902 => x"f0",
          4903 => x"78",
          4904 => x"56",
          4905 => x"57",
          4906 => x"79",
          4907 => x"7c",
          4908 => x"fd",
          4909 => x"8a",
          4910 => x"2e",
          4911 => x"22",
          4912 => x"fc",
          4913 => x"7b",
          4914 => x"ae",
          4915 => x"54",
          4916 => x"81",
          4917 => x"79",
          4918 => x"7b",
          4919 => x"08",
          4920 => x"8c",
          4921 => x"81",
          4922 => x"1c",
          4923 => x"5d",
          4924 => x"1c",
          4925 => x"d3",
          4926 => x"88",
          4927 => x"54",
          4928 => x"88",
          4929 => x"fe",
          4930 => x"2e",
          4931 => x"fb",
          4932 => x"07",
          4933 => x"7d",
          4934 => x"06",
          4935 => x"06",
          4936 => x"fd",
          4937 => x"7c",
          4938 => x"38",
          4939 => x"34",
          4940 => x"3d",
          4941 => x"38",
          4942 => x"ff",
          4943 => x"38",
          4944 => x"5c",
          4945 => x"5a",
          4946 => x"f6",
          4947 => x"ff",
          4948 => x"55",
          4949 => x"ff",
          4950 => x"54",
          4951 => x"74",
          4952 => x"b4",
          4953 => x"ff",
          4954 => x"80",
          4955 => x"81",
          4956 => x"56",
          4957 => x"ff",
          4958 => x"bf",
          4959 => x"7d",
          4960 => x"53",
          4961 => x"93",
          4962 => x"06",
          4963 => x"58",
          4964 => x"59",
          4965 => x"16",
          4966 => x"b3",
          4967 => x"ff",
          4968 => x"ae",
          4969 => x"1d",
          4970 => x"34",
          4971 => x"14",
          4972 => x"2b",
          4973 => x"1f",
          4974 => x"1b",
          4975 => x"72",
          4976 => x"05",
          4977 => x"5b",
          4978 => x"1d",
          4979 => x"09",
          4980 => x"39",
          4981 => x"f6",
          4982 => x"0c",
          4983 => x"67",
          4984 => x"33",
          4985 => x"7e",
          4986 => x"2e",
          4987 => x"5b",
          4988 => x"ba",
          4989 => x"75",
          4990 => x"e8",
          4991 => x"38",
          4992 => x"70",
          4993 => x"2e",
          4994 => x"81",
          4995 => x"80",
          4996 => x"ff",
          4997 => x"81",
          4998 => x"7c",
          4999 => x"34",
          5000 => x"33",
          5001 => x"33",
          5002 => x"8c",
          5003 => x"41",
          5004 => x"78",
          5005 => x"81",
          5006 => x"38",
          5007 => x"0b",
          5008 => x"81",
          5009 => x"81",
          5010 => x"3f",
          5011 => x"38",
          5012 => x"0c",
          5013 => x"17",
          5014 => x"2b",
          5015 => x"d4",
          5016 => x"26",
          5017 => x"42",
          5018 => x"84",
          5019 => x"81",
          5020 => x"33",
          5021 => x"07",
          5022 => x"81",
          5023 => x"33",
          5024 => x"07",
          5025 => x"17",
          5026 => x"90",
          5027 => x"33",
          5028 => x"71",
          5029 => x"56",
          5030 => x"33",
          5031 => x"ff",
          5032 => x"59",
          5033 => x"38",
          5034 => x"80",
          5035 => x"8a",
          5036 => x"87",
          5037 => x"61",
          5038 => x"80",
          5039 => x"56",
          5040 => x"8f",
          5041 => x"98",
          5042 => x"18",
          5043 => x"74",
          5044 => x"33",
          5045 => x"88",
          5046 => x"07",
          5047 => x"44",
          5048 => x"17",
          5049 => x"2b",
          5050 => x"2e",
          5051 => x"2a",
          5052 => x"38",
          5053 => x"ed",
          5054 => x"84",
          5055 => x"38",
          5056 => x"ff",
          5057 => x"83",
          5058 => x"75",
          5059 => x"5d",
          5060 => x"a4",
          5061 => x"0c",
          5062 => x"7c",
          5063 => x"22",
          5064 => x"e0",
          5065 => x"19",
          5066 => x"10",
          5067 => x"05",
          5068 => x"59",
          5069 => x"b8",
          5070 => x"0b",
          5071 => x"18",
          5072 => x"7c",
          5073 => x"05",
          5074 => x"86",
          5075 => x"18",
          5076 => x"58",
          5077 => x"0d",
          5078 => x"97",
          5079 => x"70",
          5080 => x"89",
          5081 => x"ff",
          5082 => x"2e",
          5083 => x"e5",
          5084 => x"5a",
          5085 => x"79",
          5086 => x"12",
          5087 => x"38",
          5088 => x"55",
          5089 => x"89",
          5090 => x"58",
          5091 => x"55",
          5092 => x"38",
          5093 => x"70",
          5094 => x"07",
          5095 => x"98",
          5096 => x"83",
          5097 => x"f9",
          5098 => x"38",
          5099 => x"58",
          5100 => x"c0",
          5101 => x"81",
          5102 => x"81",
          5103 => x"70",
          5104 => x"77",
          5105 => x"83",
          5106 => x"83",
          5107 => x"5b",
          5108 => x"16",
          5109 => x"2b",
          5110 => x"33",
          5111 => x"1b",
          5112 => x"40",
          5113 => x"0c",
          5114 => x"80",
          5115 => x"1d",
          5116 => x"71",
          5117 => x"f0",
          5118 => x"43",
          5119 => x"7a",
          5120 => x"83",
          5121 => x"7a",
          5122 => x"38",
          5123 => x"81",
          5124 => x"84",
          5125 => x"ff",
          5126 => x"84",
          5127 => x"7f",
          5128 => x"83",
          5129 => x"81",
          5130 => x"33",
          5131 => x"b7",
          5132 => x"70",
          5133 => x"7f",
          5134 => x"38",
          5135 => x"80",
          5136 => x"58",
          5137 => x"38",
          5138 => x"38",
          5139 => x"1a",
          5140 => x"fe",
          5141 => x"80",
          5142 => x"58",
          5143 => x"70",
          5144 => x"ff",
          5145 => x"2e",
          5146 => x"38",
          5147 => x"c0",
          5148 => x"5d",
          5149 => x"71",
          5150 => x"40",
          5151 => x"80",
          5152 => x"39",
          5153 => x"84",
          5154 => x"75",
          5155 => x"85",
          5156 => x"40",
          5157 => x"84",
          5158 => x"83",
          5159 => x"5c",
          5160 => x"33",
          5161 => x"71",
          5162 => x"77",
          5163 => x"2e",
          5164 => x"83",
          5165 => x"81",
          5166 => x"5c",
          5167 => x"58",
          5168 => x"38",
          5169 => x"77",
          5170 => x"81",
          5171 => x"33",
          5172 => x"07",
          5173 => x"06",
          5174 => x"5a",
          5175 => x"83",
          5176 => x"81",
          5177 => x"53",
          5178 => x"ff",
          5179 => x"80",
          5180 => x"77",
          5181 => x"79",
          5182 => x"84",
          5183 => x"57",
          5184 => x"81",
          5185 => x"11",
          5186 => x"71",
          5187 => x"72",
          5188 => x"5e",
          5189 => x"84",
          5190 => x"06",
          5191 => x"11",
          5192 => x"71",
          5193 => x"72",
          5194 => x"47",
          5195 => x"86",
          5196 => x"06",
          5197 => x"11",
          5198 => x"71",
          5199 => x"72",
          5200 => x"94",
          5201 => x"11",
          5202 => x"71",
          5203 => x"72",
          5204 => x"62",
          5205 => x"5c",
          5206 => x"77",
          5207 => x"5d",
          5208 => x"18",
          5209 => x"0c",
          5210 => x"39",
          5211 => x"7a",
          5212 => x"54",
          5213 => x"53",
          5214 => x"b3",
          5215 => x"09",
          5216 => x"8c",
          5217 => x"a8",
          5218 => x"08",
          5219 => x"60",
          5220 => x"8c",
          5221 => x"74",
          5222 => x"81",
          5223 => x"58",
          5224 => x"80",
          5225 => x"5f",
          5226 => x"88",
          5227 => x"80",
          5228 => x"33",
          5229 => x"81",
          5230 => x"75",
          5231 => x"7d",
          5232 => x"40",
          5233 => x"2e",
          5234 => x"39",
          5235 => x"3d",
          5236 => x"39",
          5237 => x"bf",
          5238 => x"18",
          5239 => x"33",
          5240 => x"39",
          5241 => x"33",
          5242 => x"5d",
          5243 => x"80",
          5244 => x"33",
          5245 => x"2e",
          5246 => x"ba",
          5247 => x"33",
          5248 => x"73",
          5249 => x"08",
          5250 => x"80",
          5251 => x"86",
          5252 => x"75",
          5253 => x"38",
          5254 => x"05",
          5255 => x"08",
          5256 => x"3d",
          5257 => x"0c",
          5258 => x"11",
          5259 => x"73",
          5260 => x"81",
          5261 => x"79",
          5262 => x"83",
          5263 => x"7e",
          5264 => x"33",
          5265 => x"9f",
          5266 => x"89",
          5267 => x"56",
          5268 => x"26",
          5269 => x"06",
          5270 => x"58",
          5271 => x"85",
          5272 => x"32",
          5273 => x"79",
          5274 => x"92",
          5275 => x"83",
          5276 => x"fe",
          5277 => x"7a",
          5278 => x"e6",
          5279 => x"fb",
          5280 => x"80",
          5281 => x"54",
          5282 => x"84",
          5283 => x"ba",
          5284 => x"80",
          5285 => x"56",
          5286 => x"0d",
          5287 => x"70",
          5288 => x"8c",
          5289 => x"2e",
          5290 => x"7c",
          5291 => x"2e",
          5292 => x"ea",
          5293 => x"bb",
          5294 => x"7a",
          5295 => x"11",
          5296 => x"07",
          5297 => x"56",
          5298 => x"0b",
          5299 => x"34",
          5300 => x"0b",
          5301 => x"8b",
          5302 => x"0b",
          5303 => x"34",
          5304 => x"a9",
          5305 => x"34",
          5306 => x"9e",
          5307 => x"7e",
          5308 => x"80",
          5309 => x"08",
          5310 => x"81",
          5311 => x"7c",
          5312 => x"79",
          5313 => x"05",
          5314 => x"80",
          5315 => x"06",
          5316 => x"fe",
          5317 => x"70",
          5318 => x"82",
          5319 => x"5e",
          5320 => x"06",
          5321 => x"2a",
          5322 => x"38",
          5323 => x"11",
          5324 => x"0c",
          5325 => x"71",
          5326 => x"40",
          5327 => x"38",
          5328 => x"11",
          5329 => x"71",
          5330 => x"72",
          5331 => x"70",
          5332 => x"51",
          5333 => x"1a",
          5334 => x"34",
          5335 => x"9c",
          5336 => x"55",
          5337 => x"80",
          5338 => x"0c",
          5339 => x"52",
          5340 => x"80",
          5341 => x"92",
          5342 => x"7d",
          5343 => x"78",
          5344 => x"8c",
          5345 => x"26",
          5346 => x"08",
          5347 => x"31",
          5348 => x"33",
          5349 => x"82",
          5350 => x"fc",
          5351 => x"fb",
          5352 => x"fb",
          5353 => x"fb",
          5354 => x"84",
          5355 => x"57",
          5356 => x"7a",
          5357 => x"39",
          5358 => x"98",
          5359 => x"5d",
          5360 => x"7c",
          5361 => x"79",
          5362 => x"8c",
          5363 => x"2e",
          5364 => x"81",
          5365 => x"08",
          5366 => x"74",
          5367 => x"84",
          5368 => x"17",
          5369 => x"56",
          5370 => x"81",
          5371 => x"81",
          5372 => x"55",
          5373 => x"d9",
          5374 => x"0b",
          5375 => x"16",
          5376 => x"71",
          5377 => x"5b",
          5378 => x"8f",
          5379 => x"80",
          5380 => x"a0",
          5381 => x"5e",
          5382 => x"9b",
          5383 => x"2e",
          5384 => x"a9",
          5385 => x"57",
          5386 => x"38",
          5387 => x"09",
          5388 => x"53",
          5389 => x"ff",
          5390 => x"80",
          5391 => x"76",
          5392 => x"1d",
          5393 => x"fb",
          5394 => x"39",
          5395 => x"16",
          5396 => x"ff",
          5397 => x"7d",
          5398 => x"84",
          5399 => x"16",
          5400 => x"8c",
          5401 => x"27",
          5402 => x"74",
          5403 => x"38",
          5404 => x"08",
          5405 => x"51",
          5406 => x"ec",
          5407 => x"f8",
          5408 => x"f8",
          5409 => x"79",
          5410 => x"19",
          5411 => x"5a",
          5412 => x"1a",
          5413 => x"05",
          5414 => x"38",
          5415 => x"76",
          5416 => x"0c",
          5417 => x"80",
          5418 => x"8c",
          5419 => x"39",
          5420 => x"f0",
          5421 => x"40",
          5422 => x"79",
          5423 => x"75",
          5424 => x"74",
          5425 => x"84",
          5426 => x"84",
          5427 => x"55",
          5428 => x"55",
          5429 => x"81",
          5430 => x"81",
          5431 => x"08",
          5432 => x"81",
          5433 => x"38",
          5434 => x"7a",
          5435 => x"05",
          5436 => x"38",
          5437 => x"55",
          5438 => x"ff",
          5439 => x"0c",
          5440 => x"9c",
          5441 => x"60",
          5442 => x"70",
          5443 => x"56",
          5444 => x"15",
          5445 => x"2e",
          5446 => x"75",
          5447 => x"77",
          5448 => x"33",
          5449 => x"8c",
          5450 => x"33",
          5451 => x"b4",
          5452 => x"27",
          5453 => x"1e",
          5454 => x"81",
          5455 => x"59",
          5456 => x"77",
          5457 => x"08",
          5458 => x"08",
          5459 => x"5c",
          5460 => x"84",
          5461 => x"74",
          5462 => x"04",
          5463 => x"08",
          5464 => x"71",
          5465 => x"38",
          5466 => x"77",
          5467 => x"33",
          5468 => x"09",
          5469 => x"76",
          5470 => x"51",
          5471 => x"08",
          5472 => x"5b",
          5473 => x"38",
          5474 => x"11",
          5475 => x"59",
          5476 => x"70",
          5477 => x"05",
          5478 => x"2e",
          5479 => x"56",
          5480 => x"ff",
          5481 => x"39",
          5482 => x"19",
          5483 => x"ff",
          5484 => x"8c",
          5485 => x"9c",
          5486 => x"34",
          5487 => x"84",
          5488 => x"1a",
          5489 => x"33",
          5490 => x"fe",
          5491 => x"a0",
          5492 => x"19",
          5493 => x"5b",
          5494 => x"94",
          5495 => x"1a",
          5496 => x"3f",
          5497 => x"39",
          5498 => x"3f",
          5499 => x"74",
          5500 => x"57",
          5501 => x"34",
          5502 => x"3d",
          5503 => x"82",
          5504 => x"0d",
          5505 => x"66",
          5506 => x"89",
          5507 => x"08",
          5508 => x"33",
          5509 => x"16",
          5510 => x"78",
          5511 => x"41",
          5512 => x"1a",
          5513 => x"1a",
          5514 => x"58",
          5515 => x"38",
          5516 => x"7b",
          5517 => x"7a",
          5518 => x"ff",
          5519 => x"8a",
          5520 => x"06",
          5521 => x"9e",
          5522 => x"2e",
          5523 => x"a1",
          5524 => x"74",
          5525 => x"38",
          5526 => x"16",
          5527 => x"38",
          5528 => x"08",
          5529 => x"85",
          5530 => x"29",
          5531 => x"80",
          5532 => x"89",
          5533 => x"98",
          5534 => x"85",
          5535 => x"7b",
          5536 => x"ff",
          5537 => x"85",
          5538 => x"31",
          5539 => x"84",
          5540 => x"1f",
          5541 => x"56",
          5542 => x"ff",
          5543 => x"75",
          5544 => x"7a",
          5545 => x"79",
          5546 => x"94",
          5547 => x"57",
          5548 => x"74",
          5549 => x"85",
          5550 => x"c0",
          5551 => x"56",
          5552 => x"0d",
          5553 => x"3d",
          5554 => x"82",
          5555 => x"60",
          5556 => x"ff",
          5557 => x"7a",
          5558 => x"57",
          5559 => x"80",
          5560 => x"5f",
          5561 => x"d5",
          5562 => x"52",
          5563 => x"3f",
          5564 => x"38",
          5565 => x"0c",
          5566 => x"08",
          5567 => x"05",
          5568 => x"95",
          5569 => x"75",
          5570 => x"56",
          5571 => x"83",
          5572 => x"b4",
          5573 => x"81",
          5574 => x"3f",
          5575 => x"2e",
          5576 => x"ba",
          5577 => x"08",
          5578 => x"08",
          5579 => x"fe",
          5580 => x"82",
          5581 => x"81",
          5582 => x"05",
          5583 => x"ff",
          5584 => x"39",
          5585 => x"77",
          5586 => x"7f",
          5587 => x"0c",
          5588 => x"9c",
          5589 => x"1a",
          5590 => x"3f",
          5591 => x"8c",
          5592 => x"58",
          5593 => x"ff",
          5594 => x"55",
          5595 => x"e4",
          5596 => x"b8",
          5597 => x"57",
          5598 => x"08",
          5599 => x"83",
          5600 => x"08",
          5601 => x"fd",
          5602 => x"82",
          5603 => x"81",
          5604 => x"05",
          5605 => x"ff",
          5606 => x"39",
          5607 => x"3f",
          5608 => x"74",
          5609 => x"57",
          5610 => x"08",
          5611 => x"33",
          5612 => x"ba",
          5613 => x"8c",
          5614 => x"a8",
          5615 => x"08",
          5616 => x"58",
          5617 => x"8b",
          5618 => x"17",
          5619 => x"33",
          5620 => x"b4",
          5621 => x"fd",
          5622 => x"81",
          5623 => x"0d",
          5624 => x"0b",
          5625 => x"04",
          5626 => x"77",
          5627 => x"75",
          5628 => x"74",
          5629 => x"84",
          5630 => x"83",
          5631 => x"56",
          5632 => x"70",
          5633 => x"80",
          5634 => x"08",
          5635 => x"ac",
          5636 => x"bc",
          5637 => x"52",
          5638 => x"3f",
          5639 => x"38",
          5640 => x"0c",
          5641 => x"8b",
          5642 => x"8b",
          5643 => x"70",
          5644 => x"7a",
          5645 => x"79",
          5646 => x"96",
          5647 => x"81",
          5648 => x"7b",
          5649 => x"18",
          5650 => x"18",
          5651 => x"18",
          5652 => x"18",
          5653 => x"cc",
          5654 => x"18",
          5655 => x"5b",
          5656 => x"ff",
          5657 => x"90",
          5658 => x"79",
          5659 => x"0c",
          5660 => x"17",
          5661 => x"18",
          5662 => x"81",
          5663 => x"38",
          5664 => x"b4",
          5665 => x"ba",
          5666 => x"08",
          5667 => x"55",
          5668 => x"81",
          5669 => x"18",
          5670 => x"33",
          5671 => x"fd",
          5672 => x"94",
          5673 => x"95",
          5674 => x"7b",
          5675 => x"18",
          5676 => x"18",
          5677 => x"18",
          5678 => x"18",
          5679 => x"cc",
          5680 => x"18",
          5681 => x"5b",
          5682 => x"ff",
          5683 => x"90",
          5684 => x"79",
          5685 => x"16",
          5686 => x"ba",
          5687 => x"ba",
          5688 => x"b4",
          5689 => x"55",
          5690 => x"54",
          5691 => x"56",
          5692 => x"53",
          5693 => x"52",
          5694 => x"22",
          5695 => x"2e",
          5696 => x"54",
          5697 => x"84",
          5698 => x"81",
          5699 => x"84",
          5700 => x"da",
          5701 => x"39",
          5702 => x"57",
          5703 => x"70",
          5704 => x"52",
          5705 => x"ee",
          5706 => x"d1",
          5707 => x"38",
          5708 => x"84",
          5709 => x"8b",
          5710 => x"0d",
          5711 => x"ff",
          5712 => x"91",
          5713 => x"d0",
          5714 => x"f5",
          5715 => x"58",
          5716 => x"81",
          5717 => x"57",
          5718 => x"70",
          5719 => x"81",
          5720 => x"51",
          5721 => x"70",
          5722 => x"70",
          5723 => x"09",
          5724 => x"38",
          5725 => x"07",
          5726 => x"76",
          5727 => x"1b",
          5728 => x"38",
          5729 => x"24",
          5730 => x"c3",
          5731 => x"3d",
          5732 => x"94",
          5733 => x"ba",
          5734 => x"84",
          5735 => x"7a",
          5736 => x"51",
          5737 => x"55",
          5738 => x"02",
          5739 => x"58",
          5740 => x"02",
          5741 => x"06",
          5742 => x"7a",
          5743 => x"71",
          5744 => x"5b",
          5745 => x"76",
          5746 => x"0c",
          5747 => x"08",
          5748 => x"38",
          5749 => x"3d",
          5750 => x"33",
          5751 => x"79",
          5752 => x"39",
          5753 => x"84",
          5754 => x"ff",
          5755 => x"80",
          5756 => x"34",
          5757 => x"05",
          5758 => x"3f",
          5759 => x"8c",
          5760 => x"3d",
          5761 => x"dd",
          5762 => x"5b",
          5763 => x"80",
          5764 => x"52",
          5765 => x"ba",
          5766 => x"83",
          5767 => x"58",
          5768 => x"38",
          5769 => x"5f",
          5770 => x"76",
          5771 => x"51",
          5772 => x"08",
          5773 => x"59",
          5774 => x"38",
          5775 => x"9a",
          5776 => x"70",
          5777 => x"83",
          5778 => x"3d",
          5779 => x"b7",
          5780 => x"ba",
          5781 => x"7a",
          5782 => x"8c",
          5783 => x"38",
          5784 => x"9a",
          5785 => x"70",
          5786 => x"83",
          5787 => x"a4",
          5788 => x"51",
          5789 => x"08",
          5790 => x"ff",
          5791 => x"38",
          5792 => x"fd",
          5793 => x"89",
          5794 => x"57",
          5795 => x"56",
          5796 => x"57",
          5797 => x"75",
          5798 => x"2e",
          5799 => x"ff",
          5800 => x"19",
          5801 => x"33",
          5802 => x"80",
          5803 => x"7e",
          5804 => x"fd",
          5805 => x"38",
          5806 => x"10",
          5807 => x"70",
          5808 => x"7a",
          5809 => x"70",
          5810 => x"82",
          5811 => x"80",
          5812 => x"16",
          5813 => x"5e",
          5814 => x"ee",
          5815 => x"34",
          5816 => x"df",
          5817 => x"84",
          5818 => x"04",
          5819 => x"98",
          5820 => x"59",
          5821 => x"33",
          5822 => x"90",
          5823 => x"0c",
          5824 => x"a0",
          5825 => x"84",
          5826 => x"38",
          5827 => x"08",
          5828 => x"33",
          5829 => x"59",
          5830 => x"84",
          5831 => x"16",
          5832 => x"8c",
          5833 => x"27",
          5834 => x"74",
          5835 => x"38",
          5836 => x"08",
          5837 => x"51",
          5838 => x"dd",
          5839 => x"11",
          5840 => x"84",
          5841 => x"e5",
          5842 => x"59",
          5843 => x"81",
          5844 => x"80",
          5845 => x"5a",
          5846 => x"34",
          5847 => x"e5",
          5848 => x"79",
          5849 => x"7f",
          5850 => x"82",
          5851 => x"8c",
          5852 => x"3d",
          5853 => x"74",
          5854 => x"73",
          5855 => x"72",
          5856 => x"84",
          5857 => x"83",
          5858 => x"53",
          5859 => x"53",
          5860 => x"56",
          5861 => x"15",
          5862 => x"81",
          5863 => x"89",
          5864 => x"81",
          5865 => x"fd",
          5866 => x"ff",
          5867 => x"fd",
          5868 => x"73",
          5869 => x"06",
          5870 => x"98",
          5871 => x"2e",
          5872 => x"d9",
          5873 => x"17",
          5874 => x"81",
          5875 => x"80",
          5876 => x"51",
          5877 => x"08",
          5878 => x"81",
          5879 => x"81",
          5880 => x"73",
          5881 => x"73",
          5882 => x"0b",
          5883 => x"ba",
          5884 => x"15",
          5885 => x"58",
          5886 => x"08",
          5887 => x"09",
          5888 => x"16",
          5889 => x"27",
          5890 => x"15",
          5891 => x"16",
          5892 => x"80",
          5893 => x"2e",
          5894 => x"0b",
          5895 => x"04",
          5896 => x"08",
          5897 => x"73",
          5898 => x"c2",
          5899 => x"08",
          5900 => x"0c",
          5901 => x"2e",
          5902 => x"08",
          5903 => x"27",
          5904 => x"71",
          5905 => x"2a",
          5906 => x"80",
          5907 => x"e9",
          5908 => x"b7",
          5909 => x"8a",
          5910 => x"a2",
          5911 => x"53",
          5912 => x"54",
          5913 => x"51",
          5914 => x"08",
          5915 => x"98",
          5916 => x"fd",
          5917 => x"16",
          5918 => x"39",
          5919 => x"84",
          5920 => x"f6",
          5921 => x"80",
          5922 => x"fc",
          5923 => x"c5",
          5924 => x"84",
          5925 => x"80",
          5926 => x"8c",
          5927 => x"0c",
          5928 => x"3f",
          5929 => x"8c",
          5930 => x"70",
          5931 => x"af",
          5932 => x"81",
          5933 => x"c5",
          5934 => x"9a",
          5935 => x"70",
          5936 => x"83",
          5937 => x"7a",
          5938 => x"74",
          5939 => x"84",
          5940 => x"8d",
          5941 => x"80",
          5942 => x"80",
          5943 => x"33",
          5944 => x"90",
          5945 => x"5a",
          5946 => x"78",
          5947 => x"38",
          5948 => x"38",
          5949 => x"38",
          5950 => x"52",
          5951 => x"71",
          5952 => x"73",
          5953 => x"04",
          5954 => x"3f",
          5955 => x"71",
          5956 => x"d7",
          5957 => x"55",
          5958 => x"74",
          5959 => x"73",
          5960 => x"86",
          5961 => x"72",
          5962 => x"72",
          5963 => x"76",
          5964 => x"74",
          5965 => x"8c",
          5966 => x"2e",
          5967 => x"38",
          5968 => x"3f",
          5969 => x"3f",
          5970 => x"30",
          5971 => x"8c",
          5972 => x"ba",
          5973 => x"77",
          5974 => x"3f",
          5975 => x"3f",
          5976 => x"30",
          5977 => x"8c",
          5978 => x"75",
          5979 => x"84",
          5980 => x"8a",
          5981 => x"fe",
          5982 => x"81",
          5983 => x"75",
          5984 => x"3d",
          5985 => x"70",
          5986 => x"3f",
          5987 => x"8c",
          5988 => x"ba",
          5989 => x"52",
          5990 => x"ba",
          5991 => x"e5",
          5992 => x"98",
          5993 => x"38",
          5994 => x"75",
          5995 => x"ba",
          5996 => x"0b",
          5997 => x"04",
          5998 => x"80",
          5999 => x"3d",
          6000 => x"08",
          6001 => x"7f",
          6002 => x"fe",
          6003 => x"57",
          6004 => x"0c",
          6005 => x"0d",
          6006 => x"5a",
          6007 => x"77",
          6008 => x"5a",
          6009 => x"81",
          6010 => x"08",
          6011 => x"33",
          6012 => x"81",
          6013 => x"17",
          6014 => x"ba",
          6015 => x"5a",
          6016 => x"7e",
          6017 => x"33",
          6018 => x"77",
          6019 => x"12",
          6020 => x"07",
          6021 => x"2b",
          6022 => x"80",
          6023 => x"63",
          6024 => x"62",
          6025 => x"52",
          6026 => x"f2",
          6027 => x"0c",
          6028 => x"84",
          6029 => x"95",
          6030 => x"08",
          6031 => x"33",
          6032 => x"5e",
          6033 => x"84",
          6034 => x"17",
          6035 => x"8c",
          6036 => x"27",
          6037 => x"74",
          6038 => x"38",
          6039 => x"08",
          6040 => x"51",
          6041 => x"97",
          6042 => x"56",
          6043 => x"3f",
          6044 => x"e8",
          6045 => x"80",
          6046 => x"70",
          6047 => x"7c",
          6048 => x"5c",
          6049 => x"7a",
          6050 => x"17",
          6051 => x"34",
          6052 => x"81",
          6053 => x"07",
          6054 => x"1d",
          6055 => x"5f",
          6056 => x"38",
          6057 => x"39",
          6058 => x"7a",
          6059 => x"07",
          6060 => x"39",
          6061 => x"3d",
          6062 => x"2e",
          6063 => x"2e",
          6064 => x"2e",
          6065 => x"22",
          6066 => x"38",
          6067 => x"38",
          6068 => x"38",
          6069 => x"06",
          6070 => x"80",
          6071 => x"8c",
          6072 => x"d5",
          6073 => x"54",
          6074 => x"08",
          6075 => x"0b",
          6076 => x"18",
          6077 => x"90",
          6078 => x"75",
          6079 => x"ba",
          6080 => x"54",
          6081 => x"52",
          6082 => x"ba",
          6083 => x"80",
          6084 => x"08",
          6085 => x"8c",
          6086 => x"53",
          6087 => x"3f",
          6088 => x"9c",
          6089 => x"57",
          6090 => x"38",
          6091 => x"33",
          6092 => x"78",
          6093 => x"9c",
          6094 => x"e2",
          6095 => x"54",
          6096 => x"55",
          6097 => x"18",
          6098 => x"88",
          6099 => x"08",
          6100 => x"84",
          6101 => x"38",
          6102 => x"be",
          6103 => x"84",
          6104 => x"81",
          6105 => x"18",
          6106 => x"0b",
          6107 => x"38",
          6108 => x"27",
          6109 => x"38",
          6110 => x"83",
          6111 => x"84",
          6112 => x"52",
          6113 => x"ba",
          6114 => x"80",
          6115 => x"08",
          6116 => x"8c",
          6117 => x"53",
          6118 => x"3f",
          6119 => x"9c",
          6120 => x"57",
          6121 => x"81",
          6122 => x"81",
          6123 => x"54",
          6124 => x"55",
          6125 => x"f3",
          6126 => x"0b",
          6127 => x"39",
          6128 => x"18",
          6129 => x"ba",
          6130 => x"fd",
          6131 => x"59",
          6132 => x"08",
          6133 => x"39",
          6134 => x"ff",
          6135 => x"b7",
          6136 => x"84",
          6137 => x"75",
          6138 => x"04",
          6139 => x"3d",
          6140 => x"84",
          6141 => x"08",
          6142 => x"70",
          6143 => x"56",
          6144 => x"80",
          6145 => x"05",
          6146 => x"56",
          6147 => x"08",
          6148 => x"88",
          6149 => x"57",
          6150 => x"76",
          6151 => x"2e",
          6152 => x"08",
          6153 => x"7a",
          6154 => x"3d",
          6155 => x"84",
          6156 => x"08",
          6157 => x"52",
          6158 => x"ba",
          6159 => x"a0",
          6160 => x"a7",
          6161 => x"17",
          6162 => x"07",
          6163 => x"39",
          6164 => x"38",
          6165 => x"78",
          6166 => x"57",
          6167 => x"52",
          6168 => x"ba",
          6169 => x"80",
          6170 => x"07",
          6171 => x"9a",
          6172 => x"79",
          6173 => x"38",
          6174 => x"38",
          6175 => x"51",
          6176 => x"08",
          6177 => x"04",
          6178 => x"80",
          6179 => x"b9",
          6180 => x"74",
          6181 => x"38",
          6182 => x"81",
          6183 => x"84",
          6184 => x"ff",
          6185 => x"77",
          6186 => x"58",
          6187 => x"34",
          6188 => x"38",
          6189 => x"3f",
          6190 => x"8c",
          6191 => x"84",
          6192 => x"82",
          6193 => x"17",
          6194 => x"51",
          6195 => x"ba",
          6196 => x"ff",
          6197 => x"18",
          6198 => x"31",
          6199 => x"a0",
          6200 => x"17",
          6201 => x"06",
          6202 => x"08",
          6203 => x"81",
          6204 => x"79",
          6205 => x"78",
          6206 => x"51",
          6207 => x"08",
          6208 => x"80",
          6209 => x"2e",
          6210 => x"ff",
          6211 => x"52",
          6212 => x"ba",
          6213 => x"fe",
          6214 => x"75",
          6215 => x"94",
          6216 => x"5c",
          6217 => x"7a",
          6218 => x"a2",
          6219 => x"ba",
          6220 => x"56",
          6221 => x"53",
          6222 => x"3d",
          6223 => x"8c",
          6224 => x"2e",
          6225 => x"9f",
          6226 => x"93",
          6227 => x"3f",
          6228 => x"8c",
          6229 => x"8c",
          6230 => x"8c",
          6231 => x"38",
          6232 => x"2a",
          6233 => x"ff",
          6234 => x"3d",
          6235 => x"84",
          6236 => x"ba",
          6237 => x"ba",
          6238 => x"84",
          6239 => x"38",
          6240 => x"8c",
          6241 => x"7a",
          6242 => x"08",
          6243 => x"79",
          6244 => x"71",
          6245 => x"7a",
          6246 => x"80",
          6247 => x"05",
          6248 => x"38",
          6249 => x"75",
          6250 => x"1b",
          6251 => x"fe",
          6252 => x"81",
          6253 => x"82",
          6254 => x"17",
          6255 => x"18",
          6256 => x"81",
          6257 => x"84",
          6258 => x"17",
          6259 => x"a0",
          6260 => x"17",
          6261 => x"06",
          6262 => x"08",
          6263 => x"81",
          6264 => x"fe",
          6265 => x"58",
          6266 => x"7b",
          6267 => x"74",
          6268 => x"84",
          6269 => x"08",
          6270 => x"8c",
          6271 => x"ba",
          6272 => x"80",
          6273 => x"b0",
          6274 => x"38",
          6275 => x"08",
          6276 => x"38",
          6277 => x"33",
          6278 => x"79",
          6279 => x"75",
          6280 => x"04",
          6281 => x"ff",
          6282 => x"09",
          6283 => x"b8",
          6284 => x"05",
          6285 => x"38",
          6286 => x"7d",
          6287 => x"7d",
          6288 => x"80",
          6289 => x"1a",
          6290 => x"34",
          6291 => x"56",
          6292 => x"2a",
          6293 => x"33",
          6294 => x"7d",
          6295 => x"1b",
          6296 => x"56",
          6297 => x"ff",
          6298 => x"ae",
          6299 => x"71",
          6300 => x"78",
          6301 => x"5b",
          6302 => x"55",
          6303 => x"5b",
          6304 => x"ff",
          6305 => x"56",
          6306 => x"69",
          6307 => x"34",
          6308 => x"a1",
          6309 => x"99",
          6310 => x"9a",
          6311 => x"9b",
          6312 => x"2e",
          6313 => x"8b",
          6314 => x"18",
          6315 => x"84",
          6316 => x"8c",
          6317 => x"2a",
          6318 => x"88",
          6319 => x"fe",
          6320 => x"80",
          6321 => x"74",
          6322 => x"0b",
          6323 => x"56",
          6324 => x"77",
          6325 => x"7b",
          6326 => x"8b",
          6327 => x"18",
          6328 => x"84",
          6329 => x"d1",
          6330 => x"70",
          6331 => x"38",
          6332 => x"9f",
          6333 => x"b8",
          6334 => x"81",
          6335 => x"fc",
          6336 => x"b4",
          6337 => x"ba",
          6338 => x"84",
          6339 => x"7f",
          6340 => x"a5",
          6341 => x"3f",
          6342 => x"8c",
          6343 => x"33",
          6344 => x"ce",
          6345 => x"08",
          6346 => x"57",
          6347 => x"ff",
          6348 => x"58",
          6349 => x"70",
          6350 => x"05",
          6351 => x"38",
          6352 => x"9e",
          6353 => x"84",
          6354 => x"a8",
          6355 => x"0b",
          6356 => x"04",
          6357 => x"06",
          6358 => x"38",
          6359 => x"05",
          6360 => x"38",
          6361 => x"08",
          6362 => x"70",
          6363 => x"05",
          6364 => x"56",
          6365 => x"70",
          6366 => x"17",
          6367 => x"17",
          6368 => x"30",
          6369 => x"2e",
          6370 => x"be",
          6371 => x"72",
          6372 => x"55",
          6373 => x"84",
          6374 => x"c2",
          6375 => x"96",
          6376 => x"79",
          6377 => x"fc",
          6378 => x"e4",
          6379 => x"ba",
          6380 => x"39",
          6381 => x"06",
          6382 => x"a8",
          6383 => x"ba",
          6384 => x"93",
          6385 => x"cd",
          6386 => x"05",
          6387 => x"34",
          6388 => x"80",
          6389 => x"18",
          6390 => x"56",
          6391 => x"76",
          6392 => x"83",
          6393 => x"2a",
          6394 => x"81",
          6395 => x"81",
          6396 => x"1a",
          6397 => x"41",
          6398 => x"e0",
          6399 => x"05",
          6400 => x"38",
          6401 => x"19",
          6402 => x"82",
          6403 => x"17",
          6404 => x"33",
          6405 => x"75",
          6406 => x"51",
          6407 => x"08",
          6408 => x"5c",
          6409 => x"80",
          6410 => x"38",
          6411 => x"09",
          6412 => x"ff",
          6413 => x"18",
          6414 => x"f3",
          6415 => x"2e",
          6416 => x"2a",
          6417 => x"88",
          6418 => x"7f",
          6419 => x"08",
          6420 => x"5c",
          6421 => x"52",
          6422 => x"ba",
          6423 => x"80",
          6424 => x"08",
          6425 => x"2e",
          6426 => x"5f",
          6427 => x"a8",
          6428 => x"52",
          6429 => x"3f",
          6430 => x"38",
          6431 => x"0c",
          6432 => x"08",
          6433 => x"17",
          6434 => x"38",
          6435 => x"3f",
          6436 => x"8c",
          6437 => x"56",
          6438 => x"56",
          6439 => x"e5",
          6440 => x"ba",
          6441 => x"0b",
          6442 => x"04",
          6443 => x"98",
          6444 => x"58",
          6445 => x"8c",
          6446 => x"ba",
          6447 => x"75",
          6448 => x"04",
          6449 => x"52",
          6450 => x"3f",
          6451 => x"2e",
          6452 => x"ba",
          6453 => x"08",
          6454 => x"08",
          6455 => x"fe",
          6456 => x"82",
          6457 => x"81",
          6458 => x"05",
          6459 => x"fe",
          6460 => x"39",
          6461 => x"17",
          6462 => x"fe",
          6463 => x"8c",
          6464 => x"08",
          6465 => x"18",
          6466 => x"55",
          6467 => x"38",
          6468 => x"09",
          6469 => x"b4",
          6470 => x"7a",
          6471 => x"eb",
          6472 => x"3d",
          6473 => x"84",
          6474 => x"82",
          6475 => x"3d",
          6476 => x"8c",
          6477 => x"2e",
          6478 => x"96",
          6479 => x"96",
          6480 => x"3f",
          6481 => x"8c",
          6482 => x"33",
          6483 => x"d2",
          6484 => x"8b",
          6485 => x"07",
          6486 => x"34",
          6487 => x"78",
          6488 => x"8c",
          6489 => x"0d",
          6490 => x"53",
          6491 => x"51",
          6492 => x"08",
          6493 => x"8a",
          6494 => x"3d",
          6495 => x"3d",
          6496 => x"84",
          6497 => x"08",
          6498 => x"81",
          6499 => x"38",
          6500 => x"71",
          6501 => x"96",
          6502 => x"97",
          6503 => x"98",
          6504 => x"99",
          6505 => x"18",
          6506 => x"84",
          6507 => x"96",
          6508 => x"6d",
          6509 => x"05",
          6510 => x"3f",
          6511 => x"08",
          6512 => x"80",
          6513 => x"8b",
          6514 => x"78",
          6515 => x"07",
          6516 => x"81",
          6517 => x"58",
          6518 => x"a4",
          6519 => x"16",
          6520 => x"16",
          6521 => x"09",
          6522 => x"76",
          6523 => x"51",
          6524 => x"08",
          6525 => x"59",
          6526 => x"bd",
          6527 => x"c3",
          6528 => x"e4",
          6529 => x"56",
          6530 => x"82",
          6531 => x"2b",
          6532 => x"88",
          6533 => x"5f",
          6534 => x"ba",
          6535 => x"5e",
          6536 => x"52",
          6537 => x"8c",
          6538 => x"2e",
          6539 => x"81",
          6540 => x"80",
          6541 => x"16",
          6542 => x"17",
          6543 => x"77",
          6544 => x"09",
          6545 => x"8c",
          6546 => x"a8",
          6547 => x"5a",
          6548 => x"ad",
          6549 => x"2e",
          6550 => x"54",
          6551 => x"53",
          6552 => x"db",
          6553 => x"53",
          6554 => x"fe",
          6555 => x"80",
          6556 => x"75",
          6557 => x"84",
          6558 => x"08",
          6559 => x"84",
          6560 => x"79",
          6561 => x"56",
          6562 => x"8a",
          6563 => x"57",
          6564 => x"fc",
          6565 => x"33",
          6566 => x"38",
          6567 => x"39",
          6568 => x"ff",
          6569 => x"9c",
          6570 => x"84",
          6571 => x"3d",
          6572 => x"70",
          6573 => x"74",
          6574 => x"33",
          6575 => x"5a",
          6576 => x"3d",
          6577 => x"06",
          6578 => x"38",
          6579 => x"26",
          6580 => x"3f",
          6581 => x"51",
          6582 => x"83",
          6583 => x"81",
          6584 => x"e7",
          6585 => x"56",
          6586 => x"74",
          6587 => x"18",
          6588 => x"57",
          6589 => x"77",
          6590 => x"81",
          6591 => x"81",
          6592 => x"89",
          6593 => x"27",
          6594 => x"7b",
          6595 => x"5a",
          6596 => x"81",
          6597 => x"81",
          6598 => x"9f",
          6599 => x"57",
          6600 => x"38",
          6601 => x"05",
          6602 => x"7a",
          6603 => x"ff",
          6604 => x"80",
          6605 => x"56",
          6606 => x"08",
          6607 => x"b4",
          6608 => x"0c",
          6609 => x"74",
          6610 => x"08",
          6611 => x"f8",
          6612 => x"0c",
          6613 => x"33",
          6614 => x"51",
          6615 => x"08",
          6616 => x"38",
          6617 => x"6c",
          6618 => x"05",
          6619 => x"34",
          6620 => x"5d",
          6621 => x"fe",
          6622 => x"55",
          6623 => x"27",
          6624 => x"39",
          6625 => x"81",
          6626 => x"75",
          6627 => x"53",
          6628 => x"84",
          6629 => x"08",
          6630 => x"38",
          6631 => x"5a",
          6632 => x"18",
          6633 => x"33",
          6634 => x"81",
          6635 => x"18",
          6636 => x"c4",
          6637 => x"85",
          6638 => x"19",
          6639 => x"9c",
          6640 => x"74",
          6641 => x"30",
          6642 => x"74",
          6643 => x"5a",
          6644 => x"75",
          6645 => x"8c",
          6646 => x"2e",
          6647 => x"2e",
          6648 => x"b9",
          6649 => x"70",
          6650 => x"74",
          6651 => x"17",
          6652 => x"76",
          6653 => x"81",
          6654 => x"80",
          6655 => x"05",
          6656 => x"34",
          6657 => x"d6",
          6658 => x"5d",
          6659 => x"fe",
          6660 => x"55",
          6661 => x"39",
          6662 => x"52",
          6663 => x"3f",
          6664 => x"81",
          6665 => x"08",
          6666 => x"19",
          6667 => x"27",
          6668 => x"82",
          6669 => x"59",
          6670 => x"75",
          6671 => x"8c",
          6672 => x"2e",
          6673 => x"70",
          6674 => x"38",
          6675 => x"08",
          6676 => x"81",
          6677 => x"fd",
          6678 => x"02",
          6679 => x"5b",
          6680 => x"38",
          6681 => x"38",
          6682 => x"38",
          6683 => x"59",
          6684 => x"54",
          6685 => x"17",
          6686 => x"80",
          6687 => x"81",
          6688 => x"2a",
          6689 => x"81",
          6690 => x"89",
          6691 => x"59",
          6692 => x"06",
          6693 => x"84",
          6694 => x"79",
          6695 => x"27",
          6696 => x"83",
          6697 => x"80",
          6698 => x"87",
          6699 => x"14",
          6700 => x"84",
          6701 => x"38",
          6702 => x"d8",
          6703 => x"38",
          6704 => x"38",
          6705 => x"38",
          6706 => x"8c",
          6707 => x"84",
          6708 => x"81",
          6709 => x"84",
          6710 => x"fe",
          6711 => x"fe",
          6712 => x"38",
          6713 => x"ab",
          6714 => x"80",
          6715 => x"51",
          6716 => x"08",
          6717 => x"38",
          6718 => x"5e",
          6719 => x"0c",
          6720 => x"7a",
          6721 => x"90",
          6722 => x"90",
          6723 => x"94",
          6724 => x"fe",
          6725 => x"0c",
          6726 => x"84",
          6727 => x"ff",
          6728 => x"59",
          6729 => x"39",
          6730 => x"5e",
          6731 => x"e3",
          6732 => x"08",
          6733 => x"44",
          6734 => x"70",
          6735 => x"8a",
          6736 => x"70",
          6737 => x"85",
          6738 => x"2e",
          6739 => x"56",
          6740 => x"10",
          6741 => x"56",
          6742 => x"75",
          6743 => x"33",
          6744 => x"5d",
          6745 => x"3f",
          6746 => x"70",
          6747 => x"84",
          6748 => x"40",
          6749 => x"3d",
          6750 => x"fe",
          6751 => x"84",
          6752 => x"84",
          6753 => x"84",
          6754 => x"74",
          6755 => x"38",
          6756 => x"7e",
          6757 => x"ff",
          6758 => x"38",
          6759 => x"2a",
          6760 => x"5b",
          6761 => x"30",
          6762 => x"91",
          6763 => x"2e",
          6764 => x"60",
          6765 => x"81",
          6766 => x"38",
          6767 => x"fe",
          6768 => x"56",
          6769 => x"09",
          6770 => x"29",
          6771 => x"58",
          6772 => x"b6",
          6773 => x"71",
          6774 => x"14",
          6775 => x"33",
          6776 => x"33",
          6777 => x"88",
          6778 => x"07",
          6779 => x"a2",
          6780 => x"3d",
          6781 => x"41",
          6782 => x"ff",
          6783 => x"7a",
          6784 => x"81",
          6785 => x"80",
          6786 => x"45",
          6787 => x"06",
          6788 => x"70",
          6789 => x"83",
          6790 => x"78",
          6791 => x"b0",
          6792 => x"38",
          6793 => x"b0",
          6794 => x"57",
          6795 => x"76",
          6796 => x"51",
          6797 => x"08",
          6798 => x"08",
          6799 => x"84",
          6800 => x"08",
          6801 => x"57",
          6802 => x"5d",
          6803 => x"11",
          6804 => x"6b",
          6805 => x"62",
          6806 => x"5d",
          6807 => x"56",
          6808 => x"78",
          6809 => x"68",
          6810 => x"84",
          6811 => x"89",
          6812 => x"06",
          6813 => x"84",
          6814 => x"7a",
          6815 => x"80",
          6816 => x"fe",
          6817 => x"8c",
          6818 => x"0c",
          6819 => x"0b",
          6820 => x"84",
          6821 => x"11",
          6822 => x"74",
          6823 => x"81",
          6824 => x"7a",
          6825 => x"e5",
          6826 => x"5b",
          6827 => x"70",
          6828 => x"45",
          6829 => x"e0",
          6830 => x"ff",
          6831 => x"38",
          6832 => x"46",
          6833 => x"76",
          6834 => x"78",
          6835 => x"30",
          6836 => x"5d",
          6837 => x"38",
          6838 => x"7c",
          6839 => x"e0",
          6840 => x"52",
          6841 => x"57",
          6842 => x"61",
          6843 => x"08",
          6844 => x"6c",
          6845 => x"9c",
          6846 => x"39",
          6847 => x"24",
          6848 => x"0c",
          6849 => x"48",
          6850 => x"38",
          6851 => x"fc",
          6852 => x"f5",
          6853 => x"18",
          6854 => x"38",
          6855 => x"9f",
          6856 => x"80",
          6857 => x"9f",
          6858 => x"06",
          6859 => x"84",
          6860 => x"81",
          6861 => x"f4",
          6862 => x"57",
          6863 => x"76",
          6864 => x"55",
          6865 => x"74",
          6866 => x"77",
          6867 => x"ff",
          6868 => x"6a",
          6869 => x"34",
          6870 => x"32",
          6871 => x"05",
          6872 => x"68",
          6873 => x"83",
          6874 => x"83",
          6875 => x"05",
          6876 => x"94",
          6877 => x"bf",
          6878 => x"05",
          6879 => x"61",
          6880 => x"34",
          6881 => x"05",
          6882 => x"9e",
          6883 => x"98",
          6884 => x"05",
          6885 => x"80",
          6886 => x"05",
          6887 => x"cc",
          6888 => x"ff",
          6889 => x"74",
          6890 => x"34",
          6891 => x"61",
          6892 => x"83",
          6893 => x"81",
          6894 => x"58",
          6895 => x"60",
          6896 => x"34",
          6897 => x"6b",
          6898 => x"79",
          6899 => x"84",
          6900 => x"17",
          6901 => x"69",
          6902 => x"05",
          6903 => x"38",
          6904 => x"86",
          6905 => x"62",
          6906 => x"61",
          6907 => x"74",
          6908 => x"90",
          6909 => x"46",
          6910 => x"34",
          6911 => x"83",
          6912 => x"60",
          6913 => x"84",
          6914 => x"80",
          6915 => x"05",
          6916 => x"38",
          6917 => x"76",
          6918 => x"80",
          6919 => x"83",
          6920 => x"75",
          6921 => x"54",
          6922 => x"c4",
          6923 => x"9b",
          6924 => x"5b",
          6925 => x"2e",
          6926 => x"ff",
          6927 => x"2e",
          6928 => x"38",
          6929 => x"81",
          6930 => x"80",
          6931 => x"19",
          6932 => x"34",
          6933 => x"05",
          6934 => x"05",
          6935 => x"67",
          6936 => x"34",
          6937 => x"1f",
          6938 => x"85",
          6939 => x"2a",
          6940 => x"34",
          6941 => x"34",
          6942 => x"61",
          6943 => x"c8",
          6944 => x"83",
          6945 => x"05",
          6946 => x"83",
          6947 => x"77",
          6948 => x"2a",
          6949 => x"81",
          6950 => x"fe",
          6951 => x"8c",
          6952 => x"52",
          6953 => x"57",
          6954 => x"84",
          6955 => x"9f",
          6956 => x"62",
          6957 => x"16",
          6958 => x"38",
          6959 => x"e7",
          6960 => x"9d",
          6961 => x"e7",
          6962 => x"22",
          6963 => x"38",
          6964 => x"78",
          6965 => x"8c",
          6966 => x"89",
          6967 => x"84",
          6968 => x"58",
          6969 => x"f5",
          6970 => x"84",
          6971 => x"f8",
          6972 => x"81",
          6973 => x"57",
          6974 => x"63",
          6975 => x"f4",
          6976 => x"75",
          6977 => x"34",
          6978 => x"05",
          6979 => x"a3",
          6980 => x"80",
          6981 => x"05",
          6982 => x"80",
          6983 => x"61",
          6984 => x"7b",
          6985 => x"59",
          6986 => x"2a",
          6987 => x"61",
          6988 => x"34",
          6989 => x"af",
          6990 => x"80",
          6991 => x"05",
          6992 => x"80",
          6993 => x"80",
          6994 => x"05",
          6995 => x"70",
          6996 => x"05",
          6997 => x"2e",
          6998 => x"58",
          6999 => x"ff",
          7000 => x"39",
          7001 => x"51",
          7002 => x"ba",
          7003 => x"29",
          7004 => x"05",
          7005 => x"53",
          7006 => x"3f",
          7007 => x"8c",
          7008 => x"0c",
          7009 => x"6a",
          7010 => x"70",
          7011 => x"ff",
          7012 => x"05",
          7013 => x"61",
          7014 => x"34",
          7015 => x"8a",
          7016 => x"f9",
          7017 => x"60",
          7018 => x"84",
          7019 => x"81",
          7020 => x"f4",
          7021 => x"81",
          7022 => x"75",
          7023 => x"75",
          7024 => x"75",
          7025 => x"34",
          7026 => x"80",
          7027 => x"e1",
          7028 => x"05",
          7029 => x"7a",
          7030 => x"05",
          7031 => x"83",
          7032 => x"7f",
          7033 => x"83",
          7034 => x"05",
          7035 => x"76",
          7036 => x"69",
          7037 => x"87",
          7038 => x"bd",
          7039 => x"60",
          7040 => x"69",
          7041 => x"3d",
          7042 => x"61",
          7043 => x"25",
          7044 => x"f8",
          7045 => x"51",
          7046 => x"09",
          7047 => x"55",
          7048 => x"70",
          7049 => x"74",
          7050 => x"cd",
          7051 => x"83",
          7052 => x"0c",
          7053 => x"7b",
          7054 => x"57",
          7055 => x"17",
          7056 => x"88",
          7057 => x"59",
          7058 => x"bb",
          7059 => x"81",
          7060 => x"04",
          7061 => x"8c",
          7062 => x"d1",
          7063 => x"72",
          7064 => x"0c",
          7065 => x"56",
          7066 => x"94",
          7067 => x"02",
          7068 => x"58",
          7069 => x"70",
          7070 => x"74",
          7071 => x"77",
          7072 => x"80",
          7073 => x"17",
          7074 => x"81",
          7075 => x"74",
          7076 => x"0c",
          7077 => x"9f",
          7078 => x"c0",
          7079 => x"c9",
          7080 => x"7c",
          7081 => x"ba",
          7082 => x"3d",
          7083 => x"05",
          7084 => x"3f",
          7085 => x"07",
          7086 => x"56",
          7087 => x"fd",
          7088 => x"ba",
          7089 => x"3d",
          7090 => x"22",
          7091 => x"26",
          7092 => x"52",
          7093 => x"0d",
          7094 => x"70",
          7095 => x"38",
          7096 => x"d0",
          7097 => x"81",
          7098 => x"54",
          7099 => x"10",
          7100 => x"51",
          7101 => x"ff",
          7102 => x"3d",
          7103 => x"05",
          7104 => x"53",
          7105 => x"8c",
          7106 => x"0c",
          7107 => x"2e",
          7108 => x"ff",
          7109 => x"d0",
          7110 => x"51",
          7111 => x"77",
          7112 => x"e1",
          7113 => x"e9",
          7114 => x"80",
          7115 => x"22",
          7116 => x"7a",
          7117 => x"b7",
          7118 => x"72",
          7119 => x"06",
          7120 => x"b1",
          7121 => x"70",
          7122 => x"30",
          7123 => x"53",
          7124 => x"75",
          7125 => x"3d",
          7126 => x"a2",
          7127 => x"10",
          7128 => x"08",
          7129 => x"ff",
          7130 => x"ff",
          7131 => x"57",
          7132 => x"ff",
          7133 => x"16",
          7134 => x"db",
          7135 => x"06",
          7136 => x"83",
          7137 => x"f0",
          7138 => x"51",
          7139 => x"06",
          7140 => x"06",
          7141 => x"73",
          7142 => x"52",
          7143 => x"ff",
          7144 => x"ff",
          7145 => x"8b",
          7146 => x"75",
          7147 => x"5f",
          7148 => x"49",
          7149 => x"33",
          7150 => x"1d",
          7151 => x"07",
          7152 => x"f1",
          7153 => x"db",
          7154 => x"c5",
          7155 => x"bf",
          7156 => x"59",
          7157 => x"59",
          7158 => x"59",
          7159 => x"59",
          7160 => x"59",
          7161 => x"59",
          7162 => x"59",
          7163 => x"59",
          7164 => x"59",
          7165 => x"59",
          7166 => x"59",
          7167 => x"59",
          7168 => x"59",
          7169 => x"59",
          7170 => x"59",
          7171 => x"59",
          7172 => x"59",
          7173 => x"59",
          7174 => x"59",
          7175 => x"59",
          7176 => x"59",
          7177 => x"59",
          7178 => x"59",
          7179 => x"59",
          7180 => x"59",
          7181 => x"59",
          7182 => x"59",
          7183 => x"59",
          7184 => x"59",
          7185 => x"11",
          7186 => x"59",
          7187 => x"b2",
          7188 => x"36",
          7189 => x"59",
          7190 => x"59",
          7191 => x"59",
          7192 => x"59",
          7193 => x"59",
          7194 => x"59",
          7195 => x"59",
          7196 => x"59",
          7197 => x"59",
          7198 => x"59",
          7199 => x"59",
          7200 => x"59",
          7201 => x"59",
          7202 => x"59",
          7203 => x"59",
          7204 => x"59",
          7205 => x"59",
          7206 => x"59",
          7207 => x"59",
          7208 => x"59",
          7209 => x"59",
          7210 => x"59",
          7211 => x"59",
          7212 => x"59",
          7213 => x"59",
          7214 => x"59",
          7215 => x"b5",
          7216 => x"59",
          7217 => x"59",
          7218 => x"59",
          7219 => x"59",
          7220 => x"6d",
          7221 => x"59",
          7222 => x"59",
          7223 => x"51",
          7224 => x"1c",
          7225 => x"40",
          7226 => x"58",
          7227 => x"91",
          7228 => x"fb",
          7229 => x"1b",
          7230 => x"95",
          7231 => x"c5",
          7232 => x"0c",
          7233 => x"d8",
          7234 => x"05",
          7235 => x"d8",
          7236 => x"0c",
          7237 => x"6e",
          7238 => x"76",
          7239 => x"b4",
          7240 => x"36",
          7241 => x"4f",
          7242 => x"5c",
          7243 => x"5c",
          7244 => x"5c",
          7245 => x"35",
          7246 => x"5c",
          7247 => x"5c",
          7248 => x"5c",
          7249 => x"5c",
          7250 => x"5c",
          7251 => x"5c",
          7252 => x"5c",
          7253 => x"5c",
          7254 => x"5c",
          7255 => x"5c",
          7256 => x"5c",
          7257 => x"62",
          7258 => x"3c",
          7259 => x"2a",
          7260 => x"7f",
          7261 => x"7f",
          7262 => x"84",
          7263 => x"8e",
          7264 => x"e3",
          7265 => x"c2",
          7266 => x"66",
          7267 => x"71",
          7268 => x"9a",
          7269 => x"56",
          7270 => x"fc",
          7271 => x"d6",
          7272 => x"83",
          7273 => x"83",
          7274 => x"83",
          7275 => x"9f",
          7276 => x"64",
          7277 => x"83",
          7278 => x"83",
          7279 => x"83",
          7280 => x"83",
          7281 => x"83",
          7282 => x"83",
          7283 => x"83",
          7284 => x"83",
          7285 => x"83",
          7286 => x"21",
          7287 => x"83",
          7288 => x"c4",
          7289 => x"75",
          7290 => x"83",
          7291 => x"83",
          7292 => x"83",
          7293 => x"a6",
          7294 => x"1b",
          7295 => x"1b",
          7296 => x"1b",
          7297 => x"1b",
          7298 => x"1b",
          7299 => x"1b",
          7300 => x"1b",
          7301 => x"1b",
          7302 => x"1b",
          7303 => x"1b",
          7304 => x"1b",
          7305 => x"1b",
          7306 => x"1b",
          7307 => x"1b",
          7308 => x"b8",
          7309 => x"ed",
          7310 => x"c8",
          7311 => x"78",
          7312 => x"1b",
          7313 => x"48",
          7314 => x"24",
          7315 => x"83",
          7316 => x"61",
          7317 => x"1b",
          7318 => x"75",
          7319 => x"d1",
          7320 => x"d1",
          7321 => x"d1",
          7322 => x"d1",
          7323 => x"d1",
          7324 => x"d1",
          7325 => x"f3",
          7326 => x"d1",
          7327 => x"d1",
          7328 => x"d1",
          7329 => x"d1",
          7330 => x"4a",
          7331 => x"61",
          7332 => x"33",
          7333 => x"1b",
          7334 => x"04",
          7335 => x"ee",
          7336 => x"d7",
          7337 => x"01",
          7338 => x"fd",
          7339 => x"fd",
          7340 => x"fd",
          7341 => x"fd",
          7342 => x"fd",
          7343 => x"fd",
          7344 => x"0d",
          7345 => x"fd",
          7346 => x"fd",
          7347 => x"fd",
          7348 => x"fd",
          7349 => x"fd",
          7350 => x"fd",
          7351 => x"fd",
          7352 => x"fd",
          7353 => x"fd",
          7354 => x"fd",
          7355 => x"fd",
          7356 => x"fd",
          7357 => x"fd",
          7358 => x"fd",
          7359 => x"fd",
          7360 => x"fd",
          7361 => x"fd",
          7362 => x"fd",
          7363 => x"fd",
          7364 => x"fd",
          7365 => x"17",
          7366 => x"fd",
          7367 => x"fd",
          7368 => x"fd",
          7369 => x"fd",
          7370 => x"fd",
          7371 => x"e1",
          7372 => x"b8",
          7373 => x"fd",
          7374 => x"fd",
          7375 => x"ff",
          7376 => x"fd",
          7377 => x"0f",
          7378 => x"fd",
          7379 => x"fd",
          7380 => x"fd",
          7381 => x"17",
          7382 => x"00",
          7383 => x"00",
          7384 => x"00",
          7385 => x"00",
          7386 => x"00",
          7387 => x"00",
          7388 => x"00",
          7389 => x"00",
          7390 => x"00",
          7391 => x"00",
          7392 => x"00",
          7393 => x"00",
          7394 => x"6c",
          7395 => x"00",
          7396 => x"00",
          7397 => x"00",
          7398 => x"00",
          7399 => x"00",
          7400 => x"00",
          7401 => x"00",
          7402 => x"00",
          7403 => x"00",
          7404 => x"6e",
          7405 => x"6f",
          7406 => x"61",
          7407 => x"69",
          7408 => x"74",
          7409 => x"20",
          7410 => x"65",
          7411 => x"2e",
          7412 => x"75",
          7413 => x"74",
          7414 => x"2e",
          7415 => x"65",
          7416 => x"6b",
          7417 => x"65",
          7418 => x"65",
          7419 => x"63",
          7420 => x"64",
          7421 => x"6d",
          7422 => x"74",
          7423 => x"63",
          7424 => x"6c",
          7425 => x"79",
          7426 => x"75",
          7427 => x"69",
          7428 => x"6b",
          7429 => x"61",
          7430 => x"00",
          7431 => x"75",
          7432 => x"20",
          7433 => x"2e",
          7434 => x"69",
          7435 => x"20",
          7436 => x"65",
          7437 => x"65",
          7438 => x"20",
          7439 => x"2e",
          7440 => x"65",
          7441 => x"79",
          7442 => x"2e",
          7443 => x"65",
          7444 => x"65",
          7445 => x"61",
          7446 => x"65",
          7447 => x"00",
          7448 => x"20",
          7449 => x"00",
          7450 => x"20",
          7451 => x"00",
          7452 => x"74",
          7453 => x"00",
          7454 => x"6c",
          7455 => x"00",
          7456 => x"72",
          7457 => x"63",
          7458 => x"00",
          7459 => x"74",
          7460 => x"74",
          7461 => x"74",
          7462 => x"0a",
          7463 => x"64",
          7464 => x"6c",
          7465 => x"00",
          7466 => x"00",
          7467 => x"00",
          7468 => x"58",
          7469 => x"20",
          7470 => x"00",
          7471 => x"25",
          7472 => x"31",
          7473 => x"00",
          7474 => x"00",
          7475 => x"65",
          7476 => x"20",
          7477 => x"2a",
          7478 => x"20",
          7479 => x"70",
          7480 => x"65",
          7481 => x"54",
          7482 => x"74",
          7483 => x"00",
          7484 => x"58",
          7485 => x"75",
          7486 => x"54",
          7487 => x"74",
          7488 => x"00",
          7489 => x"58",
          7490 => x"75",
          7491 => x"54",
          7492 => x"74",
          7493 => x"00",
          7494 => x"44",
          7495 => x"75",
          7496 => x"20",
          7497 => x"70",
          7498 => x"65",
          7499 => x"72",
          7500 => x"74",
          7501 => x"74",
          7502 => x"00",
          7503 => x"67",
          7504 => x"2e",
          7505 => x"6f",
          7506 => x"74",
          7507 => x"5f",
          7508 => x"00",
          7509 => x"74",
          7510 => x"61",
          7511 => x"20",
          7512 => x"20",
          7513 => x"69",
          7514 => x"75",
          7515 => x"00",
          7516 => x"5c",
          7517 => x"6b",
          7518 => x"6c",
          7519 => x"00",
          7520 => x"20",
          7521 => x"2e",
          7522 => x"00",
          7523 => x"5c",
          7524 => x"73",
          7525 => x"64",
          7526 => x"69",
          7527 => x"00",
          7528 => x"69",
          7529 => x"69",
          7530 => x"2e",
          7531 => x"6c",
          7532 => x"65",
          7533 => x"78",
          7534 => x"00",
          7535 => x"74",
          7536 => x"6f",
          7537 => x"2e",
          7538 => x"63",
          7539 => x"6f",
          7540 => x"38",
          7541 => x"00",
          7542 => x"30",
          7543 => x"00",
          7544 => x"30",
          7545 => x"70",
          7546 => x"2e",
          7547 => x"6c",
          7548 => x"2d",
          7549 => x"25",
          7550 => x"00",
          7551 => x"2e",
          7552 => x"6c",
          7553 => x"00",
          7554 => x"67",
          7555 => x"00",
          7556 => x"6d",
          7557 => x"6d",
          7558 => x"00",
          7559 => x"25",
          7560 => x"6f",
          7561 => x"75",
          7562 => x"61",
          7563 => x"6f",
          7564 => x"6d",
          7565 => x"00",
          7566 => x"25",
          7567 => x"3a",
          7568 => x"64",
          7569 => x"20",
          7570 => x"72",
          7571 => x"00",
          7572 => x"65",
          7573 => x"6d",
          7574 => x"00",
          7575 => x"65",
          7576 => x"20",
          7577 => x"65",
          7578 => x"72",
          7579 => x"73",
          7580 => x"0a",
          7581 => x"20",
          7582 => x"6f",
          7583 => x"74",
          7584 => x"73",
          7585 => x"0a",
          7586 => x"20",
          7587 => x"74",
          7588 => x"72",
          7589 => x"20",
          7590 => x"0a",
          7591 => x"63",
          7592 => x"20",
          7593 => x"20",
          7594 => x"20",
          7595 => x"20",
          7596 => x"0a",
          7597 => x"20",
          7598 => x"43",
          7599 => x"65",
          7600 => x"20",
          7601 => x"30",
          7602 => x"00",
          7603 => x"68",
          7604 => x"52",
          7605 => x"6b",
          7606 => x"25",
          7607 => x"48",
          7608 => x"20",
          7609 => x"6c",
          7610 => x"71",
          7611 => x"20",
          7612 => x"30",
          7613 => x"00",
          7614 => x"00",
          7615 => x"00",
          7616 => x"54",
          7617 => x"20",
          7618 => x"00",
          7619 => x"48",
          7620 => x"53",
          7621 => x"20",
          7622 => x"52",
          7623 => x"6e",
          7624 => x"64",
          7625 => x"20",
          7626 => x"20",
          7627 => x"72",
          7628 => x"64",
          7629 => x"20",
          7630 => x"20",
          7631 => x"63",
          7632 => x"64",
          7633 => x"20",
          7634 => x"20",
          7635 => x"3a",
          7636 => x"00",
          7637 => x"4d",
          7638 => x"25",
          7639 => x"58",
          7640 => x"20",
          7641 => x"41",
          7642 => x"3a",
          7643 => x"00",
          7644 => x"41",
          7645 => x"25",
          7646 => x"58",
          7647 => x"20",
          7648 => x"4d",
          7649 => x"3a",
          7650 => x"00",
          7651 => x"53",
          7652 => x"69",
          7653 => x"6e",
          7654 => x"6d",
          7655 => x"6c",
          7656 => x"69",
          7657 => x"78",
          7658 => x"00",
          7659 => x"00",
          7660 => x"b0",
          7661 => x"03",
          7662 => x"00",
          7663 => x"a8",
          7664 => x"05",
          7665 => x"00",
          7666 => x"a0",
          7667 => x"07",
          7668 => x"00",
          7669 => x"98",
          7670 => x"08",
          7671 => x"00",
          7672 => x"90",
          7673 => x"09",
          7674 => x"00",
          7675 => x"88",
          7676 => x"0d",
          7677 => x"00",
          7678 => x"80",
          7679 => x"0e",
          7680 => x"00",
          7681 => x"78",
          7682 => x"0f",
          7683 => x"00",
          7684 => x"70",
          7685 => x"11",
          7686 => x"00",
          7687 => x"68",
          7688 => x"13",
          7689 => x"00",
          7690 => x"60",
          7691 => x"15",
          7692 => x"00",
          7693 => x"00",
          7694 => x"7e",
          7695 => x"00",
          7696 => x"7e",
          7697 => x"00",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"00",
          7703 => x"6f",
          7704 => x"61",
          7705 => x"6f",
          7706 => x"2c",
          7707 => x"69",
          7708 => x"74",
          7709 => x"74",
          7710 => x"00",
          7711 => x"25",
          7712 => x"6c",
          7713 => x"65",
          7714 => x"20",
          7715 => x"20",
          7716 => x"20",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"00",
          7721 => x"00",
          7722 => x"00",
          7723 => x"00",
          7724 => x"00",
          7725 => x"00",
          7726 => x"00",
          7727 => x"00",
          7728 => x"00",
          7729 => x"00",
          7730 => x"00",
          7731 => x"00",
          7732 => x"00",
          7733 => x"00",
          7734 => x"7e",
          7735 => x"7e",
          7736 => x"64",
          7737 => x"25",
          7738 => x"3a",
          7739 => x"00",
          7740 => x"2d",
          7741 => x"64",
          7742 => x"00",
          7743 => x"64",
          7744 => x"78",
          7745 => x"25",
          7746 => x"00",
          7747 => x"43",
          7748 => x"00",
          7749 => x"20",
          7750 => x"00",
          7751 => x"20",
          7752 => x"00",
          7753 => x"20",
          7754 => x"20",
          7755 => x"44",
          7756 => x"00",
          7757 => x"74",
          7758 => x"61",
          7759 => x"20",
          7760 => x"44",
          7761 => x"00",
          7762 => x"20",
          7763 => x"2e",
          7764 => x"00",
          7765 => x"7f",
          7766 => x"3d",
          7767 => x"00",
          7768 => x"00",
          7769 => x"53",
          7770 => x"4e",
          7771 => x"46",
          7772 => x"00",
          7773 => x"20",
          7774 => x"32",
          7775 => x"a4",
          7776 => x"00",
          7777 => x"07",
          7778 => x"1c",
          7779 => x"41",
          7780 => x"49",
          7781 => x"4f",
          7782 => x"9b",
          7783 => x"55",
          7784 => x"ab",
          7785 => x"b3",
          7786 => x"bb",
          7787 => x"c3",
          7788 => x"cb",
          7789 => x"d3",
          7790 => x"db",
          7791 => x"e3",
          7792 => x"eb",
          7793 => x"f3",
          7794 => x"fb",
          7795 => x"3b",
          7796 => x"3a",
          7797 => x"00",
          7798 => x"40",
          7799 => x"00",
          7800 => x"08",
          7801 => x"00",
          7802 => x"e2",
          7803 => x"e7",
          7804 => x"ef",
          7805 => x"c5",
          7806 => x"f4",
          7807 => x"f9",
          7808 => x"a2",
          7809 => x"92",
          7810 => x"fa",
          7811 => x"ba",
          7812 => x"bd",
          7813 => x"bb",
          7814 => x"02",
          7815 => x"56",
          7816 => x"57",
          7817 => x"10",
          7818 => x"1c",
          7819 => x"5f",
          7820 => x"66",
          7821 => x"67",
          7822 => x"59",
          7823 => x"6b",
          7824 => x"88",
          7825 => x"80",
          7826 => x"c0",
          7827 => x"c4",
          7828 => x"b4",
          7829 => x"29",
          7830 => x"64",
          7831 => x"48",
          7832 => x"1a",
          7833 => x"a0",
          7834 => x"17",
          7835 => x"01",
          7836 => x"32",
          7837 => x"4a",
          7838 => x"80",
          7839 => x"82",
          7840 => x"86",
          7841 => x"8a",
          7842 => x"8e",
          7843 => x"91",
          7844 => x"96",
          7845 => x"3d",
          7846 => x"20",
          7847 => x"a2",
          7848 => x"a6",
          7849 => x"aa",
          7850 => x"ae",
          7851 => x"b2",
          7852 => x"b5",
          7853 => x"ba",
          7854 => x"be",
          7855 => x"c2",
          7856 => x"c4",
          7857 => x"ca",
          7858 => x"10",
          7859 => x"de",
          7860 => x"f1",
          7861 => x"28",
          7862 => x"09",
          7863 => x"3d",
          7864 => x"41",
          7865 => x"53",
          7866 => x"55",
          7867 => x"8f",
          7868 => x"5d",
          7869 => x"61",
          7870 => x"65",
          7871 => x"96",
          7872 => x"6d",
          7873 => x"71",
          7874 => x"9f",
          7875 => x"79",
          7876 => x"64",
          7877 => x"81",
          7878 => x"85",
          7879 => x"44",
          7880 => x"8d",
          7881 => x"91",
          7882 => x"fd",
          7883 => x"04",
          7884 => x"8a",
          7885 => x"02",
          7886 => x"08",
          7887 => x"8e",
          7888 => x"f2",
          7889 => x"f4",
          7890 => x"f7",
          7891 => x"30",
          7892 => x"60",
          7893 => x"c1",
          7894 => x"c0",
          7895 => x"26",
          7896 => x"01",
          7897 => x"a0",
          7898 => x"10",
          7899 => x"30",
          7900 => x"51",
          7901 => x"5b",
          7902 => x"5f",
          7903 => x"0e",
          7904 => x"c9",
          7905 => x"db",
          7906 => x"eb",
          7907 => x"08",
          7908 => x"08",
          7909 => x"b9",
          7910 => x"01",
          7911 => x"e0",
          7912 => x"ec",
          7913 => x"4e",
          7914 => x"10",
          7915 => x"d0",
          7916 => x"60",
          7917 => x"75",
          7918 => x"00",
          7919 => x"00",
          7920 => x"b0",
          7921 => x"00",
          7922 => x"b8",
          7923 => x"00",
          7924 => x"c0",
          7925 => x"00",
          7926 => x"c8",
          7927 => x"00",
          7928 => x"d0",
          7929 => x"00",
          7930 => x"d8",
          7931 => x"00",
          7932 => x"e0",
          7933 => x"00",
          7934 => x"e8",
          7935 => x"00",
          7936 => x"f0",
          7937 => x"00",
          7938 => x"f8",
          7939 => x"00",
          7940 => x"fc",
          7941 => x"00",
          7942 => x"00",
          7943 => x"00",
          7944 => x"04",
          7945 => x"00",
          7946 => x"08",
          7947 => x"00",
          7948 => x"0c",
          7949 => x"00",
          7950 => x"10",
          7951 => x"00",
          7952 => x"14",
          7953 => x"00",
          7954 => x"1c",
          7955 => x"00",
          7956 => x"20",
          7957 => x"00",
          7958 => x"28",
          7959 => x"00",
          7960 => x"30",
          7961 => x"00",
          7962 => x"38",
          7963 => x"00",
          7964 => x"40",
          7965 => x"00",
          7966 => x"44",
          7967 => x"00",
          7968 => x"48",
          7969 => x"00",
          7970 => x"50",
          7971 => x"00",
          7972 => x"58",
          7973 => x"00",
          7974 => x"60",
          7975 => x"00",
          7976 => x"00",
          7977 => x"ff",
          7978 => x"ff",
          7979 => x"ff",
          7980 => x"00",
          7981 => x"ff",
          7982 => x"00",
          7983 => x"00",
          7984 => x"00",
          7985 => x"00",
          7986 => x"01",
          7987 => x"00",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"00",
          7996 => x"00",
          7997 => x"00",
          7998 => x"00",
          7999 => x"00",
          8000 => x"00",
          8001 => x"00",
          8002 => x"00",
          8003 => x"fd",
          8004 => x"5b",
          8005 => x"74",
          8006 => x"6c",
          8007 => x"64",
          8008 => x"34",
          8009 => x"20",
          8010 => x"f4",
          8011 => x"f0",
          8012 => x"83",
          8013 => x"fd",
          8014 => x"5b",
          8015 => x"54",
          8016 => x"4c",
          8017 => x"44",
          8018 => x"34",
          8019 => x"20",
          8020 => x"f4",
          8021 => x"f0",
          8022 => x"83",
          8023 => x"fd",
          8024 => x"7b",
          8025 => x"54",
          8026 => x"4c",
          8027 => x"44",
          8028 => x"24",
          8029 => x"20",
          8030 => x"e1",
          8031 => x"f0",
          8032 => x"88",
          8033 => x"fa",
          8034 => x"1b",
          8035 => x"14",
          8036 => x"0c",
          8037 => x"04",
          8038 => x"f0",
          8039 => x"f0",
          8040 => x"f0",
          8041 => x"f0",
          8042 => x"83",
          8043 => x"c9",
          8044 => x"b3",
          8045 => x"31",
          8046 => x"56",
          8047 => x"48",
          8048 => x"3b",
          8049 => x"00",
          8050 => x"c1",
          8051 => x"f0",
          8052 => x"83",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"38",
          8068 => x"40",
          8069 => x"44",
          8070 => x"48",
          8071 => x"4c",
          8072 => x"50",
          8073 => x"58",
          8074 => x"60",
          8075 => x"68",
          8076 => x"70",
          8077 => x"78",
          8078 => x"80",
          8079 => x"88",
          8080 => x"90",
          8081 => x"98",
          8082 => x"a0",
          8083 => x"a8",
          8084 => x"b0",
          8085 => x"b4",
          8086 => x"bc",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"19",
          9088 => x"00",
          9089 => x"f7",
          9090 => x"ff",
          9091 => x"e2",
          9092 => x"f4",
          9093 => x"67",
          9094 => x"2d",
          9095 => x"27",
          9096 => x"49",
          9097 => x"07",
          9098 => x"0f",
          9099 => x"17",
          9100 => x"3c",
          9101 => x"87",
          9102 => x"8f",
          9103 => x"97",
          9104 => x"c0",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"00",
          9113 => x"00",
          9114 => x"00",
          9115 => x"00",
          9116 => x"00",
          9117 => x"00",
          9118 => x"00",
          9119 => x"00",
          9120 => x"01",
          9121 => x"01",
        others => X"00"
    );

    shared variable RAM5 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"88",
             5 => x"88",
             6 => x"00",
             7 => x"00",
             8 => x"06",
             9 => x"2a",
            10 => x"00",
            11 => x"00",
            12 => x"ff",
            13 => x"05",
            14 => x"ff",
            15 => x"04",
            16 => x"73",
            17 => x"73",
            18 => x"04",
            19 => x"00",
            20 => x"07",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"81",
            25 => x"0a",
            26 => x"81",
            27 => x"00",
            28 => x"07",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"00",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"51",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"05",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"06",
            49 => x"ff",
            50 => x"00",
            51 => x"00",
            52 => x"73",
            53 => x"83",
            54 => x"0c",
            55 => x"00",
            56 => x"09",
            57 => x"06",
            58 => x"00",
            59 => x"00",
            60 => x"09",
            61 => x"81",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"53",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"09",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"06",
            77 => x"10",
            78 => x"00",
            79 => x"00",
            80 => x"83",
            81 => x"05",
            82 => x"04",
            83 => x"00",
            84 => x"75",
            85 => x"50",
            86 => x"0c",
            87 => x"00",
            88 => x"75",
            89 => x"50",
            90 => x"0c",
            91 => x"00",
            92 => x"06",
            93 => x"71",
            94 => x"05",
            95 => x"00",
            96 => x"06",
            97 => x"54",
            98 => x"ff",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"05",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"53",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"0b",
           134 => x"a6",
           135 => x"0b",
           136 => x"0b",
           137 => x"e6",
           138 => x"0b",
           139 => x"0b",
           140 => x"a6",
           141 => x"0b",
           142 => x"0b",
           143 => x"e8",
           144 => x"0b",
           145 => x"0b",
           146 => x"ac",
           147 => x"0b",
           148 => x"0b",
           149 => x"f0",
           150 => x"0b",
           151 => x"0b",
           152 => x"b4",
           153 => x"0b",
           154 => x"0b",
           155 => x"f8",
           156 => x"0b",
           157 => x"0b",
           158 => x"bc",
           159 => x"0b",
           160 => x"0b",
           161 => x"80",
           162 => x"0b",
           163 => x"0b",
           164 => x"c4",
           165 => x"0b",
           166 => x"0b",
           167 => x"88",
           168 => x"0b",
           169 => x"0b",
           170 => x"cb",
           171 => x"0b",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"ba",
           193 => x"ba",
           194 => x"84",
           195 => x"ba",
           196 => x"84",
           197 => x"ba",
           198 => x"84",
           199 => x"ba",
           200 => x"84",
           201 => x"ba",
           202 => x"84",
           203 => x"ba",
           204 => x"84",
           205 => x"ba",
           206 => x"84",
           207 => x"ba",
           208 => x"84",
           209 => x"ba",
           210 => x"84",
           211 => x"ba",
           212 => x"84",
           213 => x"ba",
           214 => x"84",
           215 => x"ba",
           216 => x"84",
           217 => x"84",
           218 => x"04",
           219 => x"2d",
           220 => x"90",
           221 => x"97",
           222 => x"80",
           223 => x"d3",
           224 => x"c0",
           225 => x"82",
           226 => x"80",
           227 => x"0c",
           228 => x"08",
           229 => x"98",
           230 => x"98",
           231 => x"ba",
           232 => x"ba",
           233 => x"84",
           234 => x"84",
           235 => x"04",
           236 => x"2d",
           237 => x"90",
           238 => x"d0",
           239 => x"80",
           240 => x"f2",
           241 => x"c0",
           242 => x"82",
           243 => x"80",
           244 => x"0c",
           245 => x"08",
           246 => x"98",
           247 => x"98",
           248 => x"ba",
           249 => x"ba",
           250 => x"84",
           251 => x"84",
           252 => x"04",
           253 => x"2d",
           254 => x"90",
           255 => x"c6",
           256 => x"80",
           257 => x"95",
           258 => x"c0",
           259 => x"82",
           260 => x"80",
           261 => x"0c",
           262 => x"08",
           263 => x"98",
           264 => x"98",
           265 => x"ba",
           266 => x"ba",
           267 => x"84",
           268 => x"84",
           269 => x"04",
           270 => x"2d",
           271 => x"90",
           272 => x"b2",
           273 => x"80",
           274 => x"c7",
           275 => x"c0",
           276 => x"83",
           277 => x"80",
           278 => x"0c",
           279 => x"08",
           280 => x"98",
           281 => x"98",
           282 => x"ba",
           283 => x"ba",
           284 => x"84",
           285 => x"84",
           286 => x"04",
           287 => x"2d",
           288 => x"90",
           289 => x"99",
           290 => x"80",
           291 => x"d1",
           292 => x"c0",
           293 => x"80",
           294 => x"80",
           295 => x"0c",
           296 => x"80",
           297 => x"0c",
           298 => x"08",
           299 => x"98",
           300 => x"98",
           301 => x"ba",
           302 => x"ba",
           303 => x"84",
           304 => x"84",
           305 => x"04",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"81",
           311 => x"05",
           312 => x"72",
           313 => x"72",
           314 => x"72",
           315 => x"10",
           316 => x"53",
           317 => x"d5",
           318 => x"84",
           319 => x"ec",
           320 => x"04",
           321 => x"70",
           322 => x"52",
           323 => x"3f",
           324 => x"78",
           325 => x"81",
           326 => x"55",
           327 => x"81",
           328 => x"74",
           329 => x"9f",
           330 => x"74",
           331 => x"38",
           332 => x"8c",
           333 => x"2e",
           334 => x"70",
           335 => x"8a",
           336 => x"2a",
           337 => x"cb",
           338 => x"84",
           339 => x"80",
           340 => x"0d",
           341 => x"02",
           342 => x"fe",
           343 => x"7e",
           344 => x"3f",
           345 => x"3d",
           346 => x"88",
           347 => x"3f",
           348 => x"61",
           349 => x"8c",
           350 => x"2a",
           351 => x"ff",
           352 => x"80",
           353 => x"2e",
           354 => x"06",
           355 => x"38",
           356 => x"a3",
           357 => x"80",
           358 => x"72",
           359 => x"70",
           360 => x"80",
           361 => x"5b",
           362 => x"8c",
           363 => x"0c",
           364 => x"54",
           365 => x"70",
           366 => x"81",
           367 => x"98",
           368 => x"79",
           369 => x"53",
           370 => x"58",
           371 => x"39",
           372 => x"38",
           373 => x"7c",
           374 => x"ff",
           375 => x"af",
           376 => x"38",
           377 => x"81",
           378 => x"70",
           379 => x"e0",
           380 => x"38",
           381 => x"54",
           382 => x"59",
           383 => x"52",
           384 => x"33",
           385 => x"c7",
           386 => x"88",
           387 => x"7d",
           388 => x"54",
           389 => x"51",
           390 => x"81",
           391 => x"df",
           392 => x"38",
           393 => x"74",
           394 => x"52",
           395 => x"8c",
           396 => x"38",
           397 => x"7b",
           398 => x"8f",
           399 => x"80",
           400 => x"7a",
           401 => x"73",
           402 => x"80",
           403 => x"90",
           404 => x"29",
           405 => x"2c",
           406 => x"54",
           407 => x"98",
           408 => x"78",
           409 => x"ff",
           410 => x"2a",
           411 => x"73",
           412 => x"31",
           413 => x"80",
           414 => x"85",
           415 => x"54",
           416 => x"81",
           417 => x"85",
           418 => x"38",
           419 => x"38",
           420 => x"80",
           421 => x"80",
           422 => x"2c",
           423 => x"38",
           424 => x"77",
           425 => x"80",
           426 => x"73",
           427 => x"53",
           428 => x"81",
           429 => x"70",
           430 => x"25",
           431 => x"ef",
           432 => x"81",
           433 => x"55",
           434 => x"87",
           435 => x"80",
           436 => x"2e",
           437 => x"81",
           438 => x"e2",
           439 => x"38",
           440 => x"5e",
           441 => x"2e",
           442 => x"06",
           443 => x"77",
           444 => x"80",
           445 => x"80",
           446 => x"a0",
           447 => x"90",
           448 => x"58",
           449 => x"39",
           450 => x"57",
           451 => x"7e",
           452 => x"55",
           453 => x"05",
           454 => x"33",
           455 => x"80",
           456 => x"90",
           457 => x"5f",
           458 => x"55",
           459 => x"80",
           460 => x"90",
           461 => x"fe",
           462 => x"f7",
           463 => x"ff",
           464 => x"ff",
           465 => x"70",
           466 => x"3f",
           467 => x"ff",
           468 => x"2e",
           469 => x"81",
           470 => x"e2",
           471 => x"0a",
           472 => x"80",
           473 => x"56",
           474 => x"06",
           475 => x"fe",
           476 => x"08",
           477 => x"24",
           478 => x"06",
           479 => x"39",
           480 => x"76",
           481 => x"88",
           482 => x"76",
           483 => x"60",
           484 => x"56",
           485 => x"75",
           486 => x"08",
           487 => x"90",
           488 => x"fe",
           489 => x"33",
           490 => x"ff",
           491 => x"77",
           492 => x"81",
           493 => x"84",
           494 => x"78",
           495 => x"39",
           496 => x"5b",
           497 => x"77",
           498 => x"80",
           499 => x"80",
           500 => x"a0",
           501 => x"52",
           502 => x"2e",
           503 => x"52",
           504 => x"2a",
           505 => x"8c",
           506 => x"78",
           507 => x"7d",
           508 => x"73",
           509 => x"52",
           510 => x"06",
           511 => x"ff",
           512 => x"51",
           513 => x"7a",
           514 => x"39",
           515 => x"2c",
           516 => x"ab",
           517 => x"52",
           518 => x"39",
           519 => x"84",
           520 => x"78",
           521 => x"f3",
           522 => x"83",
           523 => x"99",
           524 => x"08",
           525 => x"3f",
           526 => x"78",
           527 => x"85",
           528 => x"70",
           529 => x"ff",
           530 => x"80",
           531 => x"33",
           532 => x"d5",
           533 => x"08",
           534 => x"80",
           535 => x"81",
           536 => x"88",
           537 => x"39",
           538 => x"f0",
           539 => x"55",
           540 => x"2e",
           541 => x"84",
           542 => x"fa",
           543 => x"0b",
           544 => x"32",
           545 => x"ff",
           546 => x"92",
           547 => x"53",
           548 => x"38",
           549 => x"88",
           550 => x"55",
           551 => x"74",
           552 => x"72",
           553 => x"e3",
           554 => x"33",
           555 => x"ff",
           556 => x"73",
           557 => x"fa",
           558 => x"70",
           559 => x"56",
           560 => x"73",
           561 => x"2e",
           562 => x"88",
           563 => x"56",
           564 => x"75",
           565 => x"8c",
           566 => x"8c",
           567 => x"76",
           568 => x"54",
           569 => x"08",
           570 => x"8c",
           571 => x"3d",
           572 => x"ff",
           573 => x"55",
           574 => x"72",
           575 => x"38",
           576 => x"80",
           577 => x"33",
           578 => x"38",
           579 => x"81",
           580 => x"06",
           581 => x"3d",
           582 => x"72",
           583 => x"05",
           584 => x"ba",
           585 => x"51",
           586 => x"ba",
           587 => x"80",
           588 => x"70",
           589 => x"08",
           590 => x"53",
           591 => x"84",
           592 => x"74",
           593 => x"ff",
           594 => x"77",
           595 => x"05",
           596 => x"12",
           597 => x"51",
           598 => x"70",
           599 => x"85",
           600 => x"79",
           601 => x"80",
           602 => x"38",
           603 => x"81",
           604 => x"55",
           605 => x"73",
           606 => x"04",
           607 => x"38",
           608 => x"ff",
           609 => x"ff",
           610 => x"ff",
           611 => x"73",
           612 => x"c7",
           613 => x"53",
           614 => x"70",
           615 => x"84",
           616 => x"04",
           617 => x"54",
           618 => x"51",
           619 => x"70",
           620 => x"85",
           621 => x"78",
           622 => x"80",
           623 => x"53",
           624 => x"ff",
           625 => x"ba",
           626 => x"3d",
           627 => x"72",
           628 => x"70",
           629 => x"71",
           630 => x"14",
           631 => x"13",
           632 => x"84",
           633 => x"72",
           634 => x"ff",
           635 => x"15",
           636 => x"de",
           637 => x"0c",
           638 => x"8c",
           639 => x"0d",
           640 => x"c1",
           641 => x"8c",
           642 => x"b3",
           643 => x"ba",
           644 => x"ba",
           645 => x"74",
           646 => x"51",
           647 => x"54",
           648 => x"0d",
           649 => x"71",
           650 => x"9f",
           651 => x"51",
           652 => x"52",
           653 => x"38",
           654 => x"70",
           655 => x"04",
           656 => x"55",
           657 => x"38",
           658 => x"ff",
           659 => x"ba",
           660 => x"3d",
           661 => x"76",
           662 => x"f5",
           663 => x"12",
           664 => x"51",
           665 => x"08",
           666 => x"80",
           667 => x"80",
           668 => x"a0",
           669 => x"54",
           670 => x"38",
           671 => x"10",
           672 => x"9f",
           673 => x"75",
           674 => x"52",
           675 => x"73",
           676 => x"8c",
           677 => x"0d",
           678 => x"30",
           679 => x"2b",
           680 => x"83",
           681 => x"25",
           682 => x"2a",
           683 => x"80",
           684 => x"71",
           685 => x"8c",
           686 => x"82",
           687 => x"2a",
           688 => x"82",
           689 => x"ba",
           690 => x"54",
           691 => x"56",
           692 => x"52",
           693 => x"75",
           694 => x"81",
           695 => x"29",
           696 => x"53",
           697 => x"78",
           698 => x"2e",
           699 => x"84",
           700 => x"73",
           701 => x"bd",
           702 => x"52",
           703 => x"38",
           704 => x"81",
           705 => x"76",
           706 => x"56",
           707 => x"74",
           708 => x"78",
           709 => x"81",
           710 => x"ff",
           711 => x"55",
           712 => x"8c",
           713 => x"0d",
           714 => x"9f",
           715 => x"32",
           716 => x"72",
           717 => x"56",
           718 => x"75",
           719 => x"88",
           720 => x"7d",
           721 => x"08",
           722 => x"2e",
           723 => x"70",
           724 => x"a0",
           725 => x"f5",
           726 => x"d0",
           727 => x"80",
           728 => x"74",
           729 => x"27",
           730 => x"06",
           731 => x"06",
           732 => x"f9",
           733 => x"89",
           734 => x"27",
           735 => x"81",
           736 => x"56",
           737 => x"78",
           738 => x"75",
           739 => x"8c",
           740 => x"16",
           741 => x"59",
           742 => x"ff",
           743 => x"33",
           744 => x"38",
           745 => x"38",
           746 => x"d0",
           747 => x"73",
           748 => x"8c",
           749 => x"81",
           750 => x"55",
           751 => x"84",
           752 => x"f7",
           753 => x"70",
           754 => x"56",
           755 => x"8f",
           756 => x"33",
           757 => x"73",
           758 => x"2e",
           759 => x"56",
           760 => x"58",
           761 => x"38",
           762 => x"14",
           763 => x"14",
           764 => x"73",
           765 => x"ff",
           766 => x"89",
           767 => x"77",
           768 => x"0c",
           769 => x"26",
           770 => x"38",
           771 => x"56",
           772 => x"0d",
           773 => x"70",
           774 => x"09",
           775 => x"70",
           776 => x"80",
           777 => x"80",
           778 => x"74",
           779 => x"56",
           780 => x"38",
           781 => x"0d",
           782 => x"0c",
           783 => x"ca",
           784 => x"8b",
           785 => x"84",
           786 => x"ba",
           787 => x"52",
           788 => x"10",
           789 => x"04",
           790 => x"83",
           791 => x"ef",
           792 => x"cf",
           793 => x"0d",
           794 => x"3f",
           795 => x"51",
           796 => x"83",
           797 => x"3d",
           798 => x"fc",
           799 => x"fc",
           800 => x"04",
           801 => x"83",
           802 => x"ee",
           803 => x"d0",
           804 => x"0d",
           805 => x"3f",
           806 => x"51",
           807 => x"83",
           808 => x"3d",
           809 => x"a4",
           810 => x"c0",
           811 => x"04",
           812 => x"83",
           813 => x"ee",
           814 => x"d1",
           815 => x"0d",
           816 => x"3f",
           817 => x"51",
           818 => x"ec",
           819 => x"e3",
           820 => x"30",
           821 => x"57",
           822 => x"83",
           823 => x"81",
           824 => x"80",
           825 => x"3d",
           826 => x"84",
           827 => x"08",
           828 => x"82",
           829 => x"07",
           830 => x"72",
           831 => x"2e",
           832 => x"55",
           833 => x"74",
           834 => x"8e",
           835 => x"d2",
           836 => x"51",
           837 => x"0c",
           838 => x"08",
           839 => x"8c",
           840 => x"84",
           841 => x"9e",
           842 => x"84",
           843 => x"55",
           844 => x"19",
           845 => x"e8",
           846 => x"ba",
           847 => x"3f",
           848 => x"bc",
           849 => x"de",
           850 => x"0d",
           851 => x"58",
           852 => x"7a",
           853 => x"08",
           854 => x"76",
           855 => x"8c",
           856 => x"84",
           857 => x"84",
           858 => x"78",
           859 => x"8c",
           860 => x"0d",
           861 => x"cf",
           862 => x"5f",
           863 => x"2e",
           864 => x"c4",
           865 => x"51",
           866 => x"27",
           867 => x"38",
           868 => x"18",
           869 => x"72",
           870 => x"d1",
           871 => x"53",
           872 => x"74",
           873 => x"dd",
           874 => x"80",
           875 => x"53",
           876 => x"81",
           877 => x"38",
           878 => x"ff",
           879 => x"38",
           880 => x"84",
           881 => x"df",
           882 => x"c2",
           883 => x"3f",
           884 => x"51",
           885 => x"98",
           886 => x"a0",
           887 => x"82",
           888 => x"26",
           889 => x"8c",
           890 => x"e0",
           891 => x"d5",
           892 => x"87",
           893 => x"fe",
           894 => x"91",
           895 => x"53",
           896 => x"79",
           897 => x"72",
           898 => x"83",
           899 => x"14",
           900 => x"51",
           901 => x"38",
           902 => x"db",
           903 => x"08",
           904 => x"73",
           905 => x"53",
           906 => x"52",
           907 => x"84",
           908 => x"a0",
           909 => x"dd",
           910 => x"08",
           911 => x"16",
           912 => x"3f",
           913 => x"53",
           914 => x"38",
           915 => x"81",
           916 => x"db",
           917 => x"ba",
           918 => x"70",
           919 => x"70",
           920 => x"06",
           921 => x"72",
           922 => x"9b",
           923 => x"2b",
           924 => x"30",
           925 => x"07",
           926 => x"59",
           927 => x"a9",
           928 => x"ba",
           929 => x"3d",
           930 => x"aa",
           931 => x"83",
           932 => x"51",
           933 => x"81",
           934 => x"72",
           935 => x"71",
           936 => x"81",
           937 => x"72",
           938 => x"71",
           939 => x"81",
           940 => x"72",
           941 => x"71",
           942 => x"81",
           943 => x"88",
           944 => x"a9",
           945 => x"51",
           946 => x"9c",
           947 => x"a9",
           948 => x"51",
           949 => x"9b",
           950 => x"72",
           951 => x"2e",
           952 => x"cd",
           953 => x"3f",
           954 => x"2a",
           955 => x"2e",
           956 => x"9b",
           957 => x"bd",
           958 => x"86",
           959 => x"80",
           960 => x"81",
           961 => x"51",
           962 => x"3f",
           963 => x"52",
           964 => x"bd",
           965 => x"d4",
           966 => x"9a",
           967 => x"06",
           968 => x"38",
           969 => x"3f",
           970 => x"80",
           971 => x"70",
           972 => x"fd",
           973 => x"9a",
           974 => x"b5",
           975 => x"82",
           976 => x"80",
           977 => x"ca",
           978 => x"61",
           979 => x"60",
           980 => x"8c",
           981 => x"59",
           982 => x"d5",
           983 => x"43",
           984 => x"7e",
           985 => x"51",
           986 => x"80",
           987 => x"79",
           988 => x"2e",
           989 => x"5e",
           990 => x"70",
           991 => x"38",
           992 => x"81",
           993 => x"5d",
           994 => x"5c",
           995 => x"29",
           996 => x"5b",
           997 => x"84",
           998 => x"08",
           999 => x"8c",
          1000 => x"7d",
          1001 => x"70",
          1002 => x"27",
          1003 => x"80",
          1004 => x"7e",
          1005 => x"08",
          1006 => x"8d",
          1007 => x"b8",
          1008 => x"3f",
          1009 => x"5c",
          1010 => x"84",
          1011 => x"84",
          1012 => x"38",
          1013 => x"82",
          1014 => x"8c",
          1015 => x"38",
          1016 => x"52",
          1017 => x"c8",
          1018 => x"67",
          1019 => x"90",
          1020 => x"3f",
          1021 => x"08",
          1022 => x"25",
          1023 => x"83",
          1024 => x"06",
          1025 => x"1b",
          1026 => x"ff",
          1027 => x"32",
          1028 => x"ff",
          1029 => x"95",
          1030 => x"d1",
          1031 => x"52",
          1032 => x"83",
          1033 => x"5b",
          1034 => x"83",
          1035 => x"82",
          1036 => x"80",
          1037 => x"ef",
          1038 => x"f8",
          1039 => x"84",
          1040 => x"84",
          1041 => x"0b",
          1042 => x"ff",
          1043 => x"81",
          1044 => x"d1",
          1045 => x"0b",
          1046 => x"d5",
          1047 => x"a7",
          1048 => x"fc",
          1049 => x"0c",
          1050 => x"26",
          1051 => x"bf",
          1052 => x"d5",
          1053 => x"5f",
          1054 => x"51",
          1055 => x"84",
          1056 => x"84",
          1057 => x"06",
          1058 => x"45",
          1059 => x"84",
          1060 => x"93",
          1061 => x"94",
          1062 => x"80",
          1063 => x"d2",
          1064 => x"e3",
          1065 => x"fa",
          1066 => x"94",
          1067 => x"3f",
          1068 => x"de",
          1069 => x"d6",
          1070 => x"3f",
          1071 => x"11",
          1072 => x"3f",
          1073 => x"b0",
          1074 => x"d0",
          1075 => x"ba",
          1076 => x"84",
          1077 => x"51",
          1078 => x"3d",
          1079 => x"51",
          1080 => x"80",
          1081 => x"d7",
          1082 => x"78",
          1083 => x"ff",
          1084 => x"ba",
          1085 => x"b8",
          1086 => x"05",
          1087 => x"08",
          1088 => x"53",
          1089 => x"f9",
          1090 => x"f8",
          1091 => x"48",
          1092 => x"98",
          1093 => x"64",
          1094 => x"b8",
          1095 => x"05",
          1096 => x"08",
          1097 => x"fe",
          1098 => x"e8",
          1099 => x"b0",
          1100 => x"52",
          1101 => x"84",
          1102 => x"7e",
          1103 => x"33",
          1104 => x"78",
          1105 => x"05",
          1106 => x"ff",
          1107 => x"e9",
          1108 => x"2e",
          1109 => x"11",
          1110 => x"3f",
          1111 => x"80",
          1112 => x"ff",
          1113 => x"ba",
          1114 => x"83",
          1115 => x"67",
          1116 => x"38",
          1117 => x"5a",
          1118 => x"79",
          1119 => x"d7",
          1120 => x"5b",
          1121 => x"d2",
          1122 => x"ff",
          1123 => x"ba",
          1124 => x"b8",
          1125 => x"05",
          1126 => x"08",
          1127 => x"fe",
          1128 => x"e8",
          1129 => x"2e",
          1130 => x"cd",
          1131 => x"82",
          1132 => x"05",
          1133 => x"46",
          1134 => x"53",
          1135 => x"84",
          1136 => x"38",
          1137 => x"80",
          1138 => x"8c",
          1139 => x"52",
          1140 => x"84",
          1141 => x"7e",
          1142 => x"33",
          1143 => x"78",
          1144 => x"05",
          1145 => x"db",
          1146 => x"49",
          1147 => x"80",
          1148 => x"8c",
          1149 => x"59",
          1150 => x"68",
          1151 => x"11",
          1152 => x"3f",
          1153 => x"f5",
          1154 => x"53",
          1155 => x"84",
          1156 => x"38",
          1157 => x"80",
          1158 => x"8c",
          1159 => x"3d",
          1160 => x"51",
          1161 => x"86",
          1162 => x"d8",
          1163 => x"5b",
          1164 => x"5b",
          1165 => x"79",
          1166 => x"e7",
          1167 => x"80",
          1168 => x"8c",
          1169 => x"59",
          1170 => x"8c",
          1171 => x"84",
          1172 => x"38",
          1173 => x"3f",
          1174 => x"11",
          1175 => x"3f",
          1176 => x"f3",
          1177 => x"c0",
          1178 => x"3d",
          1179 => x"51",
          1180 => x"91",
          1181 => x"80",
          1182 => x"08",
          1183 => x"ff",
          1184 => x"ba",
          1185 => x"66",
          1186 => x"81",
          1187 => x"72",
          1188 => x"5d",
          1189 => x"2e",
          1190 => x"51",
          1191 => x"65",
          1192 => x"3f",
          1193 => x"f2",
          1194 => x"64",
          1195 => x"11",
          1196 => x"3f",
          1197 => x"d0",
          1198 => x"84",
          1199 => x"53",
          1200 => x"84",
          1201 => x"39",
          1202 => x"7e",
          1203 => x"b8",
          1204 => x"05",
          1205 => x"08",
          1206 => x"02",
          1207 => x"05",
          1208 => x"f0",
          1209 => x"b3",
          1210 => x"38",
          1211 => x"11",
          1212 => x"3f",
          1213 => x"dc",
          1214 => x"33",
          1215 => x"9b",
          1216 => x"ff",
          1217 => x"ba",
          1218 => x"64",
          1219 => x"70",
          1220 => x"2e",
          1221 => x"55",
          1222 => x"d8",
          1223 => x"f3",
          1224 => x"80",
          1225 => x"51",
          1226 => x"3d",
          1227 => x"51",
          1228 => x"80",
          1229 => x"ce",
          1230 => x"23",
          1231 => x"91",
          1232 => x"38",
          1233 => x"39",
          1234 => x"2e",
          1235 => x"fc",
          1236 => x"cc",
          1237 => x"d8",
          1238 => x"f6",
          1239 => x"78",
          1240 => x"08",
          1241 => x"51",
          1242 => x"f3",
          1243 => x"38",
          1244 => x"39",
          1245 => x"2e",
          1246 => x"fb",
          1247 => x"7d",
          1248 => x"08",
          1249 => x"33",
          1250 => x"f2",
          1251 => x"f3",
          1252 => x"38",
          1253 => x"39",
          1254 => x"49",
          1255 => x"88",
          1256 => x"0d",
          1257 => x"c0",
          1258 => x"84",
          1259 => x"84",
          1260 => x"57",
          1261 => x"da",
          1262 => x"07",
          1263 => x"08",
          1264 => x"51",
          1265 => x"90",
          1266 => x"80",
          1267 => x"84",
          1268 => x"80",
          1269 => x"8c",
          1270 => x"0c",
          1271 => x"5d",
          1272 => x"80",
          1273 => x"70",
          1274 => x"d5",
          1275 => x"83",
          1276 => x"94",
          1277 => x"d2",
          1278 => x"fc",
          1279 => x"83",
          1280 => x"81",
          1281 => x"c3",
          1282 => x"3f",
          1283 => x"08",
          1284 => x"73",
          1285 => x"81",
          1286 => x"09",
          1287 => x"33",
          1288 => x"70",
          1289 => x"06",
          1290 => x"74",
          1291 => x"80",
          1292 => x"54",
          1293 => x"54",
          1294 => x"2e",
          1295 => x"80",
          1296 => x"a0",
          1297 => x"54",
          1298 => x"25",
          1299 => x"2e",
          1300 => x"54",
          1301 => x"84",
          1302 => x"70",
          1303 => x"ff",
          1304 => x"33",
          1305 => x"70",
          1306 => x"39",
          1307 => x"72",
          1308 => x"38",
          1309 => x"72",
          1310 => x"8c",
          1311 => x"fc",
          1312 => x"84",
          1313 => x"74",
          1314 => x"04",
          1315 => x"ff",
          1316 => x"26",
          1317 => x"05",
          1318 => x"8a",
          1319 => x"70",
          1320 => x"33",
          1321 => x"f2",
          1322 => x"74",
          1323 => x"22",
          1324 => x"80",
          1325 => x"52",
          1326 => x"81",
          1327 => x"22",
          1328 => x"33",
          1329 => x"33",
          1330 => x"33",
          1331 => x"33",
          1332 => x"33",
          1333 => x"c0",
          1334 => x"a0",
          1335 => x"0c",
          1336 => x"86",
          1337 => x"5b",
          1338 => x"0c",
          1339 => x"7b",
          1340 => x"7b",
          1341 => x"08",
          1342 => x"98",
          1343 => x"87",
          1344 => x"1c",
          1345 => x"7b",
          1346 => x"08",
          1347 => x"98",
          1348 => x"80",
          1349 => x"59",
          1350 => x"1b",
          1351 => x"1b",
          1352 => x"1b",
          1353 => x"52",
          1354 => x"3f",
          1355 => x"02",
          1356 => x"a8",
          1357 => x"84",
          1358 => x"2c",
          1359 => x"06",
          1360 => x"71",
          1361 => x"04",
          1362 => x"ba",
          1363 => x"51",
          1364 => x"df",
          1365 => x"84",
          1366 => x"2c",
          1367 => x"c7",
          1368 => x"52",
          1369 => x"e7",
          1370 => x"2b",
          1371 => x"2e",
          1372 => x"54",
          1373 => x"84",
          1374 => x"fc",
          1375 => x"f2",
          1376 => x"55",
          1377 => x"87",
          1378 => x"70",
          1379 => x"2e",
          1380 => x"06",
          1381 => x"32",
          1382 => x"38",
          1383 => x"cf",
          1384 => x"c0",
          1385 => x"38",
          1386 => x"0c",
          1387 => x"0d",
          1388 => x"51",
          1389 => x"81",
          1390 => x"71",
          1391 => x"2e",
          1392 => x"70",
          1393 => x"52",
          1394 => x"0d",
          1395 => x"9f",
          1396 => x"c4",
          1397 => x"0d",
          1398 => x"52",
          1399 => x"81",
          1400 => x"ff",
          1401 => x"80",
          1402 => x"70",
          1403 => x"52",
          1404 => x"2a",
          1405 => x"38",
          1406 => x"80",
          1407 => x"06",
          1408 => x"06",
          1409 => x"80",
          1410 => x"52",
          1411 => x"55",
          1412 => x"ba",
          1413 => x"91",
          1414 => x"98",
          1415 => x"72",
          1416 => x"81",
          1417 => x"38",
          1418 => x"2a",
          1419 => x"ce",
          1420 => x"c0",
          1421 => x"06",
          1422 => x"38",
          1423 => x"c8",
          1424 => x"f2",
          1425 => x"83",
          1426 => x"08",
          1427 => x"9c",
          1428 => x"9e",
          1429 => x"c0",
          1430 => x"87",
          1431 => x"0c",
          1432 => x"e8",
          1433 => x"f2",
          1434 => x"83",
          1435 => x"08",
          1436 => x"c4",
          1437 => x"9e",
          1438 => x"23",
          1439 => x"80",
          1440 => x"f3",
          1441 => x"83",
          1442 => x"8c",
          1443 => x"08",
          1444 => x"52",
          1445 => x"8d",
          1446 => x"08",
          1447 => x"52",
          1448 => x"71",
          1449 => x"c0",
          1450 => x"06",
          1451 => x"38",
          1452 => x"80",
          1453 => x"88",
          1454 => x"80",
          1455 => x"f3",
          1456 => x"90",
          1457 => x"52",
          1458 => x"52",
          1459 => x"87",
          1460 => x"80",
          1461 => x"83",
          1462 => x"34",
          1463 => x"70",
          1464 => x"70",
          1465 => x"83",
          1466 => x"9e",
          1467 => x"51",
          1468 => x"81",
          1469 => x"0b",
          1470 => x"80",
          1471 => x"2e",
          1472 => x"95",
          1473 => x"08",
          1474 => x"52",
          1475 => x"71",
          1476 => x"c0",
          1477 => x"51",
          1478 => x"81",
          1479 => x"c0",
          1480 => x"8a",
          1481 => x"34",
          1482 => x"70",
          1483 => x"80",
          1484 => x"f3",
          1485 => x"83",
          1486 => x"71",
          1487 => x"c0",
          1488 => x"52",
          1489 => x"52",
          1490 => x"9e",
          1491 => x"f3",
          1492 => x"52",
          1493 => x"d9",
          1494 => x"f3",
          1495 => x"83",
          1496 => x"f3",
          1497 => x"83",
          1498 => x"38",
          1499 => x"a8",
          1500 => x"84",
          1501 => x"73",
          1502 => x"56",
          1503 => x"33",
          1504 => x"99",
          1505 => x"f3",
          1506 => x"83",
          1507 => x"38",
          1508 => x"93",
          1509 => x"82",
          1510 => x"73",
          1511 => x"c2",
          1512 => x"83",
          1513 => x"83",
          1514 => x"51",
          1515 => x"08",
          1516 => x"a1",
          1517 => x"3f",
          1518 => x"c4",
          1519 => x"80",
          1520 => x"51",
          1521 => x"bd",
          1522 => x"54",
          1523 => x"ec",
          1524 => x"93",
          1525 => x"f3",
          1526 => x"51",
          1527 => x"83",
          1528 => x"52",
          1529 => x"8c",
          1530 => x"31",
          1531 => x"83",
          1532 => x"8a",
          1533 => x"04",
          1534 => x"c0",
          1535 => x"ba",
          1536 => x"71",
          1537 => x"52",
          1538 => x"3f",
          1539 => x"2e",
          1540 => x"db",
          1541 => x"b8",
          1542 => x"08",
          1543 => x"c9",
          1544 => x"d9",
          1545 => x"f2",
          1546 => x"ff",
          1547 => x"c0",
          1548 => x"83",
          1549 => x"83",
          1550 => x"52",
          1551 => x"8c",
          1552 => x"31",
          1553 => x"83",
          1554 => x"83",
          1555 => x"fe",
          1556 => x"f8",
          1557 => x"96",
          1558 => x"38",
          1559 => x"ff",
          1560 => x"56",
          1561 => x"39",
          1562 => x"3f",
          1563 => x"2e",
          1564 => x"98",
          1565 => x"8f",
          1566 => x"38",
          1567 => x"83",
          1568 => x"83",
          1569 => x"fc",
          1570 => x"33",
          1571 => x"e9",
          1572 => x"80",
          1573 => x"f3",
          1574 => x"ff",
          1575 => x"54",
          1576 => x"39",
          1577 => x"08",
          1578 => x"ff",
          1579 => x"56",
          1580 => x"39",
          1581 => x"08",
          1582 => x"ff",
          1583 => x"54",
          1584 => x"39",
          1585 => x"08",
          1586 => x"ff",
          1587 => x"55",
          1588 => x"39",
          1589 => x"08",
          1590 => x"ff",
          1591 => x"56",
          1592 => x"39",
          1593 => x"08",
          1594 => x"ff",
          1595 => x"54",
          1596 => x"39",
          1597 => x"3f",
          1598 => x"3f",
          1599 => x"2e",
          1600 => x"0d",
          1601 => x"26",
          1602 => x"c4",
          1603 => x"ac",
          1604 => x"0d",
          1605 => x"d9",
          1606 => x"bc",
          1607 => x"0d",
          1608 => x"c1",
          1609 => x"cc",
          1610 => x"0d",
          1611 => x"a9",
          1612 => x"80",
          1613 => x"84",
          1614 => x"c0",
          1615 => x"aa",
          1616 => x"81",
          1617 => x"f8",
          1618 => x"ba",
          1619 => x"57",
          1620 => x"55",
          1621 => x"df",
          1622 => x"a4",
          1623 => x"ba",
          1624 => x"0b",
          1625 => x"84",
          1626 => x"55",
          1627 => x"30",
          1628 => x"55",
          1629 => x"b0",
          1630 => x"08",
          1631 => x"ba",
          1632 => x"9a",
          1633 => x"3d",
          1634 => x"ad",
          1635 => x"06",
          1636 => x"a0",
          1637 => x"ab",
          1638 => x"76",
          1639 => x"ff",
          1640 => x"8c",
          1641 => x"0d",
          1642 => x"72",
          1643 => x"73",
          1644 => x"8d",
          1645 => x"83",
          1646 => x"ff",
          1647 => x"53",
          1648 => x"3f",
          1649 => x"14",
          1650 => x"38",
          1651 => x"70",
          1652 => x"27",
          1653 => x"8c",
          1654 => x"5a",
          1655 => x"80",
          1656 => x"8c",
          1657 => x"53",
          1658 => x"84",
          1659 => x"73",
          1660 => x"81",
          1661 => x"fe",
          1662 => x"77",
          1663 => x"38",
          1664 => x"55",
          1665 => x"d5",
          1666 => x"0b",
          1667 => x"73",
          1668 => x"f8",
          1669 => x"84",
          1670 => x"f3",
          1671 => x"51",
          1672 => x"08",
          1673 => x"bd",
          1674 => x"80",
          1675 => x"38",
          1676 => x"19",
          1677 => x"75",
          1678 => x"56",
          1679 => x"09",
          1680 => x"84",
          1681 => x"ce",
          1682 => x"08",
          1683 => x"0b",
          1684 => x"83",
          1685 => x"38",
          1686 => x"74",
          1687 => x"2e",
          1688 => x"5a",
          1689 => x"2e",
          1690 => x"5f",
          1691 => x"ba",
          1692 => x"5b",
          1693 => x"81",
          1694 => x"98",
          1695 => x"33",
          1696 => x"98",
          1697 => x"d8",
          1698 => x"53",
          1699 => x"59",
          1700 => x"38",
          1701 => x"81",
          1702 => x"70",
          1703 => x"81",
          1704 => x"2b",
          1705 => x"16",
          1706 => x"38",
          1707 => x"33",
          1708 => x"38",
          1709 => x"d1",
          1710 => x"81",
          1711 => x"70",
          1712 => x"98",
          1713 => x"05",
          1714 => x"33",
          1715 => x"57",
          1716 => x"84",
          1717 => x"57",
          1718 => x"0a",
          1719 => x"2c",
          1720 => x"76",
          1721 => x"16",
          1722 => x"83",
          1723 => x"61",
          1724 => x"08",
          1725 => x"2e",
          1726 => x"bc",
          1727 => x"80",
          1728 => x"81",
          1729 => x"fe",
          1730 => x"76",
          1731 => x"76",
          1732 => x"fd",
          1733 => x"dc",
          1734 => x"e0",
          1735 => x"d1",
          1736 => x"34",
          1737 => x"75",
          1738 => x"f0",
          1739 => x"3f",
          1740 => x"76",
          1741 => x"84",
          1742 => x"84",
          1743 => x"79",
          1744 => x"08",
          1745 => x"d0",
          1746 => x"ff",
          1747 => x"93",
          1748 => x"83",
          1749 => x"75",
          1750 => x"34",
          1751 => x"84",
          1752 => x"2e",
          1753 => x"88",
          1754 => x"f0",
          1755 => x"3f",
          1756 => x"ff",
          1757 => x"ff",
          1758 => x"7a",
          1759 => x"7b",
          1760 => x"d1",
          1761 => x"38",
          1762 => x"9e",
          1763 => x"05",
          1764 => x"f9",
          1765 => x"fb",
          1766 => x"3f",
          1767 => x"34",
          1768 => x"81",
          1769 => x"b8",
          1770 => x"d1",
          1771 => x"ff",
          1772 => x"88",
          1773 => x"f0",
          1774 => x"3f",
          1775 => x"ff",
          1776 => x"ff",
          1777 => x"74",
          1778 => x"d1",
          1779 => x"d1",
          1780 => x"27",
          1781 => x"52",
          1782 => x"34",
          1783 => x"b3",
          1784 => x"81",
          1785 => x"57",
          1786 => x"84",
          1787 => x"76",
          1788 => x"33",
          1789 => x"d1",
          1790 => x"d1",
          1791 => x"26",
          1792 => x"d1",
          1793 => x"56",
          1794 => x"15",
          1795 => x"98",
          1796 => x"06",
          1797 => x"ef",
          1798 => x"51",
          1799 => x"33",
          1800 => x"d1",
          1801 => x"77",
          1802 => x"08",
          1803 => x"74",
          1804 => x"05",
          1805 => x"5d",
          1806 => x"38",
          1807 => x"ff",
          1808 => x"29",
          1809 => x"84",
          1810 => x"75",
          1811 => x"7b",
          1812 => x"84",
          1813 => x"ff",
          1814 => x"29",
          1815 => x"84",
          1816 => x"79",
          1817 => x"81",
          1818 => x"08",
          1819 => x"3f",
          1820 => x"0a",
          1821 => x"33",
          1822 => x"a7",
          1823 => x"33",
          1824 => x"84",
          1825 => x"b0",
          1826 => x"05",
          1827 => x"81",
          1828 => x"cc",
          1829 => x"84",
          1830 => x"b0",
          1831 => x"51",
          1832 => x"81",
          1833 => x"84",
          1834 => x"80",
          1835 => x"10",
          1836 => x"57",
          1837 => x"82",
          1838 => x"05",
          1839 => x"e8",
          1840 => x"0c",
          1841 => x"83",
          1842 => x"41",
          1843 => x"08",
          1844 => x"f3",
          1845 => x"bc",
          1846 => x"80",
          1847 => x"ba",
          1848 => x"d1",
          1849 => x"38",
          1850 => x"ff",
          1851 => x"52",
          1852 => x"d5",
          1853 => x"ff",
          1854 => x"56",
          1855 => x"ff",
          1856 => x"b8",
          1857 => x"84",
          1858 => x"cc",
          1859 => x"80",
          1860 => x"33",
          1861 => x"d5",
          1862 => x"b7",
          1863 => x"51",
          1864 => x"08",
          1865 => x"84",
          1866 => x"84",
          1867 => x"55",
          1868 => x"ff",
          1869 => x"d0",
          1870 => x"7b",
          1871 => x"04",
          1872 => x"06",
          1873 => x"38",
          1874 => x"78",
          1875 => x"77",
          1876 => x"08",
          1877 => x"84",
          1878 => x"98",
          1879 => x"5b",
          1880 => x"84",
          1881 => x"ad",
          1882 => x"98",
          1883 => x"33",
          1884 => x"f3",
          1885 => x"88",
          1886 => x"80",
          1887 => x"98",
          1888 => x"55",
          1889 => x"d5",
          1890 => x"d7",
          1891 => x"80",
          1892 => x"cc",
          1893 => x"ff",
          1894 => x"57",
          1895 => x"f0",
          1896 => x"a7",
          1897 => x"80",
          1898 => x"cc",
          1899 => x"fe",
          1900 => x"33",
          1901 => x"76",
          1902 => x"81",
          1903 => x"70",
          1904 => x"57",
          1905 => x"fe",
          1906 => x"81",
          1907 => x"f2",
          1908 => x"76",
          1909 => x"70",
          1910 => x"a1",
          1911 => x"1c",
          1912 => x"ff",
          1913 => x"d0",
          1914 => x"e1",
          1915 => x"d0",
          1916 => x"5a",
          1917 => x"cc",
          1918 => x"81",
          1919 => x"75",
          1920 => x"80",
          1921 => x"98",
          1922 => x"5c",
          1923 => x"77",
          1924 => x"ff",
          1925 => x"f1",
          1926 => x"88",
          1927 => x"80",
          1928 => x"98",
          1929 => x"41",
          1930 => x"d5",
          1931 => x"8f",
          1932 => x"80",
          1933 => x"cc",
          1934 => x"ff",
          1935 => x"a4",
          1936 => x"38",
          1937 => x"ba",
          1938 => x"ba",
          1939 => x"53",
          1940 => x"3f",
          1941 => x"33",
          1942 => x"38",
          1943 => x"ff",
          1944 => x"52",
          1945 => x"d5",
          1946 => x"97",
          1947 => x"5b",
          1948 => x"ff",
          1949 => x"e1",
          1950 => x"f3",
          1951 => x"a5",
          1952 => x"ef",
          1953 => x"f0",
          1954 => x"58",
          1955 => x"0a",
          1956 => x"2c",
          1957 => x"76",
          1958 => x"33",
          1959 => x"81",
          1960 => x"7a",
          1961 => x"83",
          1962 => x"38",
          1963 => x"08",
          1964 => x"18",
          1965 => x"80",
          1966 => x"f8",
          1967 => x"38",
          1968 => x"f3",
          1969 => x"80",
          1970 => x"b4",
          1971 => x"51",
          1972 => x"ff",
          1973 => x"25",
          1974 => x"51",
          1975 => x"08",
          1976 => x"08",
          1977 => x"52",
          1978 => x"0b",
          1979 => x"33",
          1980 => x"97",
          1981 => x"51",
          1982 => x"08",
          1983 => x"84",
          1984 => x"a6",
          1985 => x"05",
          1986 => x"81",
          1987 => x"34",
          1988 => x"0b",
          1989 => x"8c",
          1990 => x"ff",
          1991 => x"84",
          1992 => x"81",
          1993 => x"7b",
          1994 => x"70",
          1995 => x"84",
          1996 => x"74",
          1997 => x"f0",
          1998 => x"3f",
          1999 => x"ff",
          2000 => x"52",
          2001 => x"d1",
          2002 => x"d1",
          2003 => x"c7",
          2004 => x"84",
          2005 => x"84",
          2006 => x"05",
          2007 => x"ab",
          2008 => x"84",
          2009 => x"58",
          2010 => x"a7",
          2011 => x"51",
          2012 => x"08",
          2013 => x"84",
          2014 => x"a4",
          2015 => x"05",
          2016 => x"81",
          2017 => x"80",
          2018 => x"70",
          2019 => x"a4",
          2020 => x"56",
          2021 => x"08",
          2022 => x"10",
          2023 => x"57",
          2024 => x"38",
          2025 => x"a8",
          2026 => x"05",
          2027 => x"79",
          2028 => x"fc",
          2029 => x"f8",
          2030 => x"51",
          2031 => x"08",
          2032 => x"83",
          2033 => x"3f",
          2034 => x"0b",
          2035 => x"8c",
          2036 => x"77",
          2037 => x"ca",
          2038 => x"a5",
          2039 => x"5c",
          2040 => x"f8",
          2041 => x"84",
          2042 => x"08",
          2043 => x"38",
          2044 => x"c1",
          2045 => x"0b",
          2046 => x"38",
          2047 => x"1b",
          2048 => x"ff",
          2049 => x"10",
          2050 => x"40",
          2051 => x"82",
          2052 => x"05",
          2053 => x"db",
          2054 => x"0c",
          2055 => x"83",
          2056 => x"41",
          2057 => x"ff",
          2058 => x"38",
          2059 => x"06",
          2060 => x"f9",
          2061 => x"51",
          2062 => x"33",
          2063 => x"57",
          2064 => x"0b",
          2065 => x"74",
          2066 => x"fc",
          2067 => x"83",
          2068 => x"52",
          2069 => x"ba",
          2070 => x"33",
          2071 => x"70",
          2072 => x"ff",
          2073 => x"f3",
          2074 => x"f3",
          2075 => x"b8",
          2076 => x"eb",
          2077 => x"02",
          2078 => x"80",
          2079 => x"26",
          2080 => x"8b",
          2081 => x"72",
          2082 => x"a0",
          2083 => x"5e",
          2084 => x"76",
          2085 => x"34",
          2086 => x"f9",
          2087 => x"98",
          2088 => x"2b",
          2089 => x"56",
          2090 => x"74",
          2091 => x"70",
          2092 => x"ee",
          2093 => x"f9",
          2094 => x"78",
          2095 => x"e0",
          2096 => x"56",
          2097 => x"90",
          2098 => x"0b",
          2099 => x"11",
          2100 => x"11",
          2101 => x"87",
          2102 => x"33",
          2103 => x"33",
          2104 => x"22",
          2105 => x"29",
          2106 => x"5d",
          2107 => x"31",
          2108 => x"7e",
          2109 => x"7a",
          2110 => x"06",
          2111 => x"57",
          2112 => x"83",
          2113 => x"70",
          2114 => x"06",
          2115 => x"78",
          2116 => x"c1",
          2117 => x"34",
          2118 => x"05",
          2119 => x"80",
          2120 => x"b8",
          2121 => x"b7",
          2122 => x"f9",
          2123 => x"5d",
          2124 => x"27",
          2125 => x"73",
          2126 => x"5a",
          2127 => x"38",
          2128 => x"0b",
          2129 => x"33",
          2130 => x"71",
          2131 => x"56",
          2132 => x"ae",
          2133 => x"38",
          2134 => x"06",
          2135 => x"33",
          2136 => x"80",
          2137 => x"87",
          2138 => x"80",
          2139 => x"ff",
          2140 => x"ba",
          2141 => x"75",
          2142 => x"58",
          2143 => x"8b",
          2144 => x"29",
          2145 => x"74",
          2146 => x"83",
          2147 => x"70",
          2148 => x"55",
          2149 => x"29",
          2150 => x"06",
          2151 => x"83",
          2152 => x"f2",
          2153 => x"fe",
          2154 => x"80",
          2155 => x"b0",
          2156 => x"80",
          2157 => x"80",
          2158 => x"34",
          2159 => x"8c",
          2160 => x"34",
          2161 => x"52",
          2162 => x"87",
          2163 => x"56",
          2164 => x"84",
          2165 => x"08",
          2166 => x"51",
          2167 => x"cc",
          2168 => x"53",
          2169 => x"08",
          2170 => x"75",
          2171 => x"34",
          2172 => x"3d",
          2173 => x"ba",
          2174 => x"af",
          2175 => x"33",
          2176 => x"81",
          2177 => x"84",
          2178 => x"83",
          2179 => x"87",
          2180 => x"22",
          2181 => x"05",
          2182 => x"92",
          2183 => x"2e",
          2184 => x"76",
          2185 => x"83",
          2186 => x"ff",
          2187 => x"55",
          2188 => x"19",
          2189 => x"f9",
          2190 => x"84",
          2191 => x"74",
          2192 => x"33",
          2193 => x"72",
          2194 => x"de",
          2195 => x"33",
          2196 => x"05",
          2197 => x"34",
          2198 => x"27",
          2199 => x"38",
          2200 => x"15",
          2201 => x"34",
          2202 => x"81",
          2203 => x"38",
          2204 => x"75",
          2205 => x"81",
          2206 => x"54",
          2207 => x"72",
          2208 => x"33",
          2209 => x"55",
          2210 => x"b0",
          2211 => x"ff",
          2212 => x"54",
          2213 => x"98",
          2214 => x"53",
          2215 => x"81",
          2216 => x"55",
          2217 => x"81",
          2218 => x"ff",
          2219 => x"5a",
          2220 => x"53",
          2221 => x"0d",
          2222 => x"f9",
          2223 => x"84",
          2224 => x"7a",
          2225 => x"fe",
          2226 => x"05",
          2227 => x"75",
          2228 => x"73",
          2229 => x"33",
          2230 => x"56",
          2231 => x"ae",
          2232 => x"de",
          2233 => x"a0",
          2234 => x"70",
          2235 => x"72",
          2236 => x"e0",
          2237 => x"05",
          2238 => x"38",
          2239 => x"80",
          2240 => x"f9",
          2241 => x"19",
          2242 => x"59",
          2243 => x"02",
          2244 => x"70",
          2245 => x"83",
          2246 => x"84",
          2247 => x"86",
          2248 => x"0b",
          2249 => x"04",
          2250 => x"f9",
          2251 => x"52",
          2252 => x"51",
          2253 => x"84",
          2254 => x"83",
          2255 => x"09",
          2256 => x"53",
          2257 => x"39",
          2258 => x"b7",
          2259 => x"70",
          2260 => x"83",
          2261 => x"8c",
          2262 => x"bd",
          2263 => x"9f",
          2264 => x"70",
          2265 => x"ba",
          2266 => x"f9",
          2267 => x"33",
          2268 => x"25",
          2269 => x"bd",
          2270 => x"86",
          2271 => x"bd",
          2272 => x"ff",
          2273 => x"25",
          2274 => x"83",
          2275 => x"3d",
          2276 => x"b1",
          2277 => x"c4",
          2278 => x"f9",
          2279 => x"84",
          2280 => x"2a",
          2281 => x"f0",
          2282 => x"f2",
          2283 => x"84",
          2284 => x"83",
          2285 => x"07",
          2286 => x"0b",
          2287 => x"04",
          2288 => x"51",
          2289 => x"83",
          2290 => x"07",
          2291 => x"39",
          2292 => x"80",
          2293 => x"0d",
          2294 => x"06",
          2295 => x"34",
          2296 => x"87",
          2297 => x"ff",
          2298 => x"fd",
          2299 => x"b8",
          2300 => x"33",
          2301 => x"83",
          2302 => x"f9",
          2303 => x"51",
          2304 => x"39",
          2305 => x"51",
          2306 => x"39",
          2307 => x"80",
          2308 => x"34",
          2309 => x"81",
          2310 => x"f9",
          2311 => x"b8",
          2312 => x"51",
          2313 => x"39",
          2314 => x"80",
          2315 => x"34",
          2316 => x"81",
          2317 => x"f9",
          2318 => x"b8",
          2319 => x"f9",
          2320 => x"b8",
          2321 => x"70",
          2322 => x"f3",
          2323 => x"84",
          2324 => x"bc",
          2325 => x"bd",
          2326 => x"5f",
          2327 => x"a1",
          2328 => x"81",
          2329 => x"82",
          2330 => x"7a",
          2331 => x"ba",
          2332 => x"3d",
          2333 => x"06",
          2334 => x"34",
          2335 => x"0b",
          2336 => x"f9",
          2337 => x"23",
          2338 => x"84",
          2339 => x"33",
          2340 => x"83",
          2341 => x"7d",
          2342 => x"b8",
          2343 => x"7b",
          2344 => x"bd",
          2345 => x"84",
          2346 => x"84",
          2347 => x"a8",
          2348 => x"83",
          2349 => x"58",
          2350 => x"8d",
          2351 => x"53",
          2352 => x"81",
          2353 => x"33",
          2354 => x"79",
          2355 => x"53",
          2356 => x"e1",
          2357 => x"84",
          2358 => x"7a",
          2359 => x"ff",
          2360 => x"34",
          2361 => x"83",
          2362 => x"23",
          2363 => x"0d",
          2364 => x"81",
          2365 => x"83",
          2366 => x"bd",
          2367 => x"83",
          2368 => x"84",
          2369 => x"51",
          2370 => x"f7",
          2371 => x"84",
          2372 => x"83",
          2373 => x"84",
          2374 => x"70",
          2375 => x"f9",
          2376 => x"05",
          2377 => x"bd",
          2378 => x"29",
          2379 => x"f9",
          2380 => x"7c",
          2381 => x"83",
          2382 => x"57",
          2383 => x"75",
          2384 => x"24",
          2385 => x"85",
          2386 => x"84",
          2387 => x"83",
          2388 => x"55",
          2389 => x"87",
          2390 => x"80",
          2391 => x"ba",
          2392 => x"56",
          2393 => x"83",
          2394 => x"58",
          2395 => x"b0",
          2396 => x"70",
          2397 => x"83",
          2398 => x"57",
          2399 => x"33",
          2400 => x"70",
          2401 => x"26",
          2402 => x"58",
          2403 => x"72",
          2404 => x"33",
          2405 => x"b8",
          2406 => x"fb",
          2407 => x"89",
          2408 => x"38",
          2409 => x"8a",
          2410 => x"81",
          2411 => x"0b",
          2412 => x"83",
          2413 => x"88",
          2414 => x"09",
          2415 => x"76",
          2416 => x"13",
          2417 => x"83",
          2418 => x"51",
          2419 => x"ff",
          2420 => x"38",
          2421 => x"34",
          2422 => x"f9",
          2423 => x"0c",
          2424 => x"2e",
          2425 => x"f9",
          2426 => x"ff",
          2427 => x"72",
          2428 => x"51",
          2429 => x"70",
          2430 => x"73",
          2431 => x"f9",
          2432 => x"83",
          2433 => x"ef",
          2434 => x"75",
          2435 => x"e6",
          2436 => x"84",
          2437 => x"2e",
          2438 => x"82",
          2439 => x"78",
          2440 => x"2e",
          2441 => x"8f",
          2442 => x"bc",
          2443 => x"29",
          2444 => x"19",
          2445 => x"84",
          2446 => x"83",
          2447 => x"5a",
          2448 => x"18",
          2449 => x"29",
          2450 => x"33",
          2451 => x"84",
          2452 => x"83",
          2453 => x"72",
          2454 => x"59",
          2455 => x"1f",
          2456 => x"42",
          2457 => x"84",
          2458 => x"38",
          2459 => x"34",
          2460 => x"3d",
          2461 => x"38",
          2462 => x"b8",
          2463 => x"2e",
          2464 => x"88",
          2465 => x"bc",
          2466 => x"29",
          2467 => x"19",
          2468 => x"84",
          2469 => x"83",
          2470 => x"41",
          2471 => x"1f",
          2472 => x"29",
          2473 => x"87",
          2474 => x"80",
          2475 => x"ba",
          2476 => x"29",
          2477 => x"f9",
          2478 => x"34",
          2479 => x"41",
          2480 => x"83",
          2481 => x"8c",
          2482 => x"2e",
          2483 => x"81",
          2484 => x"fd",
          2485 => x"34",
          2486 => x"3d",
          2487 => x"38",
          2488 => x"d0",
          2489 => x"59",
          2490 => x"84",
          2491 => x"06",
          2492 => x"34",
          2493 => x"3d",
          2494 => x"38",
          2495 => x"b8",
          2496 => x"f9",
          2497 => x"40",
          2498 => x"a3",
          2499 => x"33",
          2500 => x"22",
          2501 => x"56",
          2502 => x"f9",
          2503 => x"57",
          2504 => x"80",
          2505 => x"81",
          2506 => x"f9",
          2507 => x"42",
          2508 => x"60",
          2509 => x"58",
          2510 => x"ea",
          2511 => x"34",
          2512 => x"83",
          2513 => x"83",
          2514 => x"87",
          2515 => x"22",
          2516 => x"70",
          2517 => x"33",
          2518 => x"2e",
          2519 => x"ff",
          2520 => x"76",
          2521 => x"90",
          2522 => x"80",
          2523 => x"84",
          2524 => x"8f",
          2525 => x"80",
          2526 => x"0d",
          2527 => x"f4",
          2528 => x"f5",
          2529 => x"f6",
          2530 => x"80",
          2531 => x"0d",
          2532 => x"06",
          2533 => x"84",
          2534 => x"83",
          2535 => x"72",
          2536 => x"05",
          2537 => x"7b",
          2538 => x"83",
          2539 => x"42",
          2540 => x"38",
          2541 => x"56",
          2542 => x"f9",
          2543 => x"81",
          2544 => x"72",
          2545 => x"a8",
          2546 => x"84",
          2547 => x"83",
          2548 => x"5a",
          2549 => x"be",
          2550 => x"71",
          2551 => x"b8",
          2552 => x"84",
          2553 => x"83",
          2554 => x"72",
          2555 => x"59",
          2556 => x"de",
          2557 => x"06",
          2558 => x"38",
          2559 => x"d0",
          2560 => x"bd",
          2561 => x"ff",
          2562 => x"39",
          2563 => x"bd",
          2564 => x"95",
          2565 => x"7e",
          2566 => x"75",
          2567 => x"10",
          2568 => x"04",
          2569 => x"52",
          2570 => x"84",
          2571 => x"83",
          2572 => x"70",
          2573 => x"70",
          2574 => x"87",
          2575 => x"22",
          2576 => x"83",
          2577 => x"46",
          2578 => x"81",
          2579 => x"81",
          2580 => x"81",
          2581 => x"58",
          2582 => x"a0",
          2583 => x"83",
          2584 => x"72",
          2585 => x"a0",
          2586 => x"f9",
          2587 => x"5e",
          2588 => x"80",
          2589 => x"81",
          2590 => x"f9",
          2591 => x"44",
          2592 => x"84",
          2593 => x"70",
          2594 => x"26",
          2595 => x"58",
          2596 => x"75",
          2597 => x"81",
          2598 => x"f7",
          2599 => x"b8",
          2600 => x"81",
          2601 => x"81",
          2602 => x"5b",
          2603 => x"33",
          2604 => x"b8",
          2605 => x"f9",
          2606 => x"41",
          2607 => x"1c",
          2608 => x"29",
          2609 => x"87",
          2610 => x"80",
          2611 => x"ba",
          2612 => x"29",
          2613 => x"f9",
          2614 => x"60",
          2615 => x"58",
          2616 => x"83",
          2617 => x"0b",
          2618 => x"ba",
          2619 => x"f9",
          2620 => x"19",
          2621 => x"70",
          2622 => x"f9",
          2623 => x"34",
          2624 => x"3d",
          2625 => x"5b",
          2626 => x"83",
          2627 => x"83",
          2628 => x"5c",
          2629 => x"9c",
          2630 => x"ff",
          2631 => x"80",
          2632 => x"33",
          2633 => x"8d",
          2634 => x"02",
          2635 => x"e0",
          2636 => x"be",
          2637 => x"33",
          2638 => x"b8",
          2639 => x"5b",
          2640 => x"33",
          2641 => x"33",
          2642 => x"84",
          2643 => x"a0",
          2644 => x"83",
          2645 => x"72",
          2646 => x"78",
          2647 => x"bc",
          2648 => x"83",
          2649 => x"80",
          2650 => x"81",
          2651 => x"f9",
          2652 => x"5f",
          2653 => x"84",
          2654 => x"81",
          2655 => x"90",
          2656 => x"77",
          2657 => x"83",
          2658 => x"88",
          2659 => x"80",
          2660 => x"33",
          2661 => x"81",
          2662 => x"ba",
          2663 => x"b9",
          2664 => x"b9",
          2665 => x"b9",
          2666 => x"23",
          2667 => x"84",
          2668 => x"84",
          2669 => x"84",
          2670 => x"b9",
          2671 => x"93",
          2672 => x"86",
          2673 => x"83",
          2674 => x"f9",
          2675 => x"83",
          2676 => x"57",
          2677 => x"fe",
          2678 => x"ff",
          2679 => x"05",
          2680 => x"76",
          2681 => x"c3",
          2682 => x"b9",
          2683 => x"06",
          2684 => x"77",
          2685 => x"33",
          2686 => x"38",
          2687 => x"5f",
          2688 => x"5e",
          2689 => x"f9",
          2690 => x"71",
          2691 => x"06",
          2692 => x"f9",
          2693 => x"8d",
          2694 => x"38",
          2695 => x"81",
          2696 => x"57",
          2697 => x"75",
          2698 => x"80",
          2699 => x"bc",
          2700 => x"7b",
          2701 => x"56",
          2702 => x"39",
          2703 => x"f9",
          2704 => x"05",
          2705 => x"38",
          2706 => x"34",
          2707 => x"40",
          2708 => x"f9",
          2709 => x"71",
          2710 => x"06",
          2711 => x"f9",
          2712 => x"8d",
          2713 => x"38",
          2714 => x"2e",
          2715 => x"b8",
          2716 => x"f9",
          2717 => x"a3",
          2718 => x"43",
          2719 => x"70",
          2720 => x"08",
          2721 => x"5d",
          2722 => x"bf",
          2723 => x"fb",
          2724 => x"79",
          2725 => x"e0",
          2726 => x"06",
          2727 => x"91",
          2728 => x"33",
          2729 => x"84",
          2730 => x"5d",
          2731 => x"11",
          2732 => x"38",
          2733 => x"fb",
          2734 => x"76",
          2735 => x"e1",
          2736 => x"05",
          2737 => x"41",
          2738 => x"57",
          2739 => x"39",
          2740 => x"3f",
          2741 => x"57",
          2742 => x"10",
          2743 => x"5a",
          2744 => x"3f",
          2745 => x"b9",
          2746 => x"82",
          2747 => x"7d",
          2748 => x"22",
          2749 => x"57",
          2750 => x"d5",
          2751 => x"8d",
          2752 => x"38",
          2753 => x"81",
          2754 => x"05",
          2755 => x"33",
          2756 => x"43",
          2757 => x"27",
          2758 => x"ba",
          2759 => x"58",
          2760 => x"57",
          2761 => x"80",
          2762 => x"27",
          2763 => x"f9",
          2764 => x"8d",
          2765 => x"38",
          2766 => x"33",
          2767 => x"38",
          2768 => x"33",
          2769 => x"33",
          2770 => x"80",
          2771 => x"71",
          2772 => x"06",
          2773 => x"59",
          2774 => x"38",
          2775 => x"31",
          2776 => x"38",
          2777 => x"27",
          2778 => x"83",
          2779 => x"70",
          2780 => x"8e",
          2781 => x"76",
          2782 => x"56",
          2783 => x"ff",
          2784 => x"80",
          2785 => x"77",
          2786 => x"71",
          2787 => x"87",
          2788 => x"80",
          2789 => x"06",
          2790 => x"5c",
          2791 => x"98",
          2792 => x"5f",
          2793 => x"81",
          2794 => x"58",
          2795 => x"81",
          2796 => x"ff",
          2797 => x"5e",
          2798 => x"e0",
          2799 => x"1f",
          2800 => x"76",
          2801 => x"81",
          2802 => x"80",
          2803 => x"29",
          2804 => x"26",
          2805 => x"b9",
          2806 => x"e0",
          2807 => x"51",
          2808 => x"0b",
          2809 => x"b9",
          2810 => x"78",
          2811 => x"56",
          2812 => x"be",
          2813 => x"81",
          2814 => x"43",
          2815 => x"38",
          2816 => x"26",
          2817 => x"56",
          2818 => x"76",
          2819 => x"f5",
          2820 => x"90",
          2821 => x"11",
          2822 => x"80",
          2823 => x"75",
          2824 => x"76",
          2825 => x"70",
          2826 => x"88",
          2827 => x"52",
          2828 => x"80",
          2829 => x"76",
          2830 => x"26",
          2831 => x"b7",
          2832 => x"06",
          2833 => x"22",
          2834 => x"59",
          2835 => x"78",
          2836 => x"57",
          2837 => x"76",
          2838 => x"33",
          2839 => x"0b",
          2840 => x"81",
          2841 => x"76",
          2842 => x"e0",
          2843 => x"5a",
          2844 => x"d6",
          2845 => x"81",
          2846 => x"83",
          2847 => x"71",
          2848 => x"2a",
          2849 => x"2e",
          2850 => x"0b",
          2851 => x"81",
          2852 => x"83",
          2853 => x"88",
          2854 => x"33",
          2855 => x"22",
          2856 => x"5d",
          2857 => x"87",
          2858 => x"81",
          2859 => x"f4",
          2860 => x"fd",
          2861 => x"b8",
          2862 => x"81",
          2863 => x"f9",
          2864 => x"33",
          2865 => x"83",
          2866 => x"b8",
          2867 => x"75",
          2868 => x"80",
          2869 => x"18",
          2870 => x"a4",
          2871 => x"06",
          2872 => x"8f",
          2873 => x"06",
          2874 => x"34",
          2875 => x"81",
          2876 => x"83",
          2877 => x"f9",
          2878 => x"07",
          2879 => x"d7",
          2880 => x"06",
          2881 => x"34",
          2882 => x"81",
          2883 => x"f9",
          2884 => x"b8",
          2885 => x"75",
          2886 => x"83",
          2887 => x"07",
          2888 => x"8f",
          2889 => x"06",
          2890 => x"ff",
          2891 => x"07",
          2892 => x"ef",
          2893 => x"07",
          2894 => x"df",
          2895 => x"06",
          2896 => x"b8",
          2897 => x"33",
          2898 => x"83",
          2899 => x"0b",
          2900 => x"51",
          2901 => x"b9",
          2902 => x"b9",
          2903 => x"b9",
          2904 => x"23",
          2905 => x"c7",
          2906 => x"80",
          2907 => x"0d",
          2908 => x"f9",
          2909 => x"ff",
          2910 => x"90",
          2911 => x"05",
          2912 => x"8c",
          2913 => x"84",
          2914 => x"8c",
          2915 => x"9c",
          2916 => x"34",
          2917 => x"81",
          2918 => x"34",
          2919 => x"80",
          2920 => x"23",
          2921 => x"39",
          2922 => x"52",
          2923 => x"bd",
          2924 => x"05",
          2925 => x"f9",
          2926 => x"fb",
          2927 => x"eb",
          2928 => x"bd",
          2929 => x"2c",
          2930 => x"39",
          2931 => x"b8",
          2932 => x"eb",
          2933 => x"e3",
          2934 => x"70",
          2935 => x"40",
          2936 => x"33",
          2937 => x"11",
          2938 => x"c0",
          2939 => x"b7",
          2940 => x"5c",
          2941 => x"f9",
          2942 => x"81",
          2943 => x"74",
          2944 => x"83",
          2945 => x"29",
          2946 => x"f8",
          2947 => x"5d",
          2948 => x"83",
          2949 => x"80",
          2950 => x"ff",
          2951 => x"38",
          2952 => x"23",
          2953 => x"57",
          2954 => x"b7",
          2955 => x"ec",
          2956 => x"bc",
          2957 => x"ba",
          2958 => x"26",
          2959 => x"7e",
          2960 => x"5e",
          2961 => x"5b",
          2962 => x"06",
          2963 => x"1d",
          2964 => x"ec",
          2965 => x"e0",
          2966 => x"1e",
          2967 => x"76",
          2968 => x"81",
          2969 => x"80",
          2970 => x"29",
          2971 => x"27",
          2972 => x"5e",
          2973 => x"81",
          2974 => x"58",
          2975 => x"81",
          2976 => x"ff",
          2977 => x"5d",
          2978 => x"eb",
          2979 => x"5c",
          2980 => x"83",
          2981 => x"83",
          2982 => x"5f",
          2983 => x"eb",
          2984 => x"81",
          2985 => x"76",
          2986 => x"83",
          2987 => x"ff",
          2988 => x"38",
          2989 => x"84",
          2990 => x"ff",
          2991 => x"eb",
          2992 => x"bd",
          2993 => x"33",
          2994 => x"11",
          2995 => x"ca",
          2996 => x"81",
          2997 => x"83",
          2998 => x"83",
          2999 => x"57",
          3000 => x"b8",
          3001 => x"75",
          3002 => x"ff",
          3003 => x"fc",
          3004 => x"83",
          3005 => x"7d",
          3006 => x"38",
          3007 => x"83",
          3008 => x"59",
          3009 => x"80",
          3010 => x"f9",
          3011 => x"34",
          3012 => x"39",
          3013 => x"ba",
          3014 => x"f9",
          3015 => x"f9",
          3016 => x"83",
          3017 => x"0b",
          3018 => x"83",
          3019 => x"88",
          3020 => x"f8",
          3021 => x"0d",
          3022 => x"33",
          3023 => x"73",
          3024 => x"ba",
          3025 => x"52",
          3026 => x"84",
          3027 => x"f3",
          3028 => x"ff",
          3029 => x"ff",
          3030 => x"55",
          3031 => x"38",
          3032 => x"34",
          3033 => x"8f",
          3034 => x"54",
          3035 => x"73",
          3036 => x"09",
          3037 => x"72",
          3038 => x"54",
          3039 => x"38",
          3040 => x"70",
          3041 => x"79",
          3042 => x"80",
          3043 => x"bc",
          3044 => x"a0",
          3045 => x"59",
          3046 => x"ff",
          3047 => x"59",
          3048 => x"38",
          3049 => x"80",
          3050 => x"0c",
          3051 => x"80",
          3052 => x"08",
          3053 => x"81",
          3054 => x"81",
          3055 => x"83",
          3056 => x"06",
          3057 => x"55",
          3058 => x"81",
          3059 => x"f7",
          3060 => x"5a",
          3061 => x"75",
          3062 => x"ac",
          3063 => x"81",
          3064 => x"89",
          3065 => x"b4",
          3066 => x"58",
          3067 => x"73",
          3068 => x"32",
          3069 => x"80",
          3070 => x"f7",
          3071 => x"72",
          3072 => x"83",
          3073 => x"e5",
          3074 => x"e6",
          3075 => x"f7",
          3076 => x"5e",
          3077 => x"74",
          3078 => x"d4",
          3079 => x"82",
          3080 => x"72",
          3081 => x"d4",
          3082 => x"74",
          3083 => x"2e",
          3084 => x"53",
          3085 => x"81",
          3086 => x"84",
          3087 => x"54",
          3088 => x"f7",
          3089 => x"98",
          3090 => x"83",
          3091 => x"9c",
          3092 => x"16",
          3093 => x"76",
          3094 => x"e7",
          3095 => x"9e",
          3096 => x"38",
          3097 => x"5a",
          3098 => x"54",
          3099 => x"14",
          3100 => x"7d",
          3101 => x"83",
          3102 => x"2e",
          3103 => x"92",
          3104 => x"f8",
          3105 => x"77",
          3106 => x"17",
          3107 => x"76",
          3108 => x"83",
          3109 => x"82",
          3110 => x"38",
          3111 => x"fc",
          3112 => x"80",
          3113 => x"2e",
          3114 => x"06",
          3115 => x"ed",
          3116 => x"79",
          3117 => x"75",
          3118 => x"a1",
          3119 => x"17",
          3120 => x"fe",
          3121 => x"57",
          3122 => x"e1",
          3123 => x"05",
          3124 => x"f4",
          3125 => x"78",
          3126 => x"e0",
          3127 => x"7d",
          3128 => x"ff",
          3129 => x"ff",
          3130 => x"38",
          3131 => x"54",
          3132 => x"82",
          3133 => x"07",
          3134 => x"83",
          3135 => x"78",
          3136 => x"72",
          3137 => x"70",
          3138 => x"ba",
          3139 => x"54",
          3140 => x"b8",
          3141 => x"9a",
          3142 => x"f9",
          3143 => x"82",
          3144 => x"8c",
          3145 => x"34",
          3146 => x"81",
          3147 => x"14",
          3148 => x"d4",
          3149 => x"83",
          3150 => x"f7",
          3151 => x"ca",
          3152 => x"ff",
          3153 => x"96",
          3154 => x"81",
          3155 => x"ff",
          3156 => x"06",
          3157 => x"81",
          3158 => x"54",
          3159 => x"87",
          3160 => x"0c",
          3161 => x"39",
          3162 => x"f9",
          3163 => x"73",
          3164 => x"38",
          3165 => x"83",
          3166 => x"83",
          3167 => x"33",
          3168 => x"5e",
          3169 => x"82",
          3170 => x"7a",
          3171 => x"79",
          3172 => x"38",
          3173 => x"f0",
          3174 => x"b8",
          3175 => x"81",
          3176 => x"59",
          3177 => x"82",
          3178 => x"54",
          3179 => x"f7",
          3180 => x"08",
          3181 => x"83",
          3182 => x"b7",
          3183 => x"11",
          3184 => x"38",
          3185 => x"73",
          3186 => x"80",
          3187 => x"83",
          3188 => x"70",
          3189 => x"80",
          3190 => x"83",
          3191 => x"39",
          3192 => x"3f",
          3193 => x"fc",
          3194 => x"f7",
          3195 => x"0b",
          3196 => x"33",
          3197 => x"81",
          3198 => x"04",
          3199 => x"98",
          3200 => x"82",
          3201 => x"80",
          3202 => x"98",
          3203 => x"34",
          3204 => x"87",
          3205 => x"08",
          3206 => x"c0",
          3207 => x"9c",
          3208 => x"81",
          3209 => x"57",
          3210 => x"81",
          3211 => x"a4",
          3212 => x"80",
          3213 => x"80",
          3214 => x"80",
          3215 => x"9c",
          3216 => x"56",
          3217 => x"33",
          3218 => x"71",
          3219 => x"2e",
          3220 => x"52",
          3221 => x"72",
          3222 => x"80",
          3223 => x"53",
          3224 => x"95",
          3225 => x"3d",
          3226 => x"06",
          3227 => x"83",
          3228 => x"3f",
          3229 => x"0d",
          3230 => x"05",
          3231 => x"83",
          3232 => x"fc",
          3233 => x"07",
          3234 => x"34",
          3235 => x"34",
          3236 => x"34",
          3237 => x"08",
          3238 => x"98",
          3239 => x"0b",
          3240 => x"0b",
          3241 => x"80",
          3242 => x"83",
          3243 => x"05",
          3244 => x"87",
          3245 => x"2e",
          3246 => x"98",
          3247 => x"87",
          3248 => x"87",
          3249 => x"71",
          3250 => x"72",
          3251 => x"98",
          3252 => x"87",
          3253 => x"98",
          3254 => x"38",
          3255 => x"08",
          3256 => x"72",
          3257 => x"98",
          3258 => x"27",
          3259 => x"2e",
          3260 => x"dd",
          3261 => x"fe",
          3262 => x"06",
          3263 => x"7c",
          3264 => x"74",
          3265 => x"54",
          3266 => x"73",
          3267 => x"8c",
          3268 => x"83",
          3269 => x"3f",
          3270 => x"0d",
          3271 => x"58",
          3272 => x"ff",
          3273 => x"84",
          3274 => x"0b",
          3275 => x"87",
          3276 => x"2a",
          3277 => x"16",
          3278 => x"16",
          3279 => x"16",
          3280 => x"f4",
          3281 => x"13",
          3282 => x"97",
          3283 => x"73",
          3284 => x"26",
          3285 => x"75",
          3286 => x"56",
          3287 => x"f4",
          3288 => x"16",
          3289 => x"34",
          3290 => x"98",
          3291 => x"87",
          3292 => x"98",
          3293 => x"38",
          3294 => x"08",
          3295 => x"72",
          3296 => x"98",
          3297 => x"27",
          3298 => x"2e",
          3299 => x"08",
          3300 => x"98",
          3301 => x"08",
          3302 => x"15",
          3303 => x"53",
          3304 => x"ff",
          3305 => x"08",
          3306 => x"38",
          3307 => x"76",
          3308 => x"06",
          3309 => x"81",
          3310 => x"77",
          3311 => x"04",
          3312 => x"54",
          3313 => x"06",
          3314 => x"81",
          3315 => x"d1",
          3316 => x"89",
          3317 => x"f4",
          3318 => x"85",
          3319 => x"fe",
          3320 => x"f0",
          3321 => x"08",
          3322 => x"90",
          3323 => x"52",
          3324 => x"72",
          3325 => x"c0",
          3326 => x"27",
          3327 => x"38",
          3328 => x"53",
          3329 => x"53",
          3330 => x"c0",
          3331 => x"54",
          3332 => x"c0",
          3333 => x"f6",
          3334 => x"9c",
          3335 => x"38",
          3336 => x"c0",
          3337 => x"74",
          3338 => x"2e",
          3339 => x"72",
          3340 => x"38",
          3341 => x"06",
          3342 => x"83",
          3343 => x"82",
          3344 => x"b9",
          3345 => x"70",
          3346 => x"73",
          3347 => x"8b",
          3348 => x"70",
          3349 => x"71",
          3350 => x"53",
          3351 => x"80",
          3352 => x"82",
          3353 => x"2b",
          3354 => x"33",
          3355 => x"90",
          3356 => x"56",
          3357 => x"84",
          3358 => x"2b",
          3359 => x"88",
          3360 => x"13",
          3361 => x"87",
          3362 => x"17",
          3363 => x"88",
          3364 => x"59",
          3365 => x"85",
          3366 => x"52",
          3367 => x"87",
          3368 => x"74",
          3369 => x"84",
          3370 => x"12",
          3371 => x"80",
          3372 => x"52",
          3373 => x"89",
          3374 => x"13",
          3375 => x"07",
          3376 => x"33",
          3377 => x"58",
          3378 => x"84",
          3379 => x"b9",
          3380 => x"85",
          3381 => x"2b",
          3382 => x"86",
          3383 => x"2b",
          3384 => x"52",
          3385 => x"34",
          3386 => x"81",
          3387 => x"ff",
          3388 => x"54",
          3389 => x"34",
          3390 => x"33",
          3391 => x"83",
          3392 => x"12",
          3393 => x"2b",
          3394 => x"88",
          3395 => x"57",
          3396 => x"83",
          3397 => x"17",
          3398 => x"2b",
          3399 => x"33",
          3400 => x"81",
          3401 => x"52",
          3402 => x"73",
          3403 => x"fc",
          3404 => x"12",
          3405 => x"07",
          3406 => x"71",
          3407 => x"53",
          3408 => x"80",
          3409 => x"13",
          3410 => x"80",
          3411 => x"76",
          3412 => x"b9",
          3413 => x"12",
          3414 => x"07",
          3415 => x"33",
          3416 => x"57",
          3417 => x"72",
          3418 => x"89",
          3419 => x"84",
          3420 => x"2e",
          3421 => x"77",
          3422 => x"04",
          3423 => x"0c",
          3424 => x"82",
          3425 => x"f4",
          3426 => x"fc",
          3427 => x"81",
          3428 => x"76",
          3429 => x"34",
          3430 => x"17",
          3431 => x"b9",
          3432 => x"05",
          3433 => x"ff",
          3434 => x"56",
          3435 => x"34",
          3436 => x"10",
          3437 => x"55",
          3438 => x"83",
          3439 => x"0d",
          3440 => x"72",
          3441 => x"82",
          3442 => x"51",
          3443 => x"fc",
          3444 => x"71",
          3445 => x"58",
          3446 => x"2e",
          3447 => x"17",
          3448 => x"2b",
          3449 => x"31",
          3450 => x"27",
          3451 => x"74",
          3452 => x"38",
          3453 => x"85",
          3454 => x"5a",
          3455 => x"2e",
          3456 => x"76",
          3457 => x"12",
          3458 => x"ff",
          3459 => x"59",
          3460 => x"80",
          3461 => x"78",
          3462 => x"72",
          3463 => x"70",
          3464 => x"80",
          3465 => x"56",
          3466 => x"34",
          3467 => x"2a",
          3468 => x"83",
          3469 => x"19",
          3470 => x"2b",
          3471 => x"06",
          3472 => x"70",
          3473 => x"52",
          3474 => x"ff",
          3475 => x"b9",
          3476 => x"72",
          3477 => x"70",
          3478 => x"71",
          3479 => x"05",
          3480 => x"15",
          3481 => x"fc",
          3482 => x"11",
          3483 => x"07",
          3484 => x"70",
          3485 => x"84",
          3486 => x"33",
          3487 => x"83",
          3488 => x"5a",
          3489 => x"15",
          3490 => x"55",
          3491 => x"33",
          3492 => x"54",
          3493 => x"79",
          3494 => x"18",
          3495 => x"0c",
          3496 => x"87",
          3497 => x"2b",
          3498 => x"18",
          3499 => x"2a",
          3500 => x"84",
          3501 => x"b9",
          3502 => x"85",
          3503 => x"2b",
          3504 => x"15",
          3505 => x"2a",
          3506 => x"52",
          3507 => x"34",
          3508 => x"81",
          3509 => x"ff",
          3510 => x"54",
          3511 => x"34",
          3512 => x"51",
          3513 => x"84",
          3514 => x"2e",
          3515 => x"73",
          3516 => x"04",
          3517 => x"8c",
          3518 => x"0d",
          3519 => x"fc",
          3520 => x"23",
          3521 => x"ff",
          3522 => x"b9",
          3523 => x"0b",
          3524 => x"54",
          3525 => x"15",
          3526 => x"86",
          3527 => x"84",
          3528 => x"ff",
          3529 => x"ff",
          3530 => x"55",
          3531 => x"17",
          3532 => x"10",
          3533 => x"05",
          3534 => x"0b",
          3535 => x"2e",
          3536 => x"3d",
          3537 => x"84",
          3538 => x"61",
          3539 => x"85",
          3540 => x"38",
          3541 => x"7f",
          3542 => x"83",
          3543 => x"ff",
          3544 => x"70",
          3545 => x"7a",
          3546 => x"88",
          3547 => x"ff",
          3548 => x"05",
          3549 => x"81",
          3550 => x"90",
          3551 => x"46",
          3552 => x"59",
          3553 => x"85",
          3554 => x"33",
          3555 => x"10",
          3556 => x"98",
          3557 => x"53",
          3558 => x"c9",
          3559 => x"63",
          3560 => x"38",
          3561 => x"1b",
          3562 => x"63",
          3563 => x"38",
          3564 => x"71",
          3565 => x"11",
          3566 => x"2b",
          3567 => x"52",
          3568 => x"8c",
          3569 => x"83",
          3570 => x"2b",
          3571 => x"12",
          3572 => x"07",
          3573 => x"33",
          3574 => x"59",
          3575 => x"5c",
          3576 => x"85",
          3577 => x"17",
          3578 => x"8b",
          3579 => x"86",
          3580 => x"2b",
          3581 => x"52",
          3582 => x"34",
          3583 => x"08",
          3584 => x"88",
          3585 => x"88",
          3586 => x"34",
          3587 => x"08",
          3588 => x"33",
          3589 => x"74",
          3590 => x"88",
          3591 => x"45",
          3592 => x"34",
          3593 => x"08",
          3594 => x"71",
          3595 => x"05",
          3596 => x"88",
          3597 => x"45",
          3598 => x"1a",
          3599 => x"fc",
          3600 => x"12",
          3601 => x"62",
          3602 => x"5d",
          3603 => x"a3",
          3604 => x"05",
          3605 => x"ff",
          3606 => x"81",
          3607 => x"8c",
          3608 => x"f4",
          3609 => x"0b",
          3610 => x"53",
          3611 => x"c7",
          3612 => x"60",
          3613 => x"84",
          3614 => x"34",
          3615 => x"fc",
          3616 => x"0b",
          3617 => x"84",
          3618 => x"80",
          3619 => x"88",
          3620 => x"18",
          3621 => x"f8",
          3622 => x"fc",
          3623 => x"82",
          3624 => x"84",
          3625 => x"38",
          3626 => x"54",
          3627 => x"51",
          3628 => x"84",
          3629 => x"61",
          3630 => x"2b",
          3631 => x"33",
          3632 => x"81",
          3633 => x"44",
          3634 => x"81",
          3635 => x"05",
          3636 => x"19",
          3637 => x"fc",
          3638 => x"33",
          3639 => x"8f",
          3640 => x"ff",
          3641 => x"47",
          3642 => x"05",
          3643 => x"63",
          3644 => x"1e",
          3645 => x"34",
          3646 => x"05",
          3647 => x"bc",
          3648 => x"ff",
          3649 => x"81",
          3650 => x"ff",
          3651 => x"33",
          3652 => x"10",
          3653 => x"98",
          3654 => x"53",
          3655 => x"25",
          3656 => x"78",
          3657 => x"8b",
          3658 => x"5b",
          3659 => x"8f",
          3660 => x"fc",
          3661 => x"23",
          3662 => x"ff",
          3663 => x"b9",
          3664 => x"0b",
          3665 => x"59",
          3666 => x"1a",
          3667 => x"86",
          3668 => x"84",
          3669 => x"ff",
          3670 => x"ff",
          3671 => x"57",
          3672 => x"64",
          3673 => x"70",
          3674 => x"05",
          3675 => x"05",
          3676 => x"ee",
          3677 => x"61",
          3678 => x"27",
          3679 => x"80",
          3680 => x"fb",
          3681 => x"0c",
          3682 => x"11",
          3683 => x"71",
          3684 => x"33",
          3685 => x"83",
          3686 => x"85",
          3687 => x"88",
          3688 => x"58",
          3689 => x"05",
          3690 => x"b9",
          3691 => x"85",
          3692 => x"2b",
          3693 => x"15",
          3694 => x"2a",
          3695 => x"41",
          3696 => x"87",
          3697 => x"70",
          3698 => x"07",
          3699 => x"5f",
          3700 => x"81",
          3701 => x"1f",
          3702 => x"8b",
          3703 => x"73",
          3704 => x"07",
          3705 => x"43",
          3706 => x"81",
          3707 => x"1f",
          3708 => x"2b",
          3709 => x"14",
          3710 => x"07",
          3711 => x"40",
          3712 => x"60",
          3713 => x"70",
          3714 => x"71",
          3715 => x"70",
          3716 => x"05",
          3717 => x"84",
          3718 => x"83",
          3719 => x"39",
          3720 => x"0c",
          3721 => x"82",
          3722 => x"f4",
          3723 => x"fc",
          3724 => x"81",
          3725 => x"7f",
          3726 => x"34",
          3727 => x"15",
          3728 => x"b9",
          3729 => x"05",
          3730 => x"ff",
          3731 => x"5e",
          3732 => x"34",
          3733 => x"10",
          3734 => x"5c",
          3735 => x"83",
          3736 => x"7f",
          3737 => x"87",
          3738 => x"2b",
          3739 => x"1d",
          3740 => x"2a",
          3741 => x"61",
          3742 => x"34",
          3743 => x"11",
          3744 => x"71",
          3745 => x"33",
          3746 => x"70",
          3747 => x"56",
          3748 => x"78",
          3749 => x"08",
          3750 => x"88",
          3751 => x"88",
          3752 => x"34",
          3753 => x"08",
          3754 => x"71",
          3755 => x"05",
          3756 => x"2b",
          3757 => x"06",
          3758 => x"5d",
          3759 => x"82",
          3760 => x"b9",
          3761 => x"12",
          3762 => x"07",
          3763 => x"71",
          3764 => x"70",
          3765 => x"5a",
          3766 => x"81",
          3767 => x"5b",
          3768 => x"16",
          3769 => x"07",
          3770 => x"33",
          3771 => x"5e",
          3772 => x"1e",
          3773 => x"fc",
          3774 => x"12",
          3775 => x"07",
          3776 => x"33",
          3777 => x"44",
          3778 => x"7c",
          3779 => x"05",
          3780 => x"33",
          3781 => x"81",
          3782 => x"5b",
          3783 => x"16",
          3784 => x"70",
          3785 => x"71",
          3786 => x"81",
          3787 => x"83",
          3788 => x"63",
          3789 => x"59",
          3790 => x"7b",
          3791 => x"70",
          3792 => x"8b",
          3793 => x"70",
          3794 => x"07",
          3795 => x"5d",
          3796 => x"75",
          3797 => x"b9",
          3798 => x"83",
          3799 => x"2b",
          3800 => x"12",
          3801 => x"07",
          3802 => x"33",
          3803 => x"59",
          3804 => x"5d",
          3805 => x"79",
          3806 => x"70",
          3807 => x"71",
          3808 => x"05",
          3809 => x"88",
          3810 => x"5e",
          3811 => x"16",
          3812 => x"fc",
          3813 => x"71",
          3814 => x"70",
          3815 => x"79",
          3816 => x"fc",
          3817 => x"12",
          3818 => x"07",
          3819 => x"71",
          3820 => x"5c",
          3821 => x"79",
          3822 => x"fc",
          3823 => x"33",
          3824 => x"74",
          3825 => x"71",
          3826 => x"5c",
          3827 => x"82",
          3828 => x"b9",
          3829 => x"83",
          3830 => x"57",
          3831 => x"5a",
          3832 => x"b5",
          3833 => x"84",
          3834 => x"ff",
          3835 => x"39",
          3836 => x"8b",
          3837 => x"84",
          3838 => x"2b",
          3839 => x"43",
          3840 => x"63",
          3841 => x"08",
          3842 => x"33",
          3843 => x"74",
          3844 => x"71",
          3845 => x"41",
          3846 => x"64",
          3847 => x"34",
          3848 => x"81",
          3849 => x"ff",
          3850 => x"42",
          3851 => x"34",
          3852 => x"33",
          3853 => x"83",
          3854 => x"12",
          3855 => x"2b",
          3856 => x"88",
          3857 => x"45",
          3858 => x"83",
          3859 => x"1f",
          3860 => x"2b",
          3861 => x"33",
          3862 => x"81",
          3863 => x"5f",
          3864 => x"7d",
          3865 => x"ff",
          3866 => x"60",
          3867 => x"8c",
          3868 => x"2e",
          3869 => x"ba",
          3870 => x"73",
          3871 => x"7b",
          3872 => x"f9",
          3873 => x"fc",
          3874 => x"38",
          3875 => x"ba",
          3876 => x"51",
          3877 => x"54",
          3878 => x"38",
          3879 => x"08",
          3880 => x"ba",
          3881 => x"ff",
          3882 => x"80",
          3883 => x"80",
          3884 => x"fe",
          3885 => x"55",
          3886 => x"34",
          3887 => x"15",
          3888 => x"b9",
          3889 => x"81",
          3890 => x"08",
          3891 => x"80",
          3892 => x"70",
          3893 => x"88",
          3894 => x"b9",
          3895 => x"b9",
          3896 => x"76",
          3897 => x"34",
          3898 => x"38",
          3899 => x"8f",
          3900 => x"26",
          3901 => x"52",
          3902 => x"0d",
          3903 => x"33",
          3904 => x"38",
          3905 => x"8c",
          3906 => x"38",
          3907 => x"ba",
          3908 => x"8c",
          3909 => x"0d",
          3910 => x"05",
          3911 => x"76",
          3912 => x"17",
          3913 => x"55",
          3914 => x"87",
          3915 => x"52",
          3916 => x"8c",
          3917 => x"2e",
          3918 => x"54",
          3919 => x"38",
          3920 => x"80",
          3921 => x"74",
          3922 => x"04",
          3923 => x"ff",
          3924 => x"ff",
          3925 => x"7c",
          3926 => x"33",
          3927 => x"74",
          3928 => x"33",
          3929 => x"73",
          3930 => x"c0",
          3931 => x"76",
          3932 => x"08",
          3933 => x"a7",
          3934 => x"73",
          3935 => x"74",
          3936 => x"2e",
          3937 => x"84",
          3938 => x"84",
          3939 => x"06",
          3940 => x"ac",
          3941 => x"02",
          3942 => x"05",
          3943 => x"53",
          3944 => x"88",
          3945 => x"83",
          3946 => x"c0",
          3947 => x"2e",
          3948 => x"70",
          3949 => x"84",
          3950 => x"88",
          3951 => x"8c",
          3952 => x"75",
          3953 => x"86",
          3954 => x"c0",
          3955 => x"38",
          3956 => x"51",
          3957 => x"c0",
          3958 => x"87",
          3959 => x"38",
          3960 => x"14",
          3961 => x"80",
          3962 => x"06",
          3963 => x"f6",
          3964 => x"19",
          3965 => x"2e",
          3966 => x"56",
          3967 => x"53",
          3968 => x"a3",
          3969 => x"83",
          3970 => x"0c",
          3971 => x"18",
          3972 => x"19",
          3973 => x"59",
          3974 => x"81",
          3975 => x"83",
          3976 => x"1a",
          3977 => x"8c",
          3978 => x"27",
          3979 => x"74",
          3980 => x"38",
          3981 => x"81",
          3982 => x"78",
          3983 => x"81",
          3984 => x"57",
          3985 => x"ee",
          3986 => x"56",
          3987 => x"34",
          3988 => x"d5",
          3989 => x"0b",
          3990 => x"34",
          3991 => x"e1",
          3992 => x"bb",
          3993 => x"19",
          3994 => x"34",
          3995 => x"80",
          3996 => x"18",
          3997 => x"74",
          3998 => x"34",
          3999 => x"19",
          4000 => x"a3",
          4001 => x"84",
          4002 => x"74",
          4003 => x"56",
          4004 => x"2a",
          4005 => x"18",
          4006 => x"5b",
          4007 => x"18",
          4008 => x"19",
          4009 => x"33",
          4010 => x"08",
          4011 => x"39",
          4012 => x"59",
          4013 => x"9c",
          4014 => x"58",
          4015 => x"0d",
          4016 => x"82",
          4017 => x"82",
          4018 => x"06",
          4019 => x"89",
          4020 => x"80",
          4021 => x"38",
          4022 => x"09",
          4023 => x"78",
          4024 => x"51",
          4025 => x"80",
          4026 => x"78",
          4027 => x"79",
          4028 => x"81",
          4029 => x"05",
          4030 => x"79",
          4031 => x"33",
          4032 => x"09",
          4033 => x"78",
          4034 => x"51",
          4035 => x"80",
          4036 => x"78",
          4037 => x"7a",
          4038 => x"70",
          4039 => x"71",
          4040 => x"79",
          4041 => x"84",
          4042 => x"75",
          4043 => x"b4",
          4044 => x"0b",
          4045 => x"7b",
          4046 => x"38",
          4047 => x"81",
          4048 => x"ba",
          4049 => x"59",
          4050 => x"fd",
          4051 => x"77",
          4052 => x"33",
          4053 => x"0c",
          4054 => x"83",
          4055 => x"75",
          4056 => x"b4",
          4057 => x"0b",
          4058 => x"7c",
          4059 => x"38",
          4060 => x"81",
          4061 => x"ba",
          4062 => x"59",
          4063 => x"fc",
          4064 => x"06",
          4065 => x"82",
          4066 => x"2b",
          4067 => x"88",
          4068 => x"fe",
          4069 => x"41",
          4070 => x"0d",
          4071 => x"b8",
          4072 => x"5c",
          4073 => x"8c",
          4074 => x"be",
          4075 => x"34",
          4076 => x"84",
          4077 => x"18",
          4078 => x"33",
          4079 => x"fd",
          4080 => x"a0",
          4081 => x"17",
          4082 => x"fd",
          4083 => x"53",
          4084 => x"52",
          4085 => x"08",
          4086 => x"38",
          4087 => x"b4",
          4088 => x"7c",
          4089 => x"17",
          4090 => x"38",
          4091 => x"39",
          4092 => x"17",
          4093 => x"f5",
          4094 => x"08",
          4095 => x"38",
          4096 => x"b4",
          4097 => x"ba",
          4098 => x"08",
          4099 => x"55",
          4100 => x"b8",
          4101 => x"18",
          4102 => x"33",
          4103 => x"a0",
          4104 => x"b8",
          4105 => x"5e",
          4106 => x"8c",
          4107 => x"cb",
          4108 => x"34",
          4109 => x"84",
          4110 => x"18",
          4111 => x"33",
          4112 => x"fb",
          4113 => x"a0",
          4114 => x"17",
          4115 => x"fa",
          4116 => x"a0",
          4117 => x"17",
          4118 => x"39",
          4119 => x"9f",
          4120 => x"5d",
          4121 => x"9c",
          4122 => x"38",
          4123 => x"38",
          4124 => x"81",
          4125 => x"8c",
          4126 => x"2a",
          4127 => x"b4",
          4128 => x"86",
          4129 => x"5d",
          4130 => x"fa",
          4131 => x"52",
          4132 => x"84",
          4133 => x"ff",
          4134 => x"79",
          4135 => x"83",
          4136 => x"ff",
          4137 => x"76",
          4138 => x"81",
          4139 => x"8c",
          4140 => x"2e",
          4141 => x"87",
          4142 => x"0b",
          4143 => x"2e",
          4144 => x"5b",
          4145 => x"84",
          4146 => x"19",
          4147 => x"3f",
          4148 => x"38",
          4149 => x"0c",
          4150 => x"82",
          4151 => x"11",
          4152 => x"0a",
          4153 => x"57",
          4154 => x"2a",
          4155 => x"2a",
          4156 => x"2a",
          4157 => x"83",
          4158 => x"2a",
          4159 => x"05",
          4160 => x"78",
          4161 => x"33",
          4162 => x"09",
          4163 => x"77",
          4164 => x"51",
          4165 => x"80",
          4166 => x"77",
          4167 => x"ac",
          4168 => x"05",
          4169 => x"57",
          4170 => x"7a",
          4171 => x"8f",
          4172 => x"34",
          4173 => x"2a",
          4174 => x"b4",
          4175 => x"83",
          4176 => x"19",
          4177 => x"f0",
          4178 => x"08",
          4179 => x"38",
          4180 => x"b4",
          4181 => x"a0",
          4182 => x"5c",
          4183 => x"82",
          4184 => x"e4",
          4185 => x"81",
          4186 => x"ba",
          4187 => x"56",
          4188 => x"fc",
          4189 => x"b8",
          4190 => x"8f",
          4191 => x"f0",
          4192 => x"74",
          4193 => x"fc",
          4194 => x"19",
          4195 => x"ef",
          4196 => x"08",
          4197 => x"38",
          4198 => x"b4",
          4199 => x"a0",
          4200 => x"59",
          4201 => x"38",
          4202 => x"09",
          4203 => x"76",
          4204 => x"51",
          4205 => x"39",
          4206 => x"53",
          4207 => x"3f",
          4208 => x"2e",
          4209 => x"ba",
          4210 => x"08",
          4211 => x"08",
          4212 => x"5f",
          4213 => x"19",
          4214 => x"06",
          4215 => x"53",
          4216 => x"e4",
          4217 => x"54",
          4218 => x"1a",
          4219 => x"5a",
          4220 => x"81",
          4221 => x"08",
          4222 => x"a8",
          4223 => x"ba",
          4224 => x"7d",
          4225 => x"55",
          4226 => x"fa",
          4227 => x"52",
          4228 => x"7b",
          4229 => x"1c",
          4230 => x"ec",
          4231 => x"7b",
          4232 => x"7c",
          4233 => x"76",
          4234 => x"79",
          4235 => x"58",
          4236 => x"83",
          4237 => x"11",
          4238 => x"7f",
          4239 => x"5d",
          4240 => x"56",
          4241 => x"5a",
          4242 => x"5b",
          4243 => x"f6",
          4244 => x"5c",
          4245 => x"08",
          4246 => x"76",
          4247 => x"94",
          4248 => x"2e",
          4249 => x"93",
          4250 => x"19",
          4251 => x"75",
          4252 => x"79",
          4253 => x"08",
          4254 => x"84",
          4255 => x"84",
          4256 => x"72",
          4257 => x"51",
          4258 => x"77",
          4259 => x"73",
          4260 => x"3d",
          4261 => x"84",
          4262 => x"52",
          4263 => x"74",
          4264 => x"84",
          4265 => x"08",
          4266 => x"84",
          4267 => x"57",
          4268 => x"19",
          4269 => x"75",
          4270 => x"58",
          4271 => x"a0",
          4272 => x"30",
          4273 => x"07",
          4274 => x"55",
          4275 => x"8c",
          4276 => x"08",
          4277 => x"73",
          4278 => x"73",
          4279 => x"80",
          4280 => x"52",
          4281 => x"8c",
          4282 => x"84",
          4283 => x"58",
          4284 => x"e3",
          4285 => x"08",
          4286 => x"74",
          4287 => x"1a",
          4288 => x"79",
          4289 => x"ba",
          4290 => x"0b",
          4291 => x"04",
          4292 => x"39",
          4293 => x"53",
          4294 => x"84",
          4295 => x"84",
          4296 => x"8c",
          4297 => x"2e",
          4298 => x"39",
          4299 => x"59",
          4300 => x"80",
          4301 => x"80",
          4302 => x"18",
          4303 => x"33",
          4304 => x"73",
          4305 => x"22",
          4306 => x"ac",
          4307 => x"19",
          4308 => x"72",
          4309 => x"13",
          4310 => x"17",
          4311 => x"75",
          4312 => x"04",
          4313 => x"3d",
          4314 => x"80",
          4315 => x"70",
          4316 => x"a5",
          4317 => x"fe",
          4318 => x"27",
          4319 => x"29",
          4320 => x"98",
          4321 => x"77",
          4322 => x"08",
          4323 => x"a4",
          4324 => x"27",
          4325 => x"84",
          4326 => x"38",
          4327 => x"cd",
          4328 => x"ba",
          4329 => x"3d",
          4330 => x"a0",
          4331 => x"7a",
          4332 => x"0c",
          4333 => x"80",
          4334 => x"5b",
          4335 => x"08",
          4336 => x"2a",
          4337 => x"27",
          4338 => x"79",
          4339 => x"9c",
          4340 => x"8c",
          4341 => x"18",
          4342 => x"89",
          4343 => x"52",
          4344 => x"8c",
          4345 => x"ba",
          4346 => x"84",
          4347 => x"9c",
          4348 => x"82",
          4349 => x"38",
          4350 => x"a7",
          4351 => x"56",
          4352 => x"9c",
          4353 => x"81",
          4354 => x"ba",
          4355 => x"84",
          4356 => x"58",
          4357 => x"1a",
          4358 => x"75",
          4359 => x"76",
          4360 => x"5e",
          4361 => x"84",
          4362 => x"81",
          4363 => x"f4",
          4364 => x"75",
          4365 => x"75",
          4366 => x"51",
          4367 => x"80",
          4368 => x"7a",
          4369 => x"8c",
          4370 => x"b4",
          4371 => x"81",
          4372 => x"84",
          4373 => x"ba",
          4374 => x"08",
          4375 => x"1a",
          4376 => x"33",
          4377 => x"fe",
          4378 => x"a0",
          4379 => x"19",
          4380 => x"39",
          4381 => x"ff",
          4382 => x"06",
          4383 => x"1d",
          4384 => x"80",
          4385 => x"8a",
          4386 => x"08",
          4387 => x"39",
          4388 => x"3d",
          4389 => x"41",
          4390 => x"ff",
          4391 => x"75",
          4392 => x"5f",
          4393 => x"76",
          4394 => x"78",
          4395 => x"06",
          4396 => x"b8",
          4397 => x"bd",
          4398 => x"85",
          4399 => x"1a",
          4400 => x"9c",
          4401 => x"80",
          4402 => x"bf",
          4403 => x"60",
          4404 => x"70",
          4405 => x"80",
          4406 => x"45",
          4407 => x"df",
          4408 => x"bf",
          4409 => x"81",
          4410 => x"f6",
          4411 => x"ba",
          4412 => x"08",
          4413 => x"ba",
          4414 => x"54",
          4415 => x"19",
          4416 => x"84",
          4417 => x"06",
          4418 => x"83",
          4419 => x"08",
          4420 => x"7a",
          4421 => x"82",
          4422 => x"81",
          4423 => x"19",
          4424 => x"52",
          4425 => x"77",
          4426 => x"09",
          4427 => x"2a",
          4428 => x"38",
          4429 => x"70",
          4430 => x"59",
          4431 => x"81",
          4432 => x"81",
          4433 => x"fe",
          4434 => x"0b",
          4435 => x"0c",
          4436 => x"df",
          4437 => x"2e",
          4438 => x"08",
          4439 => x"88",
          4440 => x"b7",
          4441 => x"8d",
          4442 => x"58",
          4443 => x"05",
          4444 => x"2b",
          4445 => x"80",
          4446 => x"87",
          4447 => x"42",
          4448 => x"17",
          4449 => x"33",
          4450 => x"77",
          4451 => x"26",
          4452 => x"43",
          4453 => x"ff",
          4454 => x"83",
          4455 => x"55",
          4456 => x"55",
          4457 => x"80",
          4458 => x"33",
          4459 => x"ff",
          4460 => x"74",
          4461 => x"ac",
          4462 => x"94",
          4463 => x"70",
          4464 => x"f5",
          4465 => x"84",
          4466 => x"ff",
          4467 => x"0c",
          4468 => x"80",
          4469 => x"cc",
          4470 => x"74",
          4471 => x"38",
          4472 => x"81",
          4473 => x"ba",
          4474 => x"56",
          4475 => x"5a",
          4476 => x"70",
          4477 => x"99",
          4478 => x"81",
          4479 => x"34",
          4480 => x"75",
          4481 => x"2e",
          4482 => x"75",
          4483 => x"38",
          4484 => x"81",
          4485 => x"70",
          4486 => x"70",
          4487 => x"5d",
          4488 => x"cd",
          4489 => x"76",
          4490 => x"57",
          4491 => x"70",
          4492 => x"ff",
          4493 => x"2e",
          4494 => x"38",
          4495 => x"0c",
          4496 => x"84",
          4497 => x"08",
          4498 => x"ba",
          4499 => x"54",
          4500 => x"1b",
          4501 => x"84",
          4502 => x"06",
          4503 => x"83",
          4504 => x"08",
          4505 => x"78",
          4506 => x"82",
          4507 => x"81",
          4508 => x"1b",
          4509 => x"52",
          4510 => x"77",
          4511 => x"e4",
          4512 => x"81",
          4513 => x"76",
          4514 => x"2e",
          4515 => x"bf",
          4516 => x"05",
          4517 => x"af",
          4518 => x"52",
          4519 => x"8c",
          4520 => x"2e",
          4521 => x"80",
          4522 => x"ff",
          4523 => x"8d",
          4524 => x"81",
          4525 => x"1a",
          4526 => x"07",
          4527 => x"78",
          4528 => x"05",
          4529 => x"e6",
          4530 => x"33",
          4531 => x"42",
          4532 => x"79",
          4533 => x"51",
          4534 => x"08",
          4535 => x"43",
          4536 => x"3f",
          4537 => x"81",
          4538 => x"18",
          4539 => x"78",
          4540 => x"59",
          4541 => x"2e",
          4542 => x"22",
          4543 => x"1d",
          4544 => x"ae",
          4545 => x"93",
          4546 => x"2e",
          4547 => x"94",
          4548 => x"70",
          4549 => x"5a",
          4550 => x"38",
          4551 => x"57",
          4552 => x"1d",
          4553 => x"5d",
          4554 => x"5b",
          4555 => x"75",
          4556 => x"81",
          4557 => x"ef",
          4558 => x"81",
          4559 => x"aa",
          4560 => x"81",
          4561 => x"08",
          4562 => x"57",
          4563 => x"76",
          4564 => x"55",
          4565 => x"c2",
          4566 => x"80",
          4567 => x"56",
          4568 => x"07",
          4569 => x"06",
          4570 => x"56",
          4571 => x"84",
          4572 => x"77",
          4573 => x"74",
          4574 => x"cf",
          4575 => x"06",
          4576 => x"15",
          4577 => x"19",
          4578 => x"e3",
          4579 => x"34",
          4580 => x"a0",
          4581 => x"98",
          4582 => x"88",
          4583 => x"57",
          4584 => x"38",
          4585 => x"26",
          4586 => x"05",
          4587 => x"74",
          4588 => x"38",
          4589 => x"8c",
          4590 => x"e3",
          4591 => x"7a",
          4592 => x"ba",
          4593 => x"84",
          4594 => x"02",
          4595 => x"7d",
          4596 => x"33",
          4597 => x"5f",
          4598 => x"8d",
          4599 => x"3f",
          4600 => x"52",
          4601 => x"8c",
          4602 => x"82",
          4603 => x"5e",
          4604 => x"b4",
          4605 => x"83",
          4606 => x"81",
          4607 => x"53",
          4608 => x"d4",
          4609 => x"2e",
          4610 => x"b4",
          4611 => x"9c",
          4612 => x"81",
          4613 => x"70",
          4614 => x"80",
          4615 => x"78",
          4616 => x"7d",
          4617 => x"08",
          4618 => x"ff",
          4619 => x"81",
          4620 => x"38",
          4621 => x"98",
          4622 => x"2e",
          4623 => x"40",
          4624 => x"53",
          4625 => x"d3",
          4626 => x"2e",
          4627 => x"b4",
          4628 => x"38",
          4629 => x"80",
          4630 => x"15",
          4631 => x"1f",
          4632 => x"81",
          4633 => x"59",
          4634 => x"9c",
          4635 => x"5e",
          4636 => x"83",
          4637 => x"8c",
          4638 => x"30",
          4639 => x"57",
          4640 => x"52",
          4641 => x"8c",
          4642 => x"2e",
          4643 => x"54",
          4644 => x"18",
          4645 => x"8c",
          4646 => x"bf",
          4647 => x"34",
          4648 => x"55",
          4649 => x"82",
          4650 => x"ac",
          4651 => x"9c",
          4652 => x"71",
          4653 => x"3f",
          4654 => x"8c",
          4655 => x"8c",
          4656 => x"2a",
          4657 => x"81",
          4658 => x"81",
          4659 => x"76",
          4660 => x"1d",
          4661 => x"56",
          4662 => x"83",
          4663 => x"81",
          4664 => x"53",
          4665 => x"d0",
          4666 => x"2e",
          4667 => x"b4",
          4668 => x"38",
          4669 => x"81",
          4670 => x"1c",
          4671 => x"8c",
          4672 => x"9b",
          4673 => x"76",
          4674 => x"ff",
          4675 => x"22",
          4676 => x"8c",
          4677 => x"70",
          4678 => x"56",
          4679 => x"ff",
          4680 => x"27",
          4681 => x"81",
          4682 => x"58",
          4683 => x"7c",
          4684 => x"80",
          4685 => x"ba",
          4686 => x"fc",
          4687 => x"fe",
          4688 => x"b4",
          4689 => x"81",
          4690 => x"81",
          4691 => x"38",
          4692 => x"b4",
          4693 => x"ba",
          4694 => x"08",
          4695 => x"42",
          4696 => x"bc",
          4697 => x"1d",
          4698 => x"33",
          4699 => x"a4",
          4700 => x"57",
          4701 => x"81",
          4702 => x"81",
          4703 => x"9f",
          4704 => x"07",
          4705 => x"1c",
          4706 => x"51",
          4707 => x"76",
          4708 => x"ba",
          4709 => x"08",
          4710 => x"1d",
          4711 => x"5f",
          4712 => x"8c",
          4713 => x"1c",
          4714 => x"38",
          4715 => x"e8",
          4716 => x"2e",
          4717 => x"54",
          4718 => x"53",
          4719 => x"ac",
          4720 => x"18",
          4721 => x"52",
          4722 => x"f8",
          4723 => x"71",
          4724 => x"1e",
          4725 => x"b5",
          4726 => x"d9",
          4727 => x"08",
          4728 => x"72",
          4729 => x"14",
          4730 => x"7a",
          4731 => x"70",
          4732 => x"8f",
          4733 => x"1a",
          4734 => x"5b",
          4735 => x"25",
          4736 => x"7c",
          4737 => x"18",
          4738 => x"58",
          4739 => x"18",
          4740 => x"38",
          4741 => x"89",
          4742 => x"25",
          4743 => x"38",
          4744 => x"70",
          4745 => x"74",
          4746 => x"18",
          4747 => x"7c",
          4748 => x"16",
          4749 => x"38",
          4750 => x"1e",
          4751 => x"56",
          4752 => x"08",
          4753 => x"38",
          4754 => x"53",
          4755 => x"1c",
          4756 => x"12",
          4757 => x"07",
          4758 => x"2b",
          4759 => x"97",
          4760 => x"2b",
          4761 => x"5b",
          4762 => x"33",
          4763 => x"5d",
          4764 => x"0d",
          4765 => x"77",
          4766 => x"58",
          4767 => x"2b",
          4768 => x"84",
          4769 => x"55",
          4770 => x"76",
          4771 => x"54",
          4772 => x"82",
          4773 => x"08",
          4774 => x"22",
          4775 => x"fd",
          4776 => x"78",
          4777 => x"58",
          4778 => x"7a",
          4779 => x"8c",
          4780 => x"73",
          4781 => x"80",
          4782 => x"7e",
          4783 => x"bf",
          4784 => x"38",
          4785 => x"5b",
          4786 => x"2a",
          4787 => x"2e",
          4788 => x"ff",
          4789 => x"05",
          4790 => x"19",
          4791 => x"56",
          4792 => x"39",
          4793 => x"7b",
          4794 => x"06",
          4795 => x"ef",
          4796 => x"57",
          4797 => x"53",
          4798 => x"74",
          4799 => x"80",
          4800 => x"88",
          4801 => x"3d",
          4802 => x"a7",
          4803 => x"80",
          4804 => x"33",
          4805 => x"7f",
          4806 => x"83",
          4807 => x"10",
          4808 => x"57",
          4809 => x"32",
          4810 => x"25",
          4811 => x"90",
          4812 => x"38",
          4813 => x"e5",
          4814 => x"81",
          4815 => x"2e",
          4816 => x"38",
          4817 => x"06",
          4818 => x"81",
          4819 => x"76",
          4820 => x"10",
          4821 => x"62",
          4822 => x"54",
          4823 => x"80",
          4824 => x"70",
          4825 => x"55",
          4826 => x"81",
          4827 => x"54",
          4828 => x"80",
          4829 => x"77",
          4830 => x"72",
          4831 => x"94",
          4832 => x"fe",
          4833 => x"73",
          4834 => x"8c",
          4835 => x"fe",
          4836 => x"8c",
          4837 => x"a8",
          4838 => x"7a",
          4839 => x"ff",
          4840 => x"7b",
          4841 => x"08",
          4842 => x"04",
          4843 => x"70",
          4844 => x"56",
          4845 => x"42",
          4846 => x"72",
          4847 => x"32",
          4848 => x"40",
          4849 => x"0c",
          4850 => x"81",
          4851 => x"83",
          4852 => x"2e",
          4853 => x"05",
          4854 => x"70",
          4855 => x"59",
          4856 => x"38",
          4857 => x"59",
          4858 => x"80",
          4859 => x"70",
          4860 => x"55",
          4861 => x"73",
          4862 => x"2e",
          4863 => x"38",
          4864 => x"54",
          4865 => x"18",
          4866 => x"80",
          4867 => x"5e",
          4868 => x"eb",
          4869 => x"a0",
          4870 => x"13",
          4871 => x"5e",
          4872 => x"59",
          4873 => x"ed",
          4874 => x"74",
          4875 => x"55",
          4876 => x"38",
          4877 => x"7b",
          4878 => x"32",
          4879 => x"70",
          4880 => x"80",
          4881 => x"86",
          4882 => x"79",
          4883 => x"38",
          4884 => x"2b",
          4885 => x"5d",
          4886 => x"56",
          4887 => x"33",
          4888 => x"38",
          4889 => x"8c",
          4890 => x"38",
          4891 => x"82",
          4892 => x"56",
          4893 => x"7c",
          4894 => x"5a",
          4895 => x"80",
          4896 => x"79",
          4897 => x"3f",
          4898 => x"56",
          4899 => x"81",
          4900 => x"2e",
          4901 => x"85",
          4902 => x"84",
          4903 => x"59",
          4904 => x"55",
          4905 => x"80",
          4906 => x"11",
          4907 => x"56",
          4908 => x"2e",
          4909 => x"fd",
          4910 => x"ae",
          4911 => x"77",
          4912 => x"06",
          4913 => x"80",
          4914 => x"53",
          4915 => x"a0",
          4916 => x"34",
          4917 => x"38",
          4918 => x"34",
          4919 => x"8c",
          4920 => x"ba",
          4921 => x"2a",
          4922 => x"86",
          4923 => x"56",
          4924 => x"90",
          4925 => x"80",
          4926 => x"71",
          4927 => x"54",
          4928 => x"74",
          4929 => x"56",
          4930 => x"ae",
          4931 => x"76",
          4932 => x"83",
          4933 => x"39",
          4934 => x"8c",
          4935 => x"81",
          4936 => x"5a",
          4937 => x"34",
          4938 => x"f6",
          4939 => x"1d",
          4940 => x"93",
          4941 => x"9d",
          4942 => x"38",
          4943 => x"f7",
          4944 => x"57",
          4945 => x"07",
          4946 => x"85",
          4947 => x"ff",
          4948 => x"5a",
          4949 => x"80",
          4950 => x"56",
          4951 => x"38",
          4952 => x"e5",
          4953 => x"81",
          4954 => x"2e",
          4955 => x"38",
          4956 => x"06",
          4957 => x"81",
          4958 => x"ff",
          4959 => x"38",
          4960 => x"5f",
          4961 => x"26",
          4962 => x"ff",
          4963 => x"06",
          4964 => x"05",
          4965 => x"75",
          4966 => x"fa",
          4967 => x"81",
          4968 => x"ff",
          4969 => x"7d",
          4970 => x"79",
          4971 => x"cd",
          4972 => x"98",
          4973 => x"88",
          4974 => x"7b",
          4975 => x"54",
          4976 => x"a0",
          4977 => x"1b",
          4978 => x"a0",
          4979 => x"2e",
          4980 => x"a3",
          4981 => x"7b",
          4982 => x"8c",
          4983 => x"0d",
          4984 => x"05",
          4985 => x"ff",
          4986 => x"80",
          4987 => x"05",
          4988 => x"75",
          4989 => x"38",
          4990 => x"d1",
          4991 => x"b2",
          4992 => x"05",
          4993 => x"80",
          4994 => x"7f",
          4995 => x"7b",
          4996 => x"51",
          4997 => x"08",
          4998 => x"58",
          4999 => x"77",
          5000 => x"1d",
          5001 => x"17",
          5002 => x"ba",
          5003 => x"06",
          5004 => x"38",
          5005 => x"2a",
          5006 => x"b1",
          5007 => x"ff",
          5008 => x"55",
          5009 => x"53",
          5010 => x"95",
          5011 => x"85",
          5012 => x"18",
          5013 => x"b7",
          5014 => x"88",
          5015 => x"82",
          5016 => x"81",
          5017 => x"33",
          5018 => x"75",
          5019 => x"75",
          5020 => x"17",
          5021 => x"2b",
          5022 => x"09",
          5023 => x"17",
          5024 => x"2b",
          5025 => x"dc",
          5026 => x"71",
          5027 => x"14",
          5028 => x"33",
          5029 => x"5f",
          5030 => x"17",
          5031 => x"33",
          5032 => x"40",
          5033 => x"d9",
          5034 => x"29",
          5035 => x"77",
          5036 => x"2e",
          5037 => x"42",
          5038 => x"33",
          5039 => x"07",
          5040 => x"75",
          5041 => x"82",
          5042 => x"cb",
          5043 => x"5c",
          5044 => x"11",
          5045 => x"71",
          5046 => x"72",
          5047 => x"53",
          5048 => x"c7",
          5049 => x"88",
          5050 => x"80",
          5051 => x"84",
          5052 => x"c1",
          5053 => x"fd",
          5054 => x"56",
          5055 => x"a9",
          5056 => x"ff",
          5057 => x"75",
          5058 => x"5d",
          5059 => x"81",
          5060 => x"7b",
          5061 => x"1a",
          5062 => x"59",
          5063 => x"17",
          5064 => x"80",
          5065 => x"78",
          5066 => x"78",
          5067 => x"06",
          5068 => x"2a",
          5069 => x"26",
          5070 => x"ff",
          5071 => x"84",
          5072 => x"38",
          5073 => x"81",
          5074 => x"7c",
          5075 => x"8c",
          5076 => x"80",
          5077 => x"3d",
          5078 => x"0c",
          5079 => x"11",
          5080 => x"74",
          5081 => x"81",
          5082 => x"7a",
          5083 => x"83",
          5084 => x"7f",
          5085 => x"33",
          5086 => x"9f",
          5087 => x"89",
          5088 => x"57",
          5089 => x"26",
          5090 => x"06",
          5091 => x"59",
          5092 => x"85",
          5093 => x"32",
          5094 => x"7a",
          5095 => x"87",
          5096 => x"5c",
          5097 => x"56",
          5098 => x"cf",
          5099 => x"8a",
          5100 => x"fe",
          5101 => x"75",
          5102 => x"38",
          5103 => x"30",
          5104 => x"5c",
          5105 => x"2e",
          5106 => x"5a",
          5107 => x"59",
          5108 => x"81",
          5109 => x"90",
          5110 => x"19",
          5111 => x"fe",
          5112 => x"40",
          5113 => x"5c",
          5114 => x"78",
          5115 => x"81",
          5116 => x"72",
          5117 => x"05",
          5118 => x"52",
          5119 => x"56",
          5120 => x"0b",
          5121 => x"0c",
          5122 => x"a5",
          5123 => x"52",
          5124 => x"3f",
          5125 => x"38",
          5126 => x"0c",
          5127 => x"33",
          5128 => x"5e",
          5129 => x"09",
          5130 => x"18",
          5131 => x"82",
          5132 => x"30",
          5133 => x"42",
          5134 => x"b6",
          5135 => x"56",
          5136 => x"5d",
          5137 => x"83",
          5138 => x"bd",
          5139 => x"81",
          5140 => x"27",
          5141 => x"0b",
          5142 => x"5d",
          5143 => x"7e",
          5144 => x"31",
          5145 => x"80",
          5146 => x"e1",
          5147 => x"e5",
          5148 => x"05",
          5149 => x"33",
          5150 => x"42",
          5151 => x"75",
          5152 => x"f3",
          5153 => x"77",
          5154 => x"04",
          5155 => x"38",
          5156 => x"c0",
          5157 => x"0b",
          5158 => x"04",
          5159 => x"bc",
          5160 => x"5a",
          5161 => x"71",
          5162 => x"5f",
          5163 => x"80",
          5164 => x"18",
          5165 => x"70",
          5166 => x"05",
          5167 => x"5b",
          5168 => x"91",
          5169 => x"3d",
          5170 => x"39",
          5171 => x"17",
          5172 => x"2b",
          5173 => x"81",
          5174 => x"80",
          5175 => x"38",
          5176 => x"09",
          5177 => x"77",
          5178 => x"51",
          5179 => x"08",
          5180 => x"5a",
          5181 => x"38",
          5182 => x"33",
          5183 => x"07",
          5184 => x"09",
          5185 => x"83",
          5186 => x"2b",
          5187 => x"70",
          5188 => x"07",
          5189 => x"77",
          5190 => x"81",
          5191 => x"83",
          5192 => x"2b",
          5193 => x"70",
          5194 => x"07",
          5195 => x"60",
          5196 => x"81",
          5197 => x"83",
          5198 => x"2b",
          5199 => x"70",
          5200 => x"07",
          5201 => x"83",
          5202 => x"2b",
          5203 => x"70",
          5204 => x"07",
          5205 => x"46",
          5206 => x"7c",
          5207 => x"05",
          5208 => x"86",
          5209 => x"18",
          5210 => x"cf",
          5211 => x"7b",
          5212 => x"75",
          5213 => x"70",
          5214 => x"af",
          5215 => x"2e",
          5216 => x"ba",
          5217 => x"08",
          5218 => x"18",
          5219 => x"41",
          5220 => x"ba",
          5221 => x"56",
          5222 => x"0b",
          5223 => x"5a",
          5224 => x"33",
          5225 => x"07",
          5226 => x"38",
          5227 => x"38",
          5228 => x"12",
          5229 => x"07",
          5230 => x"2b",
          5231 => x"5a",
          5232 => x"59",
          5233 => x"80",
          5234 => x"e3",
          5235 => x"93",
          5236 => x"f2",
          5237 => x"fc",
          5238 => x"a0",
          5239 => x"17",
          5240 => x"85",
          5241 => x"05",
          5242 => x"57",
          5243 => x"2e",
          5244 => x"5a",
          5245 => x"ba",
          5246 => x"74",
          5247 => x"e8",
          5248 => x"38",
          5249 => x"70",
          5250 => x"38",
          5251 => x"2e",
          5252 => x"73",
          5253 => x"92",
          5254 => x"84",
          5255 => x"8c",
          5256 => x"92",
          5257 => x"8c",
          5258 => x"d0",
          5259 => x"57",
          5260 => x"77",
          5261 => x"77",
          5262 => x"08",
          5263 => x"08",
          5264 => x"5b",
          5265 => x"ff",
          5266 => x"26",
          5267 => x"06",
          5268 => x"99",
          5269 => x"ff",
          5270 => x"2a",
          5271 => x"06",
          5272 => x"79",
          5273 => x"2a",
          5274 => x"2e",
          5275 => x"5b",
          5276 => x"54",
          5277 => x"38",
          5278 => x"39",
          5279 => x"80",
          5280 => x"78",
          5281 => x"70",
          5282 => x"3d",
          5283 => x"84",
          5284 => x"08",
          5285 => x"76",
          5286 => x"3d",
          5287 => x"3d",
          5288 => x"ba",
          5289 => x"80",
          5290 => x"5d",
          5291 => x"80",
          5292 => x"83",
          5293 => x"ff",
          5294 => x"5b",
          5295 => x"9b",
          5296 => x"2b",
          5297 => x"5e",
          5298 => x"80",
          5299 => x"17",
          5300 => x"cc",
          5301 => x"0b",
          5302 => x"80",
          5303 => x"17",
          5304 => x"84",
          5305 => x"1c",
          5306 => x"0b",
          5307 => x"34",
          5308 => x"7b",
          5309 => x"11",
          5310 => x"57",
          5311 => x"08",
          5312 => x"80",
          5313 => x"e7",
          5314 => x"7b",
          5315 => x"9c",
          5316 => x"76",
          5317 => x"33",
          5318 => x"7b",
          5319 => x"06",
          5320 => x"81",
          5321 => x"83",
          5322 => x"86",
          5323 => x"b4",
          5324 => x"1b",
          5325 => x"33",
          5326 => x"5e",
          5327 => x"f1",
          5328 => x"83",
          5329 => x"2b",
          5330 => x"70",
          5331 => x"07",
          5332 => x"0c",
          5333 => x"86",
          5334 => x"1a",
          5335 => x"0b",
          5336 => x"06",
          5337 => x"75",
          5338 => x"1a",
          5339 => x"7c",
          5340 => x"07",
          5341 => x"84",
          5342 => x"5b",
          5343 => x"52",
          5344 => x"ba",
          5345 => x"81",
          5346 => x"8c",
          5347 => x"7a",
          5348 => x"05",
          5349 => x"77",
          5350 => x"2e",
          5351 => x"0c",
          5352 => x"0c",
          5353 => x"0c",
          5354 => x"3f",
          5355 => x"59",
          5356 => x"39",
          5357 => x"f3",
          5358 => x"71",
          5359 => x"07",
          5360 => x"55",
          5361 => x"52",
          5362 => x"ba",
          5363 => x"80",
          5364 => x"08",
          5365 => x"8c",
          5366 => x"53",
          5367 => x"3f",
          5368 => x"9c",
          5369 => x"58",
          5370 => x"38",
          5371 => x"33",
          5372 => x"7c",
          5373 => x"80",
          5374 => x"80",
          5375 => x"95",
          5376 => x"2b",
          5377 => x"56",
          5378 => x"0b",
          5379 => x"34",
          5380 => x"56",
          5381 => x"57",
          5382 => x"0b",
          5383 => x"83",
          5384 => x"ff",
          5385 => x"59",
          5386 => x"ae",
          5387 => x"2e",
          5388 => x"7d",
          5389 => x"51",
          5390 => x"08",
          5391 => x"5b",
          5392 => x"ff",
          5393 => x"2e",
          5394 => x"97",
          5395 => x"b8",
          5396 => x"5a",
          5397 => x"08",
          5398 => x"38",
          5399 => x"b4",
          5400 => x"ba",
          5401 => x"08",
          5402 => x"55",
          5403 => x"85",
          5404 => x"17",
          5405 => x"33",
          5406 => x"fe",
          5407 => x"56",
          5408 => x"76",
          5409 => x"5a",
          5410 => x"fe",
          5411 => x"59",
          5412 => x"8a",
          5413 => x"08",
          5414 => x"cd",
          5415 => x"0c",
          5416 => x"1a",
          5417 => x"57",
          5418 => x"ba",
          5419 => x"cf",
          5420 => x"39",
          5421 => x"40",
          5422 => x"57",
          5423 => x"56",
          5424 => x"55",
          5425 => x"22",
          5426 => x"2e",
          5427 => x"76",
          5428 => x"33",
          5429 => x"33",
          5430 => x"2e",
          5431 => x"1b",
          5432 => x"26",
          5433 => x"d5",
          5434 => x"5b",
          5435 => x"ff",
          5436 => x"9b",
          5437 => x"08",
          5438 => x"74",
          5439 => x"1b",
          5440 => x"05",
          5441 => x"76",
          5442 => x"22",
          5443 => x"56",
          5444 => x"7a",
          5445 => x"80",
          5446 => x"75",
          5447 => x"58",
          5448 => x"19",
          5449 => x"ba",
          5450 => x"11",
          5451 => x"38",
          5452 => x"78",
          5453 => x"29",
          5454 => x"70",
          5455 => x"05",
          5456 => x"38",
          5457 => x"7e",
          5458 => x"1c",
          5459 => x"5e",
          5460 => x"75",
          5461 => x"04",
          5462 => x"0d",
          5463 => x"1a",
          5464 => x"80",
          5465 => x"83",
          5466 => x"08",
          5467 => x"1a",
          5468 => x"2e",
          5469 => x"54",
          5470 => x"33",
          5471 => x"8c",
          5472 => x"81",
          5473 => x"dc",
          5474 => x"06",
          5475 => x"56",
          5476 => x"74",
          5477 => x"81",
          5478 => x"80",
          5479 => x"05",
          5480 => x"34",
          5481 => x"bc",
          5482 => x"b8",
          5483 => x"40",
          5484 => x"ba",
          5485 => x"ff",
          5486 => x"1a",
          5487 => x"31",
          5488 => x"a0",
          5489 => x"19",
          5490 => x"06",
          5491 => x"08",
          5492 => x"81",
          5493 => x"7e",
          5494 => x"0c",
          5495 => x"98",
          5496 => x"98",
          5497 => x"a1",
          5498 => x"83",
          5499 => x"55",
          5500 => x"56",
          5501 => x"1b",
          5502 => x"92",
          5503 => x"34",
          5504 => x"3d",
          5505 => x"67",
          5506 => x"0c",
          5507 => x"79",
          5508 => x"75",
          5509 => x"86",
          5510 => x"78",
          5511 => x"74",
          5512 => x"91",
          5513 => x"90",
          5514 => x"58",
          5515 => x"a1",
          5516 => x"57",
          5517 => x"5b",
          5518 => x"83",
          5519 => x"60",
          5520 => x"2a",
          5521 => x"84",
          5522 => x"80",
          5523 => x"86",
          5524 => x"38",
          5525 => x"85",
          5526 => x"b4",
          5527 => x"d3",
          5528 => x"17",
          5529 => x"27",
          5530 => x"79",
          5531 => x"74",
          5532 => x"7b",
          5533 => x"83",
          5534 => x"27",
          5535 => x"54",
          5536 => x"51",
          5537 => x"08",
          5538 => x"7d",
          5539 => x"38",
          5540 => x"29",
          5541 => x"05",
          5542 => x"34",
          5543 => x"59",
          5544 => x"59",
          5545 => x"0c",
          5546 => x"71",
          5547 => x"5a",
          5548 => x"38",
          5549 => x"fe",
          5550 => x"80",
          5551 => x"80",
          5552 => x"3d",
          5553 => x"92",
          5554 => x"74",
          5555 => x"39",
          5556 => x"83",
          5557 => x"5c",
          5558 => x"77",
          5559 => x"38",
          5560 => x"41",
          5561 => x"80",
          5562 => x"16",
          5563 => x"cd",
          5564 => x"85",
          5565 => x"17",
          5566 => x"1b",
          5567 => x"b8",
          5568 => x"2e",
          5569 => x"33",
          5570 => x"16",
          5571 => x"0b",
          5572 => x"54",
          5573 => x"53",
          5574 => x"f4",
          5575 => x"7f",
          5576 => x"84",
          5577 => x"16",
          5578 => x"8c",
          5579 => x"27",
          5580 => x"74",
          5581 => x"38",
          5582 => x"08",
          5583 => x"51",
          5584 => x"ca",
          5585 => x"08",
          5586 => x"40",
          5587 => x"12",
          5588 => x"7c",
          5589 => x"98",
          5590 => x"e7",
          5591 => x"ba",
          5592 => x"33",
          5593 => x"51",
          5594 => x"08",
          5595 => x"38",
          5596 => x"53",
          5597 => x"52",
          5598 => x"8c",
          5599 => x"08",
          5600 => x"17",
          5601 => x"27",
          5602 => x"7b",
          5603 => x"38",
          5604 => x"08",
          5605 => x"51",
          5606 => x"89",
          5607 => x"9b",
          5608 => x"55",
          5609 => x"56",
          5610 => x"16",
          5611 => x"17",
          5612 => x"84",
          5613 => x"ba",
          5614 => x"08",
          5615 => x"17",
          5616 => x"33",
          5617 => x"fe",
          5618 => x"a0",
          5619 => x"16",
          5620 => x"7c",
          5621 => x"56",
          5622 => x"34",
          5623 => x"3d",
          5624 => x"82",
          5625 => x"0d",
          5626 => x"5a",
          5627 => x"56",
          5628 => x"55",
          5629 => x"22",
          5630 => x"2e",
          5631 => x"79",
          5632 => x"33",
          5633 => x"7a",
          5634 => x"19",
          5635 => x"2e",
          5636 => x"81",
          5637 => x"17",
          5638 => x"f5",
          5639 => x"85",
          5640 => x"18",
          5641 => x"08",
          5642 => x"78",
          5643 => x"08",
          5644 => x"56",
          5645 => x"5a",
          5646 => x"33",
          5647 => x"2e",
          5648 => x"74",
          5649 => x"9d",
          5650 => x"9e",
          5651 => x"9f",
          5652 => x"97",
          5653 => x"80",
          5654 => x"92",
          5655 => x"7b",
          5656 => x"51",
          5657 => x"08",
          5658 => x"56",
          5659 => x"8c",
          5660 => x"b4",
          5661 => x"81",
          5662 => x"3f",
          5663 => x"c9",
          5664 => x"34",
          5665 => x"84",
          5666 => x"18",
          5667 => x"33",
          5668 => x"fe",
          5669 => x"a0",
          5670 => x"17",
          5671 => x"56",
          5672 => x"74",
          5673 => x"75",
          5674 => x"74",
          5675 => x"9d",
          5676 => x"9e",
          5677 => x"9f",
          5678 => x"97",
          5679 => x"80",
          5680 => x"92",
          5681 => x"7b",
          5682 => x"51",
          5683 => x"08",
          5684 => x"56",
          5685 => x"81",
          5686 => x"84",
          5687 => x"fc",
          5688 => x"fc",
          5689 => x"52",
          5690 => x"08",
          5691 => x"89",
          5692 => x"08",
          5693 => x"33",
          5694 => x"13",
          5695 => x"77",
          5696 => x"75",
          5697 => x"73",
          5698 => x"04",
          5699 => x"3f",
          5700 => x"72",
          5701 => x"d5",
          5702 => x"5b",
          5703 => x"75",
          5704 => x"26",
          5705 => x"70",
          5706 => x"84",
          5707 => x"90",
          5708 => x"0b",
          5709 => x"04",
          5710 => x"3d",
          5711 => x"81",
          5712 => x"26",
          5713 => x"06",
          5714 => x"80",
          5715 => x"5b",
          5716 => x"70",
          5717 => x"05",
          5718 => x"52",
          5719 => x"70",
          5720 => x"13",
          5721 => x"13",
          5722 => x"30",
          5723 => x"2e",
          5724 => x"be",
          5725 => x"72",
          5726 => x"52",
          5727 => x"84",
          5728 => x"99",
          5729 => x"83",
          5730 => x"fe",
          5731 => x"98",
          5732 => x"d1",
          5733 => x"84",
          5734 => x"74",
          5735 => x"04",
          5736 => x"05",
          5737 => x"08",
          5738 => x"38",
          5739 => x"2b",
          5740 => x"38",
          5741 => x"81",
          5742 => x"38",
          5743 => x"33",
          5744 => x"5a",
          5745 => x"38",
          5746 => x"8c",
          5747 => x"8c",
          5748 => x"8f",
          5749 => x"98",
          5750 => x"17",
          5751 => x"07",
          5752 => x"cc",
          5753 => x"74",
          5754 => x"04",
          5755 => x"08",
          5756 => x"7c",
          5757 => x"b4",
          5758 => x"c5",
          5759 => x"ba",
          5760 => x"d9",
          5761 => x"80",
          5762 => x"08",
          5763 => x"38",
          5764 => x"a0",
          5765 => x"84",
          5766 => x"08",
          5767 => x"08",
          5768 => x"b1",
          5769 => x"33",
          5770 => x"54",
          5771 => x"33",
          5772 => x"8c",
          5773 => x"81",
          5774 => x"d4",
          5775 => x"33",
          5776 => x"63",
          5777 => x"78",
          5778 => x"db",
          5779 => x"a3",
          5780 => x"84",
          5781 => x"52",
          5782 => x"ba",
          5783 => x"bb",
          5784 => x"33",
          5785 => x"63",
          5786 => x"7d",
          5787 => x"2e",
          5788 => x"7a",
          5789 => x"8c",
          5790 => x"2e",
          5791 => x"d8",
          5792 => x"3d",
          5793 => x"bd",
          5794 => x"5b",
          5795 => x"1f",
          5796 => x"5f",
          5797 => x"56",
          5798 => x"80",
          5799 => x"56",
          5800 => x"ff",
          5801 => x"75",
          5802 => x"18",
          5803 => x"af",
          5804 => x"79",
          5805 => x"8a",
          5806 => x"70",
          5807 => x"08",
          5808 => x"7e",
          5809 => x"17",
          5810 => x"38",
          5811 => x"38",
          5812 => x"76",
          5813 => x"05",
          5814 => x"26",
          5815 => x"5e",
          5816 => x"81",
          5817 => x"78",
          5818 => x"0d",
          5819 => x"71",
          5820 => x"07",
          5821 => x"16",
          5822 => x"71",
          5823 => x"3d",
          5824 => x"ff",
          5825 => x"59",
          5826 => x"96",
          5827 => x"16",
          5828 => x"17",
          5829 => x"81",
          5830 => x"38",
          5831 => x"b4",
          5832 => x"ba",
          5833 => x"08",
          5834 => x"55",
          5835 => x"f6",
          5836 => x"17",
          5837 => x"33",
          5838 => x"fb",
          5839 => x"08",
          5840 => x"0b",
          5841 => x"83",
          5842 => x"43",
          5843 => x"09",
          5844 => x"39",
          5845 => x"59",
          5846 => x"5e",
          5847 => x"80",
          5848 => x"5a",
          5849 => x"34",
          5850 => x"39",
          5851 => x"ba",
          5852 => x"f7",
          5853 => x"56",
          5854 => x"54",
          5855 => x"53",
          5856 => x"22",
          5857 => x"2e",
          5858 => x"75",
          5859 => x"33",
          5860 => x"08",
          5861 => x"94",
          5862 => x"2e",
          5863 => x"70",
          5864 => x"2e",
          5865 => x"51",
          5866 => x"08",
          5867 => x"53",
          5868 => x"08",
          5869 => x"74",
          5870 => x"31",
          5871 => x"80",
          5872 => x"81",
          5873 => x"08",
          5874 => x"70",
          5875 => x"78",
          5876 => x"74",
          5877 => x"8c",
          5878 => x"2e",
          5879 => x"38",
          5880 => x"53",
          5881 => x"38",
          5882 => x"81",
          5883 => x"84",
          5884 => x"90",
          5885 => x"55",
          5886 => x"16",
          5887 => x"2e",
          5888 => x"94",
          5889 => x"74",
          5890 => x"90",
          5891 => x"90",
          5892 => x"78",
          5893 => x"78",
          5894 => x"80",
          5895 => x"0d",
          5896 => x"15",
          5897 => x"38",
          5898 => x"80",
          5899 => x"8c",
          5900 => x"16",
          5901 => x"80",
          5902 => x"12",
          5903 => x"78",
          5904 => x"74",
          5905 => x"89",
          5906 => x"2e",
          5907 => x"fe",
          5908 => x"89",
          5909 => x"fe",
          5910 => x"82",
          5911 => x"06",
          5912 => x"08",
          5913 => x"74",
          5914 => x"8c",
          5915 => x"2e",
          5916 => x"2e",
          5917 => x"88",
          5918 => x"dc",
          5919 => x"0b",
          5920 => x"04",
          5921 => x"75",
          5922 => x"3d",
          5923 => x"51",
          5924 => x"55",
          5925 => x"38",
          5926 => x"ba",
          5927 => x"76",
          5928 => x"97",
          5929 => x"ba",
          5930 => x"33",
          5931 => x"24",
          5932 => x"2a",
          5933 => x"80",
          5934 => x"33",
          5935 => x"7d",
          5936 => x"78",
          5937 => x"0c",
          5938 => x"23",
          5939 => x"3f",
          5940 => x"2e",
          5941 => x"38",
          5942 => x"55",
          5943 => x"17",
          5944 => x"71",
          5945 => x"0c",
          5946 => x"0d",
          5947 => x"9e",
          5948 => x"96",
          5949 => x"8e",
          5950 => x"57",
          5951 => x"52",
          5952 => x"0c",
          5953 => x"0d",
          5954 => x"c3",
          5955 => x"52",
          5956 => x"54",
          5957 => x"58",
          5958 => x"38",
          5959 => x"38",
          5960 => x"38",
          5961 => x"53",
          5962 => x"53",
          5963 => x"38",
          5964 => x"52",
          5965 => x"ba",
          5966 => x"84",
          5967 => x"a6",
          5968 => x"92",
          5969 => x"be",
          5970 => x"70",
          5971 => x"ba",
          5972 => x"84",
          5973 => x"75",
          5974 => x"e2",
          5975 => x"8e",
          5976 => x"70",
          5977 => x"ba",
          5978 => x"39",
          5979 => x"3f",
          5980 => x"0c",
          5981 => x"51",
          5982 => x"08",
          5983 => x"72",
          5984 => x"ed",
          5985 => x"3d",
          5986 => x"a5",
          5987 => x"ba",
          5988 => x"84",
          5989 => x"65",
          5990 => x"84",
          5991 => x"08",
          5992 => x"70",
          5993 => x"97",
          5994 => x"52",
          5995 => x"84",
          5996 => x"86",
          5997 => x"0d",
          5998 => x"5f",
          5999 => x"96",
          6000 => x"8c",
          6001 => x"38",
          6002 => x"08",
          6003 => x"59",
          6004 => x"7f",
          6005 => x"3d",
          6006 => x"33",
          6007 => x"38",
          6008 => x"08",
          6009 => x"7b",
          6010 => x"17",
          6011 => x"17",
          6012 => x"38",
          6013 => x"81",
          6014 => x"84",
          6015 => x"ff",
          6016 => x"7f",
          6017 => x"76",
          6018 => x"38",
          6019 => x"82",
          6020 => x"2b",
          6021 => x"88",
          6022 => x"fe",
          6023 => x"25",
          6024 => x"06",
          6025 => x"54",
          6026 => x"fe",
          6027 => x"18",
          6028 => x"77",
          6029 => x"0c",
          6030 => x"17",
          6031 => x"18",
          6032 => x"81",
          6033 => x"38",
          6034 => x"b4",
          6035 => x"ba",
          6036 => x"08",
          6037 => x"55",
          6038 => x"b0",
          6039 => x"18",
          6040 => x"33",
          6041 => x"fe",
          6042 => x"59",
          6043 => x"80",
          6044 => x"80",
          6045 => x"2e",
          6046 => x"30",
          6047 => x"25",
          6048 => x"5c",
          6049 => x"38",
          6050 => x"84",
          6051 => x"18",
          6052 => x"05",
          6053 => x"2b",
          6054 => x"82",
          6055 => x"5d",
          6056 => x"83",
          6057 => x"bf",
          6058 => x"0c",
          6059 => x"81",
          6060 => x"83",
          6061 => x"f7",
          6062 => x"80",
          6063 => x"80",
          6064 => x"80",
          6065 => x"18",
          6066 => x"da",
          6067 => x"dc",
          6068 => x"d4",
          6069 => x"81",
          6070 => x"2e",
          6071 => x"73",
          6072 => x"81",
          6073 => x"57",
          6074 => x"16",
          6075 => x"80",
          6076 => x"8c",
          6077 => x"78",
          6078 => x"38",
          6079 => x"84",
          6080 => x"78",
          6081 => x"73",
          6082 => x"84",
          6083 => x"08",
          6084 => x"8c",
          6085 => x"ba",
          6086 => x"80",
          6087 => x"81",
          6088 => x"38",
          6089 => x"08",
          6090 => x"af",
          6091 => x"16",
          6092 => x"34",
          6093 => x"38",
          6094 => x"f6",
          6095 => x"06",
          6096 => x"08",
          6097 => x"90",
          6098 => x"0b",
          6099 => x"17",
          6100 => x"3f",
          6101 => x"c2",
          6102 => x"81",
          6103 => x"58",
          6104 => x"27",
          6105 => x"98",
          6106 => x"81",
          6107 => x"a1",
          6108 => x"08",
          6109 => x"97",
          6110 => x"ff",
          6111 => x"55",
          6112 => x"73",
          6113 => x"84",
          6114 => x"08",
          6115 => x"8c",
          6116 => x"ba",
          6117 => x"80",
          6118 => x"89",
          6119 => x"38",
          6120 => x"08",
          6121 => x"38",
          6122 => x"33",
          6123 => x"78",
          6124 => x"80",
          6125 => x"fc",
          6126 => x"82",
          6127 => x"e4",
          6128 => x"90",
          6129 => x"84",
          6130 => x"54",
          6131 => x"33",
          6132 => x"8c",
          6133 => x"bb",
          6134 => x"3d",
          6135 => x"ff",
          6136 => x"56",
          6137 => x"38",
          6138 => x"0d",
          6139 => x"9b",
          6140 => x"3f",
          6141 => x"8c",
          6142 => x"33",
          6143 => x"86",
          6144 => x"5b",
          6145 => x"ee",
          6146 => x"87",
          6147 => x"3d",
          6148 => x"71",
          6149 => x"5c",
          6150 => x"38",
          6151 => x"80",
          6152 => x"18",
          6153 => x"5f",
          6154 => x"8f",
          6155 => x"3f",
          6156 => x"8c",
          6157 => x"08",
          6158 => x"84",
          6159 => x"08",
          6160 => x"0c",
          6161 => x"94",
          6162 => x"2b",
          6163 => x"98",
          6164 => x"88",
          6165 => x"38",
          6166 => x"5d",
          6167 => x"74",
          6168 => x"84",
          6169 => x"08",
          6170 => x"77",
          6171 => x"2e",
          6172 => x"7a",
          6173 => x"89",
          6174 => x"fd",
          6175 => x"7d",
          6176 => x"8c",
          6177 => x"0d",
          6178 => x"56",
          6179 => x"82",
          6180 => x"55",
          6181 => x"dd",
          6182 => x"52",
          6183 => x"3f",
          6184 => x"38",
          6185 => x"0c",
          6186 => x"08",
          6187 => x"18",
          6188 => x"ec",
          6189 => x"de",
          6190 => x"ba",
          6191 => x"75",
          6192 => x"38",
          6193 => x"b4",
          6194 => x"33",
          6195 => x"84",
          6196 => x"06",
          6197 => x"83",
          6198 => x"08",
          6199 => x"74",
          6200 => x"82",
          6201 => x"81",
          6202 => x"17",
          6203 => x"52",
          6204 => x"3f",
          6205 => x"79",
          6206 => x"78",
          6207 => x"8c",
          6208 => x"2e",
          6209 => x"81",
          6210 => x"08",
          6211 => x"74",
          6212 => x"84",
          6213 => x"08",
          6214 => x"58",
          6215 => x"16",
          6216 => x"07",
          6217 => x"77",
          6218 => x"fd",
          6219 => x"84",
          6220 => x"81",
          6221 => x"82",
          6222 => x"a0",
          6223 => x"ba",
          6224 => x"80",
          6225 => x"0c",
          6226 => x"52",
          6227 => x"bf",
          6228 => x"ba",
          6229 => x"ba",
          6230 => x"ba",
          6231 => x"cb",
          6232 => x"85",
          6233 => x"74",
          6234 => x"8f",
          6235 => x"3f",
          6236 => x"84",
          6237 => x"84",
          6238 => x"38",
          6239 => x"cb",
          6240 => x"ba",
          6241 => x"57",
          6242 => x"18",
          6243 => x"75",
          6244 => x"76",
          6245 => x"58",
          6246 => x"84",
          6247 => x"81",
          6248 => x"f4",
          6249 => x"77",
          6250 => x"77",
          6251 => x"51",
          6252 => x"08",
          6253 => x"39",
          6254 => x"b4",
          6255 => x"81",
          6256 => x"3f",
          6257 => x"38",
          6258 => x"b4",
          6259 => x"74",
          6260 => x"82",
          6261 => x"81",
          6262 => x"17",
          6263 => x"52",
          6264 => x"3f",
          6265 => x"08",
          6266 => x"38",
          6267 => x"38",
          6268 => x"3f",
          6269 => x"8c",
          6270 => x"ba",
          6271 => x"84",
          6272 => x"38",
          6273 => x"f9",
          6274 => x"f3",
          6275 => x"19",
          6276 => x"90",
          6277 => x"17",
          6278 => x"34",
          6279 => x"38",
          6280 => x"0d",
          6281 => x"ff",
          6282 => x"2e",
          6283 => x"0b",
          6284 => x"81",
          6285 => x"f4",
          6286 => x"34",
          6287 => x"34",
          6288 => x"75",
          6289 => x"d0",
          6290 => x"1a",
          6291 => x"59",
          6292 => x"88",
          6293 => x"75",
          6294 => x"38",
          6295 => x"b8",
          6296 => x"05",
          6297 => x"34",
          6298 => x"56",
          6299 => x"7e",
          6300 => x"57",
          6301 => x"2a",
          6302 => x"33",
          6303 => x"7d",
          6304 => x"51",
          6305 => x"08",
          6306 => x"38",
          6307 => x"17",
          6308 => x"34",
          6309 => x"0b",
          6310 => x"77",
          6311 => x"78",
          6312 => x"83",
          6313 => x"0b",
          6314 => x"83",
          6315 => x"3f",
          6316 => x"ba",
          6317 => x"90",
          6318 => x"74",
          6319 => x"34",
          6320 => x"7a",
          6321 => x"55",
          6322 => x"a0",
          6323 => x"58",
          6324 => x"58",
          6325 => x"5c",
          6326 => x"0b",
          6327 => x"83",
          6328 => x"3f",
          6329 => x"39",
          6330 => x"08",
          6331 => x"9b",
          6332 => x"70",
          6333 => x"81",
          6334 => x"2e",
          6335 => x"fe",
          6336 => x"ab",
          6337 => x"84",
          6338 => x"75",
          6339 => x"04",
          6340 => x"52",
          6341 => x"af",
          6342 => x"ba",
          6343 => x"05",
          6344 => x"7c",
          6345 => x"3d",
          6346 => x"05",
          6347 => x"34",
          6348 => x"3d",
          6349 => x"75",
          6350 => x"81",
          6351 => x"ef",
          6352 => x"ff",
          6353 => x"56",
          6354 => x"6a",
          6355 => x"88",
          6356 => x"0d",
          6357 => x"ff",
          6358 => x"91",
          6359 => x"d0",
          6360 => x"fa",
          6361 => x"70",
          6362 => x"7a",
          6363 => x"81",
          6364 => x"58",
          6365 => x"16",
          6366 => x"9f",
          6367 => x"e0",
          6368 => x"75",
          6369 => x"77",
          6370 => x"ff",
          6371 => x"70",
          6372 => x"58",
          6373 => x"1c",
          6374 => x"fd",
          6375 => x"ff",
          6376 => x"38",
          6377 => x"fe",
          6378 => x"a8",
          6379 => x"84",
          6380 => x"b8",
          6381 => x"81",
          6382 => x"8d",
          6383 => x"84",
          6384 => x"58",
          6385 => x"80",
          6386 => x"81",
          6387 => x"57",
          6388 => x"02",
          6389 => x"8b",
          6390 => x"40",
          6391 => x"57",
          6392 => x"0b",
          6393 => x"84",
          6394 => x"2e",
          6395 => x"2e",
          6396 => x"9a",
          6397 => x"33",
          6398 => x"82",
          6399 => x"fe",
          6400 => x"c7",
          6401 => x"b0",
          6402 => x"2e",
          6403 => x"b4",
          6404 => x"17",
          6405 => x"54",
          6406 => x"33",
          6407 => x"8c",
          6408 => x"81",
          6409 => x"7b",
          6410 => x"bf",
          6411 => x"2e",
          6412 => x"83",
          6413 => x"f2",
          6414 => x"80",
          6415 => x"83",
          6416 => x"90",
          6417 => x"7d",
          6418 => x"34",
          6419 => x"78",
          6420 => x"57",
          6421 => x"74",
          6422 => x"84",
          6423 => x"08",
          6424 => x"19",
          6425 => x"77",
          6426 => x"59",
          6427 => x"81",
          6428 => x"16",
          6429 => x"bd",
          6430 => x"85",
          6431 => x"17",
          6432 => x"19",
          6433 => x"83",
          6434 => x"a5",
          6435 => x"ae",
          6436 => x"ba",
          6437 => x"82",
          6438 => x"74",
          6439 => x"fe",
          6440 => x"84",
          6441 => x"82",
          6442 => x"0d",
          6443 => x"71",
          6444 => x"07",
          6445 => x"ba",
          6446 => x"84",
          6447 => x"38",
          6448 => x"0d",
          6449 => x"7b",
          6450 => x"94",
          6451 => x"7a",
          6452 => x"84",
          6453 => x"16",
          6454 => x"8c",
          6455 => x"27",
          6456 => x"7c",
          6457 => x"38",
          6458 => x"08",
          6459 => x"51",
          6460 => x"fa",
          6461 => x"b8",
          6462 => x"5b",
          6463 => x"ba",
          6464 => x"8c",
          6465 => x"a8",
          6466 => x"5d",
          6467 => x"8e",
          6468 => x"2e",
          6469 => x"54",
          6470 => x"53",
          6471 => x"e0",
          6472 => x"ec",
          6473 => x"02",
          6474 => x"57",
          6475 => x"97",
          6476 => x"ba",
          6477 => x"80",
          6478 => x"0c",
          6479 => x"52",
          6480 => x"d7",
          6481 => x"ba",
          6482 => x"05",
          6483 => x"73",
          6484 => x"09",
          6485 => x"06",
          6486 => x"17",
          6487 => x"34",
          6488 => x"ba",
          6489 => x"3d",
          6490 => x"82",
          6491 => x"3d",
          6492 => x"8c",
          6493 => x"2e",
          6494 => x"96",
          6495 => x"96",
          6496 => x"3f",
          6497 => x"8c",
          6498 => x"33",
          6499 => x"d2",
          6500 => x"22",
          6501 => x"76",
          6502 => x"74",
          6503 => x"77",
          6504 => x"73",
          6505 => x"83",
          6506 => x"3f",
          6507 => x"0c",
          6508 => x"6b",
          6509 => x"cc",
          6510 => x"c5",
          6511 => x"8c",
          6512 => x"07",
          6513 => x"2e",
          6514 => x"56",
          6515 => x"78",
          6516 => x"2e",
          6517 => x"5a",
          6518 => x"7c",
          6519 => x"b4",
          6520 => x"83",
          6521 => x"2e",
          6522 => x"54",
          6523 => x"33",
          6524 => x"8c",
          6525 => x"81",
          6526 => x"78",
          6527 => x"80",
          6528 => x"80",
          6529 => x"a7",
          6530 => x"33",
          6531 => x"88",
          6532 => x"07",
          6533 => x"0c",
          6534 => x"84",
          6535 => x"7c",
          6536 => x"70",
          6537 => x"ba",
          6538 => x"80",
          6539 => x"09",
          6540 => x"34",
          6541 => x"b4",
          6542 => x"81",
          6543 => x"3f",
          6544 => x"2e",
          6545 => x"ba",
          6546 => x"08",
          6547 => x"08",
          6548 => x"fe",
          6549 => x"82",
          6550 => x"77",
          6551 => x"05",
          6552 => x"fe",
          6553 => x"76",
          6554 => x"51",
          6555 => x"08",
          6556 => x"39",
          6557 => x"3f",
          6558 => x"8c",
          6559 => x"08",
          6560 => x"59",
          6561 => x"59",
          6562 => x"59",
          6563 => x"1c",
          6564 => x"2e",
          6565 => x"70",
          6566 => x"ea",
          6567 => x"ba",
          6568 => x"3d",
          6569 => x"ff",
          6570 => x"56",
          6571 => x"8f",
          6572 => x"76",
          6573 => x"55",
          6574 => x"70",
          6575 => x"58",
          6576 => x"a2",
          6577 => x"ff",
          6578 => x"f5",
          6579 => x"ff",
          6580 => x"95",
          6581 => x"08",
          6582 => x"08",
          6583 => x"2e",
          6584 => x"83",
          6585 => x"5b",
          6586 => x"38",
          6587 => x"81",
          6588 => x"57",
          6589 => x"74",
          6590 => x"75",
          6591 => x"38",
          6592 => x"79",
          6593 => x"77",
          6594 => x"74",
          6595 => x"1a",
          6596 => x"34",
          6597 => x"70",
          6598 => x"77",
          6599 => x"33",
          6600 => x"bc",
          6601 => x"b7",
          6602 => x"5c",
          6603 => x"38",
          6604 => x"45",
          6605 => x"52",
          6606 => x"8c",
          6607 => x"2e",
          6608 => x"8c",
          6609 => x"52",
          6610 => x"8c",
          6611 => x"fd",
          6612 => x"8c",
          6613 => x"9c",
          6614 => x"75",
          6615 => x"8c",
          6616 => x"c1",
          6617 => x"8b",
          6618 => x"81",
          6619 => x"58",
          6620 => x"7d",
          6621 => x"51",
          6622 => x"08",
          6623 => x"7a",
          6624 => x"9c",
          6625 => x"09",
          6626 => x"79",
          6627 => x"75",
          6628 => x"3f",
          6629 => x"8c",
          6630 => x"84",
          6631 => x"5c",
          6632 => x"b4",
          6633 => x"18",
          6634 => x"06",
          6635 => x"b8",
          6636 => x"d5",
          6637 => x"2e",
          6638 => x"b4",
          6639 => x"78",
          6640 => x"57",
          6641 => x"74",
          6642 => x"5c",
          6643 => x"1a",
          6644 => x"52",
          6645 => x"ba",
          6646 => x"80",
          6647 => x"84",
          6648 => x"fd",
          6649 => x"76",
          6650 => x"55",
          6651 => x"8b",
          6652 => x"55",
          6653 => x"70",
          6654 => x"74",
          6655 => x"81",
          6656 => x"58",
          6657 => x"fd",
          6658 => x"7d",
          6659 => x"51",
          6660 => x"08",
          6661 => x"df",
          6662 => x"7a",
          6663 => x"ec",
          6664 => x"09",
          6665 => x"8c",
          6666 => x"a8",
          6667 => x"08",
          6668 => x"74",
          6669 => x"08",
          6670 => x"52",
          6671 => x"ba",
          6672 => x"80",
          6673 => x"81",
          6674 => x"e7",
          6675 => x"18",
          6676 => x"52",
          6677 => x"3f",
          6678 => x"62",
          6679 => x"5e",
          6680 => x"9f",
          6681 => x"97",
          6682 => x"8f",
          6683 => x"59",
          6684 => x"80",
          6685 => x"91",
          6686 => x"79",
          6687 => x"08",
          6688 => x"81",
          6689 => x"2e",
          6690 => x"70",
          6691 => x"5c",
          6692 => x"7a",
          6693 => x"2a",
          6694 => x"08",
          6695 => x"78",
          6696 => x"26",
          6697 => x"5b",
          6698 => x"d8",
          6699 => x"9c",
          6700 => x"55",
          6701 => x"dc",
          6702 => x"81",
          6703 => x"c5",
          6704 => x"bb",
          6705 => x"c2",
          6706 => x"ba",
          6707 => x"0b",
          6708 => x"04",
          6709 => x"3f",
          6710 => x"73",
          6711 => x"56",
          6712 => x"8e",
          6713 => x"2e",
          6714 => x"2e",
          6715 => x"7e",
          6716 => x"8c",
          6717 => x"a3",
          6718 => x"59",
          6719 => x"12",
          6720 => x"38",
          6721 => x"0c",
          6722 => x"7b",
          6723 => x"05",
          6724 => x"26",
          6725 => x"16",
          6726 => x"7c",
          6727 => x"39",
          6728 => x"80",
          6729 => x"c5",
          6730 => x"1b",
          6731 => x"08",
          6732 => x"3d",
          6733 => x"33",
          6734 => x"08",
          6735 => x"85",
          6736 => x"33",
          6737 => x"2e",
          6738 => x"ba",
          6739 => x"33",
          6740 => x"75",
          6741 => x"08",
          6742 => x"80",
          6743 => x"11",
          6744 => x"5b",
          6745 => x"a9",
          6746 => x"06",
          6747 => x"7b",
          6748 => x"06",
          6749 => x"9f",
          6750 => x"51",
          6751 => x"08",
          6752 => x"2e",
          6753 => x"26",
          6754 => x"55",
          6755 => x"88",
          6756 => x"38",
          6757 => x"38",
          6758 => x"e7",
          6759 => x"89",
          6760 => x"47",
          6761 => x"65",
          6762 => x"5f",
          6763 => x"80",
          6764 => x"53",
          6765 => x"3f",
          6766 => x"95",
          6767 => x"83",
          6768 => x"59",
          6769 => x"2e",
          6770 => x"90",
          6771 => x"44",
          6772 => x"83",
          6773 => x"33",
          6774 => x"81",
          6775 => x"75",
          6776 => x"11",
          6777 => x"71",
          6778 => x"72",
          6779 => x"5c",
          6780 => x"a3",
          6781 => x"4f",
          6782 => x"80",
          6783 => x"57",
          6784 => x"61",
          6785 => x"63",
          6786 => x"06",
          6787 => x"81",
          6788 => x"6e",
          6789 => x"62",
          6790 => x"38",
          6791 => x"e7",
          6792 => x"9d",
          6793 => x"e7",
          6794 => x"22",
          6795 => x"38",
          6796 => x"78",
          6797 => x"8c",
          6798 => x"8c",
          6799 => x"0b",
          6800 => x"8c",
          6801 => x"05",
          6802 => x"2a",
          6803 => x"7d",
          6804 => x"70",
          6805 => x"44",
          6806 => x"1d",
          6807 => x"31",
          6808 => x"38",
          6809 => x"70",
          6810 => x"3f",
          6811 => x"2e",
          6812 => x"81",
          6813 => x"0b",
          6814 => x"38",
          6815 => x"74",
          6816 => x"5b",
          6817 => x"ba",
          6818 => x"98",
          6819 => x"93",
          6820 => x"0d",
          6821 => x"d0",
          6822 => x"57",
          6823 => x"77",
          6824 => x"77",
          6825 => x"83",
          6826 => x"57",
          6827 => x"76",
          6828 => x"12",
          6829 => x"38",
          6830 => x"44",
          6831 => x"89",
          6832 => x"59",
          6833 => x"47",
          6834 => x"38",
          6835 => x"70",
          6836 => x"07",
          6837 => x"ce",
          6838 => x"83",
          6839 => x"f9",
          6840 => x"81",
          6841 => x"81",
          6842 => x"38",
          6843 => x"8c",
          6844 => x"5f",
          6845 => x"fe",
          6846 => x"fb",
          6847 => x"83",
          6848 => x"3d",
          6849 => x"06",
          6850 => x"f5",
          6851 => x"43",
          6852 => x"9f",
          6853 => x"77",
          6854 => x"f5",
          6855 => x"0c",
          6856 => x"04",
          6857 => x"38",
          6858 => x"81",
          6859 => x"38",
          6860 => x"70",
          6861 => x"74",
          6862 => x"59",
          6863 => x"33",
          6864 => x"15",
          6865 => x"45",
          6866 => x"34",
          6867 => x"ff",
          6868 => x"34",
          6869 => x"05",
          6870 => x"83",
          6871 => x"91",
          6872 => x"49",
          6873 => x"75",
          6874 => x"75",
          6875 => x"93",
          6876 => x"61",
          6877 => x"34",
          6878 => x"99",
          6879 => x"80",
          6880 => x"05",
          6881 => x"9d",
          6882 => x"61",
          6883 => x"ba",
          6884 => x"9f",
          6885 => x"38",
          6886 => x"a8",
          6887 => x"80",
          6888 => x"ff",
          6889 => x"34",
          6890 => x"05",
          6891 => x"a9",
          6892 => x"05",
          6893 => x"70",
          6894 => x"05",
          6895 => x"38",
          6896 => x"69",
          6897 => x"aa",
          6898 => x"52",
          6899 => x"57",
          6900 => x"60",
          6901 => x"38",
          6902 => x"81",
          6903 => x"f4",
          6904 => x"2e",
          6905 => x"57",
          6906 => x"76",
          6907 => x"55",
          6908 => x"76",
          6909 => x"05",
          6910 => x"64",
          6911 => x"26",
          6912 => x"53",
          6913 => x"3f",
          6914 => x"84",
          6915 => x"81",
          6916 => x"f4",
          6917 => x"5b",
          6918 => x"7f",
          6919 => x"62",
          6920 => x"55",
          6921 => x"74",
          6922 => x"fe",
          6923 => x"85",
          6924 => x"57",
          6925 => x"83",
          6926 => x"ff",
          6927 => x"82",
          6928 => x"c1",
          6929 => x"7d",
          6930 => x"59",
          6931 => x"ff",
          6932 => x"69",
          6933 => x"be",
          6934 => x"81",
          6935 => x"78",
          6936 => x"05",
          6937 => x"62",
          6938 => x"67",
          6939 => x"82",
          6940 => x"05",
          6941 => x"05",
          6942 => x"67",
          6943 => x"83",
          6944 => x"61",
          6945 => x"ca",
          6946 => x"61",
          6947 => x"58",
          6948 => x"98",
          6949 => x"34",
          6950 => x"51",
          6951 => x"ba",
          6952 => x"80",
          6953 => x"81",
          6954 => x"38",
          6955 => x"0c",
          6956 => x"04",
          6957 => x"64",
          6958 => x"ae",
          6959 => x"83",
          6960 => x"2e",
          6961 => x"83",
          6962 => x"70",
          6963 => x"86",
          6964 => x"52",
          6965 => x"ba",
          6966 => x"70",
          6967 => x"0b",
          6968 => x"05",
          6969 => x"27",
          6970 => x"39",
          6971 => x"26",
          6972 => x"77",
          6973 => x"8e",
          6974 => x"44",
          6975 => x"43",
          6976 => x"34",
          6977 => x"05",
          6978 => x"a2",
          6979 => x"61",
          6980 => x"61",
          6981 => x"c4",
          6982 => x"34",
          6983 => x"7c",
          6984 => x"5c",
          6985 => x"2a",
          6986 => x"98",
          6987 => x"82",
          6988 => x"05",
          6989 => x"61",
          6990 => x"34",
          6991 => x"b2",
          6992 => x"ff",
          6993 => x"61",
          6994 => x"c7",
          6995 => x"76",
          6996 => x"81",
          6997 => x"80",
          6998 => x"05",
          6999 => x"34",
          7000 => x"b8",
          7001 => x"79",
          7002 => x"84",
          7003 => x"90",
          7004 => x"b2",
          7005 => x"08",
          7006 => x"b4",
          7007 => x"ba",
          7008 => x"98",
          7009 => x"ff",
          7010 => x"6a",
          7011 => x"34",
          7012 => x"85",
          7013 => x"ff",
          7014 => x"05",
          7015 => x"61",
          7016 => x"57",
          7017 => x"53",
          7018 => x"3f",
          7019 => x"70",
          7020 => x"76",
          7021 => x"70",
          7022 => x"d2",
          7023 => x"e1",
          7024 => x"c1",
          7025 => x"05",
          7026 => x"34",
          7027 => x"80",
          7028 => x"ff",
          7029 => x"34",
          7030 => x"e9",
          7031 => x"61",
          7032 => x"40",
          7033 => x"61",
          7034 => x"ed",
          7035 => x"34",
          7036 => x"d5",
          7037 => x"54",
          7038 => x"fe",
          7039 => x"53",
          7040 => x"3f",
          7041 => x"f4",
          7042 => x"7b",
          7043 => x"78",
          7044 => x"3d",
          7045 => x"79",
          7046 => x"2e",
          7047 => x"33",
          7048 => x"76",
          7049 => x"57",
          7050 => x"24",
          7051 => x"76",
          7052 => x"8c",
          7053 => x"0d",
          7054 => x"59",
          7055 => x"84",
          7056 => x"38",
          7057 => x"56",
          7058 => x"74",
          7059 => x"0c",
          7060 => x"0d",
          7061 => x"53",
          7062 => x"9e",
          7063 => x"70",
          7064 => x"1b",
          7065 => x"56",
          7066 => x"ff",
          7067 => x"0d",
          7068 => x"58",
          7069 => x"76",
          7070 => x"55",
          7071 => x"0c",
          7072 => x"56",
          7073 => x"77",
          7074 => x"34",
          7075 => x"38",
          7076 => x"18",
          7077 => x"38",
          7078 => x"54",
          7079 => x"9d",
          7080 => x"38",
          7081 => x"84",
          7082 => x"9f",
          7083 => x"c0",
          7084 => x"a2",
          7085 => x"72",
          7086 => x"56",
          7087 => x"51",
          7088 => x"84",
          7089 => x"fd",
          7090 => x"05",
          7091 => x"ff",
          7092 => x"06",
          7093 => x"3d",
          7094 => x"54",
          7095 => x"e9",
          7096 => x"e7",
          7097 => x"38",
          7098 => x"53",
          7099 => x"71",
          7100 => x"51",
          7101 => x"81",
          7102 => x"85",
          7103 => x"92",
          7104 => x"22",
          7105 => x"26",
          7106 => x"8c",
          7107 => x"b5",
          7108 => x"81",
          7109 => x"e5",
          7110 => x"0c",
          7111 => x"0d",
          7112 => x"80",
          7113 => x"83",
          7114 => x"26",
          7115 => x"56",
          7116 => x"73",
          7117 => x"70",
          7118 => x"22",
          7119 => x"ff",
          7120 => x"24",
          7121 => x"15",
          7122 => x"73",
          7123 => x"07",
          7124 => x"38",
          7125 => x"87",
          7126 => x"ff",
          7127 => x"71",
          7128 => x"73",
          7129 => x"ff",
          7130 => x"39",
          7131 => x"06",
          7132 => x"83",
          7133 => x"e6",
          7134 => x"51",
          7135 => x"ff",
          7136 => x"70",
          7137 => x"39",
          7138 => x"57",
          7139 => x"81",
          7140 => x"ff",
          7141 => x"75",
          7142 => x"52",
          7143 => x"ff",
          7144 => x"00",
          7145 => x"19",
          7146 => x"19",
          7147 => x"19",
          7148 => x"19",
          7149 => x"19",
          7150 => x"19",
          7151 => x"19",
          7152 => x"18",
          7153 => x"18",
          7154 => x"18",
          7155 => x"1e",
          7156 => x"1f",
          7157 => x"1f",
          7158 => x"1f",
          7159 => x"1f",
          7160 => x"1f",
          7161 => x"1f",
          7162 => x"1f",
          7163 => x"1f",
          7164 => x"1f",
          7165 => x"1f",
          7166 => x"1f",
          7167 => x"1f",
          7168 => x"1f",
          7169 => x"1f",
          7170 => x"1f",
          7171 => x"1f",
          7172 => x"1f",
          7173 => x"1f",
          7174 => x"1f",
          7175 => x"1f",
          7176 => x"1f",
          7177 => x"1f",
          7178 => x"1f",
          7179 => x"1f",
          7180 => x"1f",
          7181 => x"1f",
          7182 => x"1f",
          7183 => x"1f",
          7184 => x"1f",
          7185 => x"24",
          7186 => x"1f",
          7187 => x"24",
          7188 => x"22",
          7189 => x"1f",
          7190 => x"1f",
          7191 => x"1f",
          7192 => x"1f",
          7193 => x"1f",
          7194 => x"1f",
          7195 => x"1f",
          7196 => x"1f",
          7197 => x"1f",
          7198 => x"1f",
          7199 => x"1f",
          7200 => x"1f",
          7201 => x"1f",
          7202 => x"1f",
          7203 => x"1f",
          7204 => x"1f",
          7205 => x"1f",
          7206 => x"1f",
          7207 => x"1f",
          7208 => x"1f",
          7209 => x"1f",
          7210 => x"1f",
          7211 => x"1f",
          7212 => x"1f",
          7213 => x"1f",
          7214 => x"1f",
          7215 => x"21",
          7216 => x"1f",
          7217 => x"1f",
          7218 => x"1f",
          7219 => x"1f",
          7220 => x"21",
          7221 => x"1f",
          7222 => x"1f",
          7223 => x"21",
          7224 => x"32",
          7225 => x"32",
          7226 => x"32",
          7227 => x"3b",
          7228 => x"38",
          7229 => x"3a",
          7230 => x"37",
          7231 => x"39",
          7232 => x"37",
          7233 => x"34",
          7234 => x"38",
          7235 => x"34",
          7236 => x"37",
          7237 => x"36",
          7238 => x"46",
          7239 => x"46",
          7240 => x"46",
          7241 => x"46",
          7242 => x"47",
          7243 => x"47",
          7244 => x"47",
          7245 => x"47",
          7246 => x"47",
          7247 => x"47",
          7248 => x"47",
          7249 => x"47",
          7250 => x"47",
          7251 => x"47",
          7252 => x"47",
          7253 => x"47",
          7254 => x"47",
          7255 => x"47",
          7256 => x"47",
          7257 => x"48",
          7258 => x"48",
          7259 => x"48",
          7260 => x"47",
          7261 => x"47",
          7262 => x"48",
          7263 => x"47",
          7264 => x"47",
          7265 => x"47",
          7266 => x"47",
          7267 => x"55",
          7268 => x"54",
          7269 => x"54",
          7270 => x"55",
          7271 => x"55",
          7272 => x"52",
          7273 => x"52",
          7274 => x"52",
          7275 => x"55",
          7276 => x"56",
          7277 => x"52",
          7278 => x"52",
          7279 => x"52",
          7280 => x"52",
          7281 => x"52",
          7282 => x"52",
          7283 => x"52",
          7284 => x"52",
          7285 => x"52",
          7286 => x"55",
          7287 => x"52",
          7288 => x"54",
          7289 => x"53",
          7290 => x"52",
          7291 => x"52",
          7292 => x"52",
          7293 => x"59",
          7294 => x"59",
          7295 => x"59",
          7296 => x"59",
          7297 => x"59",
          7298 => x"59",
          7299 => x"59",
          7300 => x"59",
          7301 => x"59",
          7302 => x"59",
          7303 => x"59",
          7304 => x"59",
          7305 => x"59",
          7306 => x"59",
          7307 => x"59",
          7308 => x"59",
          7309 => x"59",
          7310 => x"59",
          7311 => x"5a",
          7312 => x"59",
          7313 => x"5a",
          7314 => x"5a",
          7315 => x"59",
          7316 => x"59",
          7317 => x"59",
          7318 => x"63",
          7319 => x"61",
          7320 => x"61",
          7321 => x"61",
          7322 => x"61",
          7323 => x"61",
          7324 => x"61",
          7325 => x"5e",
          7326 => x"61",
          7327 => x"61",
          7328 => x"61",
          7329 => x"61",
          7330 => x"63",
          7331 => x"63",
          7332 => x"63",
          7333 => x"df",
          7334 => x"df",
          7335 => x"de",
          7336 => x"de",
          7337 => x"0e",
          7338 => x"0b",
          7339 => x"0b",
          7340 => x"0b",
          7341 => x"0b",
          7342 => x"0b",
          7343 => x"0b",
          7344 => x"0f",
          7345 => x"0b",
          7346 => x"0b",
          7347 => x"0b",
          7348 => x"0b",
          7349 => x"0b",
          7350 => x"0b",
          7351 => x"0b",
          7352 => x"0b",
          7353 => x"0b",
          7354 => x"0b",
          7355 => x"0b",
          7356 => x"0b",
          7357 => x"0b",
          7358 => x"0b",
          7359 => x"0b",
          7360 => x"0b",
          7361 => x"0b",
          7362 => x"0b",
          7363 => x"0b",
          7364 => x"0b",
          7365 => x"0e",
          7366 => x"0b",
          7367 => x"0b",
          7368 => x"0b",
          7369 => x"0b",
          7370 => x"0b",
          7371 => x"0e",
          7372 => x"0e",
          7373 => x"0b",
          7374 => x"0b",
          7375 => x"0e",
          7376 => x"0b",
          7377 => x"0e",
          7378 => x"0b",
          7379 => x"0b",
          7380 => x"0b",
          7381 => x"0e",
          7382 => x"00",
          7383 => x"00",
          7384 => x"00",
          7385 => x"00",
          7386 => x"00",
          7387 => x"00",
          7388 => x"00",
          7389 => x"00",
          7390 => x"00",
          7391 => x"68",
          7392 => x"64",
          7393 => x"64",
          7394 => x"6c",
          7395 => x"70",
          7396 => x"74",
          7397 => x"00",
          7398 => x"00",
          7399 => x"00",
          7400 => x"30",
          7401 => x"00",
          7402 => x"00",
          7403 => x"00",
          7404 => x"6b",
          7405 => x"72",
          7406 => x"72",
          7407 => x"20",
          7408 => x"63",
          7409 => x"6f",
          7410 => x"70",
          7411 => x"73",
          7412 => x"73",
          7413 => x"6e",
          7414 => x"79",
          7415 => x"6c",
          7416 => x"63",
          7417 => x"6d",
          7418 => x"70",
          7419 => x"20",
          7420 => x"65",
          7421 => x"72",
          7422 => x"72",
          7423 => x"20",
          7424 => x"62",
          7425 => x"73",
          7426 => x"6f",
          7427 => x"64",
          7428 => x"73",
          7429 => x"6e",
          7430 => x"00",
          7431 => x"6e",
          7432 => x"73",
          7433 => x"64",
          7434 => x"20",
          7435 => x"65",
          7436 => x"74",
          7437 => x"6c",
          7438 => x"65",
          7439 => x"64",
          7440 => x"6c",
          7441 => x"64",
          7442 => x"73",
          7443 => x"63",
          7444 => x"69",
          7445 => x"76",
          7446 => x"6c",
          7447 => x"00",
          7448 => x"68",
          7449 => x"00",
          7450 => x"65",
          7451 => x"00",
          7452 => x"6f",
          7453 => x"2e",
          7454 => x"61",
          7455 => x"2e",
          7456 => x"72",
          7457 => x"63",
          7458 => x"00",
          7459 => x"79",
          7460 => x"61",
          7461 => x"79",
          7462 => x"2e",
          7463 => x"61",
          7464 => x"38",
          7465 => x"20",
          7466 => x"00",
          7467 => x"00",
          7468 => x"34",
          7469 => x"20",
          7470 => x"00",
          7471 => x"20",
          7472 => x"2f",
          7473 => x"00",
          7474 => x"00",
          7475 => x"72",
          7476 => x"29",
          7477 => x"2a",
          7478 => x"55",
          7479 => x"75",
          7480 => x"6c",
          7481 => x"52",
          7482 => x"6e",
          7483 => x"00",
          7484 => x"52",
          7485 => x"72",
          7486 => x"52",
          7487 => x"6e",
          7488 => x"00",
          7489 => x"52",
          7490 => x"72",
          7491 => x"43",
          7492 => x"6e",
          7493 => x"00",
          7494 => x"52",
          7495 => x"72",
          7496 => x"32",
          7497 => x"75",
          7498 => x"6d",
          7499 => x"72",
          7500 => x"74",
          7501 => x"20",
          7502 => x"2e",
          7503 => x"6e",
          7504 => x"2e",
          7505 => x"74",
          7506 => x"61",
          7507 => x"53",
          7508 => x"74",
          7509 => x"20",
          7510 => x"69",
          7511 => x"64",
          7512 => x"2c",
          7513 => x"20",
          7514 => x"6e",
          7515 => x"00",
          7516 => x"3a",
          7517 => x"73",
          7518 => x"61",
          7519 => x"00",
          7520 => x"64",
          7521 => x"64",
          7522 => x"55",
          7523 => x"3a",
          7524 => x"25",
          7525 => x"6c",
          7526 => x"74",
          7527 => x"00",
          7528 => x"74",
          7529 => x"6c",
          7530 => x"2e",
          7531 => x"6c",
          7532 => x"64",
          7533 => x"6c",
          7534 => x"00",
          7535 => x"65",
          7536 => x"63",
          7537 => x"29",
          7538 => x"65",
          7539 => x"63",
          7540 => x"30",
          7541 => x"0a",
          7542 => x"25",
          7543 => x"00",
          7544 => x"25",
          7545 => x"6d",
          7546 => x"2e",
          7547 => x"38",
          7548 => x"29",
          7549 => x"28",
          7550 => x"00",
          7551 => x"67",
          7552 => x"38",
          7553 => x"2d",
          7554 => x"6e",
          7555 => x"00",
          7556 => x"65",
          7557 => x"6f",
          7558 => x"00",
          7559 => x"5c",
          7560 => x"6d",
          7561 => x"61",
          7562 => x"63",
          7563 => x"72",
          7564 => x"6f",
          7565 => x"00",
          7566 => x"2f",
          7567 => x"64",
          7568 => x"25",
          7569 => x"43",
          7570 => x"75",
          7571 => x"00",
          7572 => x"63",
          7573 => x"65",
          7574 => x"00",
          7575 => x"73",
          7576 => x"20",
          7577 => x"73",
          7578 => x"6f",
          7579 => x"73",
          7580 => x"58",
          7581 => x"20",
          7582 => x"6d",
          7583 => x"72",
          7584 => x"73",
          7585 => x"58",
          7586 => x"20",
          7587 => x"53",
          7588 => x"64",
          7589 => x"20",
          7590 => x"58",
          7591 => x"73",
          7592 => x"20",
          7593 => x"20",
          7594 => x"20",
          7595 => x"20",
          7596 => x"58",
          7597 => x"20",
          7598 => x"20",
          7599 => x"72",
          7600 => x"20",
          7601 => x"25",
          7602 => x"00",
          7603 => x"73",
          7604 => x"44",
          7605 => x"63",
          7606 => x"20",
          7607 => x"4d",
          7608 => x"20",
          7609 => x"43",
          7610 => x"65",
          7611 => x"20",
          7612 => x"25",
          7613 => x"00",
          7614 => x"49",
          7615 => x"32",
          7616 => x"43",
          7617 => x"20",
          7618 => x"00",
          7619 => x"53",
          7620 => x"55",
          7621 => x"20",
          7622 => x"54",
          7623 => x"6e",
          7624 => x"32",
          7625 => x"20",
          7626 => x"20",
          7627 => x"65",
          7628 => x"32",
          7629 => x"20",
          7630 => x"44",
          7631 => x"69",
          7632 => x"32",
          7633 => x"20",
          7634 => x"20",
          7635 => x"58",
          7636 => x"0a",
          7637 => x"41",
          7638 => x"28",
          7639 => x"38",
          7640 => x"20",
          7641 => x"52",
          7642 => x"58",
          7643 => x"0a",
          7644 => x"52",
          7645 => x"28",
          7646 => x"38",
          7647 => x"20",
          7648 => x"41",
          7649 => x"58",
          7650 => x"0a",
          7651 => x"20",
          7652 => x"66",
          7653 => x"6b",
          7654 => x"4f",
          7655 => x"61",
          7656 => x"64",
          7657 => x"65",
          7658 => x"4f",
          7659 => x"00",
          7660 => x"f0",
          7661 => x"00",
          7662 => x"00",
          7663 => x"f0",
          7664 => x"00",
          7665 => x"00",
          7666 => x"f0",
          7667 => x"00",
          7668 => x"00",
          7669 => x"f0",
          7670 => x"00",
          7671 => x"00",
          7672 => x"f0",
          7673 => x"00",
          7674 => x"00",
          7675 => x"f0",
          7676 => x"00",
          7677 => x"00",
          7678 => x"f0",
          7679 => x"00",
          7680 => x"00",
          7681 => x"f0",
          7682 => x"00",
          7683 => x"00",
          7684 => x"f0",
          7685 => x"00",
          7686 => x"00",
          7687 => x"f0",
          7688 => x"00",
          7689 => x"00",
          7690 => x"f0",
          7691 => x"00",
          7692 => x"43",
          7693 => x"41",
          7694 => x"35",
          7695 => x"46",
          7696 => x"32",
          7697 => x"00",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"00",
          7703 => x"20",
          7704 => x"65",
          7705 => x"74",
          7706 => x"65",
          7707 => x"6c",
          7708 => x"73",
          7709 => x"73",
          7710 => x"00",
          7711 => x"20",
          7712 => x"69",
          7713 => x"72",
          7714 => x"65",
          7715 => x"79",
          7716 => x"6f",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"42",
          7721 => x"44",
          7722 => x"00",
          7723 => x"00",
          7724 => x"00",
          7725 => x"00",
          7726 => x"00",
          7727 => x"00",
          7728 => x"00",
          7729 => x"00",
          7730 => x"00",
          7731 => x"00",
          7732 => x"00",
          7733 => x"00",
          7734 => x"35",
          7735 => x"36",
          7736 => x"25",
          7737 => x"2c",
          7738 => x"64",
          7739 => x"00",
          7740 => x"64",
          7741 => x"25",
          7742 => x"3a",
          7743 => x"25",
          7744 => x"32",
          7745 => x"5b",
          7746 => x"00",
          7747 => x"20",
          7748 => x"00",
          7749 => x"78",
          7750 => x"00",
          7751 => x"78",
          7752 => x"00",
          7753 => x"78",
          7754 => x"64",
          7755 => x"53",
          7756 => x"00",
          7757 => x"69",
          7758 => x"65",
          7759 => x"64",
          7760 => x"53",
          7761 => x"00",
          7762 => x"74",
          7763 => x"64",
          7764 => x"00",
          7765 => x"7c",
          7766 => x"3b",
          7767 => x"54",
          7768 => x"00",
          7769 => x"4f",
          7770 => x"20",
          7771 => x"20",
          7772 => x"20",
          7773 => x"45",
          7774 => x"33",
          7775 => x"f2",
          7776 => x"00",
          7777 => x"05",
          7778 => x"18",
          7779 => x"45",
          7780 => x"45",
          7781 => x"92",
          7782 => x"9a",
          7783 => x"4f",
          7784 => x"aa",
          7785 => x"b2",
          7786 => x"ba",
          7787 => x"c2",
          7788 => x"ca",
          7789 => x"d2",
          7790 => x"da",
          7791 => x"e2",
          7792 => x"ea",
          7793 => x"f2",
          7794 => x"fa",
          7795 => x"2c",
          7796 => x"2a",
          7797 => x"00",
          7798 => x"00",
          7799 => x"00",
          7800 => x"00",
          7801 => x"00",
          7802 => x"00",
          7803 => x"00",
          7804 => x"00",
          7805 => x"00",
          7806 => x"00",
          7807 => x"00",
          7808 => x"00",
          7809 => x"01",
          7810 => x"00",
          7811 => x"00",
          7812 => x"00",
          7813 => x"00",
          7814 => x"25",
          7815 => x"25",
          7816 => x"25",
          7817 => x"25",
          7818 => x"25",
          7819 => x"25",
          7820 => x"25",
          7821 => x"25",
          7822 => x"25",
          7823 => x"25",
          7824 => x"25",
          7825 => x"25",
          7826 => x"03",
          7827 => x"03",
          7828 => x"03",
          7829 => x"22",
          7830 => x"22",
          7831 => x"22",
          7832 => x"22",
          7833 => x"00",
          7834 => x"03",
          7835 => x"00",
          7836 => x"01",
          7837 => x"01",
          7838 => x"01",
          7839 => x"01",
          7840 => x"01",
          7841 => x"01",
          7842 => x"01",
          7843 => x"01",
          7844 => x"01",
          7845 => x"02",
          7846 => x"02",
          7847 => x"01",
          7848 => x"01",
          7849 => x"01",
          7850 => x"01",
          7851 => x"01",
          7852 => x"01",
          7853 => x"01",
          7854 => x"01",
          7855 => x"01",
          7856 => x"01",
          7857 => x"01",
          7858 => x"01",
          7859 => x"01",
          7860 => x"01",
          7861 => x"01",
          7862 => x"00",
          7863 => x"02",
          7864 => x"02",
          7865 => x"02",
          7866 => x"02",
          7867 => x"01",
          7868 => x"02",
          7869 => x"02",
          7870 => x"02",
          7871 => x"01",
          7872 => x"02",
          7873 => x"02",
          7874 => x"01",
          7875 => x"02",
          7876 => x"2c",
          7877 => x"02",
          7878 => x"02",
          7879 => x"02",
          7880 => x"02",
          7881 => x"02",
          7882 => x"03",
          7883 => x"00",
          7884 => x"03",
          7885 => x"00",
          7886 => x"03",
          7887 => x"03",
          7888 => x"03",
          7889 => x"03",
          7890 => x"03",
          7891 => x"04",
          7892 => x"04",
          7893 => x"04",
          7894 => x"04",
          7895 => x"04",
          7896 => x"00",
          7897 => x"1e",
          7898 => x"1f",
          7899 => x"1f",
          7900 => x"1f",
          7901 => x"1f",
          7902 => x"1f",
          7903 => x"00",
          7904 => x"1f",
          7905 => x"1f",
          7906 => x"1f",
          7907 => x"06",
          7908 => x"06",
          7909 => x"1f",
          7910 => x"00",
          7911 => x"1f",
          7912 => x"1f",
          7913 => x"21",
          7914 => x"02",
          7915 => x"24",
          7916 => x"2c",
          7917 => x"2c",
          7918 => x"2d",
          7919 => x"00",
          7920 => x"e6",
          7921 => x"00",
          7922 => x"e6",
          7923 => x"00",
          7924 => x"e6",
          7925 => x"00",
          7926 => x"e6",
          7927 => x"00",
          7928 => x"e6",
          7929 => x"00",
          7930 => x"e6",
          7931 => x"00",
          7932 => x"e6",
          7933 => x"00",
          7934 => x"e6",
          7935 => x"00",
          7936 => x"e6",
          7937 => x"00",
          7938 => x"e6",
          7939 => x"00",
          7940 => x"e6",
          7941 => x"00",
          7942 => x"e7",
          7943 => x"00",
          7944 => x"e7",
          7945 => x"00",
          7946 => x"e7",
          7947 => x"00",
          7948 => x"e7",
          7949 => x"00",
          7950 => x"e7",
          7951 => x"00",
          7952 => x"e7",
          7953 => x"00",
          7954 => x"e7",
          7955 => x"00",
          7956 => x"e7",
          7957 => x"00",
          7958 => x"e7",
          7959 => x"00",
          7960 => x"e7",
          7961 => x"00",
          7962 => x"e7",
          7963 => x"00",
          7964 => x"e7",
          7965 => x"00",
          7966 => x"e7",
          7967 => x"00",
          7968 => x"e7",
          7969 => x"00",
          7970 => x"e7",
          7971 => x"00",
          7972 => x"e7",
          7973 => x"00",
          7974 => x"e7",
          7975 => x"00",
          7976 => x"00",
          7977 => x"7f",
          7978 => x"7f",
          7979 => x"7f",
          7980 => x"00",
          7981 => x"ff",
          7982 => x"00",
          7983 => x"00",
          7984 => x"e1",
          7985 => x"00",
          7986 => x"01",
          7987 => x"00",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"00",
          7996 => x"00",
          7997 => x"00",
          7998 => x"00",
          7999 => x"00",
          8000 => x"00",
          8001 => x"00",
          8002 => x"00",
          8003 => x"5f",
          8004 => x"40",
          8005 => x"73",
          8006 => x"6b",
          8007 => x"63",
          8008 => x"33",
          8009 => x"2d",
          8010 => x"f3",
          8011 => x"f0",
          8012 => x"82",
          8013 => x"58",
          8014 => x"40",
          8015 => x"53",
          8016 => x"4b",
          8017 => x"43",
          8018 => x"33",
          8019 => x"2d",
          8020 => x"f3",
          8021 => x"f0",
          8022 => x"82",
          8023 => x"58",
          8024 => x"60",
          8025 => x"53",
          8026 => x"4b",
          8027 => x"43",
          8028 => x"23",
          8029 => x"3d",
          8030 => x"e0",
          8031 => x"f0",
          8032 => x"87",
          8033 => x"1e",
          8034 => x"00",
          8035 => x"13",
          8036 => x"0b",
          8037 => x"03",
          8038 => x"f0",
          8039 => x"f0",
          8040 => x"f0",
          8041 => x"f0",
          8042 => x"82",
          8043 => x"cf",
          8044 => x"d7",
          8045 => x"41",
          8046 => x"6c",
          8047 => x"d9",
          8048 => x"7e",
          8049 => x"d1",
          8050 => x"c2",
          8051 => x"f0",
          8052 => x"82",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"f1",
          8068 => x"f1",
          8069 => x"f1",
          8070 => x"f1",
          8071 => x"f1",
          8072 => x"f1",
          8073 => x"f1",
          8074 => x"f1",
          8075 => x"f1",
          8076 => x"f1",
          8077 => x"f1",
          8078 => x"f1",
          8079 => x"f1",
          8080 => x"f1",
          8081 => x"f1",
          8082 => x"f1",
          8083 => x"f1",
          8084 => x"f1",
          8085 => x"f1",
          8086 => x"f1",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"32",
          9088 => x"00",
          9089 => x"f6",
          9090 => x"fe",
          9091 => x"c6",
          9092 => x"ef",
          9093 => x"66",
          9094 => x"2e",
          9095 => x"26",
          9096 => x"57",
          9097 => x"06",
          9098 => x"0e",
          9099 => x"16",
          9100 => x"be",
          9101 => x"86",
          9102 => x"8e",
          9103 => x"96",
          9104 => x"a5",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"00",
          9113 => x"00",
          9114 => x"00",
          9115 => x"00",
          9116 => x"00",
          9117 => x"00",
          9118 => x"00",
          9119 => x"00",
          9120 => x"01",
          9121 => x"01",
        others => X"00"
    );

    shared variable RAM6 : ramArray :=
    (
             0 => x"0d",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"83",
             9 => x"2b",
            10 => x"00",
            11 => x"00",
            12 => x"ff",
            13 => x"82",
            14 => x"83",
            15 => x"a5",
            16 => x"05",
            17 => x"09",
            18 => x"51",
            19 => x"00",
            20 => x"2e",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"10",
            26 => x"0a",
            27 => x"00",
            28 => x"2e",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"04",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"53",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"81",
            45 => x"04",
            46 => x"00",
            47 => x"00",
            48 => x"9f",
            49 => x"06",
            50 => x"00",
            51 => x"00",
            52 => x"06",
            53 => x"05",
            54 => x"06",
            55 => x"00",
            56 => x"05",
            57 => x"81",
            58 => x"00",
            59 => x"00",
            60 => x"05",
            61 => x"09",
            62 => x"00",
            63 => x"00",
            64 => x"04",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"05",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"73",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"83",
            77 => x"10",
            78 => x"00",
            79 => x"00",
            80 => x"0b",
            81 => x"10",
            82 => x"b5",
            83 => x"00",
            84 => x"08",
            85 => x"2d",
            86 => x"8c",
            87 => x"00",
            88 => x"08",
            89 => x"2d",
            90 => x"8c",
            91 => x"00",
            92 => x"09",
            93 => x"54",
            94 => x"ff",
            95 => x"00",
            96 => x"09",
            97 => x"70",
            98 => x"05",
            99 => x"04",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"10",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"04",
           133 => x"0b",
           134 => x"8c",
           135 => x"04",
           136 => x"0b",
           137 => x"8c",
           138 => x"04",
           139 => x"0b",
           140 => x"8d",
           141 => x"04",
           142 => x"0b",
           143 => x"8d",
           144 => x"04",
           145 => x"0b",
           146 => x"8e",
           147 => x"04",
           148 => x"0b",
           149 => x"8e",
           150 => x"04",
           151 => x"0b",
           152 => x"8f",
           153 => x"04",
           154 => x"0b",
           155 => x"8f",
           156 => x"04",
           157 => x"0b",
           158 => x"90",
           159 => x"04",
           160 => x"0b",
           161 => x"91",
           162 => x"04",
           163 => x"0b",
           164 => x"91",
           165 => x"04",
           166 => x"0b",
           167 => x"92",
           168 => x"04",
           169 => x"0b",
           170 => x"92",
           171 => x"04",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"84",
           193 => x"84",
           194 => x"04",
           195 => x"84",
           196 => x"04",
           197 => x"84",
           198 => x"04",
           199 => x"84",
           200 => x"04",
           201 => x"84",
           202 => x"04",
           203 => x"84",
           204 => x"04",
           205 => x"84",
           206 => x"04",
           207 => x"84",
           208 => x"04",
           209 => x"84",
           210 => x"04",
           211 => x"84",
           212 => x"04",
           213 => x"84",
           214 => x"04",
           215 => x"84",
           216 => x"04",
           217 => x"2d",
           218 => x"90",
           219 => x"c0",
           220 => x"80",
           221 => x"d2",
           222 => x"c0",
           223 => x"80",
           224 => x"80",
           225 => x"0c",
           226 => x"08",
           227 => x"98",
           228 => x"98",
           229 => x"ba",
           230 => x"ba",
           231 => x"84",
           232 => x"84",
           233 => x"04",
           234 => x"2d",
           235 => x"90",
           236 => x"ee",
           237 => x"80",
           238 => x"df",
           239 => x"c0",
           240 => x"82",
           241 => x"80",
           242 => x"0c",
           243 => x"08",
           244 => x"98",
           245 => x"98",
           246 => x"ba",
           247 => x"ba",
           248 => x"84",
           249 => x"84",
           250 => x"04",
           251 => x"2d",
           252 => x"90",
           253 => x"86",
           254 => x"80",
           255 => x"94",
           256 => x"c0",
           257 => x"83",
           258 => x"80",
           259 => x"0c",
           260 => x"08",
           261 => x"98",
           262 => x"98",
           263 => x"ba",
           264 => x"ba",
           265 => x"84",
           266 => x"84",
           267 => x"04",
           268 => x"2d",
           269 => x"90",
           270 => x"c0",
           271 => x"80",
           272 => x"a1",
           273 => x"c0",
           274 => x"82",
           275 => x"80",
           276 => x"0c",
           277 => x"08",
           278 => x"98",
           279 => x"98",
           280 => x"ba",
           281 => x"ba",
           282 => x"84",
           283 => x"84",
           284 => x"04",
           285 => x"2d",
           286 => x"90",
           287 => x"aa",
           288 => x"80",
           289 => x"d0",
           290 => x"c0",
           291 => x"80",
           292 => x"80",
           293 => x"0c",
           294 => x"08",
           295 => x"98",
           296 => x"08",
           297 => x"98",
           298 => x"98",
           299 => x"ba",
           300 => x"ba",
           301 => x"84",
           302 => x"84",
           303 => x"04",
           304 => x"2d",
           305 => x"90",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"73",
           311 => x"81",
           312 => x"07",
           313 => x"72",
           314 => x"09",
           315 => x"0a",
           316 => x"51",
           317 => x"84",
           318 => x"70",
           319 => x"93",
           320 => x"c4",
           321 => x"70",
           322 => x"74",
           323 => x"c5",
           324 => x"0d",
           325 => x"32",
           326 => x"58",
           327 => x"09",
           328 => x"77",
           329 => x"07",
           330 => x"80",
           331 => x"b2",
           332 => x"ba",
           333 => x"ff",
           334 => x"75",
           335 => x"73",
           336 => x"9f",
           337 => x"24",
           338 => x"71",
           339 => x"04",
           340 => x"3d",
           341 => x"86",
           342 => x"56",
           343 => x"53",
           344 => x"9d",
           345 => x"8d",
           346 => x"3d",
           347 => x"85",
           348 => x"0d",
           349 => x"70",
           350 => x"81",
           351 => x"5b",
           352 => x"06",
           353 => x"7b",
           354 => x"81",
           355 => x"81",
           356 => x"81",
           357 => x"70",
           358 => x"38",
           359 => x"2a",
           360 => x"7e",
           361 => x"07",
           362 => x"38",
           363 => x"8c",
           364 => x"2a",
           365 => x"05",
           366 => x"70",
           367 => x"70",
           368 => x"80",
           369 => x"06",
           370 => x"33",
           371 => x"b8",
           372 => x"93",
           373 => x"8a",
           374 => x"38",
           375 => x"8b",
           376 => x"cc",
           377 => x"70",
           378 => x"81",
           379 => x"38",
           380 => x"97",
           381 => x"05",
           382 => x"54",
           383 => x"7c",
           384 => x"7c",
           385 => x"fe",
           386 => x"39",
           387 => x"08",
           388 => x"41",
           389 => x"75",
           390 => x"08",
           391 => x"18",
           392 => x"88",
           393 => x"55",
           394 => x"79",
           395 => x"ba",
           396 => x"c5",
           397 => x"2b",
           398 => x"2e",
           399 => x"fc",
           400 => x"55",
           401 => x"5f",
           402 => x"80",
           403 => x"79",
           404 => x"80",
           405 => x"90",
           406 => x"06",
           407 => x"75",
           408 => x"54",
           409 => x"83",
           410 => x"86",
           411 => x"54",
           412 => x"79",
           413 => x"83",
           414 => x"2e",
           415 => x"06",
           416 => x"2a",
           417 => x"7a",
           418 => x"97",
           419 => x"8f",
           420 => x"7e",
           421 => x"80",
           422 => x"90",
           423 => x"9d",
           424 => x"3f",
           425 => x"80",
           426 => x"54",
           427 => x"06",
           428 => x"79",
           429 => x"05",
           430 => x"75",
           431 => x"87",
           432 => x"29",
           433 => x"5b",
           434 => x"7a",
           435 => x"7a",
           436 => x"e3",
           437 => x"2e",
           438 => x"81",
           439 => x"96",
           440 => x"52",
           441 => x"9c",
           442 => x"81",
           443 => x"38",
           444 => x"80",
           445 => x"55",
           446 => x"52",
           447 => x"7a",
           448 => x"33",
           449 => x"c8",
           450 => x"f8",
           451 => x"08",
           452 => x"42",
           453 => x"84",
           454 => x"13",
           455 => x"84",
           456 => x"70",
           457 => x"41",
           458 => x"5c",
           459 => x"84",
           460 => x"70",
           461 => x"25",
           462 => x"85",
           463 => x"83",
           464 => x"ff",
           465 => x"75",
           466 => x"d8",
           467 => x"ff",
           468 => x"ff",
           469 => x"70",
           470 => x"3f",
           471 => x"fc",
           472 => x"fc",
           473 => x"58",
           474 => x"81",
           475 => x"38",
           476 => x"71",
           477 => x"7e",
           478 => x"bf",
           479 => x"ad",
           480 => x"5b",
           481 => x"7a",
           482 => x"59",
           483 => x"7f",
           484 => x"06",
           485 => x"38",
           486 => x"8c",
           487 => x"31",
           488 => x"58",
           489 => x"7c",
           490 => x"f7",
           491 => x"08",
           492 => x"79",
           493 => x"3f",
           494 => x"06",
           495 => x"c4",
           496 => x"58",
           497 => x"39",
           498 => x"80",
           499 => x"54",
           500 => x"52",
           501 => x"7c",
           502 => x"90",
           503 => x"7c",
           504 => x"88",
           505 => x"fb",
           506 => x"2c",
           507 => x"2c",
           508 => x"53",
           509 => x"7c",
           510 => x"81",
           511 => x"38",
           512 => x"2a",
           513 => x"5b",
           514 => x"c8",
           515 => x"98",
           516 => x"52",
           517 => x"7c",
           518 => x"be",
           519 => x"3f",
           520 => x"06",
           521 => x"fd",
           522 => x"71",
           523 => x"fd",
           524 => x"ec",
           525 => x"b5",
           526 => x"0d",
           527 => x"08",
           528 => x"32",
           529 => x"57",
           530 => x"06",
           531 => x"56",
           532 => x"84",
           533 => x"14",
           534 => x"08",
           535 => x"70",
           536 => x"2e",
           537 => x"d7",
           538 => x"d5",
           539 => x"08",
           540 => x"80",
           541 => x"75",
           542 => x"04",
           543 => x"80",
           544 => x"81",
           545 => x"57",
           546 => x"06",
           547 => x"33",
           548 => x"98",
           549 => x"0c",
           550 => x"05",
           551 => x"38",
           552 => x"53",
           553 => x"2e",
           554 => x"56",
           555 => x"39",
           556 => x"52",
           557 => x"04",
           558 => x"33",
           559 => x"56",
           560 => x"38",
           561 => x"80",
           562 => x"72",
           563 => x"08",
           564 => x"05",
           565 => x"13",
           566 => x"ba",
           567 => x"52",
           568 => x"08",
           569 => x"8c",
           570 => x"05",
           571 => x"fb",
           572 => x"81",
           573 => x"55",
           574 => x"38",
           575 => x"b3",
           576 => x"71",
           577 => x"70",
           578 => x"f0",
           579 => x"08",
           580 => x"ff",
           581 => x"87",
           582 => x"53",
           583 => x"81",
           584 => x"84",
           585 => x"75",
           586 => x"84",
           587 => x"08",
           588 => x"33",
           589 => x"8c",
           590 => x"07",
           591 => x"73",
           592 => x"04",
           593 => x"34",
           594 => x"75",
           595 => x"81",
           596 => x"ff",
           597 => x"33",
           598 => x"34",
           599 => x"0c",
           600 => x"76",
           601 => x"70",
           602 => x"a1",
           603 => x"70",
           604 => x"05",
           605 => x"38",
           606 => x"0d",
           607 => x"d9",
           608 => x"13",
           609 => x"34",
           610 => x"38",
           611 => x"33",
           612 => x"38",
           613 => x"53",
           614 => x"51",
           615 => x"31",
           616 => x"0d",
           617 => x"54",
           618 => x"33",
           619 => x"34",
           620 => x"0c",
           621 => x"75",
           622 => x"70",
           623 => x"05",
           624 => x"34",
           625 => x"84",
           626 => x"fc",
           627 => x"54",
           628 => x"75",
           629 => x"71",
           630 => x"81",
           631 => x"ff",
           632 => x"70",
           633 => x"04",
           634 => x"53",
           635 => x"ff",
           636 => x"2e",
           637 => x"8c",
           638 => x"ba",
           639 => x"3d",
           640 => x"80",
           641 => x"ba",
           642 => x"b3",
           643 => x"84",
           644 => x"84",
           645 => x"34",
           646 => x"08",
           647 => x"08",
           648 => x"3d",
           649 => x"71",
           650 => x"2e",
           651 => x"33",
           652 => x"12",
           653 => x"ea",
           654 => x"52",
           655 => x"0d",
           656 => x"72",
           657 => x"8e",
           658 => x"34",
           659 => x"84",
           660 => x"fa",
           661 => x"52",
           662 => x"80",
           663 => x"e0",
           664 => x"73",
           665 => x"8c",
           666 => x"26",
           667 => x"2e",
           668 => x"2a",
           669 => x"54",
           670 => x"a8",
           671 => x"74",
           672 => x"11",
           673 => x"06",
           674 => x"52",
           675 => x"38",
           676 => x"ba",
           677 => x"3d",
           678 => x"70",
           679 => x"84",
           680 => x"70",
           681 => x"80",
           682 => x"71",
           683 => x"70",
           684 => x"74",
           685 => x"73",
           686 => x"10",
           687 => x"81",
           688 => x"30",
           689 => x"84",
           690 => x"51",
           691 => x"51",
           692 => x"54",
           693 => x"0d",
           694 => x"54",
           695 => x"73",
           696 => x"0c",
           697 => x"0d",
           698 => x"80",
           699 => x"3f",
           700 => x"52",
           701 => x"fe",
           702 => x"31",
           703 => x"c5",
           704 => x"38",
           705 => x"31",
           706 => x"80",
           707 => x"10",
           708 => x"07",
           709 => x"70",
           710 => x"31",
           711 => x"58",
           712 => x"ba",
           713 => x"3d",
           714 => x"7a",
           715 => x"7d",
           716 => x"57",
           717 => x"55",
           718 => x"08",
           719 => x"0c",
           720 => x"7b",
           721 => x"77",
           722 => x"a0",
           723 => x"15",
           724 => x"73",
           725 => x"80",
           726 => x"38",
           727 => x"26",
           728 => x"a0",
           729 => x"74",
           730 => x"ff",
           731 => x"ff",
           732 => x"38",
           733 => x"54",
           734 => x"78",
           735 => x"13",
           736 => x"56",
           737 => x"38",
           738 => x"56",
           739 => x"ba",
           740 => x"70",
           741 => x"56",
           742 => x"fe",
           743 => x"70",
           744 => x"a6",
           745 => x"a0",
           746 => x"38",
           747 => x"89",
           748 => x"ba",
           749 => x"58",
           750 => x"55",
           751 => x"0b",
           752 => x"04",
           753 => x"80",
           754 => x"56",
           755 => x"06",
           756 => x"70",
           757 => x"38",
           758 => x"b0",
           759 => x"80",
           760 => x"8a",
           761 => x"c4",
           762 => x"e0",
           763 => x"d0",
           764 => x"90",
           765 => x"81",
           766 => x"81",
           767 => x"38",
           768 => x"79",
           769 => x"a0",
           770 => x"84",
           771 => x"81",
           772 => x"3d",
           773 => x"0c",
           774 => x"2e",
           775 => x"15",
           776 => x"73",
           777 => x"73",
           778 => x"a0",
           779 => x"80",
           780 => x"e1",
           781 => x"3d",
           782 => x"78",
           783 => x"fe",
           784 => x"0c",
           785 => x"3f",
           786 => x"84",
           787 => x"73",
           788 => x"10",
           789 => x"08",
           790 => x"3f",
           791 => x"51",
           792 => x"83",
           793 => x"3d",
           794 => x"9d",
           795 => x"bc",
           796 => x"04",
           797 => x"83",
           798 => x"ee",
           799 => x"cf",
           800 => x"0d",
           801 => x"3f",
           802 => x"51",
           803 => x"83",
           804 => x"3d",
           805 => x"c5",
           806 => x"84",
           807 => x"04",
           808 => x"83",
           809 => x"ee",
           810 => x"d1",
           811 => x"0d",
           812 => x"3f",
           813 => x"51",
           814 => x"83",
           815 => x"3d",
           816 => x"ed",
           817 => x"8c",
           818 => x"04",
           819 => x"80",
           820 => x"79",
           821 => x"57",
           822 => x"26",
           823 => x"70",
           824 => x"74",
           825 => x"8c",
           826 => x"3f",
           827 => x"8c",
           828 => x"51",
           829 => x"78",
           830 => x"2a",
           831 => x"80",
           832 => x"08",
           833 => x"38",
           834 => x"f5",
           835 => x"83",
           836 => x"98",
           837 => x"8c",
           838 => x"8c",
           839 => x"ba",
           840 => x"54",
           841 => x"82",
           842 => x"57",
           843 => x"7a",
           844 => x"74",
           845 => x"87",
           846 => x"84",
           847 => x"a7",
           848 => x"d2",
           849 => x"51",
           850 => x"3d",
           851 => x"33",
           852 => x"52",
           853 => x"8c",
           854 => x"38",
           855 => x"ba",
           856 => x"04",
           857 => x"54",
           858 => x"51",
           859 => x"ba",
           860 => x"3d",
           861 => x"80",
           862 => x"41",
           863 => x"80",
           864 => x"d2",
           865 => x"cc",
           866 => x"79",
           867 => x"ed",
           868 => x"73",
           869 => x"38",
           870 => x"dd",
           871 => x"08",
           872 => x"78",
           873 => x"51",
           874 => x"27",
           875 => x"55",
           876 => x"38",
           877 => x"83",
           878 => x"81",
           879 => x"88",
           880 => x"38",
           881 => x"eb",
           882 => x"26",
           883 => x"d5",
           884 => x"80",
           885 => x"08",
           886 => x"76",
           887 => x"2e",
           888 => x"78",
           889 => x"ba",
           890 => x"d2",
           891 => x"84",
           892 => x"eb",
           893 => x"38",
           894 => x"dc",
           895 => x"08",
           896 => x"73",
           897 => x"53",
           898 => x"52",
           899 => x"82",
           900 => x"a0",
           901 => x"dd",
           902 => x"51",
           903 => x"f0",
           904 => x"3f",
           905 => x"18",
           906 => x"08",
           907 => x"3f",
           908 => x"54",
           909 => x"26",
           910 => x"f0",
           911 => x"81",
           912 => x"e3",
           913 => x"06",
           914 => x"ec",
           915 => x"09",
           916 => x"fc",
           917 => x"84",
           918 => x"2c",
           919 => x"32",
           920 => x"07",
           921 => x"53",
           922 => x"51",
           923 => x"98",
           924 => x"70",
           925 => x"72",
           926 => x"58",
           927 => x"ff",
           928 => x"84",
           929 => x"fe",
           930 => x"53",
           931 => x"3f",
           932 => x"80",
           933 => x"70",
           934 => x"38",
           935 => x"52",
           936 => x"70",
           937 => x"38",
           938 => x"52",
           939 => x"70",
           940 => x"38",
           941 => x"52",
           942 => x"70",
           943 => x"72",
           944 => x"38",
           945 => x"81",
           946 => x"51",
           947 => x"3f",
           948 => x"81",
           949 => x"51",
           950 => x"3f",
           951 => x"80",
           952 => x"9b",
           953 => x"de",
           954 => x"87",
           955 => x"80",
           956 => x"51",
           957 => x"9b",
           958 => x"72",
           959 => x"71",
           960 => x"39",
           961 => x"9c",
           962 => x"fe",
           963 => x"51",
           964 => x"ff",
           965 => x"83",
           966 => x"51",
           967 => x"81",
           968 => x"94",
           969 => x"c6",
           970 => x"3f",
           971 => x"2a",
           972 => x"2e",
           973 => x"51",
           974 => x"9a",
           975 => x"72",
           976 => x"71",
           977 => x"39",
           978 => x"ff",
           979 => x"52",
           980 => x"ba",
           981 => x"40",
           982 => x"83",
           983 => x"3d",
           984 => x"3f",
           985 => x"7e",
           986 => x"ef",
           987 => x"59",
           988 => x"81",
           989 => x"06",
           990 => x"67",
           991 => x"dc",
           992 => x"09",
           993 => x"33",
           994 => x"80",
           995 => x"90",
           996 => x"52",
           997 => x"08",
           998 => x"7b",
           999 => x"ba",
          1000 => x"5e",
          1001 => x"1c",
          1002 => x"7c",
          1003 => x"7b",
          1004 => x"52",
          1005 => x"8c",
          1006 => x"2e",
          1007 => x"48",
          1008 => x"93",
          1009 => x"06",
          1010 => x"38",
          1011 => x"3f",
          1012 => x"f3",
          1013 => x"7a",
          1014 => x"24",
          1015 => x"ee",
          1016 => x"e4",
          1017 => x"f2",
          1018 => x"56",
          1019 => x"53",
          1020 => x"ae",
          1021 => x"8c",
          1022 => x"80",
          1023 => x"7a",
          1024 => x"7a",
          1025 => x"81",
          1026 => x"7a",
          1027 => x"81",
          1028 => x"61",
          1029 => x"81",
          1030 => x"d3",
          1031 => x"80",
          1032 => x"0b",
          1033 => x"06",
          1034 => x"53",
          1035 => x"51",
          1036 => x"08",
          1037 => x"83",
          1038 => x"80",
          1039 => x"3f",
          1040 => x"38",
          1041 => x"3f",
          1042 => x"81",
          1043 => x"09",
          1044 => x"84",
          1045 => x"82",
          1046 => x"83",
          1047 => x"51",
          1048 => x"79",
          1049 => x"63",
          1050 => x"89",
          1051 => x"83",
          1052 => x"83",
          1053 => x"3d",
          1054 => x"7e",
          1055 => x"52",
          1056 => x"3f",
          1057 => x"81",
          1058 => x"3d",
          1059 => x"d6",
          1060 => x"81",
          1061 => x"d6",
          1062 => x"54",
          1063 => x"51",
          1064 => x"8c",
          1065 => x"3f",
          1066 => x"bf",
          1067 => x"95",
          1068 => x"51",
          1069 => x"83",
          1070 => x"f3",
          1071 => x"84",
          1072 => x"80",
          1073 => x"fa",
          1074 => x"51",
          1075 => x"84",
          1076 => x"38",
          1077 => x"f8",
          1078 => x"b8",
          1079 => x"05",
          1080 => x"08",
          1081 => x"83",
          1082 => x"59",
          1083 => x"53",
          1084 => x"84",
          1085 => x"38",
          1086 => x"80",
          1087 => x"8c",
          1088 => x"08",
          1089 => x"cf",
          1090 => x"80",
          1091 => x"7e",
          1092 => x"f9",
          1093 => x"38",
          1094 => x"39",
          1095 => x"80",
          1096 => x"8c",
          1097 => x"3d",
          1098 => x"51",
          1099 => x"86",
          1100 => x"78",
          1101 => x"3f",
          1102 => x"52",
          1103 => x"7e",
          1104 => x"38",
          1105 => x"82",
          1106 => x"3d",
          1107 => x"51",
          1108 => x"80",
          1109 => x"fc",
          1110 => x"d0",
          1111 => x"f8",
          1112 => x"53",
          1113 => x"84",
          1114 => x"38",
          1115 => x"68",
          1116 => x"8d",
          1117 => x"5c",
          1118 => x"55",
          1119 => x"83",
          1120 => x"66",
          1121 => x"59",
          1122 => x"53",
          1123 => x"84",
          1124 => x"38",
          1125 => x"80",
          1126 => x"8c",
          1127 => x"3d",
          1128 => x"51",
          1129 => x"80",
          1130 => x"51",
          1131 => x"27",
          1132 => x"81",
          1133 => x"05",
          1134 => x"11",
          1135 => x"3f",
          1136 => x"b9",
          1137 => x"ff",
          1138 => x"ba",
          1139 => x"54",
          1140 => x"3f",
          1141 => x"52",
          1142 => x"7e",
          1143 => x"38",
          1144 => x"81",
          1145 => x"80",
          1146 => x"05",
          1147 => x"ff",
          1148 => x"ba",
          1149 => x"68",
          1150 => x"34",
          1151 => x"fc",
          1152 => x"80",
          1153 => x"38",
          1154 => x"11",
          1155 => x"3f",
          1156 => x"99",
          1157 => x"ff",
          1158 => x"ba",
          1159 => x"b8",
          1160 => x"05",
          1161 => x"08",
          1162 => x"83",
          1163 => x"67",
          1164 => x"65",
          1165 => x"0c",
          1166 => x"d9",
          1167 => x"ff",
          1168 => x"ba",
          1169 => x"52",
          1170 => x"ba",
          1171 => x"3f",
          1172 => x"99",
          1173 => x"ec",
          1174 => x"84",
          1175 => x"c8",
          1176 => x"83",
          1177 => x"83",
          1178 => x"b8",
          1179 => x"05",
          1180 => x"08",
          1181 => x"79",
          1182 => x"cc",
          1183 => x"53",
          1184 => x"84",
          1185 => x"80",
          1186 => x"38",
          1187 => x"70",
          1188 => x"5f",
          1189 => x"a0",
          1190 => x"a0",
          1191 => x"54",
          1192 => x"9e",
          1193 => x"3f",
          1194 => x"59",
          1195 => x"f0",
          1196 => x"9c",
          1197 => x"f2",
          1198 => x"64",
          1199 => x"11",
          1200 => x"3f",
          1201 => x"b1",
          1202 => x"22",
          1203 => x"45",
          1204 => x"80",
          1205 => x"8c",
          1206 => x"5e",
          1207 => x"82",
          1208 => x"fe",
          1209 => x"e1",
          1210 => x"b9",
          1211 => x"fc",
          1212 => x"a0",
          1213 => x"81",
          1214 => x"05",
          1215 => x"fb",
          1216 => x"53",
          1217 => x"84",
          1218 => x"38",
          1219 => x"05",
          1220 => x"83",
          1221 => x"7b",
          1222 => x"83",
          1223 => x"3f",
          1224 => x"da",
          1225 => x"c4",
          1226 => x"b8",
          1227 => x"05",
          1228 => x"08",
          1229 => x"80",
          1230 => x"5b",
          1231 => x"f3",
          1232 => x"cf",
          1233 => x"ea",
          1234 => x"80",
          1235 => x"49",
          1236 => x"d3",
          1237 => x"83",
          1238 => x"59",
          1239 => x"59",
          1240 => x"d8",
          1241 => x"f0",
          1242 => x"83",
          1243 => x"9b",
          1244 => x"92",
          1245 => x"80",
          1246 => x"49",
          1247 => x"5e",
          1248 => x"e4",
          1249 => x"8e",
          1250 => x"83",
          1251 => x"83",
          1252 => x"94",
          1253 => x"ca",
          1254 => x"05",
          1255 => x"08",
          1256 => x"3d",
          1257 => x"87",
          1258 => x"87",
          1259 => x"3f",
          1260 => x"08",
          1261 => x"51",
          1262 => x"08",
          1263 => x"70",
          1264 => x"74",
          1265 => x"08",
          1266 => x"84",
          1267 => x"74",
          1268 => x"8c",
          1269 => x"0c",
          1270 => x"94",
          1271 => x"eb",
          1272 => x"34",
          1273 => x"3d",
          1274 => x"84",
          1275 => x"89",
          1276 => x"51",
          1277 => x"83",
          1278 => x"f2",
          1279 => x"3f",
          1280 => x"53",
          1281 => x"51",
          1282 => x"f8",
          1283 => x"70",
          1284 => x"74",
          1285 => x"70",
          1286 => x"2e",
          1287 => x"70",
          1288 => x"55",
          1289 => x"ff",
          1290 => x"38",
          1291 => x"38",
          1292 => x"53",
          1293 => x"81",
          1294 => x"80",
          1295 => x"39",
          1296 => x"70",
          1297 => x"81",
          1298 => x"80",
          1299 => x"80",
          1300 => x"05",
          1301 => x"70",
          1302 => x"04",
          1303 => x"2e",
          1304 => x"72",
          1305 => x"54",
          1306 => x"e0",
          1307 => x"53",
          1308 => x"f8",
          1309 => x"53",
          1310 => x"ba",
          1311 => x"3d",
          1312 => x"3f",
          1313 => x"38",
          1314 => x"0d",
          1315 => x"33",
          1316 => x"8b",
          1317 => x"ff",
          1318 => x"81",
          1319 => x"52",
          1320 => x"13",
          1321 => x"80",
          1322 => x"52",
          1323 => x"13",
          1324 => x"26",
          1325 => x"87",
          1326 => x"38",
          1327 => x"72",
          1328 => x"13",
          1329 => x"13",
          1330 => x"13",
          1331 => x"13",
          1332 => x"13",
          1333 => x"87",
          1334 => x"98",
          1335 => x"9c",
          1336 => x"0c",
          1337 => x"7f",
          1338 => x"7d",
          1339 => x"7d",
          1340 => x"5c",
          1341 => x"b4",
          1342 => x"c0",
          1343 => x"34",
          1344 => x"85",
          1345 => x"5c",
          1346 => x"a4",
          1347 => x"c0",
          1348 => x"23",
          1349 => x"06",
          1350 => x"86",
          1351 => x"84",
          1352 => x"82",
          1353 => x"06",
          1354 => x"b2",
          1355 => x"0d",
          1356 => x"2e",
          1357 => x"3f",
          1358 => x"98",
          1359 => x"81",
          1360 => x"38",
          1361 => x"0d",
          1362 => x"84",
          1363 => x"2c",
          1364 => x"06",
          1365 => x"3f",
          1366 => x"98",
          1367 => x"38",
          1368 => x"54",
          1369 => x"80",
          1370 => x"98",
          1371 => x"ff",
          1372 => x"14",
          1373 => x"71",
          1374 => x"04",
          1375 => x"83",
          1376 => x"53",
          1377 => x"38",
          1378 => x"2a",
          1379 => x"80",
          1380 => x"81",
          1381 => x"81",
          1382 => x"8a",
          1383 => x"71",
          1384 => x"87",
          1385 => x"86",
          1386 => x"72",
          1387 => x"3d",
          1388 => x"06",
          1389 => x"32",
          1390 => x"38",
          1391 => x"80",
          1392 => x"08",
          1393 => x"54",
          1394 => x"3d",
          1395 => x"70",
          1396 => x"f2",
          1397 => x"3d",
          1398 => x"56",
          1399 => x"38",
          1400 => x"81",
          1401 => x"2e",
          1402 => x"08",
          1403 => x"54",
          1404 => x"91",
          1405 => x"e3",
          1406 => x"72",
          1407 => x"81",
          1408 => x"ff",
          1409 => x"70",
          1410 => x"90",
          1411 => x"33",
          1412 => x"84",
          1413 => x"71",
          1414 => x"70",
          1415 => x"53",
          1416 => x"2a",
          1417 => x"b5",
          1418 => x"96",
          1419 => x"70",
          1420 => x"87",
          1421 => x"8a",
          1422 => x"ab",
          1423 => x"f2",
          1424 => x"83",
          1425 => x"08",
          1426 => x"98",
          1427 => x"9e",
          1428 => x"c0",
          1429 => x"87",
          1430 => x"0c",
          1431 => x"e4",
          1432 => x"f2",
          1433 => x"83",
          1434 => x"08",
          1435 => x"c0",
          1436 => x"9e",
          1437 => x"c0",
          1438 => x"fc",
          1439 => x"f3",
          1440 => x"83",
          1441 => x"08",
          1442 => x"f3",
          1443 => x"90",
          1444 => x"52",
          1445 => x"f3",
          1446 => x"90",
          1447 => x"52",
          1448 => x"52",
          1449 => x"87",
          1450 => x"0a",
          1451 => x"83",
          1452 => x"34",
          1453 => x"70",
          1454 => x"70",
          1455 => x"83",
          1456 => x"9e",
          1457 => x"51",
          1458 => x"81",
          1459 => x"0b",
          1460 => x"80",
          1461 => x"2e",
          1462 => x"92",
          1463 => x"08",
          1464 => x"52",
          1465 => x"71",
          1466 => x"c0",
          1467 => x"06",
          1468 => x"38",
          1469 => x"80",
          1470 => x"81",
          1471 => x"80",
          1472 => x"f3",
          1473 => x"90",
          1474 => x"52",
          1475 => x"52",
          1476 => x"87",
          1477 => x"06",
          1478 => x"38",
          1479 => x"87",
          1480 => x"70",
          1481 => x"98",
          1482 => x"08",
          1483 => x"70",
          1484 => x"83",
          1485 => x"08",
          1486 => x"51",
          1487 => x"87",
          1488 => x"51",
          1489 => x"81",
          1490 => x"c0",
          1491 => x"83",
          1492 => x"81",
          1493 => x"83",
          1494 => x"83",
          1495 => x"38",
          1496 => x"83",
          1497 => x"38",
          1498 => x"d1",
          1499 => x"85",
          1500 => x"74",
          1501 => x"54",
          1502 => x"33",
          1503 => x"9b",
          1504 => x"f3",
          1505 => x"83",
          1506 => x"38",
          1507 => x"b1",
          1508 => x"83",
          1509 => x"75",
          1510 => x"54",
          1511 => x"51",
          1512 => x"52",
          1513 => x"3f",
          1514 => x"ec",
          1515 => x"f8",
          1516 => x"b5",
          1517 => x"85",
          1518 => x"da",
          1519 => x"f3",
          1520 => x"75",
          1521 => x"08",
          1522 => x"54",
          1523 => x"da",
          1524 => x"f3",
          1525 => x"83",
          1526 => x"8a",
          1527 => x"04",
          1528 => x"c0",
          1529 => x"ba",
          1530 => x"71",
          1531 => x"52",
          1532 => x"3f",
          1533 => x"0d",
          1534 => x"84",
          1535 => x"84",
          1536 => x"76",
          1537 => x"08",
          1538 => x"f2",
          1539 => x"80",
          1540 => x"83",
          1541 => x"d9",
          1542 => x"f0",
          1543 => x"b3",
          1544 => x"83",
          1545 => x"83",
          1546 => x"51",
          1547 => x"51",
          1548 => x"52",
          1549 => x"3f",
          1550 => x"c0",
          1551 => x"ba",
          1552 => x"71",
          1553 => x"52",
          1554 => x"3f",
          1555 => x"2e",
          1556 => x"db",
          1557 => x"f3",
          1558 => x"84",
          1559 => x"51",
          1560 => x"33",
          1561 => x"d6",
          1562 => x"9d",
          1563 => x"80",
          1564 => x"dc",
          1565 => x"f3",
          1566 => x"a9",
          1567 => x"52",
          1568 => x"3f",
          1569 => x"2e",
          1570 => x"9c",
          1571 => x"b1",
          1572 => x"74",
          1573 => x"83",
          1574 => x"51",
          1575 => x"33",
          1576 => x"cd",
          1577 => x"dc",
          1578 => x"51",
          1579 => x"33",
          1580 => x"c7",
          1581 => x"d4",
          1582 => x"51",
          1583 => x"33",
          1584 => x"c1",
          1585 => x"cc",
          1586 => x"51",
          1587 => x"33",
          1588 => x"c1",
          1589 => x"e4",
          1590 => x"51",
          1591 => x"33",
          1592 => x"c1",
          1593 => x"ec",
          1594 => x"51",
          1595 => x"33",
          1596 => x"c1",
          1597 => x"9a",
          1598 => x"fd",
          1599 => x"80",
          1600 => x"3d",
          1601 => x"85",
          1602 => x"c3",
          1603 => x"de",
          1604 => x"3d",
          1605 => x"af",
          1606 => x"de",
          1607 => x"3d",
          1608 => x"af",
          1609 => x"de",
          1610 => x"3d",
          1611 => x"af",
          1612 => x"88",
          1613 => x"96",
          1614 => x"87",
          1615 => x"0d",
          1616 => x"5a",
          1617 => x"f3",
          1618 => x"84",
          1619 => x"3d",
          1620 => x"54",
          1621 => x"d2",
          1622 => x"2e",
          1623 => x"84",
          1624 => x"80",
          1625 => x"38",
          1626 => x"18",
          1627 => x"70",
          1628 => x"55",
          1629 => x"ff",
          1630 => x"11",
          1631 => x"84",
          1632 => x"2e",
          1633 => x"a9",
          1634 => x"ff",
          1635 => x"81",
          1636 => x"c0",
          1637 => x"3f",
          1638 => x"08",
          1639 => x"51",
          1640 => x"ba",
          1641 => x"3d",
          1642 => x"71",
          1643 => x"57",
          1644 => x"0b",
          1645 => x"10",
          1646 => x"54",
          1647 => x"08",
          1648 => x"8f",
          1649 => x"84",
          1650 => x"88",
          1651 => x"16",
          1652 => x"76",
          1653 => x"ba",
          1654 => x"1a",
          1655 => x"ff",
          1656 => x"ba",
          1657 => x"1b",
          1658 => x"3f",
          1659 => x"54",
          1660 => x"70",
          1661 => x"27",
          1662 => x"33",
          1663 => x"e6",
          1664 => x"55",
          1665 => x"fe",
          1666 => x"80",
          1667 => x"39",
          1668 => x"f3",
          1669 => x"3f",
          1670 => x"83",
          1671 => x"77",
          1672 => x"8c",
          1673 => x"ff",
          1674 => x"55",
          1675 => x"9d",
          1676 => x"70",
          1677 => x"53",
          1678 => x"52",
          1679 => x"2e",
          1680 => x"0b",
          1681 => x"04",
          1682 => x"3d",
          1683 => x"80",
          1684 => x"33",
          1685 => x"9e",
          1686 => x"56",
          1687 => x"80",
          1688 => x"06",
          1689 => x"80",
          1690 => x"3d",
          1691 => x"84",
          1692 => x"2c",
          1693 => x"79",
          1694 => x"70",
          1695 => x"c4",
          1696 => x"71",
          1697 => x"de",
          1698 => x"52",
          1699 => x"5c",
          1700 => x"cd",
          1701 => x"75",
          1702 => x"05",
          1703 => x"24",
          1704 => x"82",
          1705 => x"dc",
          1706 => x"91",
          1707 => x"70",
          1708 => x"95",
          1709 => x"84",
          1710 => x"2e",
          1711 => x"2b",
          1712 => x"70",
          1713 => x"2c",
          1714 => x"11",
          1715 => x"57",
          1716 => x"76",
          1717 => x"81",
          1718 => x"80",
          1719 => x"98",
          1720 => x"41",
          1721 => x"10",
          1722 => x"0b",
          1723 => x"77",
          1724 => x"15",
          1725 => x"61",
          1726 => x"ff",
          1727 => x"76",
          1728 => x"39",
          1729 => x"76",
          1730 => x"34",
          1731 => x"34",
          1732 => x"26",
          1733 => x"c3",
          1734 => x"de",
          1735 => x"84",
          1736 => x"c4",
          1737 => x"56",
          1738 => x"d5",
          1739 => x"90",
          1740 => x"57",
          1741 => x"39",
          1742 => x"06",
          1743 => x"75",
          1744 => x"f0",
          1745 => x"d1",
          1746 => x"55",
          1747 => x"7c",
          1748 => x"10",
          1749 => x"59",
          1750 => x"cc",
          1751 => x"33",
          1752 => x"80",
          1753 => x"52",
          1754 => x"d5",
          1755 => x"90",
          1756 => x"51",
          1757 => x"33",
          1758 => x"34",
          1759 => x"38",
          1760 => x"84",
          1761 => x"8a",
          1762 => x"8d",
          1763 => x"a4",
          1764 => x"8e",
          1765 => x"2e",
          1766 => x"f2",
          1767 => x"cc",
          1768 => x"06",
          1769 => x"ff",
          1770 => x"84",
          1771 => x"2e",
          1772 => x"52",
          1773 => x"d5",
          1774 => x"f8",
          1775 => x"51",
          1776 => x"33",
          1777 => x"34",
          1778 => x"84",
          1779 => x"84",
          1780 => x"79",
          1781 => x"08",
          1782 => x"d0",
          1783 => x"ff",
          1784 => x"70",
          1785 => x"5a",
          1786 => x"38",
          1787 => x"57",
          1788 => x"70",
          1789 => x"84",
          1790 => x"84",
          1791 => x"76",
          1792 => x"84",
          1793 => x"56",
          1794 => x"ff",
          1795 => x"75",
          1796 => x"ff",
          1797 => x"80",
          1798 => x"a0",
          1799 => x"d0",
          1800 => x"84",
          1801 => x"74",
          1802 => x"f0",
          1803 => x"3f",
          1804 => x"0a",
          1805 => x"33",
          1806 => x"e2",
          1807 => x"51",
          1808 => x"0a",
          1809 => x"2c",
          1810 => x"7a",
          1811 => x"39",
          1812 => x"34",
          1813 => x"51",
          1814 => x"0a",
          1815 => x"2c",
          1816 => x"75",
          1817 => x"58",
          1818 => x"f0",
          1819 => x"90",
          1820 => x"80",
          1821 => x"cc",
          1822 => x"ff",
          1823 => x"d0",
          1824 => x"38",
          1825 => x"ff",
          1826 => x"ff",
          1827 => x"76",
          1828 => x"d1",
          1829 => x"34",
          1830 => x"ff",
          1831 => x"7b",
          1832 => x"08",
          1833 => x"38",
          1834 => x"2e",
          1835 => x"70",
          1836 => x"08",
          1837 => x"75",
          1838 => x"a4",
          1839 => x"80",
          1840 => x"7b",
          1841 => x"10",
          1842 => x"41",
          1843 => x"f8",
          1844 => x"83",
          1845 => x"8b",
          1846 => x"34",
          1847 => x"84",
          1848 => x"84",
          1849 => x"b6",
          1850 => x"51",
          1851 => x"08",
          1852 => x"84",
          1853 => x"ae",
          1854 => x"05",
          1855 => x"81",
          1856 => x"d2",
          1857 => x"0b",
          1858 => x"d1",
          1859 => x"34",
          1860 => x"d0",
          1861 => x"84",
          1862 => x"ae",
          1863 => x"a0",
          1864 => x"f0",
          1865 => x"3f",
          1866 => x"7c",
          1867 => x"06",
          1868 => x"51",
          1869 => x"d1",
          1870 => x"34",
          1871 => x"0d",
          1872 => x"ff",
          1873 => x"ca",
          1874 => x"59",
          1875 => x"58",
          1876 => x"f0",
          1877 => x"3f",
          1878 => x"70",
          1879 => x"52",
          1880 => x"38",
          1881 => x"ff",
          1882 => x"70",
          1883 => x"cc",
          1884 => x"24",
          1885 => x"52",
          1886 => x"81",
          1887 => x"70",
          1888 => x"51",
          1889 => x"84",
          1890 => x"ac",
          1891 => x"81",
          1892 => x"d1",
          1893 => x"25",
          1894 => x"16",
          1895 => x"d5",
          1896 => x"ac",
          1897 => x"81",
          1898 => x"d1",
          1899 => x"25",
          1900 => x"17",
          1901 => x"52",
          1902 => x"75",
          1903 => x"05",
          1904 => x"43",
          1905 => x"38",
          1906 => x"70",
          1907 => x"2e",
          1908 => x"55",
          1909 => x"2b",
          1910 => x"24",
          1911 => x"81",
          1912 => x"81",
          1913 => x"d1",
          1914 => x"25",
          1915 => x"d1",
          1916 => x"05",
          1917 => x"d1",
          1918 => x"38",
          1919 => x"34",
          1920 => x"81",
          1921 => x"70",
          1922 => x"58",
          1923 => x"38",
          1924 => x"81",
          1925 => x"25",
          1926 => x"52",
          1927 => x"81",
          1928 => x"70",
          1929 => x"57",
          1930 => x"84",
          1931 => x"aa",
          1932 => x"81",
          1933 => x"d1",
          1934 => x"24",
          1935 => x"f3",
          1936 => x"9d",
          1937 => x"84",
          1938 => x"84",
          1939 => x"05",
          1940 => x"c4",
          1941 => x"d0",
          1942 => x"c8",
          1943 => x"51",
          1944 => x"08",
          1945 => x"84",
          1946 => x"a9",
          1947 => x"05",
          1948 => x"81",
          1949 => x"80",
          1950 => x"83",
          1951 => x"85",
          1952 => x"77",
          1953 => x"d5",
          1954 => x"52",
          1955 => x"80",
          1956 => x"98",
          1957 => x"57",
          1958 => x"d0",
          1959 => x"79",
          1960 => x"75",
          1961 => x"39",
          1962 => x"fc",
          1963 => x"76",
          1964 => x"84",
          1965 => x"38",
          1966 => x"f3",
          1967 => x"d4",
          1968 => x"83",
          1969 => x"3f",
          1970 => x"3d",
          1971 => x"74",
          1972 => x"0c",
          1973 => x"80",
          1974 => x"75",
          1975 => x"8c",
          1976 => x"8c",
          1977 => x"75",
          1978 => x"93",
          1979 => x"d0",
          1980 => x"f2",
          1981 => x"88",
          1982 => x"f0",
          1983 => x"3f",
          1984 => x"ff",
          1985 => x"ff",
          1986 => x"79",
          1987 => x"7c",
          1988 => x"80",
          1989 => x"ba",
          1990 => x"51",
          1991 => x"08",
          1992 => x"08",
          1993 => x"52",
          1994 => x"1d",
          1995 => x"33",
          1996 => x"56",
          1997 => x"d5",
          1998 => x"f8",
          1999 => x"51",
          2000 => x"08",
          2001 => x"84",
          2002 => x"84",
          2003 => x"55",
          2004 => x"3f",
          2005 => x"34",
          2006 => x"81",
          2007 => x"a9",
          2008 => x"06",
          2009 => x"33",
          2010 => x"f0",
          2011 => x"88",
          2012 => x"f0",
          2013 => x"3f",
          2014 => x"ff",
          2015 => x"ff",
          2016 => x"60",
          2017 => x"51",
          2018 => x"33",
          2019 => x"f3",
          2020 => x"5c",
          2021 => x"8c",
          2022 => x"70",
          2023 => x"08",
          2024 => x"d5",
          2025 => x"ff",
          2026 => x"81",
          2027 => x"93",
          2028 => x"f3",
          2029 => x"fe",
          2030 => x"75",
          2031 => x"f8",
          2032 => x"3f",
          2033 => x"c2",
          2034 => x"80",
          2035 => x"ba",
          2036 => x"53",
          2037 => x"81",
          2038 => x"82",
          2039 => x"3d",
          2040 => x"80",
          2041 => x"3f",
          2042 => x"8c",
          2043 => x"ee",
          2044 => x"a6",
          2045 => x"80",
          2046 => x"e3",
          2047 => x"70",
          2048 => x"81",
          2049 => x"10",
          2050 => x"58",
          2051 => x"76",
          2052 => x"a4",
          2053 => x"80",
          2054 => x"75",
          2055 => x"10",
          2056 => x"40",
          2057 => x"81",
          2058 => x"83",
          2059 => x"81",
          2060 => x"38",
          2061 => x"74",
          2062 => x"fc",
          2063 => x"5b",
          2064 => x"80",
          2065 => x"39",
          2066 => x"f3",
          2067 => x"06",
          2068 => x"54",
          2069 => x"84",
          2070 => x"fc",
          2071 => x"05",
          2072 => x"2e",
          2073 => x"83",
          2074 => x"83",
          2075 => x"e1",
          2076 => x"e7",
          2077 => x"0d",
          2078 => x"05",
          2079 => x"83",
          2080 => x"81",
          2081 => x"38",
          2082 => x"a3",
          2083 => x"70",
          2084 => x"79",
          2085 => x"bc",
          2086 => x"83",
          2087 => x"70",
          2088 => x"88",
          2089 => x"56",
          2090 => x"80",
          2091 => x"73",
          2092 => x"26",
          2093 => x"83",
          2094 => x"79",
          2095 => x"e0",
          2096 => x"05",
          2097 => x"38",
          2098 => x"80",
          2099 => x"10",
          2100 => x"29",
          2101 => x"59",
          2102 => x"80",
          2103 => x"ff",
          2104 => x"ba",
          2105 => x"75",
          2106 => x"5b",
          2107 => x"74",
          2108 => x"06",
          2109 => x"06",
          2110 => x"ff",
          2111 => x"57",
          2112 => x"38",
          2113 => x"05",
          2114 => x"83",
          2115 => x"38",
          2116 => x"fe",
          2117 => x"55",
          2118 => x"81",
          2119 => x"a0",
          2120 => x"84",
          2121 => x"84",
          2122 => x"83",
          2123 => x"5b",
          2124 => x"78",
          2125 => x"06",
          2126 => x"18",
          2127 => x"bb",
          2128 => x"80",
          2129 => x"b8",
          2130 => x"07",
          2131 => x"7f",
          2132 => x"fd",
          2133 => x"e6",
          2134 => x"ff",
          2135 => x"bd",
          2136 => x"a0",
          2137 => x"5f",
          2138 => x"b8",
          2139 => x"b7",
          2140 => x"f9",
          2141 => x"7c",
          2142 => x"5f",
          2143 => x"26",
          2144 => x"7d",
          2145 => x"06",
          2146 => x"7d",
          2147 => x"06",
          2148 => x"5d",
          2149 => x"75",
          2150 => x"83",
          2151 => x"76",
          2152 => x"fb",
          2153 => x"56",
          2154 => x"ee",
          2155 => x"ff",
          2156 => x"53",
          2157 => x"ee",
          2158 => x"76",
          2159 => x"80",
          2160 => x"75",
          2161 => x"81",
          2162 => x"90",
          2163 => x"f8",
          2164 => x"06",
          2165 => x"73",
          2166 => x"07",
          2167 => x"87",
          2168 => x"51",
          2169 => x"73",
          2170 => x"72",
          2171 => x"80",
          2172 => x"87",
          2173 => x"84",
          2174 => x"02",
          2175 => x"05",
          2176 => x"56",
          2177 => x"38",
          2178 => x"33",
          2179 => x"12",
          2180 => x"ba",
          2181 => x"29",
          2182 => x"f8",
          2183 => x"81",
          2184 => x"22",
          2185 => x"23",
          2186 => x"81",
          2187 => x"5b",
          2188 => x"ff",
          2189 => x"83",
          2190 => x"06",
          2191 => x"79",
          2192 => x"80",
          2193 => x"54",
          2194 => x"98",
          2195 => x"13",
          2196 => x"81",
          2197 => x"57",
          2198 => x"73",
          2199 => x"a1",
          2200 => x"de",
          2201 => x"14",
          2202 => x"34",
          2203 => x"eb",
          2204 => x"56",
          2205 => x"78",
          2206 => x"06",
          2207 => x"38",
          2208 => x"80",
          2209 => x"75",
          2210 => x"a3",
          2211 => x"81",
          2212 => x"5c",
          2213 => x"84",
          2214 => x"33",
          2215 => x"70",
          2216 => x"05",
          2217 => x"34",
          2218 => x"b7",
          2219 => x"5c",
          2220 => x"80",
          2221 => x"3d",
          2222 => x"83",
          2223 => x"06",
          2224 => x"73",
          2225 => x"2e",
          2226 => x"ff",
          2227 => x"72",
          2228 => x"38",
          2229 => x"80",
          2230 => x"11",
          2231 => x"fe",
          2232 => x"98",
          2233 => x"56",
          2234 => x"75",
          2235 => x"53",
          2236 => x"0b",
          2237 => x"81",
          2238 => x"d8",
          2239 => x"b8",
          2240 => x"83",
          2241 => x"88",
          2242 => x"33",
          2243 => x"76",
          2244 => x"51",
          2245 => x"10",
          2246 => x"04",
          2247 => x"27",
          2248 => x"80",
          2249 => x"0d",
          2250 => x"83",
          2251 => x"54",
          2252 => x"12",
          2253 => x"0b",
          2254 => x"04",
          2255 => x"70",
          2256 => x"55",
          2257 => x"de",
          2258 => x"84",
          2259 => x"51",
          2260 => x"72",
          2261 => x"ba",
          2262 => x"f9",
          2263 => x"70",
          2264 => x"55",
          2265 => x"84",
          2266 => x"83",
          2267 => x"80",
          2268 => x"74",
          2269 => x"f9",
          2270 => x"0c",
          2271 => x"f9",
          2272 => x"b7",
          2273 => x"75",
          2274 => x"70",
          2275 => x"ff",
          2276 => x"70",
          2277 => x"83",
          2278 => x"83",
          2279 => x"71",
          2280 => x"84",
          2281 => x"80",
          2282 => x"80",
          2283 => x"0b",
          2284 => x"04",
          2285 => x"90",
          2286 => x"80",
          2287 => x"0d",
          2288 => x"07",
          2289 => x"39",
          2290 => x"86",
          2291 => x"d7",
          2292 => x"34",
          2293 => x"3d",
          2294 => x"fc",
          2295 => x"b8",
          2296 => x"33",
          2297 => x"34",
          2298 => x"81",
          2299 => x"f9",
          2300 => x"b8",
          2301 => x"70",
          2302 => x"83",
          2303 => x"07",
          2304 => x"ef",
          2305 => x"06",
          2306 => x"df",
          2307 => x"06",
          2308 => x"b8",
          2309 => x"33",
          2310 => x"83",
          2311 => x"f9",
          2312 => x"07",
          2313 => x"a7",
          2314 => x"06",
          2315 => x"b8",
          2316 => x"33",
          2317 => x"83",
          2318 => x"f9",
          2319 => x"83",
          2320 => x"f9",
          2321 => x"51",
          2322 => x"39",
          2323 => x"02",
          2324 => x"f9",
          2325 => x"f9",
          2326 => x"41",
          2327 => x"82",
          2328 => x"78",
          2329 => x"b8",
          2330 => x"34",
          2331 => x"f9",
          2332 => x"8f",
          2333 => x"81",
          2334 => x"82",
          2335 => x"82",
          2336 => x"83",
          2337 => x"ba",
          2338 => x"57",
          2339 => x"fe",
          2340 => x"52",
          2341 => x"3f",
          2342 => x"84",
          2343 => x"34",
          2344 => x"f9",
          2345 => x"0b",
          2346 => x"b8",
          2347 => x"34",
          2348 => x"0b",
          2349 => x"33",
          2350 => x"b9",
          2351 => x"7c",
          2352 => x"ff",
          2353 => x"8d",
          2354 => x"38",
          2355 => x"22",
          2356 => x"80",
          2357 => x"06",
          2358 => x"78",
          2359 => x"51",
          2360 => x"82",
          2361 => x"7a",
          2362 => x"ba",
          2363 => x"3d",
          2364 => x"34",
          2365 => x"0b",
          2366 => x"f9",
          2367 => x"23",
          2368 => x"3f",
          2369 => x"fc",
          2370 => x"83",
          2371 => x"78",
          2372 => x"38",
          2373 => x"e4",
          2374 => x"19",
          2375 => x"39",
          2376 => x"a7",
          2377 => x"f9",
          2378 => x"71",
          2379 => x"83",
          2380 => x"71",
          2381 => x"06",
          2382 => x"55",
          2383 => x"38",
          2384 => x"89",
          2385 => x"83",
          2386 => x"38",
          2387 => x"33",
          2388 => x"05",
          2389 => x"33",
          2390 => x"b8",
          2391 => x"f9",
          2392 => x"5a",
          2393 => x"34",
          2394 => x"16",
          2395 => x"a3",
          2396 => x"33",
          2397 => x"22",
          2398 => x"11",
          2399 => x"b8",
          2400 => x"18",
          2401 => x"78",
          2402 => x"33",
          2403 => x"53",
          2404 => x"83",
          2405 => x"84",
          2406 => x"80",
          2407 => x"0c",
          2408 => x"97",
          2409 => x"75",
          2410 => x"38",
          2411 => x"80",
          2412 => x"39",
          2413 => x"b8",
          2414 => x"2e",
          2415 => x"53",
          2416 => x"81",
          2417 => x"72",
          2418 => x"a0",
          2419 => x"81",
          2420 => x"d8",
          2421 => x"bd",
          2422 => x"51",
          2423 => x"8c",
          2424 => x"ff",
          2425 => x"83",
          2426 => x"55",
          2427 => x"53",
          2428 => x"a0",
          2429 => x"33",
          2430 => x"53",
          2431 => x"83",
          2432 => x"0b",
          2433 => x"51",
          2434 => x"52",
          2435 => x"39",
          2436 => x"33",
          2437 => x"81",
          2438 => x"83",
          2439 => x"38",
          2440 => x"88",
          2441 => x"88",
          2442 => x"f9",
          2443 => x"72",
          2444 => x"88",
          2445 => x"34",
          2446 => x"33",
          2447 => x"12",
          2448 => x"be",
          2449 => x"71",
          2450 => x"b8",
          2451 => x"34",
          2452 => x"06",
          2453 => x"33",
          2454 => x"58",
          2455 => x"de",
          2456 => x"06",
          2457 => x"38",
          2458 => x"f1",
          2459 => x"bd",
          2460 => x"9c",
          2461 => x"8a",
          2462 => x"78",
          2463 => x"db",
          2464 => x"b9",
          2465 => x"f9",
          2466 => x"72",
          2467 => x"88",
          2468 => x"34",
          2469 => x"33",
          2470 => x"12",
          2471 => x"be",
          2472 => x"71",
          2473 => x"33",
          2474 => x"b8",
          2475 => x"f9",
          2476 => x"72",
          2477 => x"83",
          2478 => x"05",
          2479 => x"06",
          2480 => x"77",
          2481 => x"ba",
          2482 => x"9b",
          2483 => x"83",
          2484 => x"06",
          2485 => x"bd",
          2486 => x"9c",
          2487 => x"aa",
          2488 => x"84",
          2489 => x"11",
          2490 => x"78",
          2491 => x"ff",
          2492 => x"1a",
          2493 => x"9c",
          2494 => x"e9",
          2495 => x"84",
          2496 => x"83",
          2497 => x"5e",
          2498 => x"87",
          2499 => x"80",
          2500 => x"ba",
          2501 => x"59",
          2502 => x"83",
          2503 => x"5b",
          2504 => x"b0",
          2505 => x"70",
          2506 => x"83",
          2507 => x"44",
          2508 => x"33",
          2509 => x"1f",
          2510 => x"51",
          2511 => x"bd",
          2512 => x"33",
          2513 => x"06",
          2514 => x"12",
          2515 => x"ba",
          2516 => x"05",
          2517 => x"92",
          2518 => x"81",
          2519 => x"06",
          2520 => x"38",
          2521 => x"fc",
          2522 => x"34",
          2523 => x"0b",
          2524 => x"b9",
          2525 => x"0c",
          2526 => x"3d",
          2527 => x"b9",
          2528 => x"b9",
          2529 => x"b9",
          2530 => x"0c",
          2531 => x"3d",
          2532 => x"81",
          2533 => x"33",
          2534 => x"06",
          2535 => x"06",
          2536 => x"80",
          2537 => x"72",
          2538 => x"06",
          2539 => x"5c",
          2540 => x"fe",
          2541 => x"58",
          2542 => x"83",
          2543 => x"7a",
          2544 => x"72",
          2545 => x"b8",
          2546 => x"34",
          2547 => x"33",
          2548 => x"12",
          2549 => x"f9",
          2550 => x"60",
          2551 => x"f9",
          2552 => x"34",
          2553 => x"06",
          2554 => x"33",
          2555 => x"5e",
          2556 => x"98",
          2557 => x"ff",
          2558 => x"ea",
          2559 => x"96",
          2560 => x"f9",
          2561 => x"81",
          2562 => x"ac",
          2563 => x"78",
          2564 => x"2e",
          2565 => x"5f",
          2566 => x"56",
          2567 => x"10",
          2568 => x"08",
          2569 => x"80",
          2570 => x"0b",
          2571 => x"04",
          2572 => x"33",
          2573 => x"33",
          2574 => x"11",
          2575 => x"ba",
          2576 => x"70",
          2577 => x"33",
          2578 => x"7f",
          2579 => x"7a",
          2580 => x"7a",
          2581 => x"5c",
          2582 => x"a3",
          2583 => x"33",
          2584 => x"22",
          2585 => x"56",
          2586 => x"83",
          2587 => x"5a",
          2588 => x"b0",
          2589 => x"70",
          2590 => x"83",
          2591 => x"5b",
          2592 => x"33",
          2593 => x"05",
          2594 => x"7a",
          2595 => x"33",
          2596 => x"56",
          2597 => x"70",
          2598 => x"26",
          2599 => x"84",
          2600 => x"72",
          2601 => x"72",
          2602 => x"54",
          2603 => x"a8",
          2604 => x"84",
          2605 => x"83",
          2606 => x"5e",
          2607 => x"be",
          2608 => x"71",
          2609 => x"33",
          2610 => x"b8",
          2611 => x"f9",
          2612 => x"72",
          2613 => x"83",
          2614 => x"34",
          2615 => x"5b",
          2616 => x"77",
          2617 => x"82",
          2618 => x"84",
          2619 => x"83",
          2620 => x"88",
          2621 => x"33",
          2622 => x"56",
          2623 => x"8e",
          2624 => x"9c",
          2625 => x"33",
          2626 => x"34",
          2627 => x"33",
          2628 => x"80",
          2629 => x"42",
          2630 => x"51",
          2631 => x"08",
          2632 => x"8d",
          2633 => x"b9",
          2634 => x"41",
          2635 => x"b9",
          2636 => x"f9",
          2637 => x"1c",
          2638 => x"84",
          2639 => x"5b",
          2640 => x"80",
          2641 => x"bd",
          2642 => x"5b",
          2643 => x"a3",
          2644 => x"33",
          2645 => x"22",
          2646 => x"56",
          2647 => x"f9",
          2648 => x"5e",
          2649 => x"b0",
          2650 => x"70",
          2651 => x"83",
          2652 => x"41",
          2653 => x"33",
          2654 => x"70",
          2655 => x"26",
          2656 => x"58",
          2657 => x"75",
          2658 => x"b9",
          2659 => x"7f",
          2660 => x"84",
          2661 => x"52",
          2662 => x"84",
          2663 => x"84",
          2664 => x"84",
          2665 => x"84",
          2666 => x"ba",
          2667 => x"33",
          2668 => x"33",
          2669 => x"33",
          2670 => x"84",
          2671 => x"ff",
          2672 => x"7c",
          2673 => x"38",
          2674 => x"83",
          2675 => x"53",
          2676 => x"52",
          2677 => x"fe",
          2678 => x"81",
          2679 => x"76",
          2680 => x"38",
          2681 => x"fd",
          2682 => x"84",
          2683 => x"ff",
          2684 => x"38",
          2685 => x"11",
          2686 => x"a5",
          2687 => x"05",
          2688 => x"33",
          2689 => x"83",
          2690 => x"71",
          2691 => x"72",
          2692 => x"83",
          2693 => x"b9",
          2694 => x"e7",
          2695 => x"70",
          2696 => x"5d",
          2697 => x"38",
          2698 => x"39",
          2699 => x"f9",
          2700 => x"57",
          2701 => x"17",
          2702 => x"9c",
          2703 => x"83",
          2704 => x"ff",
          2705 => x"84",
          2706 => x"bc",
          2707 => x"33",
          2708 => x"83",
          2709 => x"71",
          2710 => x"72",
          2711 => x"83",
          2712 => x"b9",
          2713 => x"c4",
          2714 => x"99",
          2715 => x"84",
          2716 => x"83",
          2717 => x"87",
          2718 => x"22",
          2719 => x"05",
          2720 => x"90",
          2721 => x"5a",
          2722 => x"92",
          2723 => x"34",
          2724 => x"5a",
          2725 => x"b9",
          2726 => x"81",
          2727 => x"f8",
          2728 => x"8d",
          2729 => x"38",
          2730 => x"33",
          2731 => x"ff",
          2732 => x"83",
          2733 => x"34",
          2734 => x"57",
          2735 => x"b9",
          2736 => x"61",
          2737 => x"59",
          2738 => x"75",
          2739 => x"f4",
          2740 => x"e2",
          2741 => x"57",
          2742 => x"76",
          2743 => x"53",
          2744 => x"c2",
          2745 => x"84",
          2746 => x"39",
          2747 => x"57",
          2748 => x"e0",
          2749 => x"75",
          2750 => x"51",
          2751 => x"b9",
          2752 => x"b7",
          2753 => x"70",
          2754 => x"ff",
          2755 => x"ff",
          2756 => x"40",
          2757 => x"7e",
          2758 => x"f9",
          2759 => x"18",
          2760 => x"77",
          2761 => x"b8",
          2762 => x"60",
          2763 => x"83",
          2764 => x"b9",
          2765 => x"ef",
          2766 => x"ff",
          2767 => x"94",
          2768 => x"80",
          2769 => x"bd",
          2770 => x"a0",
          2771 => x"40",
          2772 => x"ff",
          2773 => x"59",
          2774 => x"f0",
          2775 => x"7c",
          2776 => x"fe",
          2777 => x"76",
          2778 => x"75",
          2779 => x"06",
          2780 => x"24",
          2781 => x"56",
          2782 => x"16",
          2783 => x"81",
          2784 => x"57",
          2785 => x"75",
          2786 => x"06",
          2787 => x"58",
          2788 => x"b0",
          2789 => x"ff",
          2790 => x"42",
          2791 => x"84",
          2792 => x"33",
          2793 => x"70",
          2794 => x"05",
          2795 => x"34",
          2796 => x"b7",
          2797 => x"40",
          2798 => x"38",
          2799 => x"88",
          2800 => x"34",
          2801 => x"70",
          2802 => x"b8",
          2803 => x"71",
          2804 => x"78",
          2805 => x"84",
          2806 => x"87",
          2807 => x"33",
          2808 => x"80",
          2809 => x"84",
          2810 => x"79",
          2811 => x"22",
          2812 => x"8b",
          2813 => x"76",
          2814 => x"79",
          2815 => x"ed",
          2816 => x"60",
          2817 => x"06",
          2818 => x"7b",
          2819 => x"76",
          2820 => x"70",
          2821 => x"80",
          2822 => x"b0",
          2823 => x"5d",
          2824 => x"57",
          2825 => x"33",
          2826 => x"71",
          2827 => x"59",
          2828 => x"38",
          2829 => x"7d",
          2830 => x"77",
          2831 => x"84",
          2832 => x"ff",
          2833 => x"ba",
          2834 => x"59",
          2835 => x"76",
          2836 => x"05",
          2837 => x"76",
          2838 => x"b8",
          2839 => x"a0",
          2840 => x"70",
          2841 => x"76",
          2842 => x"e0",
          2843 => x"05",
          2844 => x"27",
          2845 => x"70",
          2846 => x"39",
          2847 => x"06",
          2848 => x"84",
          2849 => x"f0",
          2850 => x"f2",
          2851 => x"70",
          2852 => x"39",
          2853 => x"b8",
          2854 => x"bc",
          2855 => x"ba",
          2856 => x"5f",
          2857 => x"33",
          2858 => x"34",
          2859 => x"56",
          2860 => x"81",
          2861 => x"f9",
          2862 => x"33",
          2863 => x"83",
          2864 => x"b8",
          2865 => x"75",
          2866 => x"f9",
          2867 => x"56",
          2868 => x"39",
          2869 => x"81",
          2870 => x"f4",
          2871 => x"8f",
          2872 => x"ff",
          2873 => x"9f",
          2874 => x"b8",
          2875 => x"33",
          2876 => x"75",
          2877 => x"83",
          2878 => x"c0",
          2879 => x"fe",
          2880 => x"af",
          2881 => x"b8",
          2882 => x"33",
          2883 => x"83",
          2884 => x"f9",
          2885 => x"56",
          2886 => x"39",
          2887 => x"82",
          2888 => x"fe",
          2889 => x"f8",
          2890 => x"fd",
          2891 => x"f0",
          2892 => x"fd",
          2893 => x"f0",
          2894 => x"fd",
          2895 => x"df",
          2896 => x"f9",
          2897 => x"b8",
          2898 => x"75",
          2899 => x"80",
          2900 => x"81",
          2901 => x"84",
          2902 => x"84",
          2903 => x"84",
          2904 => x"ba",
          2905 => x"e8",
          2906 => x"34",
          2907 => x"3d",
          2908 => x"83",
          2909 => x"58",
          2910 => x"b9",
          2911 => x"d8",
          2912 => x"ba",
          2913 => x"08",
          2914 => x"b9",
          2915 => x"0c",
          2916 => x"bd",
          2917 => x"33",
          2918 => x"8d",
          2919 => x"02",
          2920 => x"1e",
          2921 => x"ca",
          2922 => x"80",
          2923 => x"f9",
          2924 => x"ff",
          2925 => x"83",
          2926 => x"d0",
          2927 => x"fe",
          2928 => x"f9",
          2929 => x"9f",
          2930 => x"a6",
          2931 => x"84",
          2932 => x"ee",
          2933 => x"ee",
          2934 => x"05",
          2935 => x"58",
          2936 => x"bc",
          2937 => x"ff",
          2938 => x"f3",
          2939 => x"84",
          2940 => x"58",
          2941 => x"83",
          2942 => x"70",
          2943 => x"71",
          2944 => x"05",
          2945 => x"7e",
          2946 => x"83",
          2947 => x"5f",
          2948 => x"79",
          2949 => x"57",
          2950 => x"b7",
          2951 => x"98",
          2952 => x"ba",
          2953 => x"57",
          2954 => x"84",
          2955 => x"82",
          2956 => x"f9",
          2957 => x"f9",
          2958 => x"76",
          2959 => x"05",
          2960 => x"5c",
          2961 => x"80",
          2962 => x"ff",
          2963 => x"29",
          2964 => x"27",
          2965 => x"57",
          2966 => x"88",
          2967 => x"34",
          2968 => x"70",
          2969 => x"b8",
          2970 => x"71",
          2971 => x"76",
          2972 => x"33",
          2973 => x"70",
          2974 => x"05",
          2975 => x"34",
          2976 => x"b7",
          2977 => x"41",
          2978 => x"38",
          2979 => x"33",
          2980 => x"34",
          2981 => x"33",
          2982 => x"33",
          2983 => x"76",
          2984 => x"70",
          2985 => x"58",
          2986 => x"79",
          2987 => x"06",
          2988 => x"83",
          2989 => x"34",
          2990 => x"06",
          2991 => x"27",
          2992 => x"f9",
          2993 => x"bd",
          2994 => x"ff",
          2995 => x"ef",
          2996 => x"75",
          2997 => x"38",
          2998 => x"06",
          2999 => x"5d",
          3000 => x"f4",
          3001 => x"56",
          3002 => x"39",
          3003 => x"23",
          3004 => x"75",
          3005 => x"77",
          3006 => x"8d",
          3007 => x"34",
          3008 => x"05",
          3009 => x"38",
          3010 => x"83",
          3011 => x"59",
          3012 => x"d3",
          3013 => x"f9",
          3014 => x"83",
          3015 => x"83",
          3016 => x"0b",
          3017 => x"80",
          3018 => x"39",
          3019 => x"b8",
          3020 => x"83",
          3021 => x"3d",
          3022 => x"82",
          3023 => x"38",
          3024 => x"84",
          3025 => x"76",
          3026 => x"0b",
          3027 => x"04",
          3028 => x"5c",
          3029 => x"81",
          3030 => x"58",
          3031 => x"d6",
          3032 => x"90",
          3033 => x"0c",
          3034 => x"08",
          3035 => x"38",
          3036 => x"70",
          3037 => x"58",
          3038 => x"80",
          3039 => x"83",
          3040 => x"30",
          3041 => x"5d",
          3042 => x"b8",
          3043 => x"f9",
          3044 => x"a3",
          3045 => x"5b",
          3046 => x"83",
          3047 => x"58",
          3048 => x"8c",
          3049 => x"80",
          3050 => x"88",
          3051 => x"75",
          3052 => x"84",
          3053 => x"34",
          3054 => x"55",
          3055 => x"54",
          3056 => x"ff",
          3057 => x"54",
          3058 => x"72",
          3059 => x"83",
          3060 => x"06",
          3061 => x"38",
          3062 => x"f7",
          3063 => x"34",
          3064 => x"5e",
          3065 => x"f7",
          3066 => x"25",
          3067 => x"34",
          3068 => x"81",
          3069 => x"72",
          3070 => x"83",
          3071 => x"53",
          3072 => x"0b",
          3073 => x"f7",
          3074 => x"f7",
          3075 => x"83",
          3076 => x"5c",
          3077 => x"55",
          3078 => x"f7",
          3079 => x"82",
          3080 => x"53",
          3081 => x"f7",
          3082 => x"38",
          3083 => x"ff",
          3084 => x"33",
          3085 => x"74",
          3086 => x"2e",
          3087 => x"33",
          3088 => x"83",
          3089 => x"c0",
          3090 => x"27",
          3091 => x"98",
          3092 => x"81",
          3093 => x"89",
          3094 => x"f7",
          3095 => x"fe",
          3096 => x"8b",
          3097 => x"05",
          3098 => x"08",
          3099 => x"f4",
          3100 => x"5e",
          3101 => x"0b",
          3102 => x"81",
          3103 => x"f8",
          3104 => x"83",
          3105 => x"58",
          3106 => x"be",
          3107 => x"33",
          3108 => x"39",
          3109 => x"2e",
          3110 => x"f4",
          3111 => x"54",
          3112 => x"39",
          3113 => x"81",
          3114 => x"81",
          3115 => x"80",
          3116 => x"38",
          3117 => x"27",
          3118 => x"25",
          3119 => x"81",
          3120 => x"81",
          3121 => x"2b",
          3122 => x"24",
          3123 => x"10",
          3124 => x"83",
          3125 => x"54",
          3126 => x"f7",
          3127 => x"59",
          3128 => x"81",
          3129 => x"59",
          3130 => x"9f",
          3131 => x"54",
          3132 => x"7b",
          3133 => x"76",
          3134 => x"7b",
          3135 => x"38",
          3136 => x"53",
          3137 => x"05",
          3138 => x"83",
          3139 => x"06",
          3140 => x"84",
          3141 => x"f9",
          3142 => x"74",
          3143 => x"52",
          3144 => x"ba",
          3145 => x"76",
          3146 => x"72",
          3147 => x"d4",
          3148 => x"f7",
          3149 => x"0b",
          3150 => x"83",
          3151 => x"f7",
          3152 => x"81",
          3153 => x"fc",
          3154 => x"55",
          3155 => x"81",
          3156 => x"81",
          3157 => x"08",
          3158 => x"08",
          3159 => x"38",
          3160 => x"e0",
          3161 => x"d7",
          3162 => x"34",
          3163 => x"34",
          3164 => x"9e",
          3165 => x"0b",
          3166 => x"08",
          3167 => x"e8",
          3168 => x"42",
          3169 => x"79",
          3170 => x"38",
          3171 => x"38",
          3172 => x"c0",
          3173 => x"81",
          3174 => x"84",
          3175 => x"38",
          3176 => x"ff",
          3177 => x"b8",
          3178 => x"81",
          3179 => x"59",
          3180 => x"ec",
          3181 => x"0b",
          3182 => x"84",
          3183 => x"ff",
          3184 => x"83",
          3185 => x"23",
          3186 => x"53",
          3187 => x"73",
          3188 => x"33",
          3189 => x"53",
          3190 => x"72",
          3191 => x"b7",
          3192 => x"a5",
          3193 => x"54",
          3194 => x"83",
          3195 => x"81",
          3196 => x"f0",
          3197 => x"0d",
          3198 => x"0d",
          3199 => x"f4",
          3200 => x"33",
          3201 => x"52",
          3202 => x"f4",
          3203 => x"16",
          3204 => x"34",
          3205 => x"98",
          3206 => x"87",
          3207 => x"98",
          3208 => x"38",
          3209 => x"08",
          3210 => x"72",
          3211 => x"98",
          3212 => x"27",
          3213 => x"2e",
          3214 => x"08",
          3215 => x"98",
          3216 => x"08",
          3217 => x"15",
          3218 => x"53",
          3219 => x"ff",
          3220 => x"08",
          3221 => x"38",
          3222 => x"76",
          3223 => x"06",
          3224 => x"2e",
          3225 => x"89",
          3226 => x"ff",
          3227 => x"0b",
          3228 => x"8d",
          3229 => x"3d",
          3230 => x"84",
          3231 => x"0b",
          3232 => x"87",
          3233 => x"2a",
          3234 => x"16",
          3235 => x"16",
          3236 => x"16",
          3237 => x"98",
          3238 => x"f4",
          3239 => x"85",
          3240 => x"fe",
          3241 => x"f0",
          3242 => x"08",
          3243 => x"90",
          3244 => x"53",
          3245 => x"73",
          3246 => x"c0",
          3247 => x"27",
          3248 => x"38",
          3249 => x"56",
          3250 => x"56",
          3251 => x"c0",
          3252 => x"54",
          3253 => x"c0",
          3254 => x"f6",
          3255 => x"9c",
          3256 => x"38",
          3257 => x"c0",
          3258 => x"74",
          3259 => x"ff",
          3260 => x"80",
          3261 => x"72",
          3262 => x"ff",
          3263 => x"15",
          3264 => x"71",
          3265 => x"05",
          3266 => x"34",
          3267 => x"ba",
          3268 => x"0b",
          3269 => x"c5",
          3270 => x"3d",
          3271 => x"06",
          3272 => x"52",
          3273 => x"02",
          3274 => x"80",
          3275 => x"2b",
          3276 => x"98",
          3277 => x"83",
          3278 => x"84",
          3279 => x"85",
          3280 => x"83",
          3281 => x"80",
          3282 => x"27",
          3283 => x"33",
          3284 => x"72",
          3285 => x"55",
          3286 => x"08",
          3287 => x"83",
          3288 => x"81",
          3289 => x"e8",
          3290 => x"f4",
          3291 => x"54",
          3292 => x"c0",
          3293 => x"f6",
          3294 => x"9c",
          3295 => x"38",
          3296 => x"c0",
          3297 => x"74",
          3298 => x"ff",
          3299 => x"9c",
          3300 => x"c0",
          3301 => x"9c",
          3302 => x"81",
          3303 => x"53",
          3304 => x"81",
          3305 => x"a4",
          3306 => x"a9",
          3307 => x"38",
          3308 => x"ff",
          3309 => x"70",
          3310 => x"38",
          3311 => x"0d",
          3312 => x"58",
          3313 => x"ff",
          3314 => x"38",
          3315 => x"fe",
          3316 => x"0c",
          3317 => x"83",
          3318 => x"34",
          3319 => x"56",
          3320 => x"86",
          3321 => x"9c",
          3322 => x"ce",
          3323 => x"08",
          3324 => x"72",
          3325 => x"87",
          3326 => x"74",
          3327 => x"db",
          3328 => x"ff",
          3329 => x"71",
          3330 => x"87",
          3331 => x"05",
          3332 => x"87",
          3333 => x"2e",
          3334 => x"98",
          3335 => x"87",
          3336 => x"87",
          3337 => x"70",
          3338 => x"ff",
          3339 => x"38",
          3340 => x"d8",
          3341 => x"ff",
          3342 => x"0d",
          3343 => x"3f",
          3344 => x"84",
          3345 => x"2a",
          3346 => x"2b",
          3347 => x"71",
          3348 => x"11",
          3349 => x"2b",
          3350 => x"53",
          3351 => x"53",
          3352 => x"16",
          3353 => x"8b",
          3354 => x"70",
          3355 => x"71",
          3356 => x"59",
          3357 => x"38",
          3358 => x"8b",
          3359 => x"76",
          3360 => x"86",
          3361 => x"73",
          3362 => x"70",
          3363 => x"71",
          3364 => x"55",
          3365 => x"71",
          3366 => x"16",
          3367 => x"0b",
          3368 => x"53",
          3369 => x"34",
          3370 => x"81",
          3371 => x"80",
          3372 => x"52",
          3373 => x"34",
          3374 => x"87",
          3375 => x"2b",
          3376 => x"17",
          3377 => x"2a",
          3378 => x"71",
          3379 => x"84",
          3380 => x"33",
          3381 => x"83",
          3382 => x"05",
          3383 => x"88",
          3384 => x"59",
          3385 => x"13",
          3386 => x"33",
          3387 => x"81",
          3388 => x"5a",
          3389 => x"13",
          3390 => x"70",
          3391 => x"71",
          3392 => x"81",
          3393 => x"83",
          3394 => x"7b",
          3395 => x"5a",
          3396 => x"73",
          3397 => x"70",
          3398 => x"8b",
          3399 => x"70",
          3400 => x"07",
          3401 => x"5f",
          3402 => x"77",
          3403 => x"b9",
          3404 => x"83",
          3405 => x"2b",
          3406 => x"33",
          3407 => x"58",
          3408 => x"70",
          3409 => x"81",
          3410 => x"80",
          3411 => x"54",
          3412 => x"84",
          3413 => x"81",
          3414 => x"2b",
          3415 => x"15",
          3416 => x"2a",
          3417 => x"53",
          3418 => x"34",
          3419 => x"79",
          3420 => x"80",
          3421 => x"38",
          3422 => x"0d",
          3423 => x"fc",
          3424 => x"23",
          3425 => x"ff",
          3426 => x"b9",
          3427 => x"0b",
          3428 => x"54",
          3429 => x"15",
          3430 => x"86",
          3431 => x"84",
          3432 => x"ff",
          3433 => x"ff",
          3434 => x"55",
          3435 => x"17",
          3436 => x"10",
          3437 => x"05",
          3438 => x"0b",
          3439 => x"3d",
          3440 => x"84",
          3441 => x"2a",
          3442 => x"51",
          3443 => x"b9",
          3444 => x"33",
          3445 => x"5a",
          3446 => x"80",
          3447 => x"10",
          3448 => x"88",
          3449 => x"79",
          3450 => x"7a",
          3451 => x"72",
          3452 => x"85",
          3453 => x"33",
          3454 => x"57",
          3455 => x"ff",
          3456 => x"80",
          3457 => x"81",
          3458 => x"81",
          3459 => x"59",
          3460 => x"59",
          3461 => x"38",
          3462 => x"38",
          3463 => x"16",
          3464 => x"80",
          3465 => x"56",
          3466 => x"15",
          3467 => x"88",
          3468 => x"75",
          3469 => x"70",
          3470 => x"88",
          3471 => x"f8",
          3472 => x"06",
          3473 => x"59",
          3474 => x"81",
          3475 => x"84",
          3476 => x"34",
          3477 => x"08",
          3478 => x"33",
          3479 => x"74",
          3480 => x"84",
          3481 => x"b9",
          3482 => x"86",
          3483 => x"2b",
          3484 => x"59",
          3485 => x"34",
          3486 => x"11",
          3487 => x"71",
          3488 => x"5c",
          3489 => x"87",
          3490 => x"16",
          3491 => x"12",
          3492 => x"2a",
          3493 => x"34",
          3494 => x"08",
          3495 => x"8c",
          3496 => x"33",
          3497 => x"83",
          3498 => x"85",
          3499 => x"88",
          3500 => x"74",
          3501 => x"84",
          3502 => x"33",
          3503 => x"83",
          3504 => x"87",
          3505 => x"88",
          3506 => x"57",
          3507 => x"1a",
          3508 => x"33",
          3509 => x"81",
          3510 => x"57",
          3511 => x"18",
          3512 => x"05",
          3513 => x"79",
          3514 => x"80",
          3515 => x"38",
          3516 => x"0d",
          3517 => x"ba",
          3518 => x"3d",
          3519 => x"b9",
          3520 => x"f8",
          3521 => x"84",
          3522 => x"84",
          3523 => x"81",
          3524 => x"08",
          3525 => x"85",
          3526 => x"76",
          3527 => x"34",
          3528 => x"22",
          3529 => x"83",
          3530 => x"51",
          3531 => x"89",
          3532 => x"10",
          3533 => x"f8",
          3534 => x"81",
          3535 => x"80",
          3536 => x"ed",
          3537 => x"70",
          3538 => x"76",
          3539 => x"2e",
          3540 => x"d7",
          3541 => x"38",
          3542 => x"70",
          3543 => x"83",
          3544 => x"2a",
          3545 => x"2b",
          3546 => x"71",
          3547 => x"83",
          3548 => x"fc",
          3549 => x"33",
          3550 => x"70",
          3551 => x"45",
          3552 => x"48",
          3553 => x"24",
          3554 => x"16",
          3555 => x"10",
          3556 => x"71",
          3557 => x"5c",
          3558 => x"85",
          3559 => x"38",
          3560 => x"a2",
          3561 => x"60",
          3562 => x"38",
          3563 => x"f7",
          3564 => x"33",
          3565 => x"7a",
          3566 => x"98",
          3567 => x"59",
          3568 => x"24",
          3569 => x"33",
          3570 => x"83",
          3571 => x"87",
          3572 => x"2b",
          3573 => x"15",
          3574 => x"2a",
          3575 => x"53",
          3576 => x"79",
          3577 => x"70",
          3578 => x"71",
          3579 => x"05",
          3580 => x"88",
          3581 => x"5e",
          3582 => x"16",
          3583 => x"fc",
          3584 => x"71",
          3585 => x"70",
          3586 => x"79",
          3587 => x"fc",
          3588 => x"12",
          3589 => x"07",
          3590 => x"71",
          3591 => x"5c",
          3592 => x"79",
          3593 => x"fc",
          3594 => x"33",
          3595 => x"74",
          3596 => x"71",
          3597 => x"5c",
          3598 => x"82",
          3599 => x"b9",
          3600 => x"83",
          3601 => x"57",
          3602 => x"5a",
          3603 => x"c4",
          3604 => x"84",
          3605 => x"ff",
          3606 => x"26",
          3607 => x"ba",
          3608 => x"ff",
          3609 => x"80",
          3610 => x"80",
          3611 => x"fe",
          3612 => x"5e",
          3613 => x"34",
          3614 => x"1e",
          3615 => x"b9",
          3616 => x"81",
          3617 => x"08",
          3618 => x"80",
          3619 => x"70",
          3620 => x"88",
          3621 => x"b9",
          3622 => x"b9",
          3623 => x"60",
          3624 => x"34",
          3625 => x"d3",
          3626 => x"7e",
          3627 => x"7f",
          3628 => x"08",
          3629 => x"04",
          3630 => x"83",
          3631 => x"70",
          3632 => x"07",
          3633 => x"48",
          3634 => x"60",
          3635 => x"08",
          3636 => x"82",
          3637 => x"b9",
          3638 => x"12",
          3639 => x"2b",
          3640 => x"83",
          3641 => x"5c",
          3642 => x"82",
          3643 => x"60",
          3644 => x"08",
          3645 => x"1c",
          3646 => x"84",
          3647 => x"fd",
          3648 => x"ff",
          3649 => x"77",
          3650 => x"83",
          3651 => x"18",
          3652 => x"10",
          3653 => x"71",
          3654 => x"5e",
          3655 => x"80",
          3656 => x"61",
          3657 => x"24",
          3658 => x"06",
          3659 => x"fe",
          3660 => x"b9",
          3661 => x"f8",
          3662 => x"84",
          3663 => x"84",
          3664 => x"81",
          3665 => x"08",
          3666 => x"85",
          3667 => x"7e",
          3668 => x"34",
          3669 => x"22",
          3670 => x"83",
          3671 => x"56",
          3672 => x"73",
          3673 => x"22",
          3674 => x"08",
          3675 => x"82",
          3676 => x"fc",
          3677 => x"38",
          3678 => x"7b",
          3679 => x"76",
          3680 => x"ea",
          3681 => x"8c",
          3682 => x"82",
          3683 => x"2b",
          3684 => x"11",
          3685 => x"71",
          3686 => x"33",
          3687 => x"70",
          3688 => x"46",
          3689 => x"84",
          3690 => x"84",
          3691 => x"33",
          3692 => x"83",
          3693 => x"87",
          3694 => x"88",
          3695 => x"5d",
          3696 => x"64",
          3697 => x"16",
          3698 => x"2b",
          3699 => x"2a",
          3700 => x"79",
          3701 => x"70",
          3702 => x"71",
          3703 => x"05",
          3704 => x"2b",
          3705 => x"40",
          3706 => x"75",
          3707 => x"70",
          3708 => x"8b",
          3709 => x"82",
          3710 => x"2b",
          3711 => x"5b",
          3712 => x"34",
          3713 => x"08",
          3714 => x"33",
          3715 => x"56",
          3716 => x"7e",
          3717 => x"3f",
          3718 => x"78",
          3719 => x"99",
          3720 => x"fc",
          3721 => x"23",
          3722 => x"ff",
          3723 => x"b9",
          3724 => x"0b",
          3725 => x"55",
          3726 => x"16",
          3727 => x"86",
          3728 => x"84",
          3729 => x"ff",
          3730 => x"ff",
          3731 => x"44",
          3732 => x"1f",
          3733 => x"10",
          3734 => x"05",
          3735 => x"0b",
          3736 => x"3f",
          3737 => x"33",
          3738 => x"83",
          3739 => x"85",
          3740 => x"88",
          3741 => x"76",
          3742 => x"05",
          3743 => x"84",
          3744 => x"2b",
          3745 => x"14",
          3746 => x"07",
          3747 => x"59",
          3748 => x"34",
          3749 => x"fc",
          3750 => x"71",
          3751 => x"70",
          3752 => x"78",
          3753 => x"fc",
          3754 => x"33",
          3755 => x"74",
          3756 => x"88",
          3757 => x"f8",
          3758 => x"5d",
          3759 => x"7f",
          3760 => x"84",
          3761 => x"81",
          3762 => x"2b",
          3763 => x"33",
          3764 => x"06",
          3765 => x"46",
          3766 => x"60",
          3767 => x"06",
          3768 => x"87",
          3769 => x"2b",
          3770 => x"19",
          3771 => x"2a",
          3772 => x"84",
          3773 => x"b9",
          3774 => x"85",
          3775 => x"2b",
          3776 => x"15",
          3777 => x"2a",
          3778 => x"56",
          3779 => x"87",
          3780 => x"70",
          3781 => x"07",
          3782 => x"5b",
          3783 => x"81",
          3784 => x"1f",
          3785 => x"2b",
          3786 => x"33",
          3787 => x"70",
          3788 => x"05",
          3789 => x"58",
          3790 => x"34",
          3791 => x"08",
          3792 => x"71",
          3793 => x"05",
          3794 => x"2b",
          3795 => x"2a",
          3796 => x"55",
          3797 => x"84",
          3798 => x"33",
          3799 => x"83",
          3800 => x"87",
          3801 => x"2b",
          3802 => x"15",
          3803 => x"2a",
          3804 => x"53",
          3805 => x"34",
          3806 => x"08",
          3807 => x"33",
          3808 => x"74",
          3809 => x"71",
          3810 => x"42",
          3811 => x"86",
          3812 => x"b9",
          3813 => x"33",
          3814 => x"06",
          3815 => x"76",
          3816 => x"b9",
          3817 => x"83",
          3818 => x"2b",
          3819 => x"33",
          3820 => x"41",
          3821 => x"79",
          3822 => x"b9",
          3823 => x"12",
          3824 => x"07",
          3825 => x"33",
          3826 => x"41",
          3827 => x"79",
          3828 => x"84",
          3829 => x"33",
          3830 => x"66",
          3831 => x"52",
          3832 => x"fe",
          3833 => x"1e",
          3834 => x"83",
          3835 => x"d5",
          3836 => x"71",
          3837 => x"05",
          3838 => x"88",
          3839 => x"5d",
          3840 => x"34",
          3841 => x"fc",
          3842 => x"12",
          3843 => x"07",
          3844 => x"33",
          3845 => x"5b",
          3846 => x"73",
          3847 => x"05",
          3848 => x"33",
          3849 => x"81",
          3850 => x"5f",
          3851 => x"16",
          3852 => x"70",
          3853 => x"71",
          3854 => x"81",
          3855 => x"83",
          3856 => x"63",
          3857 => x"5e",
          3858 => x"7b",
          3859 => x"70",
          3860 => x"8b",
          3861 => x"70",
          3862 => x"07",
          3863 => x"47",
          3864 => x"7f",
          3865 => x"83",
          3866 => x"7e",
          3867 => x"ba",
          3868 => x"80",
          3869 => x"84",
          3870 => x"3f",
          3871 => x"61",
          3872 => x"39",
          3873 => x"b9",
          3874 => x"b7",
          3875 => x"84",
          3876 => x"77",
          3877 => x"08",
          3878 => x"e6",
          3879 => x"8c",
          3880 => x"84",
          3881 => x"84",
          3882 => x"a0",
          3883 => x"80",
          3884 => x"51",
          3885 => x"08",
          3886 => x"16",
          3887 => x"84",
          3888 => x"84",
          3889 => x"34",
          3890 => x"fc",
          3891 => x"fe",
          3892 => x"06",
          3893 => x"74",
          3894 => x"84",
          3895 => x"84",
          3896 => x"55",
          3897 => x"15",
          3898 => x"c6",
          3899 => x"02",
          3900 => x"72",
          3901 => x"33",
          3902 => x"3d",
          3903 => x"05",
          3904 => x"9d",
          3905 => x"ba",
          3906 => x"87",
          3907 => x"84",
          3908 => x"ba",
          3909 => x"3d",
          3910 => x"af",
          3911 => x"54",
          3912 => x"88",
          3913 => x"83",
          3914 => x"0b",
          3915 => x"75",
          3916 => x"ba",
          3917 => x"80",
          3918 => x"08",
          3919 => x"d6",
          3920 => x"73",
          3921 => x"55",
          3922 => x"0d",
          3923 => x"81",
          3924 => x"26",
          3925 => x"0d",
          3926 => x"05",
          3927 => x"76",
          3928 => x"17",
          3929 => x"55",
          3930 => x"87",
          3931 => x"52",
          3932 => x"8c",
          3933 => x"2e",
          3934 => x"54",
          3935 => x"38",
          3936 => x"80",
          3937 => x"74",
          3938 => x"04",
          3939 => x"ff",
          3940 => x"ff",
          3941 => x"78",
          3942 => x"88",
          3943 => x"81",
          3944 => x"ba",
          3945 => x"54",
          3946 => x"87",
          3947 => x"73",
          3948 => x"38",
          3949 => x"72",
          3950 => x"04",
          3951 => x"ba",
          3952 => x"80",
          3953 => x"0c",
          3954 => x"87",
          3955 => x"cd",
          3956 => x"06",
          3957 => x"87",
          3958 => x"38",
          3959 => x"ca",
          3960 => x"8c",
          3961 => x"73",
          3962 => x"82",
          3963 => x"39",
          3964 => x"83",
          3965 => x"77",
          3966 => x"33",
          3967 => x"80",
          3968 => x"fe",
          3969 => x"2e",
          3970 => x"8c",
          3971 => x"b4",
          3972 => x"81",
          3973 => x"81",
          3974 => x"09",
          3975 => x"08",
          3976 => x"a8",
          3977 => x"ba",
          3978 => x"76",
          3979 => x"55",
          3980 => x"8e",
          3981 => x"52",
          3982 => x"76",
          3983 => x"09",
          3984 => x"33",
          3985 => x"fe",
          3986 => x"7a",
          3987 => x"57",
          3988 => x"80",
          3989 => x"aa",
          3990 => x"7a",
          3991 => x"80",
          3992 => x"0b",
          3993 => x"9c",
          3994 => x"19",
          3995 => x"34",
          3996 => x"94",
          3997 => x"34",
          3998 => x"19",
          3999 => x"a2",
          4000 => x"84",
          4001 => x"7a",
          4002 => x"55",
          4003 => x"2a",
          4004 => x"98",
          4005 => x"a4",
          4006 => x"0c",
          4007 => x"81",
          4008 => x"84",
          4009 => x"18",
          4010 => x"8c",
          4011 => x"b2",
          4012 => x"08",
          4013 => x"38",
          4014 => x"81",
          4015 => x"3d",
          4016 => x"74",
          4017 => x"24",
          4018 => x"81",
          4019 => x"70",
          4020 => x"5a",
          4021 => x"b0",
          4022 => x"2e",
          4023 => x"54",
          4024 => x"33",
          4025 => x"08",
          4026 => x"5b",
          4027 => x"38",
          4028 => x"33",
          4029 => x"08",
          4030 => x"08",
          4031 => x"18",
          4032 => x"2e",
          4033 => x"54",
          4034 => x"33",
          4035 => x"08",
          4036 => x"5a",
          4037 => x"38",
          4038 => x"33",
          4039 => x"06",
          4040 => x"5d",
          4041 => x"06",
          4042 => x"04",
          4043 => x"59",
          4044 => x"80",
          4045 => x"5b",
          4046 => x"c2",
          4047 => x"52",
          4048 => x"84",
          4049 => x"ff",
          4050 => x"79",
          4051 => x"06",
          4052 => x"71",
          4053 => x"8c",
          4054 => x"74",
          4055 => x"38",
          4056 => x"59",
          4057 => x"80",
          4058 => x"5b",
          4059 => x"81",
          4060 => x"52",
          4061 => x"84",
          4062 => x"ff",
          4063 => x"79",
          4064 => x"fc",
          4065 => x"33",
          4066 => x"88",
          4067 => x"07",
          4068 => x"ff",
          4069 => x"0c",
          4070 => x"3d",
          4071 => x"53",
          4072 => x"52",
          4073 => x"ba",
          4074 => x"fe",
          4075 => x"18",
          4076 => x"31",
          4077 => x"a0",
          4078 => x"17",
          4079 => x"06",
          4080 => x"08",
          4081 => x"81",
          4082 => x"5a",
          4083 => x"08",
          4084 => x"33",
          4085 => x"8c",
          4086 => x"81",
          4087 => x"34",
          4088 => x"5d",
          4089 => x"82",
          4090 => x"cb",
          4091 => x"de",
          4092 => x"b8",
          4093 => x"5c",
          4094 => x"8c",
          4095 => x"ff",
          4096 => x"34",
          4097 => x"84",
          4098 => x"18",
          4099 => x"33",
          4100 => x"fd",
          4101 => x"a0",
          4102 => x"17",
          4103 => x"fd",
          4104 => x"53",
          4105 => x"52",
          4106 => x"ba",
          4107 => x"fb",
          4108 => x"18",
          4109 => x"31",
          4110 => x"a0",
          4111 => x"17",
          4112 => x"06",
          4113 => x"08",
          4114 => x"81",
          4115 => x"5a",
          4116 => x"08",
          4117 => x"81",
          4118 => x"86",
          4119 => x"fa",
          4120 => x"64",
          4121 => x"27",
          4122 => x"95",
          4123 => x"96",
          4124 => x"74",
          4125 => x"ba",
          4126 => x"88",
          4127 => x"0b",
          4128 => x"2e",
          4129 => x"5b",
          4130 => x"83",
          4131 => x"19",
          4132 => x"3f",
          4133 => x"38",
          4134 => x"0c",
          4135 => x"10",
          4136 => x"ff",
          4137 => x"34",
          4138 => x"34",
          4139 => x"ba",
          4140 => x"83",
          4141 => x"75",
          4142 => x"80",
          4143 => x"78",
          4144 => x"7c",
          4145 => x"06",
          4146 => x"b8",
          4147 => x"8e",
          4148 => x"85",
          4149 => x"1a",
          4150 => x"75",
          4151 => x"b8",
          4152 => x"8f",
          4153 => x"41",
          4154 => x"88",
          4155 => x"90",
          4156 => x"98",
          4157 => x"0b",
          4158 => x"81",
          4159 => x"08",
          4160 => x"76",
          4161 => x"1a",
          4162 => x"2e",
          4163 => x"54",
          4164 => x"33",
          4165 => x"08",
          4166 => x"5c",
          4167 => x"fd",
          4168 => x"b8",
          4169 => x"5f",
          4170 => x"38",
          4171 => x"33",
          4172 => x"77",
          4173 => x"89",
          4174 => x"0b",
          4175 => x"2e",
          4176 => x"b8",
          4177 => x"57",
          4178 => x"8c",
          4179 => x"c7",
          4180 => x"34",
          4181 => x"31",
          4182 => x"5b",
          4183 => x"38",
          4184 => x"82",
          4185 => x"52",
          4186 => x"84",
          4187 => x"ff",
          4188 => x"77",
          4189 => x"19",
          4190 => x"7c",
          4191 => x"81",
          4192 => x"5c",
          4193 => x"34",
          4194 => x"b8",
          4195 => x"5d",
          4196 => x"8c",
          4197 => x"88",
          4198 => x"34",
          4199 => x"31",
          4200 => x"5d",
          4201 => x"ca",
          4202 => x"2e",
          4203 => x"54",
          4204 => x"33",
          4205 => x"aa",
          4206 => x"70",
          4207 => x"ad",
          4208 => x"7d",
          4209 => x"84",
          4210 => x"19",
          4211 => x"1b",
          4212 => x"56",
          4213 => x"82",
          4214 => x"81",
          4215 => x"1f",
          4216 => x"ed",
          4217 => x"81",
          4218 => x"81",
          4219 => x"81",
          4220 => x"09",
          4221 => x"8c",
          4222 => x"70",
          4223 => x"84",
          4224 => x"7e",
          4225 => x"33",
          4226 => x"fa",
          4227 => x"76",
          4228 => x"3f",
          4229 => x"79",
          4230 => x"51",
          4231 => x"39",
          4232 => x"05",
          4233 => x"58",
          4234 => x"5a",
          4235 => x"7e",
          4236 => x"2b",
          4237 => x"83",
          4238 => x"06",
          4239 => x"5f",
          4240 => x"2a",
          4241 => x"2a",
          4242 => x"2a",
          4243 => x"39",
          4244 => x"5b",
          4245 => x"19",
          4246 => x"38",
          4247 => x"38",
          4248 => x"80",
          4249 => x"81",
          4250 => x"9c",
          4251 => x"56",
          4252 => x"52",
          4253 => x"8c",
          4254 => x"58",
          4255 => x"38",
          4256 => x"70",
          4257 => x"51",
          4258 => x"75",
          4259 => x"38",
          4260 => x"8c",
          4261 => x"39",
          4262 => x"7a",
          4263 => x"55",
          4264 => x"38",
          4265 => x"8c",
          4266 => x"08",
          4267 => x"7a",
          4268 => x"9c",
          4269 => x"56",
          4270 => x"80",
          4271 => x"81",
          4272 => x"70",
          4273 => x"7b",
          4274 => x"51",
          4275 => x"ba",
          4276 => x"19",
          4277 => x"38",
          4278 => x"38",
          4279 => x"75",
          4280 => x"75",
          4281 => x"ba",
          4282 => x"70",
          4283 => x"56",
          4284 => x"80",
          4285 => x"19",
          4286 => x"58",
          4287 => x"94",
          4288 => x"5a",
          4289 => x"84",
          4290 => x"80",
          4291 => x"0d",
          4292 => x"da",
          4293 => x"75",
          4294 => x"3f",
          4295 => x"39",
          4296 => x"0c",
          4297 => x"81",
          4298 => x"b6",
          4299 => x"08",
          4300 => x"26",
          4301 => x"72",
          4302 => x"88",
          4303 => x"76",
          4304 => x"38",
          4305 => x"18",
          4306 => x"38",
          4307 => x"94",
          4308 => x"56",
          4309 => x"2a",
          4310 => x"06",
          4311 => x"56",
          4312 => x"0d",
          4313 => x"8a",
          4314 => x"74",
          4315 => x"22",
          4316 => x"27",
          4317 => x"15",
          4318 => x"73",
          4319 => x"71",
          4320 => x"78",
          4321 => x"52",
          4322 => x"8c",
          4323 => x"2e",
          4324 => x"08",
          4325 => x"53",
          4326 => x"91",
          4327 => x"27",
          4328 => x"84",
          4329 => x"f3",
          4330 => x"08",
          4331 => x"0a",
          4332 => x"18",
          4333 => x"74",
          4334 => x"06",
          4335 => x"18",
          4336 => x"85",
          4337 => x"76",
          4338 => x"0c",
          4339 => x"05",
          4340 => x"ba",
          4341 => x"98",
          4342 => x"7a",
          4343 => x"75",
          4344 => x"ba",
          4345 => x"84",
          4346 => x"56",
          4347 => x"38",
          4348 => x"26",
          4349 => x"98",
          4350 => x"f9",
          4351 => x"87",
          4352 => x"ff",
          4353 => x"08",
          4354 => x"84",
          4355 => x"38",
          4356 => x"5f",
          4357 => x"9c",
          4358 => x"5c",
          4359 => x"22",
          4360 => x"5d",
          4361 => x"58",
          4362 => x"70",
          4363 => x"74",
          4364 => x"55",
          4365 => x"54",
          4366 => x"33",
          4367 => x"08",
          4368 => x"39",
          4369 => x"ba",
          4370 => x"54",
          4371 => x"53",
          4372 => x"3f",
          4373 => x"84",
          4374 => x"19",
          4375 => x"a0",
          4376 => x"19",
          4377 => x"06",
          4378 => x"08",
          4379 => x"81",
          4380 => x"c5",
          4381 => x"ff",
          4382 => x"81",
          4383 => x"fe",
          4384 => x"56",
          4385 => x"38",
          4386 => x"1b",
          4387 => x"f8",
          4388 => x"8f",
          4389 => x"66",
          4390 => x"81",
          4391 => x"5e",
          4392 => x"19",
          4393 => x"08",
          4394 => x"33",
          4395 => x"81",
          4396 => x"53",
          4397 => x"e1",
          4398 => x"2e",
          4399 => x"b4",
          4400 => x"38",
          4401 => x"76",
          4402 => x"33",
          4403 => x"41",
          4404 => x"32",
          4405 => x"72",
          4406 => x"45",
          4407 => x"7a",
          4408 => x"81",
          4409 => x"38",
          4410 => x"fa",
          4411 => x"84",
          4412 => x"1c",
          4413 => x"84",
          4414 => x"81",
          4415 => x"81",
          4416 => x"57",
          4417 => x"81",
          4418 => x"08",
          4419 => x"1a",
          4420 => x"5b",
          4421 => x"38",
          4422 => x"09",
          4423 => x"b4",
          4424 => x"7e",
          4425 => x"3f",
          4426 => x"2e",
          4427 => x"86",
          4428 => x"93",
          4429 => x"06",
          4430 => x"0c",
          4431 => x"38",
          4432 => x"39",
          4433 => x"06",
          4434 => x"80",
          4435 => x"8c",
          4436 => x"fd",
          4437 => x"77",
          4438 => x"19",
          4439 => x"71",
          4440 => x"ff",
          4441 => x"06",
          4442 => x"76",
          4443 => x"78",
          4444 => x"88",
          4445 => x"2e",
          4446 => x"ff",
          4447 => x"5c",
          4448 => x"81",
          4449 => x"77",
          4450 => x"57",
          4451 => x"fe",
          4452 => x"05",
          4453 => x"81",
          4454 => x"75",
          4455 => x"ff",
          4456 => x"7c",
          4457 => x"81",
          4458 => x"5a",
          4459 => x"06",
          4460 => x"38",
          4461 => x"0b",
          4462 => x"0c",
          4463 => x"63",
          4464 => x"51",
          4465 => x"5a",
          4466 => x"81",
          4467 => x"1d",
          4468 => x"56",
          4469 => x"82",
          4470 => x"55",
          4471 => x"df",
          4472 => x"52",
          4473 => x"84",
          4474 => x"ff",
          4475 => x"76",
          4476 => x"08",
          4477 => x"84",
          4478 => x"70",
          4479 => x"1d",
          4480 => x"38",
          4481 => x"8f",
          4482 => x"38",
          4483 => x"aa",
          4484 => x"74",
          4485 => x"78",
          4486 => x"05",
          4487 => x"56",
          4488 => x"80",
          4489 => x"57",
          4490 => x"59",
          4491 => x"78",
          4492 => x"31",
          4493 => x"80",
          4494 => x"e1",
          4495 => x"1d",
          4496 => x"3f",
          4497 => x"8c",
          4498 => x"84",
          4499 => x"81",
          4500 => x"81",
          4501 => x"57",
          4502 => x"81",
          4503 => x"08",
          4504 => x"1c",
          4505 => x"59",
          4506 => x"38",
          4507 => x"09",
          4508 => x"b4",
          4509 => x"7d",
          4510 => x"3f",
          4511 => x"fd",
          4512 => x"2a",
          4513 => x"38",
          4514 => x"80",
          4515 => x"81",
          4516 => x"ac",
          4517 => x"2e",
          4518 => x"80",
          4519 => x"ba",
          4520 => x"80",
          4521 => x"75",
          4522 => x"5d",
          4523 => x"39",
          4524 => x"09",
          4525 => x"9b",
          4526 => x"2b",
          4527 => x"38",
          4528 => x"f3",
          4529 => x"83",
          4530 => x"11",
          4531 => x"52",
          4532 => x"38",
          4533 => x"76",
          4534 => x"8c",
          4535 => x"53",
          4536 => x"f6",
          4537 => x"09",
          4538 => x"81",
          4539 => x"38",
          4540 => x"56",
          4541 => x"80",
          4542 => x"70",
          4543 => x"ff",
          4544 => x"fe",
          4545 => x"0c",
          4546 => x"ff",
          4547 => x"fe",
          4548 => x"08",
          4549 => x"58",
          4550 => x"b5",
          4551 => x"57",
          4552 => x"81",
          4553 => x"56",
          4554 => x"1f",
          4555 => x"55",
          4556 => x"70",
          4557 => x"74",
          4558 => x"70",
          4559 => x"82",
          4560 => x"34",
          4561 => x"1c",
          4562 => x"5a",
          4563 => x"33",
          4564 => x"15",
          4565 => x"80",
          4566 => x"74",
          4567 => x"5a",
          4568 => x"10",
          4569 => x"ff",
          4570 => x"58",
          4571 => x"76",
          4572 => x"58",
          4573 => x"55",
          4574 => x"80",
          4575 => x"bf",
          4576 => x"87",
          4577 => x"ff",
          4578 => x"76",
          4579 => x"79",
          4580 => x"27",
          4581 => x"2e",
          4582 => x"27",
          4583 => x"56",
          4584 => x"ea",
          4585 => x"87",
          4586 => x"ec",
          4587 => x"41",
          4588 => x"f4",
          4589 => x"ba",
          4590 => x"80",
          4591 => x"56",
          4592 => x"84",
          4593 => x"08",
          4594 => x"38",
          4595 => x"34",
          4596 => x"05",
          4597 => x"06",
          4598 => x"38",
          4599 => x"e7",
          4600 => x"80",
          4601 => x"ba",
          4602 => x"81",
          4603 => x"19",
          4604 => x"57",
          4605 => x"38",
          4606 => x"09",
          4607 => x"75",
          4608 => x"51",
          4609 => x"80",
          4610 => x"75",
          4611 => x"38",
          4612 => x"74",
          4613 => x"30",
          4614 => x"74",
          4615 => x"59",
          4616 => x"52",
          4617 => x"8c",
          4618 => x"2e",
          4619 => x"2e",
          4620 => x"83",
          4621 => x"38",
          4622 => x"77",
          4623 => x"57",
          4624 => x"76",
          4625 => x"51",
          4626 => x"80",
          4627 => x"76",
          4628 => x"c3",
          4629 => x"55",
          4630 => x"ff",
          4631 => x"9c",
          4632 => x"70",
          4633 => x"05",
          4634 => x"38",
          4635 => x"06",
          4636 => x"0b",
          4637 => x"ba",
          4638 => x"75",
          4639 => x"40",
          4640 => x"81",
          4641 => x"ba",
          4642 => x"80",
          4643 => x"81",
          4644 => x"81",
          4645 => x"ba",
          4646 => x"83",
          4647 => x"19",
          4648 => x"31",
          4649 => x"38",
          4650 => x"84",
          4651 => x"fd",
          4652 => x"08",
          4653 => x"e9",
          4654 => x"ba",
          4655 => x"ba",
          4656 => x"81",
          4657 => x"70",
          4658 => x"70",
          4659 => x"5d",
          4660 => x"b8",
          4661 => x"80",
          4662 => x"38",
          4663 => x"09",
          4664 => x"76",
          4665 => x"51",
          4666 => x"80",
          4667 => x"76",
          4668 => x"83",
          4669 => x"61",
          4670 => x"8d",
          4671 => x"75",
          4672 => x"75",
          4673 => x"05",
          4674 => x"ff",
          4675 => x"70",
          4676 => x"e6",
          4677 => x"75",
          4678 => x"2a",
          4679 => x"83",
          4680 => x"78",
          4681 => x"2e",
          4682 => x"22",
          4683 => x"38",
          4684 => x"34",
          4685 => x"84",
          4686 => x"08",
          4687 => x"7f",
          4688 => x"54",
          4689 => x"53",
          4690 => x"3f",
          4691 => x"83",
          4692 => x"34",
          4693 => x"84",
          4694 => x"1d",
          4695 => x"33",
          4696 => x"fb",
          4697 => x"a0",
          4698 => x"1c",
          4699 => x"fb",
          4700 => x"33",
          4701 => x"09",
          4702 => x"39",
          4703 => x"fa",
          4704 => x"c0",
          4705 => x"b4",
          4706 => x"33",
          4707 => x"08",
          4708 => x"84",
          4709 => x"1c",
          4710 => x"a0",
          4711 => x"33",
          4712 => x"ba",
          4713 => x"ff",
          4714 => x"98",
          4715 => x"f7",
          4716 => x"80",
          4717 => x"81",
          4718 => x"05",
          4719 => x"ce",
          4720 => x"b4",
          4721 => x"7c",
          4722 => x"3f",
          4723 => x"61",
          4724 => x"96",
          4725 => x"82",
          4726 => x"80",
          4727 => x"05",
          4728 => x"58",
          4729 => x"74",
          4730 => x"56",
          4731 => x"14",
          4732 => x"76",
          4733 => x"79",
          4734 => x"55",
          4735 => x"80",
          4736 => x"5e",
          4737 => x"82",
          4738 => x"57",
          4739 => x"81",
          4740 => x"b2",
          4741 => x"75",
          4742 => x"80",
          4743 => x"90",
          4744 => x"77",
          4745 => x"58",
          4746 => x"81",
          4747 => x"38",
          4748 => x"81",
          4749 => x"a5",
          4750 => x"96",
          4751 => x"05",
          4752 => x"1c",
          4753 => x"89",
          4754 => x"08",
          4755 => x"9c",
          4756 => x"82",
          4757 => x"2b",
          4758 => x"88",
          4759 => x"59",
          4760 => x"88",
          4761 => x"56",
          4762 => x"15",
          4763 => x"07",
          4764 => x"3d",
          4765 => x"39",
          4766 => x"31",
          4767 => x"90",
          4768 => x"3f",
          4769 => x"06",
          4770 => x"81",
          4771 => x"2a",
          4772 => x"34",
          4773 => x"1f",
          4774 => x"70",
          4775 => x"38",
          4776 => x"70",
          4777 => x"07",
          4778 => x"74",
          4779 => x"0b",
          4780 => x"72",
          4781 => x"77",
          4782 => x"1e",
          4783 => x"ff",
          4784 => x"a4",
          4785 => x"54",
          4786 => x"84",
          4787 => x"80",
          4788 => x"ff",
          4789 => x"81",
          4790 => x"81",
          4791 => x"59",
          4792 => x"b4",
          4793 => x"80",
          4794 => x"73",
          4795 => x"39",
          4796 => x"42",
          4797 => x"55",
          4798 => x"53",
          4799 => x"72",
          4800 => x"08",
          4801 => x"94",
          4802 => x"82",
          4803 => x"58",
          4804 => x"52",
          4805 => x"72",
          4806 => x"38",
          4807 => x"76",
          4808 => x"17",
          4809 => x"af",
          4810 => x"80",
          4811 => x"82",
          4812 => x"89",
          4813 => x"83",
          4814 => x"70",
          4815 => x"80",
          4816 => x"8f",
          4817 => x"ff",
          4818 => x"72",
          4819 => x"38",
          4820 => x"76",
          4821 => x"17",
          4822 => x"56",
          4823 => x"38",
          4824 => x"32",
          4825 => x"51",
          4826 => x"38",
          4827 => x"33",
          4828 => x"72",
          4829 => x"25",
          4830 => x"38",
          4831 => x"3d",
          4832 => x"26",
          4833 => x"52",
          4834 => x"ba",
          4835 => x"73",
          4836 => x"ba",
          4837 => x"e5",
          4838 => x"53",
          4839 => x"39",
          4840 => x"52",
          4841 => x"8c",
          4842 => x"0d",
          4843 => x"30",
          4844 => x"5a",
          4845 => x"14",
          4846 => x"56",
          4847 => x"dc",
          4848 => x"07",
          4849 => x"61",
          4850 => x"76",
          4851 => x"2e",
          4852 => x"80",
          4853 => x"fe",
          4854 => x"30",
          4855 => x"56",
          4856 => x"89",
          4857 => x"76",
          4858 => x"76",
          4859 => x"22",
          4860 => x"5d",
          4861 => x"38",
          4862 => x"ae",
          4863 => x"aa",
          4864 => x"5a",
          4865 => x"10",
          4866 => x"76",
          4867 => x"22",
          4868 => x"06",
          4869 => x"53",
          4870 => x"ff",
          4871 => x"5c",
          4872 => x"19",
          4873 => x"80",
          4874 => x"38",
          4875 => x"25",
          4876 => x"ce",
          4877 => x"7c",
          4878 => x"77",
          4879 => x"25",
          4880 => x"72",
          4881 => x"2e",
          4882 => x"38",
          4883 => x"9e",
          4884 => x"82",
          4885 => x"5f",
          4886 => x"58",
          4887 => x"1c",
          4888 => x"84",
          4889 => x"7d",
          4890 => x"ed",
          4891 => x"2e",
          4892 => x"06",
          4893 => x"5d",
          4894 => x"07",
          4895 => x"7d",
          4896 => x"5a",
          4897 => x"ec",
          4898 => x"33",
          4899 => x"2e",
          4900 => x"84",
          4901 => x"74",
          4902 => x"2e",
          4903 => x"06",
          4904 => x"65",
          4905 => x"58",
          4906 => x"70",
          4907 => x"56",
          4908 => x"80",
          4909 => x"5a",
          4910 => x"75",
          4911 => x"38",
          4912 => x"81",
          4913 => x"5b",
          4914 => x"56",
          4915 => x"38",
          4916 => x"57",
          4917 => x"e9",
          4918 => x"1d",
          4919 => x"ba",
          4920 => x"84",
          4921 => x"82",
          4922 => x"38",
          4923 => x"06",
          4924 => x"38",
          4925 => x"05",
          4926 => x"33",
          4927 => x"57",
          4928 => x"38",
          4929 => x"55",
          4930 => x"74",
          4931 => x"59",
          4932 => x"79",
          4933 => x"81",
          4934 => x"70",
          4935 => x"09",
          4936 => x"07",
          4937 => x"1d",
          4938 => x"fc",
          4939 => x"ab",
          4940 => x"0c",
          4941 => x"26",
          4942 => x"c9",
          4943 => x"81",
          4944 => x"18",
          4945 => x"82",
          4946 => x"81",
          4947 => x"83",
          4948 => x"06",
          4949 => x"74",
          4950 => x"33",
          4951 => x"b9",
          4952 => x"83",
          4953 => x"70",
          4954 => x"80",
          4955 => x"8f",
          4956 => x"ff",
          4957 => x"72",
          4958 => x"38",
          4959 => x"8a",
          4960 => x"06",
          4961 => x"99",
          4962 => x"81",
          4963 => x"ff",
          4964 => x"a0",
          4965 => x"5b",
          4966 => x"53",
          4967 => x"70",
          4968 => x"2e",
          4969 => x"07",
          4970 => x"74",
          4971 => x"80",
          4972 => x"71",
          4973 => x"07",
          4974 => x"39",
          4975 => x"54",
          4976 => x"11",
          4977 => x"81",
          4978 => x"07",
          4979 => x"e5",
          4980 => x"fd",
          4981 => x"5c",
          4982 => x"ba",
          4983 => x"3d",
          4984 => x"e7",
          4985 => x"0c",
          4986 => x"79",
          4987 => x"81",
          4988 => x"56",
          4989 => x"ed",
          4990 => x"84",
          4991 => x"85",
          4992 => x"d4",
          4993 => x"76",
          4994 => x"0c",
          4995 => x"59",
          4996 => x"33",
          4997 => x"8c",
          4998 => x"5e",
          4999 => x"80",
          5000 => x"80",
          5001 => x"81",
          5002 => x"84",
          5003 => x"81",
          5004 => x"c2",
          5005 => x"82",
          5006 => x"84",
          5007 => x"34",
          5008 => x"5a",
          5009 => x"70",
          5010 => x"bb",
          5011 => x"2e",
          5012 => x"b4",
          5013 => x"84",
          5014 => x"71",
          5015 => x"74",
          5016 => x"75",
          5017 => x"1d",
          5018 => x"58",
          5019 => x"58",
          5020 => x"c4",
          5021 => x"88",
          5022 => x"2e",
          5023 => x"cf",
          5024 => x"88",
          5025 => x"80",
          5026 => x"33",
          5027 => x"81",
          5028 => x"75",
          5029 => x"5e",
          5030 => x"c8",
          5031 => x"17",
          5032 => x"5f",
          5033 => x"82",
          5034 => x"71",
          5035 => x"5a",
          5036 => x"80",
          5037 => x"06",
          5038 => x"17",
          5039 => x"2b",
          5040 => x"74",
          5041 => x"7c",
          5042 => x"80",
          5043 => x"56",
          5044 => x"83",
          5045 => x"2b",
          5046 => x"70",
          5047 => x"07",
          5048 => x"80",
          5049 => x"71",
          5050 => x"7b",
          5051 => x"7a",
          5052 => x"81",
          5053 => x"51",
          5054 => x"08",
          5055 => x"81",
          5056 => x"ff",
          5057 => x"5d",
          5058 => x"82",
          5059 => x"38",
          5060 => x"0c",
          5061 => x"a8",
          5062 => x"57",
          5063 => x"88",
          5064 => x"2e",
          5065 => x"0c",
          5066 => x"38",
          5067 => x"81",
          5068 => x"89",
          5069 => x"08",
          5070 => x"0c",
          5071 => x"0b",
          5072 => x"96",
          5073 => x"22",
          5074 => x"23",
          5075 => x"0b",
          5076 => x"0c",
          5077 => x"97",
          5078 => x"8c",
          5079 => x"d0",
          5080 => x"58",
          5081 => x"78",
          5082 => x"78",
          5083 => x"08",
          5084 => x"08",
          5085 => x"5c",
          5086 => x"ff",
          5087 => x"26",
          5088 => x"06",
          5089 => x"99",
          5090 => x"ff",
          5091 => x"2a",
          5092 => x"06",
          5093 => x"7a",
          5094 => x"2a",
          5095 => x"2e",
          5096 => x"5e",
          5097 => x"61",
          5098 => x"fe",
          5099 => x"5e",
          5100 => x"58",
          5101 => x"59",
          5102 => x"83",
          5103 => x"70",
          5104 => x"5b",
          5105 => x"e8",
          5106 => x"57",
          5107 => x"70",
          5108 => x"84",
          5109 => x"71",
          5110 => x"ff",
          5111 => x"83",
          5112 => x"5b",
          5113 => x"05",
          5114 => x"59",
          5115 => x"ba",
          5116 => x"2a",
          5117 => x"10",
          5118 => x"5d",
          5119 => x"83",
          5120 => x"80",
          5121 => x"18",
          5122 => x"2e",
          5123 => x"17",
          5124 => x"86",
          5125 => x"85",
          5126 => x"18",
          5127 => x"1f",
          5128 => x"5d",
          5129 => x"2e",
          5130 => x"b8",
          5131 => x"2e",
          5132 => x"70",
          5133 => x"42",
          5134 => x"2e",
          5135 => x"06",
          5136 => x"33",
          5137 => x"06",
          5138 => x"f8",
          5139 => x"38",
          5140 => x"7a",
          5141 => x"83",
          5142 => x"40",
          5143 => x"33",
          5144 => x"71",
          5145 => x"77",
          5146 => x"2e",
          5147 => x"83",
          5148 => x"81",
          5149 => x"40",
          5150 => x"58",
          5151 => x"38",
          5152 => x"fe",
          5153 => x"38",
          5154 => x"0d",
          5155 => x"dc",
          5156 => x"e5",
          5157 => x"8d",
          5158 => x"0d",
          5159 => x"e5",
          5160 => x"05",
          5161 => x"33",
          5162 => x"5f",
          5163 => x"74",
          5164 => x"8a",
          5165 => x"78",
          5166 => x"81",
          5167 => x"1b",
          5168 => x"84",
          5169 => x"93",
          5170 => x"83",
          5171 => x"e9",
          5172 => x"88",
          5173 => x"09",
          5174 => x"58",
          5175 => x"b1",
          5176 => x"2e",
          5177 => x"54",
          5178 => x"33",
          5179 => x"8c",
          5180 => x"81",
          5181 => x"99",
          5182 => x"17",
          5183 => x"2b",
          5184 => x"2e",
          5185 => x"17",
          5186 => x"90",
          5187 => x"33",
          5188 => x"71",
          5189 => x"59",
          5190 => x"09",
          5191 => x"17",
          5192 => x"90",
          5193 => x"33",
          5194 => x"71",
          5195 => x"5e",
          5196 => x"09",
          5197 => x"17",
          5198 => x"90",
          5199 => x"33",
          5200 => x"71",
          5201 => x"1c",
          5202 => x"90",
          5203 => x"33",
          5204 => x"71",
          5205 => x"49",
          5206 => x"5a",
          5207 => x"81",
          5208 => x"7c",
          5209 => x"8c",
          5210 => x"f7",
          5211 => x"38",
          5212 => x"39",
          5213 => x"17",
          5214 => x"ff",
          5215 => x"7a",
          5216 => x"84",
          5217 => x"17",
          5218 => x"a0",
          5219 => x"33",
          5220 => x"84",
          5221 => x"74",
          5222 => x"85",
          5223 => x"5c",
          5224 => x"17",
          5225 => x"2b",
          5226 => x"d2",
          5227 => x"ca",
          5228 => x"82",
          5229 => x"2b",
          5230 => x"88",
          5231 => x"0c",
          5232 => x"40",
          5233 => x"75",
          5234 => x"f9",
          5235 => x"38",
          5236 => x"f7",
          5237 => x"38",
          5238 => x"08",
          5239 => x"81",
          5240 => x"fc",
          5241 => x"d3",
          5242 => x"41",
          5243 => x"80",
          5244 => x"05",
          5245 => x"74",
          5246 => x"38",
          5247 => x"d1",
          5248 => x"c4",
          5249 => x"05",
          5250 => x"84",
          5251 => x"80",
          5252 => x"54",
          5253 => x"2e",
          5254 => x"53",
          5255 => x"ba",
          5256 => x"0c",
          5257 => x"ba",
          5258 => x"33",
          5259 => x"56",
          5260 => x"16",
          5261 => x"58",
          5262 => x"7f",
          5263 => x"7b",
          5264 => x"05",
          5265 => x"33",
          5266 => x"99",
          5267 => x"ff",
          5268 => x"76",
          5269 => x"81",
          5270 => x"9f",
          5271 => x"81",
          5272 => x"77",
          5273 => x"9f",
          5274 => x"80",
          5275 => x"5d",
          5276 => x"7f",
          5277 => x"f7",
          5278 => x"8b",
          5279 => x"05",
          5280 => x"56",
          5281 => x"06",
          5282 => x"9e",
          5283 => x"3f",
          5284 => x"8c",
          5285 => x"0c",
          5286 => x"9c",
          5287 => x"90",
          5288 => x"84",
          5289 => x"08",
          5290 => x"06",
          5291 => x"76",
          5292 => x"2e",
          5293 => x"76",
          5294 => x"06",
          5295 => x"66",
          5296 => x"88",
          5297 => x"5e",
          5298 => x"38",
          5299 => x"8f",
          5300 => x"80",
          5301 => x"a0",
          5302 => x"5e",
          5303 => x"9b",
          5304 => x"2e",
          5305 => x"9c",
          5306 => x"80",
          5307 => x"1c",
          5308 => x"34",
          5309 => x"b4",
          5310 => x"5f",
          5311 => x"17",
          5312 => x"57",
          5313 => x"80",
          5314 => x"5b",
          5315 => x"78",
          5316 => x"38",
          5317 => x"05",
          5318 => x"56",
          5319 => x"81",
          5320 => x"75",
          5321 => x"77",
          5322 => x"2e",
          5323 => x"7e",
          5324 => x"a4",
          5325 => x"12",
          5326 => x"40",
          5327 => x"81",
          5328 => x"16",
          5329 => x"90",
          5330 => x"33",
          5331 => x"71",
          5332 => x"60",
          5333 => x"5e",
          5334 => x"90",
          5335 => x"80",
          5336 => x"81",
          5337 => x"38",
          5338 => x"94",
          5339 => x"2b",
          5340 => x"78",
          5341 => x"27",
          5342 => x"5f",
          5343 => x"77",
          5344 => x"84",
          5345 => x"08",
          5346 => x"ba",
          5347 => x"75",
          5348 => x"c2",
          5349 => x"38",
          5350 => x"80",
          5351 => x"79",
          5352 => x"79",
          5353 => x"79",
          5354 => x"ca",
          5355 => x"07",
          5356 => x"8b",
          5357 => x"fe",
          5358 => x"33",
          5359 => x"7d",
          5360 => x"7c",
          5361 => x"74",
          5362 => x"84",
          5363 => x"08",
          5364 => x"8c",
          5365 => x"ba",
          5366 => x"80",
          5367 => x"82",
          5368 => x"38",
          5369 => x"08",
          5370 => x"af",
          5371 => x"17",
          5372 => x"34",
          5373 => x"38",
          5374 => x"34",
          5375 => x"39",
          5376 => x"98",
          5377 => x"5e",
          5378 => x"80",
          5379 => x"17",
          5380 => x"66",
          5381 => x"67",
          5382 => x"80",
          5383 => x"7c",
          5384 => x"38",
          5385 => x"5e",
          5386 => x"2e",
          5387 => x"7d",
          5388 => x"54",
          5389 => x"33",
          5390 => x"8c",
          5391 => x"81",
          5392 => x"7a",
          5393 => x"80",
          5394 => x"f9",
          5395 => x"53",
          5396 => x"52",
          5397 => x"8c",
          5398 => x"aa",
          5399 => x"34",
          5400 => x"84",
          5401 => x"17",
          5402 => x"33",
          5403 => x"ff",
          5404 => x"a0",
          5405 => x"16",
          5406 => x"5b",
          5407 => x"76",
          5408 => x"0c",
          5409 => x"06",
          5410 => x"7e",
          5411 => x"5f",
          5412 => x"38",
          5413 => x"1c",
          5414 => x"f9",
          5415 => x"1a",
          5416 => x"94",
          5417 => x"81",
          5418 => x"84",
          5419 => x"f7",
          5420 => x"9f",
          5421 => x"66",
          5422 => x"89",
          5423 => x"08",
          5424 => x"33",
          5425 => x"16",
          5426 => x"78",
          5427 => x"41",
          5428 => x"1a",
          5429 => x"1a",
          5430 => x"80",
          5431 => x"8c",
          5432 => x"75",
          5433 => x"81",
          5434 => x"06",
          5435 => x"22",
          5436 => x"7a",
          5437 => x"1a",
          5438 => x"38",
          5439 => x"98",
          5440 => x"fe",
          5441 => x"57",
          5442 => x"19",
          5443 => x"05",
          5444 => x"38",
          5445 => x"77",
          5446 => x"55",
          5447 => x"31",
          5448 => x"81",
          5449 => x"84",
          5450 => x"83",
          5451 => x"a9",
          5452 => x"75",
          5453 => x"71",
          5454 => x"75",
          5455 => x"81",
          5456 => x"ef",
          5457 => x"31",
          5458 => x"94",
          5459 => x"0c",
          5460 => x"56",
          5461 => x"0d",
          5462 => x"3d",
          5463 => x"9c",
          5464 => x"84",
          5465 => x"27",
          5466 => x"19",
          5467 => x"83",
          5468 => x"7f",
          5469 => x"81",
          5470 => x"19",
          5471 => x"ba",
          5472 => x"56",
          5473 => x"81",
          5474 => x"ff",
          5475 => x"05",
          5476 => x"38",
          5477 => x"70",
          5478 => x"75",
          5479 => x"81",
          5480 => x"59",
          5481 => x"fe",
          5482 => x"53",
          5483 => x"52",
          5484 => x"84",
          5485 => x"06",
          5486 => x"83",
          5487 => x"08",
          5488 => x"74",
          5489 => x"82",
          5490 => x"81",
          5491 => x"19",
          5492 => x"52",
          5493 => x"3f",
          5494 => x"1b",
          5495 => x"39",
          5496 => x"a3",
          5497 => x"fc",
          5498 => x"9c",
          5499 => x"06",
          5500 => x"08",
          5501 => x"91",
          5502 => x"0c",
          5503 => x"1b",
          5504 => x"92",
          5505 => x"65",
          5506 => x"7e",
          5507 => x"38",
          5508 => x"38",
          5509 => x"38",
          5510 => x"59",
          5511 => x"55",
          5512 => x"38",
          5513 => x"38",
          5514 => x"06",
          5515 => x"82",
          5516 => x"5d",
          5517 => x"09",
          5518 => x"76",
          5519 => x"38",
          5520 => x"89",
          5521 => x"76",
          5522 => x"74",
          5523 => x"2e",
          5524 => x"8c",
          5525 => x"08",
          5526 => x"56",
          5527 => x"81",
          5528 => x"9c",
          5529 => x"77",
          5530 => x"70",
          5531 => x"57",
          5532 => x"15",
          5533 => x"2e",
          5534 => x"7f",
          5535 => x"77",
          5536 => x"33",
          5537 => x"8c",
          5538 => x"08",
          5539 => x"a5",
          5540 => x"72",
          5541 => x"81",
          5542 => x"59",
          5543 => x"60",
          5544 => x"2b",
          5545 => x"7f",
          5546 => x"70",
          5547 => x"5a",
          5548 => x"83",
          5549 => x"7a",
          5550 => x"77",
          5551 => x"34",
          5552 => x"92",
          5553 => x"0c",
          5554 => x"55",
          5555 => x"a2",
          5556 => x"76",
          5557 => x"5a",
          5558 => x"59",
          5559 => x"b6",
          5560 => x"5e",
          5561 => x"06",
          5562 => x"b8",
          5563 => x"98",
          5564 => x"2e",
          5565 => x"b4",
          5566 => x"94",
          5567 => x"58",
          5568 => x"80",
          5569 => x"58",
          5570 => x"ff",
          5571 => x"81",
          5572 => x"81",
          5573 => x"70",
          5574 => x"98",
          5575 => x"08",
          5576 => x"38",
          5577 => x"b4",
          5578 => x"ba",
          5579 => x"08",
          5580 => x"55",
          5581 => x"e3",
          5582 => x"17",
          5583 => x"33",
          5584 => x"fe",
          5585 => x"1a",
          5586 => x"33",
          5587 => x"b4",
          5588 => x"7b",
          5589 => x"39",
          5590 => x"ab",
          5591 => x"84",
          5592 => x"1a",
          5593 => x"79",
          5594 => x"8c",
          5595 => x"bd",
          5596 => x"08",
          5597 => x"33",
          5598 => x"ba",
          5599 => x"8c",
          5600 => x"a8",
          5601 => x"08",
          5602 => x"5c",
          5603 => x"fc",
          5604 => x"17",
          5605 => x"33",
          5606 => x"fb",
          5607 => x"95",
          5608 => x"06",
          5609 => x"08",
          5610 => x"b4",
          5611 => x"81",
          5612 => x"3f",
          5613 => x"84",
          5614 => x"16",
          5615 => x"a0",
          5616 => x"16",
          5617 => x"06",
          5618 => x"08",
          5619 => x"81",
          5620 => x"60",
          5621 => x"58",
          5622 => x"1b",
          5623 => x"92",
          5624 => x"34",
          5625 => x"3d",
          5626 => x"89",
          5627 => x"08",
          5628 => x"33",
          5629 => x"16",
          5630 => x"77",
          5631 => x"5c",
          5632 => x"18",
          5633 => x"57",
          5634 => x"a0",
          5635 => x"79",
          5636 => x"7a",
          5637 => x"b8",
          5638 => x"93",
          5639 => x"2e",
          5640 => x"b4",
          5641 => x"18",
          5642 => x"57",
          5643 => x"19",
          5644 => x"5a",
          5645 => x"2a",
          5646 => x"76",
          5647 => x"83",
          5648 => x"55",
          5649 => x"7a",
          5650 => x"75",
          5651 => x"78",
          5652 => x"0b",
          5653 => x"34",
          5654 => x"0b",
          5655 => x"34",
          5656 => x"7b",
          5657 => x"8c",
          5658 => x"5b",
          5659 => x"ba",
          5660 => x"54",
          5661 => x"53",
          5662 => x"b5",
          5663 => x"fe",
          5664 => x"18",
          5665 => x"31",
          5666 => x"a0",
          5667 => x"17",
          5668 => x"06",
          5669 => x"08",
          5670 => x"81",
          5671 => x"79",
          5672 => x"55",
          5673 => x"56",
          5674 => x"55",
          5675 => x"7a",
          5676 => x"75",
          5677 => x"78",
          5678 => x"0b",
          5679 => x"34",
          5680 => x"0b",
          5681 => x"34",
          5682 => x"7b",
          5683 => x"8c",
          5684 => x"5b",
          5685 => x"39",
          5686 => x"3f",
          5687 => x"74",
          5688 => x"5a",
          5689 => x"70",
          5690 => x"8c",
          5691 => x"38",
          5692 => x"74",
          5693 => x"72",
          5694 => x"86",
          5695 => x"71",
          5696 => x"58",
          5697 => x"0c",
          5698 => x"0d",
          5699 => x"bc",
          5700 => x"53",
          5701 => x"56",
          5702 => x"70",
          5703 => x"38",
          5704 => x"9f",
          5705 => x"38",
          5706 => x"38",
          5707 => x"24",
          5708 => x"80",
          5709 => x"0d",
          5710 => x"8c",
          5711 => x"70",
          5712 => x"89",
          5713 => x"ff",
          5714 => x"2e",
          5715 => x"fc",
          5716 => x"76",
          5717 => x"81",
          5718 => x"54",
          5719 => x"12",
          5720 => x"9f",
          5721 => x"e0",
          5722 => x"71",
          5723 => x"73",
          5724 => x"ff",
          5725 => x"70",
          5726 => x"52",
          5727 => x"18",
          5728 => x"ff",
          5729 => x"77",
          5730 => x"51",
          5731 => x"53",
          5732 => x"51",
          5733 => x"55",
          5734 => x"38",
          5735 => x"0d",
          5736 => x"d0",
          5737 => x"8c",
          5738 => x"c6",
          5739 => x"98",
          5740 => x"e2",
          5741 => x"2a",
          5742 => x"b2",
          5743 => x"12",
          5744 => x"5e",
          5745 => x"a4",
          5746 => x"ba",
          5747 => x"ba",
          5748 => x"ff",
          5749 => x"0c",
          5750 => x"94",
          5751 => x"2b",
          5752 => x"54",
          5753 => x"58",
          5754 => x"0d",
          5755 => x"3d",
          5756 => x"80",
          5757 => x"fd",
          5758 => x"cf",
          5759 => x"84",
          5760 => x"80",
          5761 => x"08",
          5762 => x"3d",
          5763 => x"cc",
          5764 => x"5b",
          5765 => x"3f",
          5766 => x"8c",
          5767 => x"3d",
          5768 => x"2e",
          5769 => x"17",
          5770 => x"81",
          5771 => x"16",
          5772 => x"ba",
          5773 => x"57",
          5774 => x"82",
          5775 => x"11",
          5776 => x"07",
          5777 => x"56",
          5778 => x"80",
          5779 => x"ff",
          5780 => x"59",
          5781 => x"80",
          5782 => x"84",
          5783 => x"08",
          5784 => x"11",
          5785 => x"07",
          5786 => x"56",
          5787 => x"7a",
          5788 => x"52",
          5789 => x"ba",
          5790 => x"80",
          5791 => x"83",
          5792 => x"e4",
          5793 => x"ff",
          5794 => x"33",
          5795 => x"82",
          5796 => x"33",
          5797 => x"17",
          5798 => x"76",
          5799 => x"05",
          5800 => x"11",
          5801 => x"58",
          5802 => x"ff",
          5803 => x"58",
          5804 => x"5a",
          5805 => x"82",
          5806 => x"33",
          5807 => x"70",
          5808 => x"5a",
          5809 => x"70",
          5810 => x"f5",
          5811 => x"ab",
          5812 => x"38",
          5813 => x"81",
          5814 => x"77",
          5815 => x"05",
          5816 => x"06",
          5817 => x"34",
          5818 => x"3d",
          5819 => x"33",
          5820 => x"79",
          5821 => x"95",
          5822 => x"2b",
          5823 => x"dd",
          5824 => x"51",
          5825 => x"08",
          5826 => x"fd",
          5827 => x"b4",
          5828 => x"81",
          5829 => x"3f",
          5830 => x"be",
          5831 => x"34",
          5832 => x"84",
          5833 => x"17",
          5834 => x"33",
          5835 => x"fb",
          5836 => x"a0",
          5837 => x"16",
          5838 => x"59",
          5839 => x"3d",
          5840 => x"80",
          5841 => x"10",
          5842 => x"33",
          5843 => x"2e",
          5844 => x"f1",
          5845 => x"19",
          5846 => x"05",
          5847 => x"38",
          5848 => x"59",
          5849 => x"5e",
          5850 => x"f5",
          5851 => x"84",
          5852 => x"04",
          5853 => x"89",
          5854 => x"08",
          5855 => x"33",
          5856 => x"14",
          5857 => x"78",
          5858 => x"5a",
          5859 => x"15",
          5860 => x"15",
          5861 => x"38",
          5862 => x"78",
          5863 => x"22",
          5864 => x"78",
          5865 => x"17",
          5866 => x"8c",
          5867 => x"55",
          5868 => x"8c",
          5869 => x"30",
          5870 => x"71",
          5871 => x"73",
          5872 => x"27",
          5873 => x"16",
          5874 => x"33",
          5875 => x"57",
          5876 => x"52",
          5877 => x"ba",
          5878 => x"80",
          5879 => x"98",
          5880 => x"79",
          5881 => x"aa",
          5882 => x"39",
          5883 => x"72",
          5884 => x"04",
          5885 => x"06",
          5886 => x"94",
          5887 => x"78",
          5888 => x"77",
          5889 => x"75",
          5890 => x"0c",
          5891 => x"76",
          5892 => x"59",
          5893 => x"08",
          5894 => x"0c",
          5895 => x"3d",
          5896 => x"88",
          5897 => x"fe",
          5898 => x"2e",
          5899 => x"ba",
          5900 => x"94",
          5901 => x"75",
          5902 => x"9c",
          5903 => x"73",
          5904 => x"22",
          5905 => x"78",
          5906 => x"80",
          5907 => x"56",
          5908 => x"ff",
          5909 => x"54",
          5910 => x"ff",
          5911 => x"81",
          5912 => x"75",
          5913 => x"52",
          5914 => x"ba",
          5915 => x"81",
          5916 => x"ff",
          5917 => x"08",
          5918 => x"fe",
          5919 => x"82",
          5920 => x"0d",
          5921 => x"54",
          5922 => x"8c",
          5923 => x"05",
          5924 => x"08",
          5925 => x"8f",
          5926 => x"84",
          5927 => x"7a",
          5928 => x"b9",
          5929 => x"84",
          5930 => x"16",
          5931 => x"78",
          5932 => x"84",
          5933 => x"2e",
          5934 => x"11",
          5935 => x"07",
          5936 => x"57",
          5937 => x"17",
          5938 => x"17",
          5939 => x"b9",
          5940 => x"84",
          5941 => x"84",
          5942 => x"85",
          5943 => x"95",
          5944 => x"2b",
          5945 => x"19",
          5946 => x"3d",
          5947 => x"2e",
          5948 => x"2e",
          5949 => x"2e",
          5950 => x"22",
          5951 => x"80",
          5952 => x"75",
          5953 => x"3d",
          5954 => x"ff",
          5955 => x"06",
          5956 => x"53",
          5957 => x"7c",
          5958 => x"9f",
          5959 => x"97",
          5960 => x"8f",
          5961 => x"59",
          5962 => x"80",
          5963 => x"c7",
          5964 => x"75",
          5965 => x"84",
          5966 => x"08",
          5967 => x"08",
          5968 => x"b2",
          5969 => x"99",
          5970 => x"32",
          5971 => x"84",
          5972 => x"72",
          5973 => x"04",
          5974 => x"b1",
          5975 => x"99",
          5976 => x"32",
          5977 => x"84",
          5978 => x"cf",
          5979 => x"f9",
          5980 => x"8c",
          5981 => x"33",
          5982 => x"8c",
          5983 => x"38",
          5984 => x"39",
          5985 => x"89",
          5986 => x"c1",
          5987 => x"84",
          5988 => x"74",
          5989 => x"04",
          5990 => x"3f",
          5991 => x"8c",
          5992 => x"33",
          5993 => x"24",
          5994 => x"76",
          5995 => x"74",
          5996 => x"04",
          5997 => x"3d",
          5998 => x"56",
          5999 => x"52",
          6000 => x"ba",
          6001 => x"9a",
          6002 => x"11",
          6003 => x"57",
          6004 => x"75",
          6005 => x"95",
          6006 => x"77",
          6007 => x"93",
          6008 => x"8c",
          6009 => x"38",
          6010 => x"b4",
          6011 => x"83",
          6012 => x"8d",
          6013 => x"52",
          6014 => x"3f",
          6015 => x"38",
          6016 => x"0c",
          6017 => x"38",
          6018 => x"8d",
          6019 => x"33",
          6020 => x"88",
          6021 => x"07",
          6022 => x"ff",
          6023 => x"80",
          6024 => x"ff",
          6025 => x"53",
          6026 => x"78",
          6027 => x"94",
          6028 => x"58",
          6029 => x"8c",
          6030 => x"b4",
          6031 => x"81",
          6032 => x"3f",
          6033 => x"f8",
          6034 => x"34",
          6035 => x"84",
          6036 => x"18",
          6037 => x"33",
          6038 => x"fe",
          6039 => x"a0",
          6040 => x"17",
          6041 => x"5e",
          6042 => x"3d",
          6043 => x"81",
          6044 => x"2e",
          6045 => x"81",
          6046 => x"08",
          6047 => x"80",
          6048 => x"58",
          6049 => x"ca",
          6050 => x"0c",
          6051 => x"84",
          6052 => x"b8",
          6053 => x"88",
          6054 => x"1f",
          6055 => x"5f",
          6056 => x"fd",
          6057 => x"fd",
          6058 => x"7f",
          6059 => x"33",
          6060 => x"fe",
          6061 => x"39",
          6062 => x"76",
          6063 => x"74",
          6064 => x"73",
          6065 => x"84",
          6066 => x"81",
          6067 => x"80",
          6068 => x"80",
          6069 => x"2a",
          6070 => x"80",
          6071 => x"54",
          6072 => x"73",
          6073 => x"08",
          6074 => x"9c",
          6075 => x"56",
          6076 => x"08",
          6077 => x"59",
          6078 => x"85",
          6079 => x"74",
          6080 => x"04",
          6081 => x"38",
          6082 => x"3f",
          6083 => x"8c",
          6084 => x"ba",
          6085 => x"84",
          6086 => x"38",
          6087 => x"85",
          6088 => x"c8",
          6089 => x"18",
          6090 => x"ff",
          6091 => x"84",
          6092 => x"17",
          6093 => x"a0",
          6094 => x"fe",
          6095 => x"81",
          6096 => x"77",
          6097 => x"0b",
          6098 => x"80",
          6099 => x"98",
          6100 => x"b9",
          6101 => x"81",
          6102 => x"2e",
          6103 => x"79",
          6104 => x"08",
          6105 => x"08",
          6106 => x"54",
          6107 => x"81",
          6108 => x"17",
          6109 => x"2e",
          6110 => x"51",
          6111 => x"08",
          6112 => x"38",
          6113 => x"3f",
          6114 => x"8c",
          6115 => x"ba",
          6116 => x"84",
          6117 => x"38",
          6118 => x"83",
          6119 => x"e6",
          6120 => x"18",
          6121 => x"90",
          6122 => x"16",
          6123 => x"34",
          6124 => x"38",
          6125 => x"58",
          6126 => x"39",
          6127 => x"fc",
          6128 => x"0b",
          6129 => x"39",
          6130 => x"59",
          6131 => x"18",
          6132 => x"ba",
          6133 => x"ff",
          6134 => x"a7",
          6135 => x"51",
          6136 => x"08",
          6137 => x"8a",
          6138 => x"3d",
          6139 => x"52",
          6140 => x"f8",
          6141 => x"ba",
          6142 => x"05",
          6143 => x"57",
          6144 => x"2b",
          6145 => x"80",
          6146 => x"57",
          6147 => x"a3",
          6148 => x"33",
          6149 => x"5e",
          6150 => x"d5",
          6151 => x"76",
          6152 => x"98",
          6153 => x"77",
          6154 => x"52",
          6155 => x"f9",
          6156 => x"ba",
          6157 => x"8c",
          6158 => x"3f",
          6159 => x"8c",
          6160 => x"8c",
          6161 => x"33",
          6162 => x"90",
          6163 => x"ff",
          6164 => x"2e",
          6165 => x"a1",
          6166 => x"57",
          6167 => x"38",
          6168 => x"3f",
          6169 => x"8c",
          6170 => x"70",
          6171 => x"80",
          6172 => x"38",
          6173 => x"27",
          6174 => x"81",
          6175 => x"38",
          6176 => x"ba",
          6177 => x"3d",
          6178 => x"08",
          6179 => x"2e",
          6180 => x"59",
          6181 => x"80",
          6182 => x"17",
          6183 => x"ee",
          6184 => x"85",
          6185 => x"18",
          6186 => x"19",
          6187 => x"83",
          6188 => x"fe",
          6189 => x"8b",
          6190 => x"84",
          6191 => x"38",
          6192 => x"cd",
          6193 => x"54",
          6194 => x"17",
          6195 => x"58",
          6196 => x"81",
          6197 => x"08",
          6198 => x"18",
          6199 => x"55",
          6200 => x"38",
          6201 => x"09",
          6202 => x"b4",
          6203 => x"7c",
          6204 => x"c5",
          6205 => x"55",
          6206 => x"52",
          6207 => x"ba",
          6208 => x"80",
          6209 => x"08",
          6210 => x"8c",
          6211 => x"53",
          6212 => x"3f",
          6213 => x"17",
          6214 => x"5c",
          6215 => x"81",
          6216 => x"81",
          6217 => x"55",
          6218 => x"56",
          6219 => x"39",
          6220 => x"39",
          6221 => x"0d",
          6222 => x"52",
          6223 => x"84",
          6224 => x"08",
          6225 => x"8c",
          6226 => x"6f",
          6227 => x"a6",
          6228 => x"84",
          6229 => x"84",
          6230 => x"84",
          6231 => x"06",
          6232 => x"70",
          6233 => x"56",
          6234 => x"52",
          6235 => x"c0",
          6236 => x"5c",
          6237 => x"56",
          6238 => x"f9",
          6239 => x"81",
          6240 => x"84",
          6241 => x"5a",
          6242 => x"9c",
          6243 => x"5b",
          6244 => x"22",
          6245 => x"5c",
          6246 => x"59",
          6247 => x"70",
          6248 => x"74",
          6249 => x"55",
          6250 => x"54",
          6251 => x"33",
          6252 => x"8c",
          6253 => x"dc",
          6254 => x"54",
          6255 => x"53",
          6256 => x"a5",
          6257 => x"be",
          6258 => x"34",
          6259 => x"55",
          6260 => x"38",
          6261 => x"09",
          6262 => x"b4",
          6263 => x"77",
          6264 => x"e5",
          6265 => x"7d",
          6266 => x"b4",
          6267 => x"ac",
          6268 => x"f9",
          6269 => x"ba",
          6270 => x"84",
          6271 => x"38",
          6272 => x"84",
          6273 => x"fe",
          6274 => x"fc",
          6275 => x"94",
          6276 => x"27",
          6277 => x"84",
          6278 => x"18",
          6279 => x"a1",
          6280 => x"3d",
          6281 => x"83",
          6282 => x"78",
          6283 => x"8b",
          6284 => x"70",
          6285 => x"75",
          6286 => x"18",
          6287 => x"19",
          6288 => x"34",
          6289 => x"80",
          6290 => x"d1",
          6291 => x"06",
          6292 => x"77",
          6293 => x"34",
          6294 => x"cc",
          6295 => x"1a",
          6296 => x"81",
          6297 => x"59",
          6298 => x"7d",
          6299 => x"64",
          6300 => x"57",
          6301 => x"88",
          6302 => x"75",
          6303 => x"38",
          6304 => x"79",
          6305 => x"8c",
          6306 => x"b6",
          6307 => x"96",
          6308 => x"17",
          6309 => x"cc",
          6310 => x"5d",
          6311 => x"59",
          6312 => x"79",
          6313 => x"90",
          6314 => x"0b",
          6315 => x"80",
          6316 => x"84",
          6317 => x"76",
          6318 => x"34",
          6319 => x"17",
          6320 => x"5b",
          6321 => x"2a",
          6322 => x"59",
          6323 => x"57",
          6324 => x"2a",
          6325 => x"2a",
          6326 => x"90",
          6327 => x"0b",
          6328 => x"98",
          6329 => x"96",
          6330 => x"3d",
          6331 => x"2e",
          6332 => x"33",
          6333 => x"2e",
          6334 => x"ba",
          6335 => x"3d",
          6336 => x"ff",
          6337 => x"56",
          6338 => x"38",
          6339 => x"0d",
          6340 => x"08",
          6341 => x"9f",
          6342 => x"84",
          6343 => x"bb",
          6344 => x"56",
          6345 => x"ae",
          6346 => x"81",
          6347 => x"59",
          6348 => x"99",
          6349 => x"55",
          6350 => x"70",
          6351 => x"74",
          6352 => x"51",
          6353 => x"08",
          6354 => x"38",
          6355 => x"38",
          6356 => x"3d",
          6357 => x"81",
          6358 => x"26",
          6359 => x"06",
          6360 => x"80",
          6361 => x"fc",
          6362 => x"5c",
          6363 => x"70",
          6364 => x"5a",
          6365 => x"e0",
          6366 => x"ff",
          6367 => x"38",
          6368 => x"55",
          6369 => x"75",
          6370 => x"77",
          6371 => x"30",
          6372 => x"5d",
          6373 => x"81",
          6374 => x"24",
          6375 => x"5b",
          6376 => x"b4",
          6377 => x"3d",
          6378 => x"ff",
          6379 => x"56",
          6380 => x"fd",
          6381 => x"09",
          6382 => x"ff",
          6383 => x"56",
          6384 => x"6f",
          6385 => x"05",
          6386 => x"70",
          6387 => x"05",
          6388 => x"38",
          6389 => x"34",
          6390 => x"06",
          6391 => x"07",
          6392 => x"81",
          6393 => x"70",
          6394 => x"80",
          6395 => x"6b",
          6396 => x"33",
          6397 => x"72",
          6398 => x"2e",
          6399 => x"08",
          6400 => x"82",
          6401 => x"29",
          6402 => x"80",
          6403 => x"58",
          6404 => x"83",
          6405 => x"81",
          6406 => x"17",
          6407 => x"ba",
          6408 => x"58",
          6409 => x"57",
          6410 => x"fb",
          6411 => x"ae",
          6412 => x"70",
          6413 => x"80",
          6414 => x"77",
          6415 => x"7a",
          6416 => x"75",
          6417 => x"34",
          6418 => x"18",
          6419 => x"34",
          6420 => x"08",
          6421 => x"38",
          6422 => x"3f",
          6423 => x"8c",
          6424 => x"98",
          6425 => x"08",
          6426 => x"7a",
          6427 => x"06",
          6428 => x"b8",
          6429 => x"e2",
          6430 => x"2e",
          6431 => x"b4",
          6432 => x"9c",
          6433 => x"0b",
          6434 => x"27",
          6435 => x"fc",
          6436 => x"84",
          6437 => x"38",
          6438 => x"38",
          6439 => x"51",
          6440 => x"08",
          6441 => x"04",
          6442 => x"3d",
          6443 => x"33",
          6444 => x"78",
          6445 => x"84",
          6446 => x"38",
          6447 => x"a0",
          6448 => x"3d",
          6449 => x"53",
          6450 => x"e2",
          6451 => x"08",
          6452 => x"38",
          6453 => x"b4",
          6454 => x"ba",
          6455 => x"08",
          6456 => x"5d",
          6457 => x"93",
          6458 => x"17",
          6459 => x"33",
          6460 => x"fd",
          6461 => x"53",
          6462 => x"52",
          6463 => x"84",
          6464 => x"ba",
          6465 => x"08",
          6466 => x"08",
          6467 => x"fc",
          6468 => x"82",
          6469 => x"81",
          6470 => x"05",
          6471 => x"fe",
          6472 => x"39",
          6473 => x"33",
          6474 => x"56",
          6475 => x"52",
          6476 => x"84",
          6477 => x"08",
          6478 => x"8c",
          6479 => x"66",
          6480 => x"96",
          6481 => x"84",
          6482 => x"cf",
          6483 => x"56",
          6484 => x"71",
          6485 => x"74",
          6486 => x"8b",
          6487 => x"16",
          6488 => x"84",
          6489 => x"96",
          6490 => x"57",
          6491 => x"97",
          6492 => x"ba",
          6493 => x"80",
          6494 => x"0c",
          6495 => x"52",
          6496 => x"d8",
          6497 => x"ba",
          6498 => x"05",
          6499 => x"75",
          6500 => x"19",
          6501 => x"56",
          6502 => x"55",
          6503 => x"58",
          6504 => x"54",
          6505 => x"0b",
          6506 => x"88",
          6507 => x"8c",
          6508 => x"0d",
          6509 => x"3d",
          6510 => x"a0",
          6511 => x"ba",
          6512 => x"08",
          6513 => x"80",
          6514 => x"5a",
          6515 => x"70",
          6516 => x"80",
          6517 => x"06",
          6518 => x"38",
          6519 => x"5a",
          6520 => x"38",
          6521 => x"7a",
          6522 => x"81",
          6523 => x"16",
          6524 => x"ba",
          6525 => x"57",
          6526 => x"57",
          6527 => x"58",
          6528 => x"38",
          6529 => x"38",
          6530 => x"11",
          6531 => x"71",
          6532 => x"72",
          6533 => x"62",
          6534 => x"76",
          6535 => x"04",
          6536 => x"3d",
          6537 => x"84",
          6538 => x"08",
          6539 => x"2e",
          6540 => x"7b",
          6541 => x"54",
          6542 => x"53",
          6543 => x"ad",
          6544 => x"7a",
          6545 => x"84",
          6546 => x"16",
          6547 => x"8c",
          6548 => x"27",
          6549 => x"74",
          6550 => x"38",
          6551 => x"08",
          6552 => x"51",
          6553 => x"54",
          6554 => x"33",
          6555 => x"8c",
          6556 => x"86",
          6557 => x"bb",
          6558 => x"ba",
          6559 => x"8c",
          6560 => x"59",
          6561 => x"57",
          6562 => x"19",
          6563 => x"70",
          6564 => x"80",
          6565 => x"11",
          6566 => x"2e",
          6567 => x"fd",
          6568 => x"a1",
          6569 => x"51",
          6570 => x"08",
          6571 => x"38",
          6572 => x"a0",
          6573 => x"15",
          6574 => x"08",
          6575 => x"58",
          6576 => x"38",
          6577 => x"81",
          6578 => x"81",
          6579 => x"ff",
          6580 => x"a1",
          6581 => x"8c",
          6582 => x"8c",
          6583 => x"80",
          6584 => x"0b",
          6585 => x"06",
          6586 => x"d6",
          6587 => x"38",
          6588 => x"06",
          6589 => x"38",
          6590 => x"38",
          6591 => x"a3",
          6592 => x"38",
          6593 => x"ff",
          6594 => x"55",
          6595 => x"81",
          6596 => x"5d",
          6597 => x"33",
          6598 => x"5a",
          6599 => x"3d",
          6600 => x"2e",
          6601 => x"02",
          6602 => x"5c",
          6603 => x"87",
          6604 => x"7d",
          6605 => x"70",
          6606 => x"ba",
          6607 => x"80",
          6608 => x"ba",
          6609 => x"b5",
          6610 => x"ba",
          6611 => x"74",
          6612 => x"ba",
          6613 => x"e7",
          6614 => x"52",
          6615 => x"ba",
          6616 => x"80",
          6617 => x"38",
          6618 => x"70",
          6619 => x"05",
          6620 => x"38",
          6621 => x"7d",
          6622 => x"8c",
          6623 => x"8a",
          6624 => x"ff",
          6625 => x"2e",
          6626 => x"55",
          6627 => x"08",
          6628 => x"b1",
          6629 => x"ba",
          6630 => x"81",
          6631 => x"19",
          6632 => x"59",
          6633 => x"83",
          6634 => x"81",
          6635 => x"53",
          6636 => x"fe",
          6637 => x"80",
          6638 => x"76",
          6639 => x"38",
          6640 => x"5a",
          6641 => x"38",
          6642 => x"56",
          6643 => x"81",
          6644 => x"81",
          6645 => x"84",
          6646 => x"08",
          6647 => x"76",
          6648 => x"76",
          6649 => x"80",
          6650 => x"15",
          6651 => x"0b",
          6652 => x"57",
          6653 => x"76",
          6654 => x"55",
          6655 => x"70",
          6656 => x"05",
          6657 => x"38",
          6658 => x"34",
          6659 => x"7d",
          6660 => x"8c",
          6661 => x"fe",
          6662 => x"53",
          6663 => x"d4",
          6664 => x"2e",
          6665 => x"ba",
          6666 => x"08",
          6667 => x"19",
          6668 => x"55",
          6669 => x"8c",
          6670 => x"81",
          6671 => x"84",
          6672 => x"08",
          6673 => x"39",
          6674 => x"fd",
          6675 => x"b4",
          6676 => x"7a",
          6677 => x"fd",
          6678 => x"60",
          6679 => x"33",
          6680 => x"2e",
          6681 => x"2e",
          6682 => x"2e",
          6683 => x"22",
          6684 => x"38",
          6685 => x"38",
          6686 => x"38",
          6687 => x"17",
          6688 => x"70",
          6689 => x"80",
          6690 => x"22",
          6691 => x"57",
          6692 => x"15",
          6693 => x"9f",
          6694 => x"1c",
          6695 => x"81",
          6696 => x"78",
          6697 => x"56",
          6698 => x"fe",
          6699 => x"55",
          6700 => x"82",
          6701 => x"81",
          6702 => x"2e",
          6703 => x"81",
          6704 => x"2e",
          6705 => x"06",
          6706 => x"84",
          6707 => x"87",
          6708 => x"0d",
          6709 => x"ac",
          6710 => x"54",
          6711 => x"55",
          6712 => x"81",
          6713 => x"80",
          6714 => x"81",
          6715 => x"52",
          6716 => x"ba",
          6717 => x"ff",
          6718 => x"57",
          6719 => x"90",
          6720 => x"8c",
          6721 => x"18",
          6722 => x"5c",
          6723 => x"fe",
          6724 => x"7a",
          6725 => x"94",
          6726 => x"5d",
          6727 => x"d6",
          6728 => x"5b",
          6729 => x"fe",
          6730 => x"ff",
          6731 => x"98",
          6732 => x"a5",
          6733 => x"05",
          6734 => x"3d",
          6735 => x"2e",
          6736 => x"5b",
          6737 => x"ba",
          6738 => x"75",
          6739 => x"e8",
          6740 => x"38",
          6741 => x"70",
          6742 => x"38",
          6743 => x"80",
          6744 => x"40",
          6745 => x"ce",
          6746 => x"ff",
          6747 => x"57",
          6748 => x"81",
          6749 => x"38",
          6750 => x"79",
          6751 => x"8c",
          6752 => x"80",
          6753 => x"80",
          6754 => x"06",
          6755 => x"2e",
          6756 => x"f8",
          6757 => x"f0",
          6758 => x"83",
          6759 => x"08",
          6760 => x"4c",
          6761 => x"38",
          6762 => x"56",
          6763 => x"7d",
          6764 => x"74",
          6765 => x"be",
          6766 => x"83",
          6767 => x"61",
          6768 => x"07",
          6769 => x"d5",
          6770 => x"7d",
          6771 => x"33",
          6772 => x"38",
          6773 => x"12",
          6774 => x"07",
          6775 => x"2b",
          6776 => x"83",
          6777 => x"2b",
          6778 => x"70",
          6779 => x"07",
          6780 => x"0c",
          6781 => x"59",
          6782 => x"57",
          6783 => x"93",
          6784 => x"38",
          6785 => x"49",
          6786 => x"87",
          6787 => x"61",
          6788 => x"83",
          6789 => x"58",
          6790 => x"ae",
          6791 => x"83",
          6792 => x"2e",
          6793 => x"83",
          6794 => x"70",
          6795 => x"86",
          6796 => x"52",
          6797 => x"ba",
          6798 => x"ba",
          6799 => x"81",
          6800 => x"ba",
          6801 => x"83",
          6802 => x"89",
          6803 => x"1f",
          6804 => x"05",
          6805 => x"57",
          6806 => x"74",
          6807 => x"60",
          6808 => x"f2",
          6809 => x"53",
          6810 => x"cf",
          6811 => x"83",
          6812 => x"09",
          6813 => x"f5",
          6814 => x"ac",
          6815 => x"55",
          6816 => x"74",
          6817 => x"84",
          6818 => x"ba",
          6819 => x"39",
          6820 => x"3d",
          6821 => x"33",
          6822 => x"57",
          6823 => x"1d",
          6824 => x"58",
          6825 => x"0b",
          6826 => x"7d",
          6827 => x"33",
          6828 => x"9f",
          6829 => x"89",
          6830 => x"58",
          6831 => x"26",
          6832 => x"06",
          6833 => x"5a",
          6834 => x"85",
          6835 => x"32",
          6836 => x"7b",
          6837 => x"80",
          6838 => x"5c",
          6839 => x"56",
          6840 => x"53",
          6841 => x"3f",
          6842 => x"b6",
          6843 => x"ba",
          6844 => x"bf",
          6845 => x"26",
          6846 => x"fb",
          6847 => x"7b",
          6848 => x"a3",
          6849 => x"81",
          6850 => x"fd",
          6851 => x"46",
          6852 => x"08",
          6853 => x"38",
          6854 => x"fb",
          6855 => x"8c",
          6856 => x"0c",
          6857 => x"99",
          6858 => x"74",
          6859 => x"ae",
          6860 => x"76",
          6861 => x"55",
          6862 => x"c8",
          6863 => x"58",
          6864 => x"ff",
          6865 => x"05",
          6866 => x"05",
          6867 => x"83",
          6868 => x"05",
          6869 => x"8f",
          6870 => x"62",
          6871 => x"61",
          6872 => x"06",
          6873 => x"56",
          6874 => x"38",
          6875 => x"61",
          6876 => x"6b",
          6877 => x"05",
          6878 => x"61",
          6879 => x"34",
          6880 => x"9c",
          6881 => x"61",
          6882 => x"6b",
          6883 => x"84",
          6884 => x"61",
          6885 => x"f7",
          6886 => x"61",
          6887 => x"34",
          6888 => x"83",
          6889 => x"05",
          6890 => x"97",
          6891 => x"34",
          6892 => x"ab",
          6893 => x"76",
          6894 => x"81",
          6895 => x"ef",
          6896 => x"d5",
          6897 => x"ff",
          6898 => x"60",
          6899 => x"81",
          6900 => x"38",
          6901 => x"9c",
          6902 => x"70",
          6903 => x"74",
          6904 => x"83",
          6905 => x"f8",
          6906 => x"57",
          6907 => x"45",
          6908 => x"34",
          6909 => x"81",
          6910 => x"75",
          6911 => x"66",
          6912 => x"7a",
          6913 => x"9d",
          6914 => x"38",
          6915 => x"70",
          6916 => x"74",
          6917 => x"58",
          6918 => x"40",
          6919 => x"56",
          6920 => x"65",
          6921 => x"55",
          6922 => x"51",
          6923 => x"08",
          6924 => x"31",
          6925 => x"62",
          6926 => x"83",
          6927 => x"62",
          6928 => x"84",
          6929 => x"5e",
          6930 => x"56",
          6931 => x"34",
          6932 => x"d5",
          6933 => x"83",
          6934 => x"67",
          6935 => x"34",
          6936 => x"84",
          6937 => x"52",
          6938 => x"fe",
          6939 => x"08",
          6940 => x"86",
          6941 => x"87",
          6942 => x"34",
          6943 => x"61",
          6944 => x"08",
          6945 => x"83",
          6946 => x"64",
          6947 => x"2a",
          6948 => x"62",
          6949 => x"05",
          6950 => x"79",
          6951 => x"84",
          6952 => x"53",
          6953 => x"3f",
          6954 => x"b6",
          6955 => x"8c",
          6956 => x"0c",
          6957 => x"1c",
          6958 => x"7a",
          6959 => x"0b",
          6960 => x"80",
          6961 => x"38",
          6962 => x"17",
          6963 => x"2e",
          6964 => x"77",
          6965 => x"84",
          6966 => x"05",
          6967 => x"80",
          6968 => x"8a",
          6969 => x"77",
          6970 => x"e4",
          6971 => x"f5",
          6972 => x"38",
          6973 => x"38",
          6974 => x"06",
          6975 => x"83",
          6976 => x"05",
          6977 => x"a1",
          6978 => x"61",
          6979 => x"76",
          6980 => x"80",
          6981 => x"80",
          6982 => x"05",
          6983 => x"34",
          6984 => x"2a",
          6985 => x"90",
          6986 => x"7c",
          6987 => x"34",
          6988 => x"ad",
          6989 => x"80",
          6990 => x"05",
          6991 => x"61",
          6992 => x"34",
          6993 => x"a9",
          6994 => x"80",
          6995 => x"55",
          6996 => x"70",
          6997 => x"74",
          6998 => x"81",
          6999 => x"58",
          7000 => x"f9",
          7001 => x"52",
          7002 => x"57",
          7003 => x"7d",
          7004 => x"83",
          7005 => x"8c",
          7006 => x"bf",
          7007 => x"84",
          7008 => x"ba",
          7009 => x"4a",
          7010 => x"ff",
          7011 => x"6a",
          7012 => x"61",
          7013 => x"34",
          7014 => x"88",
          7015 => x"ff",
          7016 => x"7c",
          7017 => x"1f",
          7018 => x"d5",
          7019 => x"75",
          7020 => x"57",
          7021 => x"7c",
          7022 => x"80",
          7023 => x"80",
          7024 => x"80",
          7025 => x"e4",
          7026 => x"05",
          7027 => x"34",
          7028 => x"7f",
          7029 => x"05",
          7030 => x"83",
          7031 => x"75",
          7032 => x"2a",
          7033 => x"82",
          7034 => x"83",
          7035 => x"05",
          7036 => x"80",
          7037 => x"81",
          7038 => x"51",
          7039 => x"1f",
          7040 => x"a5",
          7041 => x"39",
          7042 => x"80",
          7043 => x"76",
          7044 => x"8e",
          7045 => x"52",
          7046 => x"81",
          7047 => x"3d",
          7048 => x"74",
          7049 => x"17",
          7050 => x"77",
          7051 => x"55",
          7052 => x"ba",
          7053 => x"3d",
          7054 => x"33",
          7055 => x"38",
          7056 => x"9e",
          7057 => x"05",
          7058 => x"55",
          7059 => x"18",
          7060 => x"3d",
          7061 => x"74",
          7062 => x"ff",
          7063 => x"30",
          7064 => x"84",
          7065 => x"5a",
          7066 => x"51",
          7067 => x"3d",
          7068 => x"3d",
          7069 => x"80",
          7070 => x"15",
          7071 => x"77",
          7072 => x"7c",
          7073 => x"7d",
          7074 => x"75",
          7075 => x"b8",
          7076 => x"88",
          7077 => x"9e",
          7078 => x"75",
          7079 => x"ff",
          7080 => x"86",
          7081 => x"0b",
          7082 => x"04",
          7083 => x"54",
          7084 => x"9d",
          7085 => x"70",
          7086 => x"5a",
          7087 => x"76",
          7088 => x"7d",
          7089 => x"04",
          7090 => x"9a",
          7091 => x"80",
          7092 => x"ff",
          7093 => x"85",
          7094 => x"27",
          7095 => x"06",
          7096 => x"83",
          7097 => x"9c",
          7098 => x"06",
          7099 => x"38",
          7100 => x"22",
          7101 => x"70",
          7102 => x"53",
          7103 => x"02",
          7104 => x"05",
          7105 => x"ff",
          7106 => x"ba",
          7107 => x"83",
          7108 => x"70",
          7109 => x"83",
          7110 => x"8c",
          7111 => x"3d",
          7112 => x"26",
          7113 => x"06",
          7114 => x"ff",
          7115 => x"05",
          7116 => x"25",
          7117 => x"53",
          7118 => x"53",
          7119 => x"81",
          7120 => x"76",
          7121 => x"10",
          7122 => x"54",
          7123 => x"26",
          7124 => x"cb",
          7125 => x"0c",
          7126 => x"55",
          7127 => x"38",
          7128 => x"54",
          7129 => x"83",
          7130 => x"d3",
          7131 => x"ff",
          7132 => x"70",
          7133 => x"39",
          7134 => x"57",
          7135 => x"ff",
          7136 => x"16",
          7137 => x"c5",
          7138 => x"06",
          7139 => x"31",
          7140 => x"ff",
          7141 => x"39",
          7142 => x"22",
          7143 => x"ff",
          7144 => x"ff",
          7145 => x"00",
          7146 => x"00",
          7147 => x"00",
          7148 => x"00",
          7149 => x"00",
          7150 => x"00",
          7151 => x"00",
          7152 => x"00",
          7153 => x"00",
          7154 => x"00",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"00",
          7372 => x"00",
          7373 => x"00",
          7374 => x"00",
          7375 => x"00",
          7376 => x"00",
          7377 => x"00",
          7378 => x"00",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"00",
          7383 => x"6c",
          7384 => x"00",
          7385 => x"00",
          7386 => x"00",
          7387 => x"72",
          7388 => x"00",
          7389 => x"00",
          7390 => x"00",
          7391 => x"65",
          7392 => x"69",
          7393 => x"66",
          7394 => x"61",
          7395 => x"6d",
          7396 => x"72",
          7397 => x"00",
          7398 => x"00",
          7399 => x"00",
          7400 => x"38",
          7401 => x"63",
          7402 => x"63",
          7403 => x"00",
          7404 => x"6e",
          7405 => x"72",
          7406 => x"61",
          7407 => x"73",
          7408 => x"65",
          7409 => x"6f",
          7410 => x"6f",
          7411 => x"65",
          7412 => x"6e",
          7413 => x"65",
          7414 => x"72",
          7415 => x"69",
          7416 => x"6f",
          7417 => x"69",
          7418 => x"6f",
          7419 => x"6e",
          7420 => x"6c",
          7421 => x"6f",
          7422 => x"6f",
          7423 => x"6f",
          7424 => x"69",
          7425 => x"65",
          7426 => x"66",
          7427 => x"20",
          7428 => x"69",
          7429 => x"65",
          7430 => x"00",
          7431 => x"20",
          7432 => x"69",
          7433 => x"69",
          7434 => x"44",
          7435 => x"74",
          7436 => x"63",
          7437 => x"69",
          7438 => x"6c",
          7439 => x"69",
          7440 => x"69",
          7441 => x"61",
          7442 => x"74",
          7443 => x"63",
          7444 => x"6e",
          7445 => x"6e",
          7446 => x"69",
          7447 => x"00",
          7448 => x"74",
          7449 => x"2e",
          7450 => x"6c",
          7451 => x"2e",
          7452 => x"6e",
          7453 => x"79",
          7454 => x"6e",
          7455 => x"72",
          7456 => x"45",
          7457 => x"75",
          7458 => x"00",
          7459 => x"62",
          7460 => x"20",
          7461 => x"62",
          7462 => x"63",
          7463 => x"65",
          7464 => x"30",
          7465 => x"20",
          7466 => x"00",
          7467 => x"00",
          7468 => x"30",
          7469 => x"20",
          7470 => x"00",
          7471 => x"2a",
          7472 => x"31",
          7473 => x"30",
          7474 => x"00",
          7475 => x"20",
          7476 => x"78",
          7477 => x"20",
          7478 => x"50",
          7479 => x"72",
          7480 => x"64",
          7481 => x"41",
          7482 => x"69",
          7483 => x"74",
          7484 => x"20",
          7485 => x"72",
          7486 => x"41",
          7487 => x"69",
          7488 => x"74",
          7489 => x"20",
          7490 => x"72",
          7491 => x"4f",
          7492 => x"69",
          7493 => x"74",
          7494 => x"20",
          7495 => x"72",
          7496 => x"53",
          7497 => x"72",
          7498 => x"69",
          7499 => x"65",
          7500 => x"65",
          7501 => x"70",
          7502 => x"2e",
          7503 => x"69",
          7504 => x"72",
          7505 => x"75",
          7506 => x"62",
          7507 => x"4f",
          7508 => x"73",
          7509 => x"64",
          7510 => x"74",
          7511 => x"73",
          7512 => x"30",
          7513 => x"65",
          7514 => x"61",
          7515 => x"00",
          7516 => x"64",
          7517 => x"69",
          7518 => x"69",
          7519 => x"00",
          7520 => x"61",
          7521 => x"6e",
          7522 => x"50",
          7523 => x"64",
          7524 => x"2e",
          7525 => x"6f",
          7526 => x"6f",
          7527 => x"00",
          7528 => x"72",
          7529 => x"70",
          7530 => x"6e",
          7531 => x"61",
          7532 => x"6f",
          7533 => x"38",
          7534 => x"00",
          7535 => x"72",
          7536 => x"20",
          7537 => x"64",
          7538 => x"78",
          7539 => x"20",
          7540 => x"25",
          7541 => x"2e",
          7542 => x"20",
          7543 => x"00",
          7544 => x"20",
          7545 => x"6f",
          7546 => x"2e",
          7547 => x"30",
          7548 => x"78",
          7549 => x"78",
          7550 => x"00",
          7551 => x"6e",
          7552 => x"30",
          7553 => x"58",
          7554 => x"69",
          7555 => x"00",
          7556 => x"4d",
          7557 => x"43",
          7558 => x"2e",
          7559 => x"73",
          7560 => x"65",
          7561 => x"68",
          7562 => x"20",
          7563 => x"70",
          7564 => x"63",
          7565 => x"00",
          7566 => x"64",
          7567 => x"25",
          7568 => x"2e",
          7569 => x"6f",
          7570 => x"67",
          7571 => x"00",
          7572 => x"69",
          7573 => x"6c",
          7574 => x"3a",
          7575 => x"73",
          7576 => x"20",
          7577 => x"65",
          7578 => x"74",
          7579 => x"65",
          7580 => x"38",
          7581 => x"20",
          7582 => x"65",
          7583 => x"61",
          7584 => x"65",
          7585 => x"38",
          7586 => x"20",
          7587 => x"20",
          7588 => x"64",
          7589 => x"20",
          7590 => x"38",
          7591 => x"69",
          7592 => x"20",
          7593 => x"64",
          7594 => x"20",
          7595 => x"20",
          7596 => x"34",
          7597 => x"20",
          7598 => x"6d",
          7599 => x"46",
          7600 => x"20",
          7601 => x"2e",
          7602 => x"0a",
          7603 => x"69",
          7604 => x"53",
          7605 => x"6f",
          7606 => x"3d",
          7607 => x"64",
          7608 => x"20",
          7609 => x"20",
          7610 => x"72",
          7611 => x"20",
          7612 => x"2e",
          7613 => x"0a",
          7614 => x"50",
          7615 => x"53",
          7616 => x"4f",
          7617 => x"20",
          7618 => x"43",
          7619 => x"49",
          7620 => x"42",
          7621 => x"20",
          7622 => x"43",
          7623 => x"61",
          7624 => x"30",
          7625 => x"20",
          7626 => x"31",
          7627 => x"6d",
          7628 => x"30",
          7629 => x"20",
          7630 => x"52",
          7631 => x"76",
          7632 => x"30",
          7633 => x"20",
          7634 => x"20",
          7635 => x"38",
          7636 => x"2e",
          7637 => x"52",
          7638 => x"20",
          7639 => x"30",
          7640 => x"20",
          7641 => x"42",
          7642 => x"38",
          7643 => x"2e",
          7644 => x"44",
          7645 => x"20",
          7646 => x"30",
          7647 => x"20",
          7648 => x"52",
          7649 => x"38",
          7650 => x"2e",
          7651 => x"6d",
          7652 => x"6e",
          7653 => x"6e",
          7654 => x"56",
          7655 => x"6d",
          7656 => x"65",
          7657 => x"6c",
          7658 => x"56",
          7659 => x"00",
          7660 => x"00",
          7661 => x"00",
          7662 => x"00",
          7663 => x"00",
          7664 => x"00",
          7665 => x"00",
          7666 => x"00",
          7667 => x"00",
          7668 => x"00",
          7669 => x"00",
          7670 => x"00",
          7671 => x"00",
          7672 => x"00",
          7673 => x"00",
          7674 => x"00",
          7675 => x"00",
          7676 => x"00",
          7677 => x"00",
          7678 => x"00",
          7679 => x"00",
          7680 => x"00",
          7681 => x"00",
          7682 => x"00",
          7683 => x"00",
          7684 => x"00",
          7685 => x"00",
          7686 => x"00",
          7687 => x"00",
          7688 => x"00",
          7689 => x"00",
          7690 => x"00",
          7691 => x"00",
          7692 => x"5b",
          7693 => x"5b",
          7694 => x"5b",
          7695 => x"30",
          7696 => x"5b",
          7697 => x"00",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"00",
          7703 => x"74",
          7704 => x"72",
          7705 => x"73",
          7706 => x"6c",
          7707 => x"62",
          7708 => x"69",
          7709 => x"69",
          7710 => x"00",
          7711 => x"20",
          7712 => x"61",
          7713 => x"20",
          7714 => x"68",
          7715 => x"72",
          7716 => x"74",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"5b",
          7721 => x"5b",
          7722 => x"00",
          7723 => x"00",
          7724 => x"00",
          7725 => x"00",
          7726 => x"00",
          7727 => x"00",
          7728 => x"00",
          7729 => x"00",
          7730 => x"00",
          7731 => x"00",
          7732 => x"00",
          7733 => x"00",
          7734 => x"5b",
          7735 => x"5b",
          7736 => x"3a",
          7737 => x"64",
          7738 => x"25",
          7739 => x"00",
          7740 => x"25",
          7741 => x"3a",
          7742 => x"64",
          7743 => x"3a",
          7744 => x"30",
          7745 => x"63",
          7746 => x"00",
          7747 => x"74",
          7748 => x"3a",
          7749 => x"32",
          7750 => x"00",
          7751 => x"32",
          7752 => x"00",
          7753 => x"32",
          7754 => x"61",
          7755 => x"20",
          7756 => x"00",
          7757 => x"78",
          7758 => x"52",
          7759 => x"61",
          7760 => x"20",
          7761 => x"65",
          7762 => x"73",
          7763 => x"65",
          7764 => x"44",
          7765 => x"3f",
          7766 => x"2c",
          7767 => x"41",
          7768 => x"00",
          7769 => x"44",
          7770 => x"4f",
          7771 => x"20",
          7772 => x"20",
          7773 => x"4d",
          7774 => x"54",
          7775 => x"00",
          7776 => x"00",
          7777 => x"03",
          7778 => x"16",
          7779 => x"9a",
          7780 => x"45",
          7781 => x"92",
          7782 => x"99",
          7783 => x"49",
          7784 => x"a9",
          7785 => x"b1",
          7786 => x"b9",
          7787 => x"c1",
          7788 => x"c9",
          7789 => x"d1",
          7790 => x"d9",
          7791 => x"e1",
          7792 => x"e9",
          7793 => x"f1",
          7794 => x"f9",
          7795 => x"2e",
          7796 => x"22",
          7797 => x"00",
          7798 => x"10",
          7799 => x"00",
          7800 => x"04",
          7801 => x"00",
          7802 => x"e9",
          7803 => x"e5",
          7804 => x"e8",
          7805 => x"c4",
          7806 => x"c6",
          7807 => x"fb",
          7808 => x"dc",
          7809 => x"a7",
          7810 => x"f3",
          7811 => x"aa",
          7812 => x"ac",
          7813 => x"ab",
          7814 => x"93",
          7815 => x"62",
          7816 => x"51",
          7817 => x"5b",
          7818 => x"2c",
          7819 => x"5e",
          7820 => x"69",
          7821 => x"6c",
          7822 => x"65",
          7823 => x"53",
          7824 => x"0c",
          7825 => x"90",
          7826 => x"93",
          7827 => x"b5",
          7828 => x"a9",
          7829 => x"b5",
          7830 => x"65",
          7831 => x"f7",
          7832 => x"b7",
          7833 => x"a0",
          7834 => x"e0",
          7835 => x"ff",
          7836 => x"30",
          7837 => x"10",
          7838 => x"06",
          7839 => x"81",
          7840 => x"84",
          7841 => x"89",
          7842 => x"8d",
          7843 => x"91",
          7844 => x"f6",
          7845 => x"98",
          7846 => x"9d",
          7847 => x"a0",
          7848 => x"a4",
          7849 => x"a9",
          7850 => x"ac",
          7851 => x"b1",
          7852 => x"b5",
          7853 => x"b8",
          7854 => x"bc",
          7855 => x"c1",
          7856 => x"c5",
          7857 => x"c7",
          7858 => x"cd",
          7859 => x"8e",
          7860 => x"03",
          7861 => x"f8",
          7862 => x"3a",
          7863 => x"3b",
          7864 => x"40",
          7865 => x"0a",
          7866 => x"86",
          7867 => x"58",
          7868 => x"5c",
          7869 => x"93",
          7870 => x"64",
          7871 => x"97",
          7872 => x"6c",
          7873 => x"70",
          7874 => x"74",
          7875 => x"78",
          7876 => x"7c",
          7877 => x"a6",
          7878 => x"84",
          7879 => x"ae",
          7880 => x"45",
          7881 => x"90",
          7882 => x"03",
          7883 => x"ac",
          7884 => x"89",
          7885 => x"c2",
          7886 => x"c4",
          7887 => x"8c",
          7888 => x"18",
          7889 => x"f3",
          7890 => x"f7",
          7891 => x"fa",
          7892 => x"10",
          7893 => x"36",
          7894 => x"01",
          7895 => x"61",
          7896 => x"7d",
          7897 => x"96",
          7898 => x"08",
          7899 => x"08",
          7900 => x"06",
          7901 => x"52",
          7902 => x"56",
          7903 => x"70",
          7904 => x"c8",
          7905 => x"da",
          7906 => x"ea",
          7907 => x"80",
          7908 => x"a0",
          7909 => x"b8",
          7910 => x"cc",
          7911 => x"02",
          7912 => x"01",
          7913 => x"fc",
          7914 => x"70",
          7915 => x"83",
          7916 => x"2f",
          7917 => x"06",
          7918 => x"64",
          7919 => x"1a",
          7920 => x"00",
          7921 => x"00",
          7922 => x"00",
          7923 => x"00",
          7924 => x"00",
          7925 => x"00",
          7926 => x"00",
          7927 => x"00",
          7928 => x"00",
          7929 => x"00",
          7930 => x"00",
          7931 => x"00",
          7932 => x"00",
          7933 => x"00",
          7934 => x"00",
          7935 => x"00",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"00",
          7940 => x"00",
          7941 => x"00",
          7942 => x"00",
          7943 => x"00",
          7944 => x"00",
          7945 => x"00",
          7946 => x"00",
          7947 => x"00",
          7948 => x"00",
          7949 => x"00",
          7950 => x"00",
          7951 => x"00",
          7952 => x"00",
          7953 => x"00",
          7954 => x"00",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"00",
          7959 => x"00",
          7960 => x"00",
          7961 => x"00",
          7962 => x"00",
          7963 => x"00",
          7964 => x"00",
          7965 => x"00",
          7966 => x"00",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"00",
          7980 => x"81",
          7981 => x"7f",
          7982 => x"00",
          7983 => x"00",
          7984 => x"f5",
          7985 => x"00",
          7986 => x"01",
          7987 => x"00",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"00",
          7996 => x"00",
          7997 => x"00",
          7998 => x"00",
          7999 => x"00",
          8000 => x"00",
          8001 => x"00",
          8002 => x"00",
          8003 => x"fc",
          8004 => x"7a",
          8005 => x"72",
          8006 => x"6a",
          8007 => x"62",
          8008 => x"32",
          8009 => x"f3",
          8010 => x"7f",
          8011 => x"f0",
          8012 => x"81",
          8013 => x"fc",
          8014 => x"5a",
          8015 => x"52",
          8016 => x"4a",
          8017 => x"42",
          8018 => x"32",
          8019 => x"f3",
          8020 => x"7f",
          8021 => x"f0",
          8022 => x"81",
          8023 => x"fc",
          8024 => x"5a",
          8025 => x"52",
          8026 => x"4a",
          8027 => x"42",
          8028 => x"22",
          8029 => x"7e",
          8030 => x"e2",
          8031 => x"f0",
          8032 => x"86",
          8033 => x"fe",
          8034 => x"1a",
          8035 => x"12",
          8036 => x"0a",
          8037 => x"02",
          8038 => x"f0",
          8039 => x"1e",
          8040 => x"f0",
          8041 => x"f0",
          8042 => x"81",
          8043 => x"f0",
          8044 => x"77",
          8045 => x"70",
          8046 => x"5d",
          8047 => x"6e",
          8048 => x"36",
          8049 => x"9f",
          8050 => x"c5",
          8051 => x"f0",
          8052 => x"81",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"cf",
          9090 => x"fd",
          9091 => x"c5",
          9092 => x"ee",
          9093 => x"65",
          9094 => x"2a",
          9095 => x"25",
          9096 => x"2b",
          9097 => x"05",
          9098 => x"0d",
          9099 => x"15",
          9100 => x"54",
          9101 => x"85",
          9102 => x"8d",
          9103 => x"95",
          9104 => x"40",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"00",
          9113 => x"00",
          9114 => x"00",
          9115 => x"00",
          9116 => x"00",
          9117 => x"00",
          9118 => x"00",
          9119 => x"00",
          9120 => x"04",
          9121 => x"04",
        others => X"00"
    );

    shared variable RAM7 : ramArray :=
    (
             0 => x"f8",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"90",
             5 => x"8c",
             6 => x"00",
             7 => x"00",
             8 => x"72",
             9 => x"83",
            10 => x"04",
            11 => x"00",
            12 => x"83",
            13 => x"05",
            14 => x"73",
            15 => x"83",
            16 => x"72",
            17 => x"73",
            18 => x"53",
            19 => x"00",
            20 => x"73",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"0a",
            26 => x"05",
            27 => x"04",
            28 => x"73",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"cd",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"0a",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"09",
            45 => x"05",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"81",
            50 => x"04",
            51 => x"00",
            52 => x"04",
            53 => x"82",
            54 => x"fc",
            55 => x"00",
            56 => x"72",
            57 => x"0a",
            58 => x"00",
            59 => x"00",
            60 => x"72",
            61 => x"0a",
            62 => x"00",
            63 => x"00",
            64 => x"52",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"05",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"73",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"72",
            77 => x"10",
            78 => x"04",
            79 => x"00",
            80 => x"0b",
            81 => x"10",
            82 => x"93",
            83 => x"00",
            84 => x"90",
            85 => x"cc",
            86 => x"0c",
            87 => x"00",
            88 => x"90",
            89 => x"ab",
            90 => x"0c",
            91 => x"00",
            92 => x"05",
            93 => x"70",
            94 => x"05",
            95 => x"04",
            96 => x"05",
            97 => x"05",
            98 => x"74",
            99 => x"51",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"04",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"10",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"05",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"81",
           133 => x"0b",
           134 => x"0b",
           135 => x"b6",
           136 => x"0b",
           137 => x"0b",
           138 => x"f6",
           139 => x"0b",
           140 => x"0b",
           141 => x"b6",
           142 => x"0b",
           143 => x"0b",
           144 => x"f9",
           145 => x"0b",
           146 => x"0b",
           147 => x"bd",
           148 => x"0b",
           149 => x"0b",
           150 => x"81",
           151 => x"0b",
           152 => x"0b",
           153 => x"c5",
           154 => x"0b",
           155 => x"0b",
           156 => x"89",
           157 => x"0b",
           158 => x"0b",
           159 => x"cd",
           160 => x"0b",
           161 => x"0b",
           162 => x"91",
           163 => x"0b",
           164 => x"0b",
           165 => x"d5",
           166 => x"0b",
           167 => x"0b",
           168 => x"99",
           169 => x"0b",
           170 => x"0b",
           171 => x"dc",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"04",
           193 => x"2d",
           194 => x"90",
           195 => x"2d",
           196 => x"90",
           197 => x"2d",
           198 => x"90",
           199 => x"2d",
           200 => x"90",
           201 => x"2d",
           202 => x"90",
           203 => x"2d",
           204 => x"90",
           205 => x"2d",
           206 => x"90",
           207 => x"2d",
           208 => x"90",
           209 => x"2d",
           210 => x"90",
           211 => x"2d",
           212 => x"90",
           213 => x"2d",
           214 => x"90",
           215 => x"2d",
           216 => x"90",
           217 => x"db",
           218 => x"80",
           219 => x"d5",
           220 => x"c0",
           221 => x"80",
           222 => x"80",
           223 => x"0c",
           224 => x"08",
           225 => x"98",
           226 => x"98",
           227 => x"ba",
           228 => x"ba",
           229 => x"84",
           230 => x"84",
           231 => x"04",
           232 => x"2d",
           233 => x"90",
           234 => x"e6",
           235 => x"80",
           236 => x"fa",
           237 => x"c0",
           238 => x"82",
           239 => x"80",
           240 => x"0c",
           241 => x"08",
           242 => x"98",
           243 => x"98",
           244 => x"ba",
           245 => x"ba",
           246 => x"84",
           247 => x"84",
           248 => x"04",
           249 => x"2d",
           250 => x"90",
           251 => x"cf",
           252 => x"80",
           253 => x"f6",
           254 => x"c0",
           255 => x"83",
           256 => x"80",
           257 => x"0c",
           258 => x"08",
           259 => x"98",
           260 => x"98",
           261 => x"ba",
           262 => x"ba",
           263 => x"84",
           264 => x"84",
           265 => x"04",
           266 => x"2d",
           267 => x"90",
           268 => x"e3",
           269 => x"80",
           270 => x"9a",
           271 => x"c0",
           272 => x"83",
           273 => x"80",
           274 => x"0c",
           275 => x"08",
           276 => x"98",
           277 => x"98",
           278 => x"ba",
           279 => x"ba",
           280 => x"84",
           281 => x"84",
           282 => x"04",
           283 => x"2d",
           284 => x"90",
           285 => x"ab",
           286 => x"80",
           287 => x"f6",
           288 => x"c0",
           289 => x"80",
           290 => x"80",
           291 => x"0c",
           292 => x"08",
           293 => x"98",
           294 => x"98",
           295 => x"ba",
           296 => x"98",
           297 => x"ba",
           298 => x"ba",
           299 => x"84",
           300 => x"84",
           301 => x"04",
           302 => x"2d",
           303 => x"90",
           304 => x"da",
           305 => x"80",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"00",
           311 => x"09",
           312 => x"2b",
           313 => x"04",
           314 => x"05",
           315 => x"72",
           316 => x"51",
           317 => x"70",
           318 => x"71",
           319 => x"0b",
           320 => x"ce",
           321 => x"3d",
           322 => x"53",
           323 => x"81",
           324 => x"3d",
           325 => x"81",
           326 => x"56",
           327 => x"2e",
           328 => x"14",
           329 => x"72",
           330 => x"54",
           331 => x"2e",
           332 => x"84",
           333 => x"08",
           334 => x"08",
           335 => x"14",
           336 => x"07",
           337 => x"80",
           338 => x"52",
           339 => x"0d",
           340 => x"88",
           341 => x"54",
           342 => x"73",
           343 => x"05",
           344 => x"51",
           345 => x"34",
           346 => x"86",
           347 => x"51",
           348 => x"3d",
           349 => x"80",
           350 => x"70",
           351 => x"55",
           352 => x"81",
           353 => x"76",
           354 => x"7b",
           355 => x"81",
           356 => x"26",
           357 => x"30",
           358 => x"ae",
           359 => x"83",
           360 => x"54",
           361 => x"80",
           362 => x"bd",
           363 => x"ba",
           364 => x"83",
           365 => x"10",
           366 => x"19",
           367 => x"05",
           368 => x"5f",
           369 => x"81",
           370 => x"7c",
           371 => x"ff",
           372 => x"06",
           373 => x"5b",
           374 => x"dd",
           375 => x"51",
           376 => x"fe",
           377 => x"2a",
           378 => x"38",
           379 => x"95",
           380 => x"26",
           381 => x"cc",
           382 => x"18",
           383 => x"38",
           384 => x"80",
           385 => x"38",
           386 => x"f6",
           387 => x"71",
           388 => x"58",
           389 => x"52",
           390 => x"8c",
           391 => x"08",
           392 => x"26",
           393 => x"05",
           394 => x"34",
           395 => x"84",
           396 => x"08",
           397 => x"98",
           398 => x"80",
           399 => x"29",
           400 => x"59",
           401 => x"55",
           402 => x"84",
           403 => x"53",
           404 => x"80",
           405 => x"72",
           406 => x"81",
           407 => x"38",
           408 => x"54",
           409 => x"7a",
           410 => x"71",
           411 => x"06",
           412 => x"77",
           413 => x"7c",
           414 => x"80",
           415 => x"81",
           416 => x"84",
           417 => x"38",
           418 => x"86",
           419 => x"85",
           420 => x"5f",
           421 => x"84",
           422 => x"70",
           423 => x"25",
           424 => x"a9",
           425 => x"fc",
           426 => x"40",
           427 => x"81",
           428 => x"78",
           429 => x"0a",
           430 => x"80",
           431 => x"51",
           432 => x"0a",
           433 => x"2c",
           434 => x"38",
           435 => x"55",
           436 => x"80",
           437 => x"f3",
           438 => x"2e",
           439 => x"2e",
           440 => x"33",
           441 => x"ba",
           442 => x"74",
           443 => x"a7",
           444 => x"fc",
           445 => x"40",
           446 => x"7c",
           447 => x"39",
           448 => x"7c",
           449 => x"fa",
           450 => x"80",
           451 => x"71",
           452 => x"59",
           453 => x"60",
           454 => x"83",
           455 => x"7c",
           456 => x"05",
           457 => x"57",
           458 => x"06",
           459 => x"78",
           460 => x"05",
           461 => x"7f",
           462 => x"51",
           463 => x"70",
           464 => x"83",
           465 => x"52",
           466 => x"85",
           467 => x"83",
           468 => x"ff",
           469 => x"75",
           470 => x"b9",
           471 => x"81",
           472 => x"29",
           473 => x"5a",
           474 => x"70",
           475 => x"c6",
           476 => x"05",
           477 => x"80",
           478 => x"ff",
           479 => x"fa",
           480 => x"58",
           481 => x"39",
           482 => x"58",
           483 => x"39",
           484 => x"81",
           485 => x"8a",
           486 => x"ba",
           487 => x"71",
           488 => x"2c",
           489 => x"07",
           490 => x"38",
           491 => x"71",
           492 => x"54",
           493 => x"bb",
           494 => x"ff",
           495 => x"5a",
           496 => x"33",
           497 => x"c9",
           498 => x"fc",
           499 => x"54",
           500 => x"7c",
           501 => x"39",
           502 => x"79",
           503 => x"38",
           504 => x"7a",
           505 => x"2e",
           506 => x"98",
           507 => x"90",
           508 => x"51",
           509 => x"39",
           510 => x"7e",
           511 => x"a2",
           512 => x"98",
           513 => x"06",
           514 => x"fb",
           515 => x"70",
           516 => x"7c",
           517 => x"39",
           518 => x"ff",
           519 => x"8b",
           520 => x"ff",
           521 => x"5a",
           522 => x"30",
           523 => x"5b",
           524 => x"d5",
           525 => x"f3",
           526 => x"3d",
           527 => x"f0",
           528 => x"81",
           529 => x"55",
           530 => x"81",
           531 => x"05",
           532 => x"38",
           533 => x"90",
           534 => x"8c",
           535 => x"74",
           536 => x"80",
           537 => x"54",
           538 => x"84",
           539 => x"14",
           540 => x"08",
           541 => x"56",
           542 => x"0d",
           543 => x"54",
           544 => x"2a",
           545 => x"57",
           546 => x"81",
           547 => x"55",
           548 => x"06",
           549 => x"8c",
           550 => x"81",
           551 => x"ea",
           552 => x"08",
           553 => x"80",
           554 => x"05",
           555 => x"ca",
           556 => x"08",
           557 => x"0d",
           558 => x"11",
           559 => x"06",
           560 => x"ae",
           561 => x"73",
           562 => x"53",
           563 => x"74",
           564 => x"81",
           565 => x"81",
           566 => x"84",
           567 => x"74",
           568 => x"15",
           569 => x"ba",
           570 => x"81",
           571 => x"39",
           572 => x"70",
           573 => x"06",
           574 => x"b3",
           575 => x"71",
           576 => x"52",
           577 => x"08",
           578 => x"80",
           579 => x"16",
           580 => x"81",
           581 => x"0c",
           582 => x"06",
           583 => x"08",
           584 => x"33",
           585 => x"04",
           586 => x"2d",
           587 => x"8c",
           588 => x"16",
           589 => x"ba",
           590 => x"a0",
           591 => x"54",
           592 => x"0d",
           593 => x"17",
           594 => x"0d",
           595 => x"70",
           596 => x"38",
           597 => x"54",
           598 => x"54",
           599 => x"8c",
           600 => x"0d",
           601 => x"54",
           602 => x"27",
           603 => x"71",
           604 => x"81",
           605 => x"ef",
           606 => x"3d",
           607 => x"27",
           608 => x"ff",
           609 => x"73",
           610 => x"d9",
           611 => x"71",
           612 => x"df",
           613 => x"70",
           614 => x"33",
           615 => x"74",
           616 => x"3d",
           617 => x"71",
           618 => x"54",
           619 => x"54",
           620 => x"8c",
           621 => x"0d",
           622 => x"54",
           623 => x"81",
           624 => x"55",
           625 => x"73",
           626 => x"04",
           627 => x"56",
           628 => x"33",
           629 => x"52",
           630 => x"38",
           631 => x"38",
           632 => x"51",
           633 => x"0d",
           634 => x"33",
           635 => x"38",
           636 => x"80",
           637 => x"ba",
           638 => x"84",
           639 => x"fb",
           640 => x"56",
           641 => x"84",
           642 => x"81",
           643 => x"54",
           644 => x"38",
           645 => x"74",
           646 => x"8c",
           647 => x"8c",
           648 => x"87",
           649 => x"77",
           650 => x"80",
           651 => x"54",
           652 => x"ff",
           653 => x"06",
           654 => x"52",
           655 => x"3d",
           656 => x"79",
           657 => x"2e",
           658 => x"54",
           659 => x"73",
           660 => x"04",
           661 => x"a0",
           662 => x"51",
           663 => x"52",
           664 => x"38",
           665 => x"ba",
           666 => x"9f",
           667 => x"9f",
           668 => x"71",
           669 => x"57",
           670 => x"2e",
           671 => x"07",
           672 => x"ff",
           673 => x"72",
           674 => x"56",
           675 => x"da",
           676 => x"84",
           677 => x"fc",
           678 => x"06",
           679 => x"70",
           680 => x"2a",
           681 => x"70",
           682 => x"74",
           683 => x"30",
           684 => x"31",
           685 => x"05",
           686 => x"25",
           687 => x"70",
           688 => x"70",
           689 => x"05",
           690 => x"55",
           691 => x"55",
           692 => x"56",
           693 => x"3d",
           694 => x"54",
           695 => x"08",
           696 => x"8c",
           697 => x"3d",
           698 => x"76",
           699 => x"cf",
           700 => x"13",
           701 => x"51",
           702 => x"08",
           703 => x"80",
           704 => x"be",
           705 => x"72",
           706 => x"55",
           707 => x"72",
           708 => x"77",
           709 => x"2c",
           710 => x"71",
           711 => x"55",
           712 => x"84",
           713 => x"fa",
           714 => x"2c",
           715 => x"2c",
           716 => x"31",
           717 => x"59",
           718 => x"8c",
           719 => x"8c",
           720 => x"0d",
           721 => x"0c",
           722 => x"73",
           723 => x"81",
           724 => x"55",
           725 => x"2e",
           726 => x"83",
           727 => x"89",
           728 => x"56",
           729 => x"e0",
           730 => x"81",
           731 => x"81",
           732 => x"8f",
           733 => x"54",
           734 => x"72",
           735 => x"29",
           736 => x"33",
           737 => x"be",
           738 => x"30",
           739 => x"84",
           740 => x"81",
           741 => x"56",
           742 => x"06",
           743 => x"0c",
           744 => x"2e",
           745 => x"2e",
           746 => x"c6",
           747 => x"58",
           748 => x"84",
           749 => x"82",
           750 => x"33",
           751 => x"80",
           752 => x"0d",
           753 => x"57",
           754 => x"33",
           755 => x"81",
           756 => x"0c",
           757 => x"f3",
           758 => x"73",
           759 => x"58",
           760 => x"38",
           761 => x"80",
           762 => x"38",
           763 => x"53",
           764 => x"53",
           765 => x"70",
           766 => x"27",
           767 => x"83",
           768 => x"70",
           769 => x"73",
           770 => x"2e",
           771 => x"0c",
           772 => x"8b",
           773 => x"79",
           774 => x"b0",
           775 => x"81",
           776 => x"55",
           777 => x"58",
           778 => x"56",
           779 => x"53",
           780 => x"fe",
           781 => x"8b",
           782 => x"70",
           783 => x"56",
           784 => x"8c",
           785 => x"dc",
           786 => x"06",
           787 => x"0d",
           788 => x"71",
           789 => x"71",
           790 => x"be",
           791 => x"f4",
           792 => x"04",
           793 => x"83",
           794 => x"ef",
           795 => x"cf",
           796 => x"0d",
           797 => x"3f",
           798 => x"51",
           799 => x"83",
           800 => x"3d",
           801 => x"e6",
           802 => x"b8",
           803 => x"04",
           804 => x"83",
           805 => x"ee",
           806 => x"d1",
           807 => x"0d",
           808 => x"3f",
           809 => x"51",
           810 => x"83",
           811 => x"3d",
           812 => x"8e",
           813 => x"e0",
           814 => x"04",
           815 => x"83",
           816 => x"ed",
           817 => x"d2",
           818 => x"0d",
           819 => x"05",
           820 => x"68",
           821 => x"51",
           822 => x"ff",
           823 => x"07",
           824 => x"57",
           825 => x"52",
           826 => x"a2",
           827 => x"ba",
           828 => x"77",
           829 => x"70",
           830 => x"9f",
           831 => x"77",
           832 => x"88",
           833 => x"e0",
           834 => x"51",
           835 => x"54",
           836 => x"d2",
           837 => x"ba",
           838 => x"ba",
           839 => x"84",
           840 => x"05",
           841 => x"51",
           842 => x"08",
           843 => x"38",
           844 => x"38",
           845 => x"39",
           846 => x"3f",
           847 => x"f4",
           848 => x"83",
           849 => x"98",
           850 => x"f8",
           851 => x"05",
           852 => x"7b",
           853 => x"ba",
           854 => x"91",
           855 => x"84",
           856 => x"78",
           857 => x"60",
           858 => x"7e",
           859 => x"84",
           860 => x"f3",
           861 => x"05",
           862 => x"68",
           863 => x"78",
           864 => x"83",
           865 => x"d2",
           866 => x"73",
           867 => x"81",
           868 => x"38",
           869 => x"a7",
           870 => x"51",
           871 => x"f0",
           872 => x"3f",
           873 => x"d8",
           874 => x"79",
           875 => x"33",
           876 => x"83",
           877 => x"27",
           878 => x"70",
           879 => x"2e",
           880 => x"ee",
           881 => x"51",
           882 => x"76",
           883 => x"e9",
           884 => x"58",
           885 => x"8c",
           886 => x"54",
           887 => x"9b",
           888 => x"76",
           889 => x"84",
           890 => x"83",
           891 => x"14",
           892 => x"51",
           893 => x"b8",
           894 => x"51",
           895 => x"f0",
           896 => x"3f",
           897 => x"18",
           898 => x"22",
           899 => x"3f",
           900 => x"54",
           901 => x"26",
           902 => x"ec",
           903 => x"d5",
           904 => x"a9",
           905 => x"73",
           906 => x"72",
           907 => x"ab",
           908 => x"53",
           909 => x"74",
           910 => x"d5",
           911 => x"3f",
           912 => x"ce",
           913 => x"ff",
           914 => x"fc",
           915 => x"2e",
           916 => x"59",
           917 => x"3f",
           918 => x"98",
           919 => x"9b",
           920 => x"75",
           921 => x"58",
           922 => x"80",
           923 => x"08",
           924 => x"32",
           925 => x"70",
           926 => x"55",
           927 => x"24",
           928 => x"0b",
           929 => x"04",
           930 => x"08",
           931 => x"f7",
           932 => x"3f",
           933 => x"2a",
           934 => x"b7",
           935 => x"51",
           936 => x"2a",
           937 => x"db",
           938 => x"51",
           939 => x"2a",
           940 => x"ff",
           941 => x"51",
           942 => x"2a",
           943 => x"38",
           944 => x"88",
           945 => x"04",
           946 => x"cc",
           947 => x"f7",
           948 => x"04",
           949 => x"e0",
           950 => x"df",
           951 => x"72",
           952 => x"51",
           953 => x"9b",
           954 => x"72",
           955 => x"71",
           956 => x"81",
           957 => x"51",
           958 => x"3f",
           959 => x"52",
           960 => x"be",
           961 => x"d4",
           962 => x"9a",
           963 => x"06",
           964 => x"38",
           965 => x"3f",
           966 => x"80",
           967 => x"70",
           968 => x"fe",
           969 => x"9a",
           970 => x"d7",
           971 => x"83",
           972 => x"80",
           973 => x"81",
           974 => x"51",
           975 => x"3f",
           976 => x"52",
           977 => x"bd",
           978 => x"41",
           979 => x"81",
           980 => x"84",
           981 => x"3d",
           982 => x"38",
           983 => x"98",
           984 => x"c3",
           985 => x"52",
           986 => x"83",
           987 => x"5b",
           988 => x"79",
           989 => x"ff",
           990 => x"38",
           991 => x"83",
           992 => x"2e",
           993 => x"70",
           994 => x"38",
           995 => x"7b",
           996 => x"08",
           997 => x"8c",
           998 => x"53",
           999 => x"84",
          1000 => x"33",
          1001 => x"81",
          1002 => x"9b",
          1003 => x"5c",
          1004 => x"f8",
          1005 => x"ba",
          1006 => x"80",
          1007 => x"08",
          1008 => x"91",
          1009 => x"62",
          1010 => x"84",
          1011 => x"8b",
          1012 => x"80",
          1013 => x"5b",
          1014 => x"82",
          1015 => x"82",
          1016 => x"d5",
          1017 => x"83",
          1018 => x"7d",
          1019 => x"0a",
          1020 => x"f5",
          1021 => x"ba",
          1022 => x"07",
          1023 => x"5a",
          1024 => x"78",
          1025 => x"38",
          1026 => x"5a",
          1027 => x"61",
          1028 => x"38",
          1029 => x"51",
          1030 => x"51",
          1031 => x"53",
          1032 => x"0b",
          1033 => x"ff",
          1034 => x"81",
          1035 => x"9c",
          1036 => x"8c",
          1037 => x"0b",
          1038 => x"53",
          1039 => x"91",
          1040 => x"a0",
          1041 => x"e6",
          1042 => x"70",
          1043 => x"2e",
          1044 => x"39",
          1045 => x"3f",
          1046 => x"34",
          1047 => x"7e",
          1048 => x"5a",
          1049 => x"1a",
          1050 => x"81",
          1051 => x"10",
          1052 => x"04",
          1053 => x"9a",
          1054 => x"52",
          1055 => x"7e",
          1056 => x"c3",
          1057 => x"09",
          1058 => x"9a",
          1059 => x"83",
          1060 => x"51",
          1061 => x"83",
          1062 => x"98",
          1063 => x"7c",
          1064 => x"81",
          1065 => x"dd",
          1066 => x"51",
          1067 => x"8e",
          1068 => x"ac",
          1069 => x"04",
          1070 => x"d0",
          1071 => x"ff",
          1072 => x"ec",
          1073 => x"2e",
          1074 => x"dc",
          1075 => x"2d",
          1076 => x"9a",
          1077 => x"d6",
          1078 => x"39",
          1079 => x"80",
          1080 => x"8c",
          1081 => x"52",
          1082 => x"68",
          1083 => x"11",
          1084 => x"3f",
          1085 => x"d2",
          1086 => x"ff",
          1087 => x"ba",
          1088 => x"78",
          1089 => x"51",
          1090 => x"53",
          1091 => x"3f",
          1092 => x"2e",
          1093 => x"d3",
          1094 => x"cf",
          1095 => x"ff",
          1096 => x"ba",
          1097 => x"b8",
          1098 => x"05",
          1099 => x"08",
          1100 => x"53",
          1101 => x"9b",
          1102 => x"f8",
          1103 => x"48",
          1104 => x"ba",
          1105 => x"64",
          1106 => x"b8",
          1107 => x"05",
          1108 => x"08",
          1109 => x"fe",
          1110 => x"e9",
          1111 => x"2e",
          1112 => x"11",
          1113 => x"3f",
          1114 => x"ea",
          1115 => x"3f",
          1116 => x"83",
          1117 => x"5f",
          1118 => x"7a",
          1119 => x"52",
          1120 => x"66",
          1121 => x"47",
          1122 => x"11",
          1123 => x"3f",
          1124 => x"9a",
          1125 => x"ff",
          1126 => x"ba",
          1127 => x"b8",
          1128 => x"05",
          1129 => x"08",
          1130 => x"f8",
          1131 => x"67",
          1132 => x"70",
          1133 => x"81",
          1134 => x"84",
          1135 => x"89",
          1136 => x"f6",
          1137 => x"53",
          1138 => x"84",
          1139 => x"33",
          1140 => x"e3",
          1141 => x"f8",
          1142 => x"48",
          1143 => x"82",
          1144 => x"68",
          1145 => x"02",
          1146 => x"81",
          1147 => x"53",
          1148 => x"84",
          1149 => x"38",
          1150 => x"79",
          1151 => x"fe",
          1152 => x"e7",
          1153 => x"bd",
          1154 => x"84",
          1155 => x"e9",
          1156 => x"f5",
          1157 => x"53",
          1158 => x"84",
          1159 => x"38",
          1160 => x"80",
          1161 => x"8c",
          1162 => x"46",
          1163 => x"68",
          1164 => x"38",
          1165 => x"5b",
          1166 => x"51",
          1167 => x"3d",
          1168 => x"84",
          1169 => x"05",
          1170 => x"84",
          1171 => x"f9",
          1172 => x"f4",
          1173 => x"e7",
          1174 => x"ff",
          1175 => x"e5",
          1176 => x"38",
          1177 => x"2e",
          1178 => x"49",
          1179 => x"80",
          1180 => x"8c",
          1181 => x"5a",
          1182 => x"f2",
          1183 => x"11",
          1184 => x"3f",
          1185 => x"38",
          1186 => x"83",
          1187 => x"30",
          1188 => x"5c",
          1189 => x"7a",
          1190 => x"d8",
          1191 => x"68",
          1192 => x"eb",
          1193 => x"a6",
          1194 => x"0c",
          1195 => x"fe",
          1196 => x"e2",
          1197 => x"2e",
          1198 => x"59",
          1199 => x"f0",
          1200 => x"fd",
          1201 => x"f2",
          1202 => x"05",
          1203 => x"7d",
          1204 => x"ff",
          1205 => x"ba",
          1206 => x"64",
          1207 => x"70",
          1208 => x"3d",
          1209 => x"51",
          1210 => x"ff",
          1211 => x"fe",
          1212 => x"e3",
          1213 => x"2e",
          1214 => x"db",
          1215 => x"49",
          1216 => x"11",
          1217 => x"3f",
          1218 => x"98",
          1219 => x"84",
          1220 => x"7a",
          1221 => x"38",
          1222 => x"53",
          1223 => x"eb",
          1224 => x"51",
          1225 => x"d8",
          1226 => x"39",
          1227 => x"80",
          1228 => x"8c",
          1229 => x"02",
          1230 => x"05",
          1231 => x"83",
          1232 => x"80",
          1233 => x"fc",
          1234 => x"7b",
          1235 => x"08",
          1236 => x"51",
          1237 => x"39",
          1238 => x"64",
          1239 => x"33",
          1240 => x"f2",
          1241 => x"d8",
          1242 => x"39",
          1243 => x"2e",
          1244 => x"fc",
          1245 => x"7d",
          1246 => x"08",
          1247 => x"33",
          1248 => x"f2",
          1249 => x"f3",
          1250 => x"38",
          1251 => x"39",
          1252 => x"2e",
          1253 => x"fb",
          1254 => x"80",
          1255 => x"f8",
          1256 => x"f3",
          1257 => x"34",
          1258 => x"57",
          1259 => x"c8",
          1260 => x"77",
          1261 => x"75",
          1262 => x"8c",
          1263 => x"9c",
          1264 => x"52",
          1265 => x"8c",
          1266 => x"87",
          1267 => x"3f",
          1268 => x"0c",
          1269 => x"84",
          1270 => x"94",
          1271 => x"c7",
          1272 => x"05",
          1273 => x"89",
          1274 => x"0c",
          1275 => x"3f",
          1276 => x"8d",
          1277 => x"52",
          1278 => x"83",
          1279 => x"87",
          1280 => x"90",
          1281 => x"98",
          1282 => x"ec",
          1283 => x"77",
          1284 => x"53",
          1285 => x"33",
          1286 => x"a0",
          1287 => x"15",
          1288 => x"53",
          1289 => x"81",
          1290 => x"82",
          1291 => x"e7",
          1292 => x"06",
          1293 => x"38",
          1294 => x"73",
          1295 => x"e1",
          1296 => x"54",
          1297 => x"38",
          1298 => x"70",
          1299 => x"72",
          1300 => x"81",
          1301 => x"51",
          1302 => x"0d",
          1303 => x"80",
          1304 => x"80",
          1305 => x"54",
          1306 => x"54",
          1307 => x"53",
          1308 => x"fe",
          1309 => x"76",
          1310 => x"84",
          1311 => x"86",
          1312 => x"fd",
          1313 => x"e5",
          1314 => x"3d",
          1315 => x"11",
          1316 => x"70",
          1317 => x"33",
          1318 => x"26",
          1319 => x"83",
          1320 => x"85",
          1321 => x"26",
          1322 => x"85",
          1323 => x"88",
          1324 => x"e7",
          1325 => x"54",
          1326 => x"cc",
          1327 => x"0c",
          1328 => x"82",
          1329 => x"83",
          1330 => x"84",
          1331 => x"85",
          1332 => x"86",
          1333 => x"74",
          1334 => x"c0",
          1335 => x"98",
          1336 => x"8c",
          1337 => x"0d",
          1338 => x"81",
          1339 => x"5e",
          1340 => x"08",
          1341 => x"98",
          1342 => x"87",
          1343 => x"1c",
          1344 => x"79",
          1345 => x"08",
          1346 => x"98",
          1347 => x"87",
          1348 => x"1c",
          1349 => x"ff",
          1350 => x"58",
          1351 => x"56",
          1352 => x"54",
          1353 => x"ff",
          1354 => x"bf",
          1355 => x"3d",
          1356 => x"81",
          1357 => x"b1",
          1358 => x"70",
          1359 => x"09",
          1360 => x"e3",
          1361 => x"3d",
          1362 => x"3f",
          1363 => x"98",
          1364 => x"81",
          1365 => x"f1",
          1366 => x"70",
          1367 => x"d2",
          1368 => x"70",
          1369 => x"51",
          1370 => x"08",
          1371 => x"71",
          1372 => x"81",
          1373 => x"38",
          1374 => x"0d",
          1375 => x"33",
          1376 => x"06",
          1377 => x"f4",
          1378 => x"96",
          1379 => x"70",
          1380 => x"70",
          1381 => x"72",
          1382 => x"2e",
          1383 => x"52",
          1384 => x"51",
          1385 => x"2e",
          1386 => x"74",
          1387 => x"86",
          1388 => x"81",
          1389 => x"81",
          1390 => x"cb",
          1391 => x"71",
          1392 => x"84",
          1393 => x"53",
          1394 => x"ff",
          1395 => x"30",
          1396 => x"83",
          1397 => x"fa",
          1398 => x"70",
          1399 => x"e7",
          1400 => x"70",
          1401 => x"80",
          1402 => x"94",
          1403 => x"53",
          1404 => x"71",
          1405 => x"70",
          1406 => x"53",
          1407 => x"2a",
          1408 => x"81",
          1409 => x"52",
          1410 => x"94",
          1411 => x"75",
          1412 => x"76",
          1413 => x"04",
          1414 => x"51",
          1415 => x"06",
          1416 => x"93",
          1417 => x"ff",
          1418 => x"70",
          1419 => x"52",
          1420 => x"0d",
          1421 => x"2a",
          1422 => x"84",
          1423 => x"83",
          1424 => x"08",
          1425 => x"94",
          1426 => x"9e",
          1427 => x"c0",
          1428 => x"87",
          1429 => x"0c",
          1430 => x"e0",
          1431 => x"f2",
          1432 => x"83",
          1433 => x"08",
          1434 => x"bc",
          1435 => x"9e",
          1436 => x"c0",
          1437 => x"87",
          1438 => x"f2",
          1439 => x"83",
          1440 => x"08",
          1441 => x"8c",
          1442 => x"83",
          1443 => x"9e",
          1444 => x"51",
          1445 => x"83",
          1446 => x"9e",
          1447 => x"51",
          1448 => x"81",
          1449 => x"0b",
          1450 => x"80",
          1451 => x"2e",
          1452 => x"8f",
          1453 => x"08",
          1454 => x"52",
          1455 => x"71",
          1456 => x"c0",
          1457 => x"06",
          1458 => x"38",
          1459 => x"80",
          1460 => x"90",
          1461 => x"80",
          1462 => x"f3",
          1463 => x"90",
          1464 => x"52",
          1465 => x"52",
          1466 => x"87",
          1467 => x"80",
          1468 => x"83",
          1469 => x"34",
          1470 => x"70",
          1471 => x"70",
          1472 => x"83",
          1473 => x"9e",
          1474 => x"51",
          1475 => x"81",
          1476 => x"0b",
          1477 => x"80",
          1478 => x"83",
          1479 => x"34",
          1480 => x"06",
          1481 => x"f3",
          1482 => x"90",
          1483 => x"52",
          1484 => x"71",
          1485 => x"90",
          1486 => x"53",
          1487 => x"0b",
          1488 => x"06",
          1489 => x"38",
          1490 => x"87",
          1491 => x"70",
          1492 => x"04",
          1493 => x"0d",
          1494 => x"3f",
          1495 => x"aa",
          1496 => x"3f",
          1497 => x"fa",
          1498 => x"85",
          1499 => x"75",
          1500 => x"55",
          1501 => x"33",
          1502 => x"97",
          1503 => x"f3",
          1504 => x"83",
          1505 => x"38",
          1506 => x"cf",
          1507 => x"83",
          1508 => x"74",
          1509 => x"56",
          1510 => x"33",
          1511 => x"b8",
          1512 => x"08",
          1513 => x"bb",
          1514 => x"d9",
          1515 => x"f2",
          1516 => x"ff",
          1517 => x"c2",
          1518 => x"83",
          1519 => x"83",
          1520 => x"52",
          1521 => x"8c",
          1522 => x"31",
          1523 => x"83",
          1524 => x"83",
          1525 => x"38",
          1526 => x"38",
          1527 => x"0d",
          1528 => x"84",
          1529 => x"84",
          1530 => x"76",
          1531 => x"08",
          1532 => x"a3",
          1533 => x"3d",
          1534 => x"bd",
          1535 => x"3f",
          1536 => x"29",
          1537 => x"8c",
          1538 => x"b3",
          1539 => x"74",
          1540 => x"39",
          1541 => x"83",
          1542 => x"f2",
          1543 => x"ff",
          1544 => x"52",
          1545 => x"3f",
          1546 => x"94",
          1547 => x"bc",
          1548 => x"22",
          1549 => x"9b",
          1550 => x"84",
          1551 => x"84",
          1552 => x"76",
          1553 => x"08",
          1554 => x"f3",
          1555 => x"80",
          1556 => x"83",
          1557 => x"83",
          1558 => x"fd",
          1559 => x"80",
          1560 => x"95",
          1561 => x"38",
          1562 => x"bf",
          1563 => x"74",
          1564 => x"83",
          1565 => x"83",
          1566 => x"fc",
          1567 => x"33",
          1568 => x"83",
          1569 => x"80",
          1570 => x"f3",
          1571 => x"ff",
          1572 => x"55",
          1573 => x"39",
          1574 => x"ec",
          1575 => x"9b",
          1576 => x"38",
          1577 => x"f2",
          1578 => x"8c",
          1579 => x"97",
          1580 => x"38",
          1581 => x"f2",
          1582 => x"a8",
          1583 => x"92",
          1584 => x"38",
          1585 => x"f2",
          1586 => x"c4",
          1587 => x"91",
          1588 => x"38",
          1589 => x"f2",
          1590 => x"e0",
          1591 => x"90",
          1592 => x"38",
          1593 => x"f2",
          1594 => x"fc",
          1595 => x"93",
          1596 => x"38",
          1597 => x"b0",
          1598 => x"bc",
          1599 => x"74",
          1600 => x"ff",
          1601 => x"71",
          1602 => x"83",
          1603 => x"83",
          1604 => x"83",
          1605 => x"ff",
          1606 => x"83",
          1607 => x"83",
          1608 => x"ff",
          1609 => x"83",
          1610 => x"83",
          1611 => x"ff",
          1612 => x"71",
          1613 => x"c0",
          1614 => x"08",
          1615 => x"3d",
          1616 => x"5a",
          1617 => x"83",
          1618 => x"3f",
          1619 => x"8b",
          1620 => x"08",
          1621 => x"82",
          1622 => x"80",
          1623 => x"3f",
          1624 => x"55",
          1625 => x"8e",
          1626 => x"70",
          1627 => x"09",
          1628 => x"51",
          1629 => x"73",
          1630 => x"8c",
          1631 => x"3f",
          1632 => x"76",
          1633 => x"0c",
          1634 => x"51",
          1635 => x"09",
          1636 => x"51",
          1637 => x"fb",
          1638 => x"8c",
          1639 => x"b0",
          1640 => x"84",
          1641 => x"d8",
          1642 => x"08",
          1643 => x"5a",
          1644 => x"80",
          1645 => x"10",
          1646 => x"52",
          1647 => x"8c",
          1648 => x"c0",
          1649 => x"38",
          1650 => x"81",
          1651 => x"81",
          1652 => x"82",
          1653 => x"84",
          1654 => x"81",
          1655 => x"53",
          1656 => x"84",
          1657 => x"ff",
          1658 => x"a6",
          1659 => x"06",
          1660 => x"16",
          1661 => x"76",
          1662 => x"78",
          1663 => x"fe",
          1664 => x"33",
          1665 => x"06",
          1666 => x"38",
          1667 => x"cd",
          1668 => x"83",
          1669 => x"b9",
          1670 => x"38",
          1671 => x"52",
          1672 => x"ba",
          1673 => x"51",
          1674 => x"08",
          1675 => x"25",
          1676 => x"05",
          1677 => x"77",
          1678 => x"f8",
          1679 => x"ff",
          1680 => x"81",
          1681 => x"0d",
          1682 => x"b7",
          1683 => x"5c",
          1684 => x"fc",
          1685 => x"74",
          1686 => x"56",
          1687 => x"77",
          1688 => x"77",
          1689 => x"77",
          1690 => x"b4",
          1691 => x"3f",
          1692 => x"98",
          1693 => x"38",
          1694 => x"33",
          1695 => x"d1",
          1696 => x"2c",
          1697 => x"83",
          1698 => x"33",
          1699 => x"58",
          1700 => x"80",
          1701 => x"38",
          1702 => x"0a",
          1703 => x"76",
          1704 => x"70",
          1705 => x"de",
          1706 => x"25",
          1707 => x"18",
          1708 => x"81",
          1709 => x"75",
          1710 => x"80",
          1711 => x"98",
          1712 => x"33",
          1713 => x"98",
          1714 => x"dc",
          1715 => x"5d",
          1716 => x"38",
          1717 => x"39",
          1718 => x"81",
          1719 => x"70",
          1720 => x"57",
          1721 => x"75",
          1722 => x"80",
          1723 => x"57",
          1724 => x"d8",
          1725 => x"78",
          1726 => x"2e",
          1727 => x"57",
          1728 => x"e7",
          1729 => x"57",
          1730 => x"c8",
          1731 => x"7e",
          1732 => x"95",
          1733 => x"83",
          1734 => x"83",
          1735 => x"0b",
          1736 => x"d1",
          1737 => x"33",
          1738 => x"84",
          1739 => x"b6",
          1740 => x"05",
          1741 => x"eb",
          1742 => x"ff",
          1743 => x"55",
          1744 => x"d5",
          1745 => x"84",
          1746 => x"52",
          1747 => x"39",
          1748 => x"10",
          1749 => x"57",
          1750 => x"d1",
          1751 => x"cc",
          1752 => x"74",
          1753 => x"08",
          1754 => x"84",
          1755 => x"b5",
          1756 => x"88",
          1757 => x"d0",
          1758 => x"d0",
          1759 => x"cc",
          1760 => x"75",
          1761 => x"7c",
          1762 => x"75",
          1763 => x"f3",
          1764 => x"75",
          1765 => x"80",
          1766 => x"b7",
          1767 => x"d1",
          1768 => x"ff",
          1769 => x"51",
          1770 => x"33",
          1771 => x"80",
          1772 => x"08",
          1773 => x"84",
          1774 => x"b3",
          1775 => x"88",
          1776 => x"d0",
          1777 => x"d0",
          1778 => x"39",
          1779 => x"06",
          1780 => x"75",
          1781 => x"f0",
          1782 => x"d1",
          1783 => x"55",
          1784 => x"33",
          1785 => x"33",
          1786 => x"83",
          1787 => x"15",
          1788 => x"16",
          1789 => x"3f",
          1790 => x"06",
          1791 => x"77",
          1792 => x"39",
          1793 => x"33",
          1794 => x"38",
          1795 => x"34",
          1796 => x"81",
          1797 => x"24",
          1798 => x"52",
          1799 => x"d1",
          1800 => x"2c",
          1801 => x"41",
          1802 => x"d5",
          1803 => x"91",
          1804 => x"80",
          1805 => x"cc",
          1806 => x"f8",
          1807 => x"88",
          1808 => x"80",
          1809 => x"98",
          1810 => x"5a",
          1811 => x"bb",
          1812 => x"78",
          1813 => x"33",
          1814 => x"80",
          1815 => x"98",
          1816 => x"55",
          1817 => x"16",
          1818 => x"d5",
          1819 => x"b1",
          1820 => x"81",
          1821 => x"d1",
          1822 => x"24",
          1823 => x"d1",
          1824 => x"d3",
          1825 => x"51",
          1826 => x"33",
          1827 => x"34",
          1828 => x"84",
          1829 => x"7f",
          1830 => x"51",
          1831 => x"52",
          1832 => x"8c",
          1833 => x"cf",
          1834 => x"80",
          1835 => x"33",
          1836 => x"70",
          1837 => x"38",
          1838 => x"f3",
          1839 => x"5b",
          1840 => x"08",
          1841 => x"10",
          1842 => x"57",
          1843 => x"f3",
          1844 => x"38",
          1845 => x"2e",
          1846 => x"d0",
          1847 => x"7b",
          1848 => x"04",
          1849 => x"2e",
          1850 => x"88",
          1851 => x"f0",
          1852 => x"3f",
          1853 => x"ff",
          1854 => x"ff",
          1855 => x"75",
          1856 => x"83",
          1857 => x"80",
          1858 => x"84",
          1859 => x"7c",
          1860 => x"d1",
          1861 => x"38",
          1862 => x"ff",
          1863 => x"52",
          1864 => x"d5",
          1865 => x"a1",
          1866 => x"5d",
          1867 => x"ff",
          1868 => x"b8",
          1869 => x"84",
          1870 => x"cc",
          1871 => x"3d",
          1872 => x"81",
          1873 => x"f4",
          1874 => x"05",
          1875 => x"16",
          1876 => x"d5",
          1877 => x"c1",
          1878 => x"2b",
          1879 => x"5a",
          1880 => x"ef",
          1881 => x"51",
          1882 => x"33",
          1883 => x"d1",
          1884 => x"7a",
          1885 => x"08",
          1886 => x"74",
          1887 => x"05",
          1888 => x"5b",
          1889 => x"38",
          1890 => x"ff",
          1891 => x"29",
          1892 => x"84",
          1893 => x"75",
          1894 => x"7b",
          1895 => x"84",
          1896 => x"ff",
          1897 => x"29",
          1898 => x"84",
          1899 => x"61",
          1900 => x"81",
          1901 => x"08",
          1902 => x"3f",
          1903 => x"0a",
          1904 => x"33",
          1905 => x"a7",
          1906 => x"33",
          1907 => x"60",
          1908 => x"33",
          1909 => x"98",
          1910 => x"76",
          1911 => x"33",
          1912 => x"29",
          1913 => x"84",
          1914 => x"78",
          1915 => x"84",
          1916 => x"7c",
          1917 => x"84",
          1918 => x"8b",
          1919 => x"cc",
          1920 => x"70",
          1921 => x"05",
          1922 => x"44",
          1923 => x"ef",
          1924 => x"78",
          1925 => x"7a",
          1926 => x"08",
          1927 => x"75",
          1928 => x"05",
          1929 => x"57",
          1930 => x"38",
          1931 => x"ff",
          1932 => x"29",
          1933 => x"84",
          1934 => x"76",
          1935 => x"83",
          1936 => x"f4",
          1937 => x"3f",
          1938 => x"34",
          1939 => x"81",
          1940 => x"ad",
          1941 => x"d1",
          1942 => x"f4",
          1943 => x"88",
          1944 => x"f0",
          1945 => x"3f",
          1946 => x"ff",
          1947 => x"ff",
          1948 => x"7a",
          1949 => x"51",
          1950 => x"08",
          1951 => x"08",
          1952 => x"34",
          1953 => x"84",
          1954 => x"33",
          1955 => x"81",
          1956 => x"70",
          1957 => x"57",
          1958 => x"d1",
          1959 => x"2c",
          1960 => x"58",
          1961 => x"e4",
          1962 => x"ee",
          1963 => x"56",
          1964 => x"16",
          1965 => x"f0",
          1966 => x"83",
          1967 => x"ee",
          1968 => x"3f",
          1969 => x"cd",
          1970 => x"93",
          1971 => x"39",
          1972 => x"77",
          1973 => x"75",
          1974 => x"39",
          1975 => x"ba",
          1976 => x"ba",
          1977 => x"53",
          1978 => x"3f",
          1979 => x"d1",
          1980 => x"2e",
          1981 => x"52",
          1982 => x"d5",
          1983 => x"f1",
          1984 => x"51",
          1985 => x"33",
          1986 => x"34",
          1987 => x"80",
          1988 => x"34",
          1989 => x"84",
          1990 => x"75",
          1991 => x"8c",
          1992 => x"8c",
          1993 => x"75",
          1994 => x"81",
          1995 => x"cc",
          1996 => x"5e",
          1997 => x"84",
          1998 => x"a5",
          1999 => x"a0",
          2000 => x"f0",
          2001 => x"3f",
          2002 => x"76",
          2003 => x"06",
          2004 => x"83",
          2005 => x"cc",
          2006 => x"06",
          2007 => x"ff",
          2008 => x"ff",
          2009 => x"d0",
          2010 => x"2e",
          2011 => x"52",
          2012 => x"d5",
          2013 => x"81",
          2014 => x"51",
          2015 => x"33",
          2016 => x"34",
          2017 => x"74",
          2018 => x"fc",
          2019 => x"83",
          2020 => x"52",
          2021 => x"ba",
          2022 => x"33",
          2023 => x"70",
          2024 => x"f4",
          2025 => x"51",
          2026 => x"33",
          2027 => x"56",
          2028 => x"83",
          2029 => x"3d",
          2030 => x"52",
          2031 => x"f3",
          2032 => x"d7",
          2033 => x"e0",
          2034 => x"34",
          2035 => x"84",
          2036 => x"93",
          2037 => x"51",
          2038 => x"08",
          2039 => x"96",
          2040 => x"53",
          2041 => x"c1",
          2042 => x"ba",
          2043 => x"e9",
          2044 => x"ff",
          2045 => x"56",
          2046 => x"80",
          2047 => x"05",
          2048 => x"75",
          2049 => x"70",
          2050 => x"08",
          2051 => x"38",
          2052 => x"f3",
          2053 => x"55",
          2054 => x"08",
          2055 => x"10",
          2056 => x"57",
          2057 => x"70",
          2058 => x"27",
          2059 => x"09",
          2060 => x"ed",
          2061 => x"52",
          2062 => x"f3",
          2063 => x"06",
          2064 => x"38",
          2065 => x"bd",
          2066 => x"83",
          2067 => x"fc",
          2068 => x"70",
          2069 => x"3f",
          2070 => x"f3",
          2071 => x"a4",
          2072 => x"80",
          2073 => x"76",
          2074 => x"75",
          2075 => x"83",
          2076 => x"77",
          2077 => x"3d",
          2078 => x"84",
          2079 => x"72",
          2080 => x"2e",
          2081 => x"9e",
          2082 => x"87",
          2083 => x"80",
          2084 => x"58",
          2085 => x"f9",
          2086 => x"75",
          2087 => x"33",
          2088 => x"71",
          2089 => x"56",
          2090 => x"38",
          2091 => x"74",
          2092 => x"74",
          2093 => x"38",
          2094 => x"17",
          2095 => x"0b",
          2096 => x"81",
          2097 => x"ee",
          2098 => x"a0",
          2099 => x"10",
          2100 => x"90",
          2101 => x"40",
          2102 => x"b8",
          2103 => x"b7",
          2104 => x"f9",
          2105 => x"70",
          2106 => x"57",
          2107 => x"72",
          2108 => x"ff",
          2109 => x"ff",
          2110 => x"81",
          2111 => x"42",
          2112 => x"8f",
          2113 => x"31",
          2114 => x"76",
          2115 => x"9c",
          2116 => x"26",
          2117 => x"05",
          2118 => x"70",
          2119 => x"a3",
          2120 => x"70",
          2121 => x"06",
          2122 => x"06",
          2123 => x"5d",
          2124 => x"74",
          2125 => x"ff",
          2126 => x"29",
          2127 => x"fd",
          2128 => x"34",
          2129 => x"f9",
          2130 => x"2b",
          2131 => x"7a",
          2132 => x"26",
          2133 => x"fc",
          2134 => x"81",
          2135 => x"f9",
          2136 => x"a3",
          2137 => x"56",
          2138 => x"84",
          2139 => x"84",
          2140 => x"83",
          2141 => x"06",
          2142 => x"41",
          2143 => x"73",
          2144 => x"70",
          2145 => x"ff",
          2146 => x"29",
          2147 => x"ff",
          2148 => x"5c",
          2149 => x"77",
          2150 => x"79",
          2151 => x"38",
          2152 => x"38",
          2153 => x"29",
          2154 => x"86",
          2155 => x"34",
          2156 => x"98",
          2157 => x"86",
          2158 => x"80",
          2159 => x"ee",
          2160 => x"87",
          2161 => x"34",
          2162 => x"87",
          2163 => x"81",
          2164 => x"77",
          2165 => x"34",
          2166 => x"c0",
          2167 => x"90",
          2168 => x"07",
          2169 => x"34",
          2170 => x"53",
          2171 => x"b8",
          2172 => x"0c",
          2173 => x"33",
          2174 => x"0d",
          2175 => x"b3",
          2176 => x"59",
          2177 => x"da",
          2178 => x"bd",
          2179 => x"29",
          2180 => x"f9",
          2181 => x"7c",
          2182 => x"83",
          2183 => x"72",
          2184 => x"ba",
          2185 => x"ba",
          2186 => x"70",
          2187 => x"55",
          2188 => x"38",
          2189 => x"34",
          2190 => x"ff",
          2191 => x"57",
          2192 => x"b8",
          2193 => x"80",
          2194 => x"84",
          2195 => x"e0",
          2196 => x"70",
          2197 => x"05",
          2198 => x"fd",
          2199 => x"26",
          2200 => x"98",
          2201 => x"e0",
          2202 => x"55",
          2203 => x"27",
          2204 => x"05",
          2205 => x"57",
          2206 => x"ff",
          2207 => x"fd",
          2208 => x"b8",
          2209 => x"57",
          2210 => x"87",
          2211 => x"75",
          2212 => x"5c",
          2213 => x"38",
          2214 => x"14",
          2215 => x"78",
          2216 => x"81",
          2217 => x"59",
          2218 => x"84",
          2219 => x"56",
          2220 => x"38",
          2221 => x"8b",
          2222 => x"34",
          2223 => x"ff",
          2224 => x"57",
          2225 => x"80",
          2226 => x"06",
          2227 => x"53",
          2228 => x"c8",
          2229 => x"b8",
          2230 => x"29",
          2231 => x"27",
          2232 => x"84",
          2233 => x"56",
          2234 => x"75",
          2235 => x"13",
          2236 => x"a0",
          2237 => x"70",
          2238 => x"72",
          2239 => x"84",
          2240 => x"39",
          2241 => x"b8",
          2242 => x"ff",
          2243 => x"0d",
          2244 => x"53",
          2245 => x"10",
          2246 => x"08",
          2247 => x"71",
          2248 => x"34",
          2249 => x"3d",
          2250 => x"34",
          2251 => x"06",
          2252 => x"ff",
          2253 => x"80",
          2254 => x"0d",
          2255 => x"31",
          2256 => x"54",
          2257 => x"34",
          2258 => x"05",
          2259 => x"56",
          2260 => x"53",
          2261 => x"84",
          2262 => x"83",
          2263 => x"09",
          2264 => x"53",
          2265 => x"0b",
          2266 => x"04",
          2267 => x"b8",
          2268 => x"70",
          2269 => x"83",
          2270 => x"8c",
          2271 => x"83",
          2272 => x"84",
          2273 => x"71",
          2274 => x"51",
          2275 => x"39",
          2276 => x"51",
          2277 => x"10",
          2278 => x"04",
          2279 => x"06",
          2280 => x"72",
          2281 => x"71",
          2282 => x"38",
          2283 => x"80",
          2284 => x"0d",
          2285 => x"06",
          2286 => x"34",
          2287 => x"3d",
          2288 => x"f0",
          2289 => x"e8",
          2290 => x"06",
          2291 => x"34",
          2292 => x"b8",
          2293 => x"83",
          2294 => x"81",
          2295 => x"f9",
          2296 => x"b8",
          2297 => x"b8",
          2298 => x"33",
          2299 => x"83",
          2300 => x"f9",
          2301 => x"51",
          2302 => x"39",
          2303 => x"81",
          2304 => x"fe",
          2305 => x"f8",
          2306 => x"fe",
          2307 => x"df",
          2308 => x"f9",
          2309 => x"b8",
          2310 => x"70",
          2311 => x"83",
          2312 => x"e0",
          2313 => x"fe",
          2314 => x"cf",
          2315 => x"f9",
          2316 => x"b8",
          2317 => x"70",
          2318 => x"83",
          2319 => x"70",
          2320 => x"83",
          2321 => x"07",
          2322 => x"e0",
          2323 => x"33",
          2324 => x"83",
          2325 => x"83",
          2326 => x"43",
          2327 => x"2e",
          2328 => x"38",
          2329 => x"84",
          2330 => x"84",
          2331 => x"83",
          2332 => x"34",
          2333 => x"09",
          2334 => x"b8",
          2335 => x"34",
          2336 => x"0b",
          2337 => x"f9",
          2338 => x"33",
          2339 => x"b7",
          2340 => x"7a",
          2341 => x"db",
          2342 => x"0b",
          2343 => x"bc",
          2344 => x"83",
          2345 => x"80",
          2346 => x"84",
          2347 => x"bc",
          2348 => x"80",
          2349 => x"8f",
          2350 => x"84",
          2351 => x"54",
          2352 => x"51",
          2353 => x"b9",
          2354 => x"a5",
          2355 => x"70",
          2356 => x"ff",
          2357 => x"ff",
          2358 => x"59",
          2359 => x"ec",
          2360 => x"b8",
          2361 => x"34",
          2362 => x"f9",
          2363 => x"8f",
          2364 => x"82",
          2365 => x"81",
          2366 => x"83",
          2367 => x"ba",
          2368 => x"a3",
          2369 => x"e3",
          2370 => x"59",
          2371 => x"3f",
          2372 => x"a6",
          2373 => x"83",
          2374 => x"81",
          2375 => x"d8",
          2376 => x"05",
          2377 => x"83",
          2378 => x"72",
          2379 => x"11",
          2380 => x"5c",
          2381 => x"ff",
          2382 => x"51",
          2383 => x"e9",
          2384 => x"75",
          2385 => x"2e",
          2386 => x"d5",
          2387 => x"bc",
          2388 => x"29",
          2389 => x"16",
          2390 => x"84",
          2391 => x"83",
          2392 => x"5a",
          2393 => x"18",
          2394 => x"29",
          2395 => x"87",
          2396 => x"80",
          2397 => x"ba",
          2398 => x"29",
          2399 => x"f9",
          2400 => x"81",
          2401 => x"73",
          2402 => x"81",
          2403 => x"17",
          2404 => x"b8",
          2405 => x"38",
          2406 => x"2e",
          2407 => x"8c",
          2408 => x"2e",
          2409 => x"38",
          2410 => x"c1",
          2411 => x"3f",
          2412 => x"be",
          2413 => x"84",
          2414 => x"89",
          2415 => x"80",
          2416 => x"3f",
          2417 => x"54",
          2418 => x"52",
          2419 => x"70",
          2420 => x"27",
          2421 => x"f9",
          2422 => x"83",
          2423 => x"ba",
          2424 => x"80",
          2425 => x"38",
          2426 => x"06",
          2427 => x"73",
          2428 => x"52",
          2429 => x"bd",
          2430 => x"05",
          2431 => x"72",
          2432 => x"80",
          2433 => x"81",
          2434 => x"80",
          2435 => x"86",
          2436 => x"05",
          2437 => x"75",
          2438 => x"2e",
          2439 => x"b5",
          2440 => x"78",
          2441 => x"2e",
          2442 => x"83",
          2443 => x"72",
          2444 => x"b8",
          2445 => x"17",
          2446 => x"bd",
          2447 => x"29",
          2448 => x"f9",
          2449 => x"60",
          2450 => x"f9",
          2451 => x"05",
          2452 => x"ff",
          2453 => x"bd",
          2454 => x"5d",
          2455 => x"98",
          2456 => x"ff",
          2457 => x"b8",
          2458 => x"86",
          2459 => x"f9",
          2460 => x"0c",
          2461 => x"84",
          2462 => x"38",
          2463 => x"80",
          2464 => x"84",
          2465 => x"83",
          2466 => x"72",
          2467 => x"b8",
          2468 => x"1d",
          2469 => x"bd",
          2470 => x"29",
          2471 => x"f9",
          2472 => x"76",
          2473 => x"b8",
          2474 => x"84",
          2475 => x"83",
          2476 => x"72",
          2477 => x"59",
          2478 => x"de",
          2479 => x"ff",
          2480 => x"38",
          2481 => x"84",
          2482 => x"78",
          2483 => x"24",
          2484 => x"81",
          2485 => x"f9",
          2486 => x"0c",
          2487 => x"82",
          2488 => x"26",
          2489 => x"81",
          2490 => x"34",
          2491 => x"81",
          2492 => x"90",
          2493 => x"0c",
          2494 => x"fd",
          2495 => x"0c",
          2496 => x"33",
          2497 => x"05",
          2498 => x"33",
          2499 => x"b8",
          2500 => x"f9",
          2501 => x"5f",
          2502 => x"34",
          2503 => x"19",
          2504 => x"a3",
          2505 => x"33",
          2506 => x"22",
          2507 => x"11",
          2508 => x"b8",
          2509 => x"81",
          2510 => x"81",
          2511 => x"f9",
          2512 => x"80",
          2513 => x"ff",
          2514 => x"29",
          2515 => x"f9",
          2516 => x"29",
          2517 => x"f8",
          2518 => x"75",
          2519 => x"ff",
          2520 => x"95",
          2521 => x"34",
          2522 => x"8c",
          2523 => x"80",
          2524 => x"84",
          2525 => x"88",
          2526 => x"9c",
          2527 => x"84",
          2528 => x"84",
          2529 => x"84",
          2530 => x"88",
          2531 => x"9c",
          2532 => x"09",
          2533 => x"bc",
          2534 => x"ff",
          2535 => x"ff",
          2536 => x"a0",
          2537 => x"40",
          2538 => x"ff",
          2539 => x"43",
          2540 => x"85",
          2541 => x"1a",
          2542 => x"76",
          2543 => x"06",
          2544 => x"06",
          2545 => x"84",
          2546 => x"1e",
          2547 => x"bd",
          2548 => x"29",
          2549 => x"83",
          2550 => x"33",
          2551 => x"83",
          2552 => x"1a",
          2553 => x"ff",
          2554 => x"bd",
          2555 => x"5a",
          2556 => x"84",
          2557 => x"81",
          2558 => x"95",
          2559 => x"79",
          2560 => x"83",
          2561 => x"70",
          2562 => x"fd",
          2563 => x"38",
          2564 => x"bf",
          2565 => x"33",
          2566 => x"19",
          2567 => x"75",
          2568 => x"77",
          2569 => x"34",
          2570 => x"80",
          2571 => x"0d",
          2572 => x"80",
          2573 => x"bd",
          2574 => x"29",
          2575 => x"f9",
          2576 => x"05",
          2577 => x"92",
          2578 => x"5b",
          2579 => x"5c",
          2580 => x"06",
          2581 => x"05",
          2582 => x"87",
          2583 => x"80",
          2584 => x"ba",
          2585 => x"5e",
          2586 => x"34",
          2587 => x"1e",
          2588 => x"a3",
          2589 => x"33",
          2590 => x"22",
          2591 => x"11",
          2592 => x"b8",
          2593 => x"81",
          2594 => x"7e",
          2595 => x"81",
          2596 => x"19",
          2597 => x"1c",
          2598 => x"83",
          2599 => x"33",
          2600 => x"33",
          2601 => x"06",
          2602 => x"05",
          2603 => x"b8",
          2604 => x"34",
          2605 => x"33",
          2606 => x"12",
          2607 => x"f9",
          2608 => x"76",
          2609 => x"b8",
          2610 => x"84",
          2611 => x"83",
          2612 => x"72",
          2613 => x"59",
          2614 => x"18",
          2615 => x"06",
          2616 => x"38",
          2617 => x"39",
          2618 => x"0b",
          2619 => x"04",
          2620 => x"b8",
          2621 => x"bd",
          2622 => x"05",
          2623 => x"b9",
          2624 => x"0c",
          2625 => x"17",
          2626 => x"7c",
          2627 => x"80",
          2628 => x"5b",
          2629 => x"90",
          2630 => x"05",
          2631 => x"8c",
          2632 => x"b9",
          2633 => x"84",
          2634 => x"06",
          2635 => x"84",
          2636 => x"83",
          2637 => x"88",
          2638 => x"33",
          2639 => x"33",
          2640 => x"b8",
          2641 => x"f9",
          2642 => x"5d",
          2643 => x"87",
          2644 => x"80",
          2645 => x"ba",
          2646 => x"5b",
          2647 => x"83",
          2648 => x"41",
          2649 => x"a3",
          2650 => x"33",
          2651 => x"22",
          2652 => x"11",
          2653 => x"b8",
          2654 => x"1c",
          2655 => x"7b",
          2656 => x"33",
          2657 => x"56",
          2658 => x"84",
          2659 => x"40",
          2660 => x"b8",
          2661 => x"78",
          2662 => x"0b",
          2663 => x"04",
          2664 => x"34",
          2665 => x"34",
          2666 => x"f9",
          2667 => x"bc",
          2668 => x"bd",
          2669 => x"bb",
          2670 => x"39",
          2671 => x"2e",
          2672 => x"5d",
          2673 => x"85",
          2674 => x"55",
          2675 => x"9b",
          2676 => x"70",
          2677 => x"51",
          2678 => x"08",
          2679 => x"57",
          2680 => x"cd",
          2681 => x"fe",
          2682 => x"0b",
          2683 => x"81",
          2684 => x"ad",
          2685 => x"81",
          2686 => x"8a",
          2687 => x"ec",
          2688 => x"8d",
          2689 => x"38",
          2690 => x"33",
          2691 => x"2c",
          2692 => x"75",
          2693 => x"84",
          2694 => x"8e",
          2695 => x"05",
          2696 => x"33",
          2697 => x"c5",
          2698 => x"bd",
          2699 => x"83",
          2700 => x"5d",
          2701 => x"ff",
          2702 => x"fd",
          2703 => x"34",
          2704 => x"33",
          2705 => x"fd",
          2706 => x"f9",
          2707 => x"8d",
          2708 => x"38",
          2709 => x"33",
          2710 => x"2c",
          2711 => x"75",
          2712 => x"84",
          2713 => x"fc",
          2714 => x"60",
          2715 => x"38",
          2716 => x"33",
          2717 => x"12",
          2718 => x"ba",
          2719 => x"29",
          2720 => x"f8",
          2721 => x"42",
          2722 => x"2e",
          2723 => x"91",
          2724 => x"33",
          2725 => x"84",
          2726 => x"09",
          2727 => x"83",
          2728 => x"b9",
          2729 => x"be",
          2730 => x"bd",
          2731 => x"33",
          2732 => x"25",
          2733 => x"bd",
          2734 => x"33",
          2735 => x"84",
          2736 => x"42",
          2737 => x"11",
          2738 => x"38",
          2739 => x"fa",
          2740 => x"e8",
          2741 => x"33",
          2742 => x"38",
          2743 => x"22",
          2744 => x"e8",
          2745 => x"06",
          2746 => x"da",
          2747 => x"5f",
          2748 => x"b9",
          2749 => x"38",
          2750 => x"06",
          2751 => x"84",
          2752 => x"8e",
          2753 => x"05",
          2754 => x"33",
          2755 => x"b7",
          2756 => x"11",
          2757 => x"77",
          2758 => x"83",
          2759 => x"ff",
          2760 => x"38",
          2761 => x"84",
          2762 => x"7a",
          2763 => x"75",
          2764 => x"84",
          2765 => x"8a",
          2766 => x"b7",
          2767 => x"f9",
          2768 => x"b8",
          2769 => x"f9",
          2770 => x"a3",
          2771 => x"5f",
          2772 => x"ff",
          2773 => x"52",
          2774 => x"84",
          2775 => x"70",
          2776 => x"8e",
          2777 => x"76",
          2778 => x"56",
          2779 => x"ff",
          2780 => x"60",
          2781 => x"33",
          2782 => x"ff",
          2783 => x"7e",
          2784 => x"57",
          2785 => x"38",
          2786 => x"ff",
          2787 => x"79",
          2788 => x"a3",
          2789 => x"81",
          2790 => x"58",
          2791 => x"38",
          2792 => x"17",
          2793 => x"7b",
          2794 => x"81",
          2795 => x"5e",
          2796 => x"84",
          2797 => x"43",
          2798 => x"9d",
          2799 => x"b8",
          2800 => x"5d",
          2801 => x"7c",
          2802 => x"84",
          2803 => x"71",
          2804 => x"7f",
          2805 => x"39",
          2806 => x"2e",
          2807 => x"e1",
          2808 => x"39",
          2809 => x"11",
          2810 => x"58",
          2811 => x"e0",
          2812 => x"06",
          2813 => x"58",
          2814 => x"33",
          2815 => x"81",
          2816 => x"7a",
          2817 => x"ff",
          2818 => x"38",
          2819 => x"57",
          2820 => x"1b",
          2821 => x"a0",
          2822 => x"a3",
          2823 => x"51",
          2824 => x"06",
          2825 => x"b8",
          2826 => x"07",
          2827 => x"7f",
          2828 => x"9e",
          2829 => x"0c",
          2830 => x"79",
          2831 => x"33",
          2832 => x"81",
          2833 => x"f9",
          2834 => x"59",
          2835 => x"38",
          2836 => x"62",
          2837 => x"57",
          2838 => x"f9",
          2839 => x"5a",
          2840 => x"78",
          2841 => x"57",
          2842 => x"0b",
          2843 => x"81",
          2844 => x"77",
          2845 => x"1f",
          2846 => x"8a",
          2847 => x"f0",
          2848 => x"71",
          2849 => x"80",
          2850 => x"80",
          2851 => x"18",
          2852 => x"b6",
          2853 => x"84",
          2854 => x"f9",
          2855 => x"f9",
          2856 => x"5c",
          2857 => x"b8",
          2858 => x"b8",
          2859 => x"59",
          2860 => x"33",
          2861 => x"83",
          2862 => x"b8",
          2863 => x"75",
          2864 => x"f9",
          2865 => x"56",
          2866 => x"83",
          2867 => x"07",
          2868 => x"b1",
          2869 => x"34",
          2870 => x"56",
          2871 => x"81",
          2872 => x"34",
          2873 => x"81",
          2874 => x"f9",
          2875 => x"b8",
          2876 => x"56",
          2877 => x"39",
          2878 => x"80",
          2879 => x"34",
          2880 => x"81",
          2881 => x"f9",
          2882 => x"b8",
          2883 => x"75",
          2884 => x"83",
          2885 => x"07",
          2886 => x"a1",
          2887 => x"06",
          2888 => x"34",
          2889 => x"81",
          2890 => x"34",
          2891 => x"80",
          2892 => x"34",
          2893 => x"80",
          2894 => x"34",
          2895 => x"81",
          2896 => x"83",
          2897 => x"f9",
          2898 => x"56",
          2899 => x"39",
          2900 => x"52",
          2901 => x"39",
          2902 => x"34",
          2903 => x"34",
          2904 => x"f9",
          2905 => x"0c",
          2906 => x"8f",
          2907 => x"9c",
          2908 => x"34",
          2909 => x"06",
          2910 => x"84",
          2911 => x"53",
          2912 => x"84",
          2913 => x"8c",
          2914 => x"84",
          2915 => x"8c",
          2916 => x"f9",
          2917 => x"8d",
          2918 => x"b9",
          2919 => x"5d",
          2920 => x"e0",
          2921 => x"34",
          2922 => x"34",
          2923 => x"83",
          2924 => x"58",
          2925 => x"0b",
          2926 => x"51",
          2927 => x"51",
          2928 => x"83",
          2929 => x"70",
          2930 => x"f2",
          2931 => x"39",
          2932 => x"27",
          2933 => x"34",
          2934 => x"ff",
          2935 => x"06",
          2936 => x"f9",
          2937 => x"33",
          2938 => x"25",
          2939 => x"39",
          2940 => x"06",
          2941 => x"38",
          2942 => x"33",
          2943 => x"33",
          2944 => x"80",
          2945 => x"71",
          2946 => x"06",
          2947 => x"42",
          2948 => x"38",
          2949 => x"5c",
          2950 => x"84",
          2951 => x"83",
          2952 => x"f9",
          2953 => x"11",
          2954 => x"38",
          2955 => x"27",
          2956 => x"83",
          2957 => x"83",
          2958 => x"76",
          2959 => x"81",
          2960 => x"29",
          2961 => x"a0",
          2962 => x"81",
          2963 => x"71",
          2964 => x"7e",
          2965 => x"1a",
          2966 => x"b8",
          2967 => x"5d",
          2968 => x"7d",
          2969 => x"84",
          2970 => x"71",
          2971 => x"77",
          2972 => x"17",
          2973 => x"7b",
          2974 => x"81",
          2975 => x"5f",
          2976 => x"84",
          2977 => x"59",
          2978 => x"99",
          2979 => x"17",
          2980 => x"7b",
          2981 => x"80",
          2982 => x"ff",
          2983 => x"39",
          2984 => x"33",
          2985 => x"42",
          2986 => x"5a",
          2987 => x"ff",
          2988 => x"27",
          2989 => x"bc",
          2990 => x"ff",
          2991 => x"78",
          2992 => x"83",
          2993 => x"f9",
          2994 => x"33",
          2995 => x"25",
          2996 => x"39",
          2997 => x"c0",
          2998 => x"ff",
          2999 => x"5d",
          3000 => x"06",
          3001 => x"1d",
          3002 => x"93",
          3003 => x"ba",
          3004 => x"56",
          3005 => x"39",
          3006 => x"f5",
          3007 => x"58",
          3008 => x"81",
          3009 => x"ec",
          3010 => x"34",
          3011 => x"05",
          3012 => x"f4",
          3013 => x"83",
          3014 => x"0b",
          3015 => x"7e",
          3016 => x"80",
          3017 => x"39",
          3018 => x"a7",
          3019 => x"84",
          3020 => x"0b",
          3021 => x"fd",
          3022 => x"b8",
          3023 => x"90",
          3024 => x"0b",
          3025 => x"04",
          3026 => x"80",
          3027 => x"0d",
          3028 => x"33",
          3029 => x"70",
          3030 => x"33",
          3031 => x"80",
          3032 => x"f8",
          3033 => x"8c",
          3034 => x"ec",
          3035 => x"91",
          3036 => x"07",
          3037 => x"5e",
          3038 => x"59",
          3039 => x"06",
          3040 => x"70",
          3041 => x"5c",
          3042 => x"84",
          3043 => x"83",
          3044 => x"87",
          3045 => x"22",
          3046 => x"70",
          3047 => x"33",
          3048 => x"83",
          3049 => x"ee",
          3050 => x"98",
          3051 => x"56",
          3052 => x"80",
          3053 => x"15",
          3054 => x"55",
          3055 => x"80",
          3056 => x"81",
          3057 => x"58",
          3058 => x"38",
          3059 => x"74",
          3060 => x"ff",
          3061 => x"cd",
          3062 => x"83",
          3063 => x"15",
          3064 => x"55",
          3065 => x"83",
          3066 => x"80",
          3067 => x"e4",
          3068 => x"2a",
          3069 => x"58",
          3070 => x"0b",
          3071 => x"06",
          3072 => x"81",
          3073 => x"83",
          3074 => x"83",
          3075 => x"33",
          3076 => x"5e",
          3077 => x"33",
          3078 => x"83",
          3079 => x"2e",
          3080 => x"33",
          3081 => x"83",
          3082 => x"ec",
          3083 => x"81",
          3084 => x"16",
          3085 => x"38",
          3086 => x"ff",
          3087 => x"16",
          3088 => x"38",
          3089 => x"87",
          3090 => x"73",
          3091 => x"c0",
          3092 => x"58",
          3093 => x"54",
          3094 => x"83",
          3095 => x"34",
          3096 => x"82",
          3097 => x"b4",
          3098 => x"94",
          3099 => x"83",
          3100 => x"5e",
          3101 => x"80",
          3102 => x"72",
          3103 => x"83",
          3104 => x"08",
          3105 => x"06",
          3106 => x"f9",
          3107 => x"14",
          3108 => x"a5",
          3109 => x"80",
          3110 => x"83",
          3111 => x"f0",
          3112 => x"e0",
          3113 => x"7c",
          3114 => x"09",
          3115 => x"2e",
          3116 => x"d7",
          3117 => x"77",
          3118 => x"80",
          3119 => x"38",
          3120 => x"10",
          3121 => x"98",
          3122 => x"73",
          3123 => x"79",
          3124 => x"05",
          3125 => x"56",
          3126 => x"83",
          3127 => x"80",
          3128 => x"79",
          3129 => x"82",
          3130 => x"fa",
          3131 => x"33",
          3132 => x"38",
          3133 => x"25",
          3134 => x"38",
          3135 => x"cc",
          3136 => x"80",
          3137 => x"98",
          3138 => x"2e",
          3139 => x"ff",
          3140 => x"38",
          3141 => x"2e",
          3142 => x"55",
          3143 => x"06",
          3144 => x"84",
          3145 => x"be",
          3146 => x"39",
          3147 => x"f7",
          3148 => x"83",
          3149 => x"80",
          3150 => x"0b",
          3151 => x"83",
          3152 => x"74",
          3153 => x"2e",
          3154 => x"33",
          3155 => x"77",
          3156 => x"09",
          3157 => x"e0",
          3158 => x"9c",
          3159 => x"e8",
          3160 => x"f7",
          3161 => x"fb",
          3162 => x"15",
          3163 => x"e5",
          3164 => x"fa",
          3165 => x"80",
          3166 => x"ec",
          3167 => x"f7",
          3168 => x"5d",
          3169 => x"39",
          3170 => x"cb",
          3171 => x"ce",
          3172 => x"fc",
          3173 => x"34",
          3174 => x"0b",
          3175 => x"83",
          3176 => x"34",
          3177 => x"84",
          3178 => x"38",
          3179 => x"ff",
          3180 => x"f7",
          3181 => x"84",
          3182 => x"39",
          3183 => x"06",
          3184 => x"27",
          3185 => x"ba",
          3186 => x"55",
          3187 => x"54",
          3188 => x"80",
          3189 => x"05",
          3190 => x"53",
          3191 => x"f6",
          3192 => x"ba",
          3193 => x"72",
          3194 => x"52",
          3195 => x"3f",
          3196 => x"f7",
          3197 => x"3d",
          3198 => x"3d",
          3199 => x"83",
          3200 => x"05",
          3201 => x"08",
          3202 => x"83",
          3203 => x"81",
          3204 => x"e8",
          3205 => x"f4",
          3206 => x"54",
          3207 => x"c0",
          3208 => x"f6",
          3209 => x"9c",
          3210 => x"38",
          3211 => x"c0",
          3212 => x"74",
          3213 => x"ff",
          3214 => x"9c",
          3215 => x"c0",
          3216 => x"9c",
          3217 => x"81",
          3218 => x"53",
          3219 => x"81",
          3220 => x"a4",
          3221 => x"a4",
          3222 => x"38",
          3223 => x"ff",
          3224 => x"ff",
          3225 => x"0c",
          3226 => x"81",
          3227 => x"81",
          3228 => x"d7",
          3229 => x"89",
          3230 => x"02",
          3231 => x"80",
          3232 => x"2b",
          3233 => x"98",
          3234 => x"83",
          3235 => x"84",
          3236 => x"85",
          3237 => x"f4",
          3238 => x"83",
          3239 => x"34",
          3240 => x"57",
          3241 => x"86",
          3242 => x"9c",
          3243 => x"ce",
          3244 => x"08",
          3245 => x"71",
          3246 => x"87",
          3247 => x"74",
          3248 => x"db",
          3249 => x"ff",
          3250 => x"72",
          3251 => x"87",
          3252 => x"05",
          3253 => x"87",
          3254 => x"2e",
          3255 => x"98",
          3256 => x"87",
          3257 => x"87",
          3258 => x"71",
          3259 => x"72",
          3260 => x"2e",
          3261 => x"53",
          3262 => x"81",
          3263 => x"c6",
          3264 => x"53",
          3265 => x"81",
          3266 => x"54",
          3267 => x"84",
          3268 => x"81",
          3269 => x"d4",
          3270 => x"89",
          3271 => x"ff",
          3272 => x"ff",
          3273 => x"7a",
          3274 => x"57",
          3275 => x"88",
          3276 => x"7a",
          3277 => x"76",
          3278 => x"71",
          3279 => x"72",
          3280 => x"7b",
          3281 => x"84",
          3282 => x"74",
          3283 => x"53",
          3284 => x"73",
          3285 => x"08",
          3286 => x"98",
          3287 => x"0b",
          3288 => x"0b",
          3289 => x"80",
          3290 => x"83",
          3291 => x"05",
          3292 => x"87",
          3293 => x"2e",
          3294 => x"98",
          3295 => x"87",
          3296 => x"87",
          3297 => x"71",
          3298 => x"72",
          3299 => x"98",
          3300 => x"87",
          3301 => x"98",
          3302 => x"38",
          3303 => x"08",
          3304 => x"72",
          3305 => x"98",
          3306 => x"27",
          3307 => x"a2",
          3308 => x"81",
          3309 => x"75",
          3310 => x"a1",
          3311 => x"3d",
          3312 => x"06",
          3313 => x"81",
          3314 => x"e1",
          3315 => x"58",
          3316 => x"8c",
          3317 => x"0d",
          3318 => x"71",
          3319 => x"56",
          3320 => x"0b",
          3321 => x"98",
          3322 => x"80",
          3323 => x"9c",
          3324 => x"53",
          3325 => x"33",
          3326 => x"70",
          3327 => x"2e",
          3328 => x"51",
          3329 => x"38",
          3330 => x"38",
          3331 => x"90",
          3332 => x"52",
          3333 => x"72",
          3334 => x"c0",
          3335 => x"27",
          3336 => x"38",
          3337 => x"53",
          3338 => x"71",
          3339 => x"8a",
          3340 => x"fe",
          3341 => x"81",
          3342 => x"3d",
          3343 => x"f6",
          3344 => x"0d",
          3345 => x"83",
          3346 => x"83",
          3347 => x"33",
          3348 => x"77",
          3349 => x"98",
          3350 => x"41",
          3351 => x"57",
          3352 => x"72",
          3353 => x"71",
          3354 => x"05",
          3355 => x"2b",
          3356 => x"52",
          3357 => x"9e",
          3358 => x"71",
          3359 => x"05",
          3360 => x"74",
          3361 => x"54",
          3362 => x"08",
          3363 => x"33",
          3364 => x"5c",
          3365 => x"34",
          3366 => x"08",
          3367 => x"80",
          3368 => x"08",
          3369 => x"14",
          3370 => x"33",
          3371 => x"82",
          3372 => x"58",
          3373 => x"13",
          3374 => x"33",
          3375 => x"83",
          3376 => x"85",
          3377 => x"88",
          3378 => x"58",
          3379 => x"34",
          3380 => x"11",
          3381 => x"71",
          3382 => x"72",
          3383 => x"71",
          3384 => x"55",
          3385 => x"87",
          3386 => x"70",
          3387 => x"07",
          3388 => x"5a",
          3389 => x"81",
          3390 => x"17",
          3391 => x"2b",
          3392 => x"33",
          3393 => x"70",
          3394 => x"05",
          3395 => x"5c",
          3396 => x"34",
          3397 => x"08",
          3398 => x"71",
          3399 => x"05",
          3400 => x"2b",
          3401 => x"2a",
          3402 => x"52",
          3403 => x"84",
          3404 => x"33",
          3405 => x"83",
          3406 => x"12",
          3407 => x"07",
          3408 => x"53",
          3409 => x"33",
          3410 => x"82",
          3411 => x"59",
          3412 => x"34",
          3413 => x"33",
          3414 => x"83",
          3415 => x"83",
          3416 => x"88",
          3417 => x"52",
          3418 => x"15",
          3419 => x"0d",
          3420 => x"76",
          3421 => x"86",
          3422 => x"3d",
          3423 => x"b9",
          3424 => x"f8",
          3425 => x"84",
          3426 => x"84",
          3427 => x"81",
          3428 => x"08",
          3429 => x"85",
          3430 => x"76",
          3431 => x"34",
          3432 => x"22",
          3433 => x"83",
          3434 => x"51",
          3435 => x"89",
          3436 => x"10",
          3437 => x"f8",
          3438 => x"81",
          3439 => x"f7",
          3440 => x"51",
          3441 => x"83",
          3442 => x"06",
          3443 => x"84",
          3444 => x"12",
          3445 => x"59",
          3446 => x"75",
          3447 => x"10",
          3448 => x"71",
          3449 => x"06",
          3450 => x"70",
          3451 => x"52",
          3452 => x"2e",
          3453 => x"12",
          3454 => x"07",
          3455 => x"ff",
          3456 => x"56",
          3457 => x"33",
          3458 => x"70",
          3459 => x"56",
          3460 => x"81",
          3461 => x"8d",
          3462 => x"85",
          3463 => x"74",
          3464 => x"82",
          3465 => x"5c",
          3466 => x"81",
          3467 => x"76",
          3468 => x"34",
          3469 => x"08",
          3470 => x"71",
          3471 => x"ff",
          3472 => x"ff",
          3473 => x"57",
          3474 => x"72",
          3475 => x"34",
          3476 => x"74",
          3477 => x"fc",
          3478 => x"12",
          3479 => x"07",
          3480 => x"75",
          3481 => x"84",
          3482 => x"05",
          3483 => x"88",
          3484 => x"58",
          3485 => x"15",
          3486 => x"84",
          3487 => x"2b",
          3488 => x"5a",
          3489 => x"72",
          3490 => x"70",
          3491 => x"85",
          3492 => x"88",
          3493 => x"15",
          3494 => x"fc",
          3495 => x"ba",
          3496 => x"14",
          3497 => x"71",
          3498 => x"33",
          3499 => x"70",
          3500 => x"52",
          3501 => x"34",
          3502 => x"11",
          3503 => x"71",
          3504 => x"33",
          3505 => x"70",
          3506 => x"5b",
          3507 => x"87",
          3508 => x"70",
          3509 => x"07",
          3510 => x"59",
          3511 => x"81",
          3512 => x"84",
          3513 => x"0d",
          3514 => x"76",
          3515 => x"8a",
          3516 => x"3d",
          3517 => x"84",
          3518 => x"89",
          3519 => x"84",
          3520 => x"b9",
          3521 => x"52",
          3522 => x"3f",
          3523 => x"34",
          3524 => x"fc",
          3525 => x"0b",
          3526 => x"56",
          3527 => x"17",
          3528 => x"f8",
          3529 => x"70",
          3530 => x"58",
          3531 => x"73",
          3532 => x"70",
          3533 => x"05",
          3534 => x"34",
          3535 => x"77",
          3536 => x"39",
          3537 => x"80",
          3538 => x"41",
          3539 => x"80",
          3540 => x"88",
          3541 => x"8f",
          3542 => x"05",
          3543 => x"73",
          3544 => x"83",
          3545 => x"83",
          3546 => x"33",
          3547 => x"70",
          3548 => x"10",
          3549 => x"70",
          3550 => x"07",
          3551 => x"42",
          3552 => x"5c",
          3553 => x"7a",
          3554 => x"83",
          3555 => x"10",
          3556 => x"33",
          3557 => x"53",
          3558 => x"24",
          3559 => x"f6",
          3560 => x"87",
          3561 => x"38",
          3562 => x"be",
          3563 => x"92",
          3564 => x"12",
          3565 => x"07",
          3566 => x"71",
          3567 => x"43",
          3568 => x"60",
          3569 => x"11",
          3570 => x"71",
          3571 => x"33",
          3572 => x"83",
          3573 => x"85",
          3574 => x"88",
          3575 => x"58",
          3576 => x"34",
          3577 => x"08",
          3578 => x"33",
          3579 => x"74",
          3580 => x"71",
          3581 => x"42",
          3582 => x"86",
          3583 => x"b9",
          3584 => x"33",
          3585 => x"06",
          3586 => x"76",
          3587 => x"b9",
          3588 => x"83",
          3589 => x"2b",
          3590 => x"33",
          3591 => x"41",
          3592 => x"79",
          3593 => x"b9",
          3594 => x"12",
          3595 => x"07",
          3596 => x"33",
          3597 => x"41",
          3598 => x"79",
          3599 => x"84",
          3600 => x"33",
          3601 => x"66",
          3602 => x"52",
          3603 => x"fe",
          3604 => x"1e",
          3605 => x"83",
          3606 => x"62",
          3607 => x"84",
          3608 => x"84",
          3609 => x"a0",
          3610 => x"80",
          3611 => x"51",
          3612 => x"08",
          3613 => x"1f",
          3614 => x"84",
          3615 => x"84",
          3616 => x"34",
          3617 => x"fc",
          3618 => x"fe",
          3619 => x"06",
          3620 => x"78",
          3621 => x"84",
          3622 => x"84",
          3623 => x"56",
          3624 => x"15",
          3625 => x"fa",
          3626 => x"38",
          3627 => x"38",
          3628 => x"8c",
          3629 => x"0d",
          3630 => x"71",
          3631 => x"05",
          3632 => x"2b",
          3633 => x"2a",
          3634 => x"34",
          3635 => x"fc",
          3636 => x"75",
          3637 => x"84",
          3638 => x"81",
          3639 => x"83",
          3640 => x"64",
          3641 => x"4a",
          3642 => x"63",
          3643 => x"41",
          3644 => x"fc",
          3645 => x"81",
          3646 => x"05",
          3647 => x"54",
          3648 => x"83",
          3649 => x"39",
          3650 => x"70",
          3651 => x"83",
          3652 => x"10",
          3653 => x"33",
          3654 => x"53",
          3655 => x"73",
          3656 => x"39",
          3657 => x"7a",
          3658 => x"ff",
          3659 => x"38",
          3660 => x"84",
          3661 => x"b9",
          3662 => x"52",
          3663 => x"3f",
          3664 => x"34",
          3665 => x"fc",
          3666 => x"0b",
          3667 => x"58",
          3668 => x"19",
          3669 => x"f8",
          3670 => x"70",
          3671 => x"58",
          3672 => x"34",
          3673 => x"f8",
          3674 => x"fc",
          3675 => x"61",
          3676 => x"34",
          3677 => x"de",
          3678 => x"61",
          3679 => x"39",
          3680 => x"51",
          3681 => x"ba",
          3682 => x"1e",
          3683 => x"8b",
          3684 => x"86",
          3685 => x"2b",
          3686 => x"14",
          3687 => x"07",
          3688 => x"5b",
          3689 => x"64",
          3690 => x"34",
          3691 => x"11",
          3692 => x"71",
          3693 => x"33",
          3694 => x"70",
          3695 => x"59",
          3696 => x"7a",
          3697 => x"08",
          3698 => x"88",
          3699 => x"88",
          3700 => x"34",
          3701 => x"08",
          3702 => x"33",
          3703 => x"74",
          3704 => x"88",
          3705 => x"5e",
          3706 => x"34",
          3707 => x"08",
          3708 => x"71",
          3709 => x"05",
          3710 => x"88",
          3711 => x"40",
          3712 => x"18",
          3713 => x"fc",
          3714 => x"12",
          3715 => x"62",
          3716 => x"5d",
          3717 => x"95",
          3718 => x"05",
          3719 => x"fc",
          3720 => x"b9",
          3721 => x"f8",
          3722 => x"84",
          3723 => x"84",
          3724 => x"81",
          3725 => x"08",
          3726 => x"85",
          3727 => x"7f",
          3728 => x"34",
          3729 => x"22",
          3730 => x"83",
          3731 => x"43",
          3732 => x"89",
          3733 => x"10",
          3734 => x"f8",
          3735 => x"81",
          3736 => x"bd",
          3737 => x"19",
          3738 => x"71",
          3739 => x"33",
          3740 => x"70",
          3741 => x"55",
          3742 => x"85",
          3743 => x"1e",
          3744 => x"8b",
          3745 => x"86",
          3746 => x"2b",
          3747 => x"48",
          3748 => x"05",
          3749 => x"b9",
          3750 => x"33",
          3751 => x"06",
          3752 => x"75",
          3753 => x"b9",
          3754 => x"12",
          3755 => x"07",
          3756 => x"71",
          3757 => x"ff",
          3758 => x"48",
          3759 => x"41",
          3760 => x"34",
          3761 => x"33",
          3762 => x"83",
          3763 => x"12",
          3764 => x"ff",
          3765 => x"5e",
          3766 => x"76",
          3767 => x"ff",
          3768 => x"33",
          3769 => x"83",
          3770 => x"85",
          3771 => x"88",
          3772 => x"78",
          3773 => x"84",
          3774 => x"33",
          3775 => x"83",
          3776 => x"87",
          3777 => x"88",
          3778 => x"55",
          3779 => x"60",
          3780 => x"18",
          3781 => x"2b",
          3782 => x"2a",
          3783 => x"78",
          3784 => x"70",
          3785 => x"8b",
          3786 => x"70",
          3787 => x"07",
          3788 => x"77",
          3789 => x"5f",
          3790 => x"17",
          3791 => x"fc",
          3792 => x"33",
          3793 => x"74",
          3794 => x"88",
          3795 => x"88",
          3796 => x"5d",
          3797 => x"34",
          3798 => x"11",
          3799 => x"71",
          3800 => x"33",
          3801 => x"83",
          3802 => x"85",
          3803 => x"88",
          3804 => x"59",
          3805 => x"1d",
          3806 => x"fc",
          3807 => x"12",
          3808 => x"07",
          3809 => x"33",
          3810 => x"5f",
          3811 => x"77",
          3812 => x"84",
          3813 => x"12",
          3814 => x"ff",
          3815 => x"59",
          3816 => x"84",
          3817 => x"33",
          3818 => x"83",
          3819 => x"15",
          3820 => x"2a",
          3821 => x"55",
          3822 => x"84",
          3823 => x"81",
          3824 => x"2b",
          3825 => x"15",
          3826 => x"2a",
          3827 => x"55",
          3828 => x"34",
          3829 => x"11",
          3830 => x"07",
          3831 => x"42",
          3832 => x"51",
          3833 => x"08",
          3834 => x"70",
          3835 => x"f1",
          3836 => x"33",
          3837 => x"79",
          3838 => x"71",
          3839 => x"48",
          3840 => x"05",
          3841 => x"b9",
          3842 => x"85",
          3843 => x"2b",
          3844 => x"15",
          3845 => x"2a",
          3846 => x"56",
          3847 => x"87",
          3848 => x"70",
          3849 => x"07",
          3850 => x"5c",
          3851 => x"81",
          3852 => x"1f",
          3853 => x"2b",
          3854 => x"33",
          3855 => x"70",
          3856 => x"05",
          3857 => x"58",
          3858 => x"34",
          3859 => x"08",
          3860 => x"71",
          3861 => x"05",
          3862 => x"2b",
          3863 => x"2a",
          3864 => x"5b",
          3865 => x"77",
          3866 => x"39",
          3867 => x"84",
          3868 => x"08",
          3869 => x"52",
          3870 => x"f5",
          3871 => x"5b",
          3872 => x"e9",
          3873 => x"84",
          3874 => x"2e",
          3875 => x"73",
          3876 => x"04",
          3877 => x"8c",
          3878 => x"2e",
          3879 => x"ba",
          3880 => x"73",
          3881 => x"04",
          3882 => x"0c",
          3883 => x"82",
          3884 => x"f4",
          3885 => x"fc",
          3886 => x"81",
          3887 => x"76",
          3888 => x"34",
          3889 => x"17",
          3890 => x"b9",
          3891 => x"05",
          3892 => x"ff",
          3893 => x"56",
          3894 => x"34",
          3895 => x"10",
          3896 => x"55",
          3897 => x"83",
          3898 => x"fe",
          3899 => x"0d",
          3900 => x"70",
          3901 => x"11",
          3902 => x"83",
          3903 => x"93",
          3904 => x"26",
          3905 => x"84",
          3906 => x"72",
          3907 => x"34",
          3908 => x"84",
          3909 => x"f7",
          3910 => x"05",
          3911 => x"81",
          3912 => x"ba",
          3913 => x"54",
          3914 => x"85",
          3915 => x"53",
          3916 => x"84",
          3917 => x"74",
          3918 => x"8c",
          3919 => x"26",
          3920 => x"54",
          3921 => x"73",
          3922 => x"3d",
          3923 => x"70",
          3924 => x"78",
          3925 => x"3d",
          3926 => x"af",
          3927 => x"54",
          3928 => x"88",
          3929 => x"83",
          3930 => x"0b",
          3931 => x"75",
          3932 => x"ba",
          3933 => x"80",
          3934 => x"08",
          3935 => x"d6",
          3936 => x"73",
          3937 => x"55",
          3938 => x"0d",
          3939 => x"81",
          3940 => x"26",
          3941 => x"0d",
          3942 => x"02",
          3943 => x"55",
          3944 => x"84",
          3945 => x"06",
          3946 => x"0b",
          3947 => x"70",
          3948 => x"ad",
          3949 => x"53",
          3950 => x"0d",
          3951 => x"84",
          3952 => x"81",
          3953 => x"8c",
          3954 => x"2b",
          3955 => x"70",
          3956 => x"81",
          3957 => x"38",
          3958 => x"ea",
          3959 => x"70",
          3960 => x"92",
          3961 => x"54",
          3962 => x"08",
          3963 => x"90",
          3964 => x"0b",
          3965 => x"74",
          3966 => x"77",
          3967 => x"38",
          3968 => x"51",
          3969 => x"80",
          3970 => x"ba",
          3971 => x"54",
          3972 => x"53",
          3973 => x"3f",
          3974 => x"2e",
          3975 => x"8c",
          3976 => x"70",
          3977 => x"84",
          3978 => x"74",
          3979 => x"33",
          3980 => x"ff",
          3981 => x"79",
          3982 => x"3f",
          3983 => x"2e",
          3984 => x"18",
          3985 => x"06",
          3986 => x"80",
          3987 => x"05",
          3988 => x"38",
          3989 => x"ff",
          3990 => x"d2",
          3991 => x"34",
          3992 => x"c1",
          3993 => x"84",
          3994 => x"9d",
          3995 => x"19",
          3996 => x"34",
          3997 => x"19",
          3998 => x"a1",
          3999 => x"84",
          4000 => x"7a",
          4001 => x"5b",
          4002 => x"2a",
          4003 => x"90",
          4004 => x"7a",
          4005 => x"34",
          4006 => x"1a",
          4007 => x"52",
          4008 => x"76",
          4009 => x"81",
          4010 => x"ba",
          4011 => x"fd",
          4012 => x"70",
          4013 => x"88",
          4014 => x"38",
          4015 => x"8f",
          4016 => x"58",
          4017 => x"82",
          4018 => x"09",
          4019 => x"16",
          4020 => x"5a",
          4021 => x"2e",
          4022 => x"7b",
          4023 => x"81",
          4024 => x"17",
          4025 => x"8c",
          4026 => x"81",
          4027 => x"9a",
          4028 => x"11",
          4029 => x"1b",
          4030 => x"17",
          4031 => x"83",
          4032 => x"7d",
          4033 => x"81",
          4034 => x"17",
          4035 => x"8c",
          4036 => x"81",
          4037 => x"ca",
          4038 => x"11",
          4039 => x"81",
          4040 => x"59",
          4041 => x"ff",
          4042 => x"0d",
          4043 => x"05",
          4044 => x"38",
          4045 => x"5d",
          4046 => x"81",
          4047 => x"17",
          4048 => x"3f",
          4049 => x"38",
          4050 => x"0c",
          4051 => x"fe",
          4052 => x"33",
          4053 => x"ba",
          4054 => x"04",
          4055 => x"b8",
          4056 => x"05",
          4057 => x"38",
          4058 => x"5e",
          4059 => x"82",
          4060 => x"17",
          4061 => x"3f",
          4062 => x"38",
          4063 => x"0c",
          4064 => x"83",
          4065 => x"11",
          4066 => x"71",
          4067 => x"72",
          4068 => x"ff",
          4069 => x"8c",
          4070 => x"8f",
          4071 => x"08",
          4072 => x"33",
          4073 => x"84",
          4074 => x"06",
          4075 => x"83",
          4076 => x"08",
          4077 => x"7d",
          4078 => x"82",
          4079 => x"81",
          4080 => x"17",
          4081 => x"52",
          4082 => x"7a",
          4083 => x"17",
          4084 => x"18",
          4085 => x"ba",
          4086 => x"82",
          4087 => x"18",
          4088 => x"31",
          4089 => x"38",
          4090 => x"81",
          4091 => x"fb",
          4092 => x"53",
          4093 => x"52",
          4094 => x"ba",
          4095 => x"fd",
          4096 => x"18",
          4097 => x"31",
          4098 => x"a0",
          4099 => x"17",
          4100 => x"06",
          4101 => x"08",
          4102 => x"81",
          4103 => x"5a",
          4104 => x"08",
          4105 => x"33",
          4106 => x"84",
          4107 => x"06",
          4108 => x"83",
          4109 => x"08",
          4110 => x"74",
          4111 => x"82",
          4112 => x"81",
          4113 => x"17",
          4114 => x"52",
          4115 => x"7c",
          4116 => x"17",
          4117 => x"52",
          4118 => x"fa",
          4119 => x"38",
          4120 => x"62",
          4121 => x"76",
          4122 => x"27",
          4123 => x"2e",
          4124 => x"38",
          4125 => x"84",
          4126 => x"75",
          4127 => x"80",
          4128 => x"78",
          4129 => x"7c",
          4130 => x"06",
          4131 => x"b8",
          4132 => x"87",
          4133 => x"85",
          4134 => x"1a",
          4135 => x"75",
          4136 => x"83",
          4137 => x"1f",
          4138 => x"1f",
          4139 => x"84",
          4140 => x"74",
          4141 => x"38",
          4142 => x"58",
          4143 => x"76",
          4144 => x"33",
          4145 => x"81",
          4146 => x"53",
          4147 => x"f1",
          4148 => x"2e",
          4149 => x"b4",
          4150 => x"38",
          4151 => x"05",
          4152 => x"2b",
          4153 => x"07",
          4154 => x"7d",
          4155 => x"7d",
          4156 => x"7d",
          4157 => x"81",
          4158 => x"75",
          4159 => x"1b",
          4160 => x"5a",
          4161 => x"83",
          4162 => x"7d",
          4163 => x"81",
          4164 => x"19",
          4165 => x"8c",
          4166 => x"81",
          4167 => x"7b",
          4168 => x"19",
          4169 => x"5f",
          4170 => x"8f",
          4171 => x"77",
          4172 => x"74",
          4173 => x"7d",
          4174 => x"80",
          4175 => x"76",
          4176 => x"53",
          4177 => x"52",
          4178 => x"ba",
          4179 => x"80",
          4180 => x"1a",
          4181 => x"08",
          4182 => x"08",
          4183 => x"8b",
          4184 => x"2e",
          4185 => x"76",
          4186 => x"3f",
          4187 => x"38",
          4188 => x"0c",
          4189 => x"06",
          4190 => x"56",
          4191 => x"33",
          4192 => x"56",
          4193 => x"1a",
          4194 => x"53",
          4195 => x"52",
          4196 => x"ba",
          4197 => x"fc",
          4198 => x"1a",
          4199 => x"08",
          4200 => x"08",
          4201 => x"fb",
          4202 => x"82",
          4203 => x"81",
          4204 => x"19",
          4205 => x"fb",
          4206 => x"19",
          4207 => x"ee",
          4208 => x"08",
          4209 => x"38",
          4210 => x"b4",
          4211 => x"a0",
          4212 => x"40",
          4213 => x"38",
          4214 => x"09",
          4215 => x"7d",
          4216 => x"51",
          4217 => x"39",
          4218 => x"53",
          4219 => x"3f",
          4220 => x"2e",
          4221 => x"ba",
          4222 => x"08",
          4223 => x"08",
          4224 => x"5e",
          4225 => x"19",
          4226 => x"06",
          4227 => x"53",
          4228 => x"86",
          4229 => x"54",
          4230 => x"33",
          4231 => x"8b",
          4232 => x"7a",
          4233 => x"5f",
          4234 => x"2a",
          4235 => x"39",
          4236 => x"82",
          4237 => x"11",
          4238 => x"0a",
          4239 => x"58",
          4240 => x"88",
          4241 => x"90",
          4242 => x"98",
          4243 => x"cf",
          4244 => x"08",
          4245 => x"90",
          4246 => x"f4",
          4247 => x"ec",
          4248 => x"73",
          4249 => x"2e",
          4250 => x"56",
          4251 => x"82",
          4252 => x"75",
          4253 => x"ba",
          4254 => x"80",
          4255 => x"b1",
          4256 => x"30",
          4257 => x"07",
          4258 => x"38",
          4259 => x"b5",
          4260 => x"0c",
          4261 => x"91",
          4262 => x"39",
          4263 => x"81",
          4264 => x"db",
          4265 => x"ba",
          4266 => x"19",
          4267 => x"38",
          4268 => x"56",
          4269 => x"82",
          4270 => x"3f",
          4271 => x"2e",
          4272 => x"09",
          4273 => x"70",
          4274 => x"51",
          4275 => x"84",
          4276 => x"90",
          4277 => x"a3",
          4278 => x"9b",
          4279 => x"39",
          4280 => x"53",
          4281 => x"84",
          4282 => x"30",
          4283 => x"25",
          4284 => x"74",
          4285 => x"9c",
          4286 => x"56",
          4287 => x"15",
          4288 => x"07",
          4289 => x"74",
          4290 => x"04",
          4291 => x"3d",
          4292 => x"fe",
          4293 => x"38",
          4294 => x"8b",
          4295 => x"a7",
          4296 => x"8c",
          4297 => x"74",
          4298 => x"ff",
          4299 => x"71",
          4300 => x"0a",
          4301 => x"53",
          4302 => x"0c",
          4303 => x"38",
          4304 => x"cc",
          4305 => x"88",
          4306 => x"a9",
          4307 => x"74",
          4308 => x"82",
          4309 => x"89",
          4310 => x"ff",
          4311 => x"80",
          4312 => x"3d",
          4313 => x"0c",
          4314 => x"55",
          4315 => x"17",
          4316 => x"76",
          4317 => x"fe",
          4318 => x"75",
          4319 => x"76",
          4320 => x"53",
          4321 => x"74",
          4322 => x"ba",
          4323 => x"ff",
          4324 => x"8c",
          4325 => x"08",
          4326 => x"ff",
          4327 => x"76",
          4328 => x"0b",
          4329 => x"04",
          4330 => x"12",
          4331 => x"80",
          4332 => x"98",
          4333 => x"56",
          4334 => x"ff",
          4335 => x"94",
          4336 => x"79",
          4337 => x"74",
          4338 => x"18",
          4339 => x"b8",
          4340 => x"84",
          4341 => x"77",
          4342 => x"05",
          4343 => x"38",
          4344 => x"84",
          4345 => x"0b",
          4346 => x"81",
          4347 => x"c6",
          4348 => x"08",
          4349 => x"81",
          4350 => x"51",
          4351 => x"5d",
          4352 => x"2e",
          4353 => x"8c",
          4354 => x"56",
          4355 => x"86",
          4356 => x"33",
          4357 => x"18",
          4358 => x"80",
          4359 => x"19",
          4360 => x"05",
          4361 => x"19",
          4362 => x"76",
          4363 => x"55",
          4364 => x"22",
          4365 => x"81",
          4366 => x"19",
          4367 => x"8c",
          4368 => x"dd",
          4369 => x"84",
          4370 => x"75",
          4371 => x"70",
          4372 => x"86",
          4373 => x"38",
          4374 => x"b4",
          4375 => x"74",
          4376 => x"82",
          4377 => x"81",
          4378 => x"19",
          4379 => x"52",
          4380 => x"fe",
          4381 => x"83",
          4382 => x"09",
          4383 => x"0c",
          4384 => x"5e",
          4385 => x"85",
          4386 => x"b0",
          4387 => x"fc",
          4388 => x"0c",
          4389 => x"64",
          4390 => x"5b",
          4391 => x"5e",
          4392 => x"b8",
          4393 => x"19",
          4394 => x"19",
          4395 => x"09",
          4396 => x"75",
          4397 => x"51",
          4398 => x"80",
          4399 => x"79",
          4400 => x"90",
          4401 => x"58",
          4402 => x"18",
          4403 => x"5b",
          4404 => x"e5",
          4405 => x"30",
          4406 => x"54",
          4407 => x"74",
          4408 => x"2e",
          4409 => x"86",
          4410 => x"51",
          4411 => x"5b",
          4412 => x"98",
          4413 => x"7a",
          4414 => x"04",
          4415 => x"52",
          4416 => x"81",
          4417 => x"09",
          4418 => x"8c",
          4419 => x"a8",
          4420 => x"58",
          4421 => x"b5",
          4422 => x"2e",
          4423 => x"54",
          4424 => x"53",
          4425 => x"de",
          4426 => x"8f",
          4427 => x"76",
          4428 => x"2e",
          4429 => x"bf",
          4430 => x"05",
          4431 => x"ab",
          4432 => x"cc",
          4433 => x"81",
          4434 => x"5b",
          4435 => x"ba",
          4436 => x"5b",
          4437 => x"7d",
          4438 => x"8c",
          4439 => x"33",
          4440 => x"75",
          4441 => x"bf",
          4442 => x"81",
          4443 => x"33",
          4444 => x"71",
          4445 => x"80",
          4446 => x"26",
          4447 => x"76",
          4448 => x"5a",
          4449 => x"38",
          4450 => x"59",
          4451 => x"81",
          4452 => x"61",
          4453 => x"70",
          4454 => x"39",
          4455 => x"81",
          4456 => x"38",
          4457 => x"75",
          4458 => x"05",
          4459 => x"ff",
          4460 => x"e4",
          4461 => x"ff",
          4462 => x"8c",
          4463 => x"0d",
          4464 => x"7b",
          4465 => x"08",
          4466 => x"38",
          4467 => x"ac",
          4468 => x"08",
          4469 => x"2e",
          4470 => x"58",
          4471 => x"81",
          4472 => x"1b",
          4473 => x"3f",
          4474 => x"38",
          4475 => x"0c",
          4476 => x"1c",
          4477 => x"2e",
          4478 => x"06",
          4479 => x"86",
          4480 => x"f2",
          4481 => x"75",
          4482 => x"e2",
          4483 => x"7c",
          4484 => x"57",
          4485 => x"05",
          4486 => x"76",
          4487 => x"59",
          4488 => x"2e",
          4489 => x"06",
          4490 => x"1d",
          4491 => x"33",
          4492 => x"71",
          4493 => x"76",
          4494 => x"2e",
          4495 => x"ac",
          4496 => x"c8",
          4497 => x"ba",
          4498 => x"79",
          4499 => x"04",
          4500 => x"52",
          4501 => x"81",
          4502 => x"09",
          4503 => x"8c",
          4504 => x"a8",
          4505 => x"58",
          4506 => x"ea",
          4507 => x"2e",
          4508 => x"54",
          4509 => x"53",
          4510 => x"b6",
          4511 => x"5a",
          4512 => x"86",
          4513 => x"f2",
          4514 => x"79",
          4515 => x"77",
          4516 => x"7f",
          4517 => x"7d",
          4518 => x"5d",
          4519 => x"84",
          4520 => x"08",
          4521 => x"39",
          4522 => x"ff",
          4523 => x"a2",
          4524 => x"2e",
          4525 => x"08",
          4526 => x"88",
          4527 => x"b3",
          4528 => x"29",
          4529 => x"56",
          4530 => x"81",
          4531 => x"07",
          4532 => x"ed",
          4533 => x"38",
          4534 => x"ba",
          4535 => x"22",
          4536 => x"a0",
          4537 => x"2e",
          4538 => x"56",
          4539 => x"b0",
          4540 => x"06",
          4541 => x"74",
          4542 => x"05",
          4543 => x"38",
          4544 => x"5a",
          4545 => x"8c",
          4546 => x"ff",
          4547 => x"55",
          4548 => x"70",
          4549 => x"06",
          4550 => x"85",
          4551 => x"22",
          4552 => x"38",
          4553 => x"51",
          4554 => x"a0",
          4555 => x"58",
          4556 => x"77",
          4557 => x"55",
          4558 => x"33",
          4559 => x"2e",
          4560 => x"1f",
          4561 => x"8c",
          4562 => x"61",
          4563 => x"59",
          4564 => x"ff",
          4565 => x"27",
          4566 => x"57",
          4567 => x"1a",
          4568 => x"77",
          4569 => x"ff",
          4570 => x"44",
          4571 => x"38",
          4572 => x"18",
          4573 => x"22",
          4574 => x"05",
          4575 => x"07",
          4576 => x"38",
          4577 => x"16",
          4578 => x"56",
          4579 => x"fe",
          4580 => x"78",
          4581 => x"a0",
          4582 => x"78",
          4583 => x"33",
          4584 => x"06",
          4585 => x"77",
          4586 => x"05",
          4587 => x"59",
          4588 => x"87",
          4589 => x"84",
          4590 => x"5b",
          4591 => x"87",
          4592 => x"38",
          4593 => x"8c",
          4594 => x"d6",
          4595 => x"1f",
          4596 => x"db",
          4597 => x"81",
          4598 => x"90",
          4599 => x"89",
          4600 => x"5b",
          4601 => x"84",
          4602 => x"08",
          4603 => x"b8",
          4604 => x"80",
          4605 => x"f3",
          4606 => x"2e",
          4607 => x"54",
          4608 => x"33",
          4609 => x"08",
          4610 => x"57",
          4611 => x"bc",
          4612 => x"42",
          4613 => x"74",
          4614 => x"5f",
          4615 => x"19",
          4616 => x"81",
          4617 => x"ba",
          4618 => x"80",
          4619 => x"84",
          4620 => x"81",
          4621 => x"f3",
          4622 => x"08",
          4623 => x"78",
          4624 => x"54",
          4625 => x"33",
          4626 => x"08",
          4627 => x"56",
          4628 => x"80",
          4629 => x"57",
          4630 => x"34",
          4631 => x"0b",
          4632 => x"75",
          4633 => x"81",
          4634 => x"ef",
          4635 => x"98",
          4636 => x"81",
          4637 => x"84",
          4638 => x"81",
          4639 => x"57",
          4640 => x"59",
          4641 => x"84",
          4642 => x"08",
          4643 => x"39",
          4644 => x"52",
          4645 => x"84",
          4646 => x"06",
          4647 => x"83",
          4648 => x"08",
          4649 => x"8b",
          4650 => x"2e",
          4651 => x"57",
          4652 => x"1f",
          4653 => x"e9",
          4654 => x"84",
          4655 => x"84",
          4656 => x"74",
          4657 => x"78",
          4658 => x"05",
          4659 => x"56",
          4660 => x"06",
          4661 => x"57",
          4662 => x"b2",
          4663 => x"2e",
          4664 => x"54",
          4665 => x"33",
          4666 => x"08",
          4667 => x"56",
          4668 => x"fe",
          4669 => x"08",
          4670 => x"60",
          4671 => x"34",
          4672 => x"34",
          4673 => x"f3",
          4674 => x"83",
          4675 => x"1f",
          4676 => x"83",
          4677 => x"76",
          4678 => x"88",
          4679 => x"38",
          4680 => x"8c",
          4681 => x"ff",
          4682 => x"70",
          4683 => x"a6",
          4684 => x"1d",
          4685 => x"3f",
          4686 => x"8c",
          4687 => x"40",
          4688 => x"81",
          4689 => x"70",
          4690 => x"96",
          4691 => x"fc",
          4692 => x"1d",
          4693 => x"31",
          4694 => x"a0",
          4695 => x"1c",
          4696 => x"06",
          4697 => x"08",
          4698 => x"81",
          4699 => x"56",
          4700 => x"70",
          4701 => x"2e",
          4702 => x"ff",
          4703 => x"2e",
          4704 => x"80",
          4705 => x"54",
          4706 => x"1c",
          4707 => x"8c",
          4708 => x"38",
          4709 => x"b4",
          4710 => x"74",
          4711 => x"1c",
          4712 => x"84",
          4713 => x"75",
          4714 => x"fa",
          4715 => x"57",
          4716 => x"75",
          4717 => x"39",
          4718 => x"08",
          4719 => x"51",
          4720 => x"54",
          4721 => x"53",
          4722 => x"96",
          4723 => x"7f",
          4724 => x"0b",
          4725 => x"2e",
          4726 => x"2e",
          4727 => x"8c",
          4728 => x"5c",
          4729 => x"54",
          4730 => x"55",
          4731 => x"80",
          4732 => x"5a",
          4733 => x"73",
          4734 => x"58",
          4735 => x"70",
          4736 => x"5c",
          4737 => x"0b",
          4738 => x"59",
          4739 => x"33",
          4740 => x"2e",
          4741 => x"38",
          4742 => x"07",
          4743 => x"26",
          4744 => x"ae",
          4745 => x"18",
          4746 => x"34",
          4747 => x"ba",
          4748 => x"0b",
          4749 => x"72",
          4750 => x"0b",
          4751 => x"94",
          4752 => x"9c",
          4753 => x"73",
          4754 => x"1c",
          4755 => x"34",
          4756 => x"33",
          4757 => x"88",
          4758 => x"07",
          4759 => x"0c",
          4760 => x"71",
          4761 => x"5a",
          4762 => x"99",
          4763 => x"2b",
          4764 => x"8f",
          4765 => x"c0",
          4766 => x"7a",
          4767 => x"7a",
          4768 => x"89",
          4769 => x"ff",
          4770 => x"38",
          4771 => x"88",
          4772 => x"18",
          4773 => x"8c",
          4774 => x"11",
          4775 => x"90",
          4776 => x"30",
          4777 => x"25",
          4778 => x"38",
          4779 => x"80",
          4780 => x"39",
          4781 => x"57",
          4782 => x"96",
          4783 => x"33",
          4784 => x"26",
          4785 => x"33",
          4786 => x"72",
          4787 => x"7d",
          4788 => x"83",
          4789 => x"70",
          4790 => x"16",
          4791 => x"57",
          4792 => x"fd",
          4793 => x"39",
          4794 => x"30",
          4795 => x"a9",
          4796 => x"70",
          4797 => x"57",
          4798 => x"81",
          4799 => x"38",
          4800 => x"16",
          4801 => x"3d",
          4802 => x"27",
          4803 => x"08",
          4804 => x"05",
          4805 => x"38",
          4806 => x"ec",
          4807 => x"38",
          4808 => x"81",
          4809 => x"70",
          4810 => x"71",
          4811 => x"73",
          4812 => x"82",
          4813 => x"38",
          4814 => x"33",
          4815 => x"73",
          4816 => x"2e",
          4817 => x"81",
          4818 => x"38",
          4819 => x"84",
          4820 => x"38",
          4821 => x"81",
          4822 => x"33",
          4823 => x"f0",
          4824 => x"dc",
          4825 => x"07",
          4826 => x"a1",
          4827 => x"74",
          4828 => x"38",
          4829 => x"80",
          4830 => x"e1",
          4831 => x"96",
          4832 => x"9f",
          4833 => x"b5",
          4834 => x"84",
          4835 => x"54",
          4836 => x"84",
          4837 => x"83",
          4838 => x"5c",
          4839 => x"e4",
          4840 => x"80",
          4841 => x"ba",
          4842 => x"3d",
          4843 => x"70",
          4844 => x"55",
          4845 => x"81",
          4846 => x"55",
          4847 => x"80",
          4848 => x"78",
          4849 => x"73",
          4850 => x"5a",
          4851 => x"82",
          4852 => x"76",
          4853 => x"11",
          4854 => x"70",
          4855 => x"5f",
          4856 => x"72",
          4857 => x"38",
          4858 => x"23",
          4859 => x"78",
          4860 => x"58",
          4861 => x"e6",
          4862 => x"72",
          4863 => x"2e",
          4864 => x"22",
          4865 => x"76",
          4866 => x"57",
          4867 => x"70",
          4868 => x"81",
          4869 => x"55",
          4870 => x"34",
          4871 => x"73",
          4872 => x"81",
          4873 => x"2e",
          4874 => x"d0",
          4875 => x"80",
          4876 => x"85",
          4877 => x"59",
          4878 => x"75",
          4879 => x"80",
          4880 => x"54",
          4881 => x"8b",
          4882 => x"8a",
          4883 => x"26",
          4884 => x"7e",
          4885 => x"57",
          4886 => x"18",
          4887 => x"a0",
          4888 => x"83",
          4889 => x"38",
          4890 => x"82",
          4891 => x"83",
          4892 => x"81",
          4893 => x"06",
          4894 => x"90",
          4895 => x"5e",
          4896 => x"07",
          4897 => x"e4",
          4898 => x"1d",
          4899 => x"80",
          4900 => x"08",
          4901 => x"38",
          4902 => x"80",
          4903 => x"81",
          4904 => x"08",
          4905 => x"08",
          4906 => x"16",
          4907 => x"40",
          4908 => x"75",
          4909 => x"07",
          4910 => x"56",
          4911 => x"ac",
          4912 => x"09",
          4913 => x"18",
          4914 => x"1d",
          4915 => x"83",
          4916 => x"05",
          4917 => x"27",
          4918 => x"ab",
          4919 => x"84",
          4920 => x"54",
          4921 => x"74",
          4922 => x"ce",
          4923 => x"81",
          4924 => x"cd",
          4925 => x"60",
          4926 => x"12",
          4927 => x"41",
          4928 => x"d8",
          4929 => x"65",
          4930 => x"55",
          4931 => x"17",
          4932 => x"39",
          4933 => x"fd",
          4934 => x"06",
          4935 => x"2e",
          4936 => x"82",
          4937 => x"a0",
          4938 => x"06",
          4939 => x"0b",
          4940 => x"8c",
          4941 => x"ff",
          4942 => x"80",
          4943 => x"26",
          4944 => x"77",
          4945 => x"79",
          4946 => x"51",
          4947 => x"08",
          4948 => x"81",
          4949 => x"38",
          4950 => x"11",
          4951 => x"ff",
          4952 => x"38",
          4953 => x"33",
          4954 => x"73",
          4955 => x"2e",
          4956 => x"81",
          4957 => x"38",
          4958 => x"d4",
          4959 => x"26",
          4960 => x"ff",
          4961 => x"78",
          4962 => x"70",
          4963 => x"ff",
          4964 => x"1b",
          4965 => x"1b",
          4966 => x"80",
          4967 => x"33",
          4968 => x"80",
          4969 => x"83",
          4970 => x"55",
          4971 => x"39",
          4972 => x"33",
          4973 => x"77",
          4974 => x"95",
          4975 => x"2a",
          4976 => x"7c",
          4977 => x"34",
          4978 => x"83",
          4979 => x"81",
          4980 => x"38",
          4981 => x"06",
          4982 => x"84",
          4983 => x"eb",
          4984 => x"80",
          4985 => x"61",
          4986 => x"42",
          4987 => x"70",
          4988 => x"56",
          4989 => x"74",
          4990 => x"38",
          4991 => x"24",
          4992 => x"d1",
          4993 => x"58",
          4994 => x"61",
          4995 => x"5d",
          4996 => x"17",
          4997 => x"ba",
          4998 => x"06",
          4999 => x"38",
          5000 => x"ba",
          5001 => x"52",
          5002 => x"3f",
          5003 => x"70",
          5004 => x"84",
          5005 => x"75",
          5006 => x"60",
          5007 => x"18",
          5008 => x"7b",
          5009 => x"17",
          5010 => x"ff",
          5011 => x"7b",
          5012 => x"74",
          5013 => x"38",
          5014 => x"33",
          5015 => x"56",
          5016 => x"38",
          5017 => x"81",
          5018 => x"81",
          5019 => x"8d",
          5020 => x"80",
          5021 => x"71",
          5022 => x"80",
          5023 => x"80",
          5024 => x"71",
          5025 => x"38",
          5026 => x"12",
          5027 => x"07",
          5028 => x"2b",
          5029 => x"43",
          5030 => x"80",
          5031 => x"c8",
          5032 => x"06",
          5033 => x"26",
          5034 => x"76",
          5035 => x"5f",
          5036 => x"77",
          5037 => x"78",
          5038 => x"ca",
          5039 => x"88",
          5040 => x"23",
          5041 => x"58",
          5042 => x"33",
          5043 => x"07",
          5044 => x"17",
          5045 => x"90",
          5046 => x"33",
          5047 => x"71",
          5048 => x"42",
          5049 => x"33",
          5050 => x"58",
          5051 => x"1c",
          5052 => x"26",
          5053 => x"31",
          5054 => x"8c",
          5055 => x"2e",
          5056 => x"80",
          5057 => x"83",
          5058 => x"38",
          5059 => x"eb",
          5060 => x"19",
          5061 => x"70",
          5062 => x"0c",
          5063 => x"38",
          5064 => x"80",
          5065 => x"18",
          5066 => x"8d",
          5067 => x"7a",
          5068 => x"15",
          5069 => x"18",
          5070 => x"18",
          5071 => x"80",
          5072 => x"86",
          5073 => x"e4",
          5074 => x"e4",
          5075 => x"ec",
          5076 => x"18",
          5077 => x"0c",
          5078 => x"ba",
          5079 => x"33",
          5080 => x"57",
          5081 => x"17",
          5082 => x"59",
          5083 => x"7e",
          5084 => x"7c",
          5085 => x"05",
          5086 => x"33",
          5087 => x"99",
          5088 => x"ff",
          5089 => x"77",
          5090 => x"81",
          5091 => x"9f",
          5092 => x"81",
          5093 => x"78",
          5094 => x"9f",
          5095 => x"80",
          5096 => x"1e",
          5097 => x"38",
          5098 => x"2e",
          5099 => x"06",
          5100 => x"80",
          5101 => x"57",
          5102 => x"06",
          5103 => x"32",
          5104 => x"5a",
          5105 => x"81",
          5106 => x"77",
          5107 => x"33",
          5108 => x"38",
          5109 => x"33",
          5110 => x"83",
          5111 => x"2b",
          5112 => x"59",
          5113 => x"84",
          5114 => x"57",
          5115 => x"84",
          5116 => x"9f",
          5117 => x"10",
          5118 => x"44",
          5119 => x"5b",
          5120 => x"38",
          5121 => x"b4",
          5122 => x"ff",
          5123 => x"b8",
          5124 => x"b4",
          5125 => x"2e",
          5126 => x"b4",
          5127 => x"81",
          5128 => x"07",
          5129 => x"d5",
          5130 => x"0b",
          5131 => x"e9",
          5132 => x"32",
          5133 => x"42",
          5134 => x"e8",
          5135 => x"ff",
          5136 => x"1e",
          5137 => x"81",
          5138 => x"27",
          5139 => x"b7",
          5140 => x"83",
          5141 => x"39",
          5142 => x"bc",
          5143 => x"5d",
          5144 => x"71",
          5145 => x"56",
          5146 => x"80",
          5147 => x"18",
          5148 => x"70",
          5149 => x"05",
          5150 => x"5b",
          5151 => x"8e",
          5152 => x"58",
          5153 => x"93",
          5154 => x"3d",
          5155 => x"fe",
          5156 => x"83",
          5157 => x"39",
          5158 => x"3d",
          5159 => x"83",
          5160 => x"81",
          5161 => x"5c",
          5162 => x"57",
          5163 => x"38",
          5164 => x"81",
          5165 => x"58",
          5166 => x"70",
          5167 => x"ff",
          5168 => x"2e",
          5169 => x"38",
          5170 => x"fc",
          5171 => x"80",
          5172 => x"71",
          5173 => x"2e",
          5174 => x"1b",
          5175 => x"2e",
          5176 => x"7a",
          5177 => x"81",
          5178 => x"17",
          5179 => x"ba",
          5180 => x"58",
          5181 => x"f9",
          5182 => x"b7",
          5183 => x"88",
          5184 => x"d5",
          5185 => x"b8",
          5186 => x"71",
          5187 => x"14",
          5188 => x"33",
          5189 => x"5c",
          5190 => x"2e",
          5191 => x"9c",
          5192 => x"71",
          5193 => x"14",
          5194 => x"33",
          5195 => x"5a",
          5196 => x"2e",
          5197 => x"a0",
          5198 => x"71",
          5199 => x"14",
          5200 => x"33",
          5201 => x"a4",
          5202 => x"71",
          5203 => x"14",
          5204 => x"33",
          5205 => x"44",
          5206 => x"56",
          5207 => x"22",
          5208 => x"23",
          5209 => x"0b",
          5210 => x"0c",
          5211 => x"f0",
          5212 => x"95",
          5213 => x"b8",
          5214 => x"59",
          5215 => x"08",
          5216 => x"38",
          5217 => x"b4",
          5218 => x"7f",
          5219 => x"17",
          5220 => x"38",
          5221 => x"39",
          5222 => x"38",
          5223 => x"c0",
          5224 => x"e3",
          5225 => x"88",
          5226 => x"f6",
          5227 => x"f6",
          5228 => x"33",
          5229 => x"88",
          5230 => x"07",
          5231 => x"1e",
          5232 => x"44",
          5233 => x"58",
          5234 => x"58",
          5235 => x"a8",
          5236 => x"59",
          5237 => x"da",
          5238 => x"17",
          5239 => x"52",
          5240 => x"3f",
          5241 => x"80",
          5242 => x"3d",
          5243 => x"75",
          5244 => x"81",
          5245 => x"55",
          5246 => x"ed",
          5247 => x"84",
          5248 => x"80",
          5249 => x"d4",
          5250 => x"2e",
          5251 => x"73",
          5252 => x"62",
          5253 => x"80",
          5254 => x"70",
          5255 => x"84",
          5256 => x"8c",
          5257 => x"84",
          5258 => x"75",
          5259 => x"56",
          5260 => x"82",
          5261 => x"5c",
          5262 => x"80",
          5263 => x"5b",
          5264 => x"81",
          5265 => x"5a",
          5266 => x"76",
          5267 => x"81",
          5268 => x"57",
          5269 => x"70",
          5270 => x"70",
          5271 => x"09",
          5272 => x"38",
          5273 => x"07",
          5274 => x"79",
          5275 => x"1d",
          5276 => x"38",
          5277 => x"24",
          5278 => x"fe",
          5279 => x"84",
          5280 => x"89",
          5281 => x"bf",
          5282 => x"53",
          5283 => x"9f",
          5284 => x"ba",
          5285 => x"79",
          5286 => x"0c",
          5287 => x"52",
          5288 => x"3f",
          5289 => x"8c",
          5290 => x"9c",
          5291 => x"38",
          5292 => x"84",
          5293 => x"58",
          5294 => x"81",
          5295 => x"38",
          5296 => x"71",
          5297 => x"58",
          5298 => x"e9",
          5299 => x"0b",
          5300 => x"34",
          5301 => x"56",
          5302 => x"57",
          5303 => x"0b",
          5304 => x"83",
          5305 => x"0b",
          5306 => x"34",
          5307 => x"9f",
          5308 => x"16",
          5309 => x"7e",
          5310 => x"57",
          5311 => x"9c",
          5312 => x"82",
          5313 => x"02",
          5314 => x"5d",
          5315 => x"86",
          5316 => x"b8",
          5317 => x"c2",
          5318 => x"5d",
          5319 => x"2a",
          5320 => x"38",
          5321 => x"38",
          5322 => x"80",
          5323 => x"58",
          5324 => x"67",
          5325 => x"9a",
          5326 => x"33",
          5327 => x"2e",
          5328 => x"9c",
          5329 => x"71",
          5330 => x"14",
          5331 => x"33",
          5332 => x"60",
          5333 => x"5d",
          5334 => x"77",
          5335 => x"34",
          5336 => x"2a",
          5337 => x"ac",
          5338 => x"75",
          5339 => x"89",
          5340 => x"70",
          5341 => x"76",
          5342 => x"06",
          5343 => x"38",
          5344 => x"3f",
          5345 => x"8c",
          5346 => x"84",
          5347 => x"38",
          5348 => x"80",
          5349 => x"95",
          5350 => x"74",
          5351 => x"80",
          5352 => x"80",
          5353 => x"80",
          5354 => x"cd",
          5355 => x"88",
          5356 => x"fc",
          5357 => x"57",
          5358 => x"17",
          5359 => x"07",
          5360 => x"39",
          5361 => x"38",
          5362 => x"3f",
          5363 => x"8c",
          5364 => x"ba",
          5365 => x"84",
          5366 => x"38",
          5367 => x"b2",
          5368 => x"90",
          5369 => x"19",
          5370 => x"ff",
          5371 => x"84",
          5372 => x"18",
          5373 => x"a0",
          5374 => x"17",
          5375 => x"cc",
          5376 => x"71",
          5377 => x"07",
          5378 => x"34",
          5379 => x"90",
          5380 => x"34",
          5381 => x"7e",
          5382 => x"34",
          5383 => x"5d",
          5384 => x"84",
          5385 => x"72",
          5386 => x"7e",
          5387 => x"79",
          5388 => x"81",
          5389 => x"16",
          5390 => x"ba",
          5391 => x"57",
          5392 => x"56",
          5393 => x"7a",
          5394 => x"0c",
          5395 => x"08",
          5396 => x"33",
          5397 => x"ba",
          5398 => x"81",
          5399 => x"17",
          5400 => x"31",
          5401 => x"a0",
          5402 => x"16",
          5403 => x"06",
          5404 => x"08",
          5405 => x"81",
          5406 => x"7c",
          5407 => x"0c",
          5408 => x"1a",
          5409 => x"ff",
          5410 => x"38",
          5411 => x"05",
          5412 => x"df",
          5413 => x"b0",
          5414 => x"2e",
          5415 => x"9c",
          5416 => x"75",
          5417 => x"39",
          5418 => x"39",
          5419 => x"0c",
          5420 => x"fe",
          5421 => x"67",
          5422 => x"0c",
          5423 => x"79",
          5424 => x"75",
          5425 => x"86",
          5426 => x"78",
          5427 => x"74",
          5428 => x"91",
          5429 => x"90",
          5430 => x"76",
          5431 => x"08",
          5432 => x"7b",
          5433 => x"2e",
          5434 => x"ff",
          5435 => x"19",
          5436 => x"5b",
          5437 => x"88",
          5438 => x"85",
          5439 => x"74",
          5440 => x"08",
          5441 => x"41",
          5442 => x"8a",
          5443 => x"08",
          5444 => x"d5",
          5445 => x"57",
          5446 => x"1b",
          5447 => x"7b",
          5448 => x"52",
          5449 => x"3f",
          5450 => x"60",
          5451 => x"2e",
          5452 => x"56",
          5453 => x"76",
          5454 => x"55",
          5455 => x"70",
          5456 => x"74",
          5457 => x"78",
          5458 => x"1e",
          5459 => x"1d",
          5460 => x"80",
          5461 => x"3d",
          5462 => x"92",
          5463 => x"39",
          5464 => x"06",
          5465 => x"78",
          5466 => x"b4",
          5467 => x"0b",
          5468 => x"7f",
          5469 => x"38",
          5470 => x"81",
          5471 => x"84",
          5472 => x"ff",
          5473 => x"7a",
          5474 => x"83",
          5475 => x"b8",
          5476 => x"e6",
          5477 => x"77",
          5478 => x"56",
          5479 => x"70",
          5480 => x"05",
          5481 => x"38",
          5482 => x"08",
          5483 => x"33",
          5484 => x"5b",
          5485 => x"81",
          5486 => x"08",
          5487 => x"1a",
          5488 => x"55",
          5489 => x"38",
          5490 => x"09",
          5491 => x"b4",
          5492 => x"7f",
          5493 => x"fe",
          5494 => x"9c",
          5495 => x"84",
          5496 => x"ff",
          5497 => x"55",
          5498 => x"ff",
          5499 => x"81",
          5500 => x"7a",
          5501 => x"0b",
          5502 => x"8c",
          5503 => x"91",
          5504 => x"0c",
          5505 => x"62",
          5506 => x"80",
          5507 => x"9f",
          5508 => x"97",
          5509 => x"8f",
          5510 => x"59",
          5511 => x"80",
          5512 => x"c4",
          5513 => x"bc",
          5514 => x"81",
          5515 => x"2e",
          5516 => x"11",
          5517 => x"76",
          5518 => x"38",
          5519 => x"a2",
          5520 => x"78",
          5521 => x"38",
          5522 => x"55",
          5523 => x"81",
          5524 => x"86",
          5525 => x"1a",
          5526 => x"60",
          5527 => x"2e",
          5528 => x"05",
          5529 => x"77",
          5530 => x"22",
          5531 => x"56",
          5532 => x"78",
          5533 => x"80",
          5534 => x"76",
          5535 => x"58",
          5536 => x"16",
          5537 => x"ba",
          5538 => x"11",
          5539 => x"27",
          5540 => x"76",
          5541 => x"70",
          5542 => x"05",
          5543 => x"38",
          5544 => x"89",
          5545 => x"1a",
          5546 => x"1b",
          5547 => x"08",
          5548 => x"27",
          5549 => x"0c",
          5550 => x"58",
          5551 => x"1b",
          5552 => x"0c",
          5553 => x"8c",
          5554 => x"33",
          5555 => x"fe",
          5556 => x"56",
          5557 => x"31",
          5558 => x"7a",
          5559 => x"2e",
          5560 => x"71",
          5561 => x"81",
          5562 => x"53",
          5563 => x"ff",
          5564 => x"80",
          5565 => x"76",
          5566 => x"60",
          5567 => x"7a",
          5568 => x"78",
          5569 => x"05",
          5570 => x"34",
          5571 => x"58",
          5572 => x"39",
          5573 => x"16",
          5574 => x"ff",
          5575 => x"8c",
          5576 => x"ab",
          5577 => x"34",
          5578 => x"84",
          5579 => x"17",
          5580 => x"33",
          5581 => x"fe",
          5582 => x"a0",
          5583 => x"16",
          5584 => x"5c",
          5585 => x"8c",
          5586 => x"16",
          5587 => x"7c",
          5588 => x"56",
          5589 => x"f8",
          5590 => x"ff",
          5591 => x"55",
          5592 => x"90",
          5593 => x"52",
          5594 => x"ba",
          5595 => x"fb",
          5596 => x"16",
          5597 => x"17",
          5598 => x"84",
          5599 => x"ba",
          5600 => x"08",
          5601 => x"17",
          5602 => x"33",
          5603 => x"fc",
          5604 => x"a0",
          5605 => x"16",
          5606 => x"56",
          5607 => x"ff",
          5608 => x"81",
          5609 => x"7a",
          5610 => x"54",
          5611 => x"53",
          5612 => x"c6",
          5613 => x"38",
          5614 => x"b4",
          5615 => x"74",
          5616 => x"82",
          5617 => x"81",
          5618 => x"16",
          5619 => x"52",
          5620 => x"3f",
          5621 => x"08",
          5622 => x"91",
          5623 => x"0c",
          5624 => x"1b",
          5625 => x"92",
          5626 => x"58",
          5627 => x"77",
          5628 => x"75",
          5629 => x"86",
          5630 => x"78",
          5631 => x"74",
          5632 => x"90",
          5633 => x"5c",
          5634 => x"7b",
          5635 => x"08",
          5636 => x"5b",
          5637 => x"53",
          5638 => x"ff",
          5639 => x"80",
          5640 => x"78",
          5641 => x"a4",
          5642 => x"5a",
          5643 => x"88",
          5644 => x"5d",
          5645 => x"88",
          5646 => x"17",
          5647 => x"74",
          5648 => x"08",
          5649 => x"5b",
          5650 => x"56",
          5651 => x"59",
          5652 => x"80",
          5653 => x"18",
          5654 => x"80",
          5655 => x"18",
          5656 => x"34",
          5657 => x"ba",
          5658 => x"06",
          5659 => x"84",
          5660 => x"81",
          5661 => x"70",
          5662 => x"93",
          5663 => x"08",
          5664 => x"83",
          5665 => x"08",
          5666 => x"74",
          5667 => x"82",
          5668 => x"81",
          5669 => x"17",
          5670 => x"52",
          5671 => x"3f",
          5672 => x"2a",
          5673 => x"2a",
          5674 => x"08",
          5675 => x"5b",
          5676 => x"56",
          5677 => x"59",
          5678 => x"80",
          5679 => x"18",
          5680 => x"80",
          5681 => x"18",
          5682 => x"34",
          5683 => x"ba",
          5684 => x"06",
          5685 => x"ae",
          5686 => x"a5",
          5687 => x"55",
          5688 => x"56",
          5689 => x"79",
          5690 => x"ba",
          5691 => x"b1",
          5692 => x"38",
          5693 => x"38",
          5694 => x"38",
          5695 => x"52",
          5696 => x"71",
          5697 => x"75",
          5698 => x"3d",
          5699 => x"8f",
          5700 => x"06",
          5701 => x"53",
          5702 => x"7d",
          5703 => x"b2",
          5704 => x"70",
          5705 => x"ac",
          5706 => x"a4",
          5707 => x"71",
          5708 => x"34",
          5709 => x"3d",
          5710 => x"0c",
          5711 => x"11",
          5712 => x"70",
          5713 => x"81",
          5714 => x"76",
          5715 => x"e5",
          5716 => x"57",
          5717 => x"70",
          5718 => x"53",
          5719 => x"e0",
          5720 => x"ff",
          5721 => x"38",
          5722 => x"54",
          5723 => x"71",
          5724 => x"73",
          5725 => x"30",
          5726 => x"59",
          5727 => x"81",
          5728 => x"25",
          5729 => x"39",
          5730 => x"5e",
          5731 => x"80",
          5732 => x"3d",
          5733 => x"08",
          5734 => x"8a",
          5735 => x"3d",
          5736 => x"3d",
          5737 => x"ba",
          5738 => x"80",
          5739 => x"70",
          5740 => x"80",
          5741 => x"84",
          5742 => x"2e",
          5743 => x"9a",
          5744 => x"33",
          5745 => x"2e",
          5746 => x"84",
          5747 => x"84",
          5748 => x"06",
          5749 => x"8c",
          5750 => x"33",
          5751 => x"90",
          5752 => x"5b",
          5753 => x"0c",
          5754 => x"3d",
          5755 => x"e6",
          5756 => x"40",
          5757 => x"3d",
          5758 => x"51",
          5759 => x"59",
          5760 => x"60",
          5761 => x"11",
          5762 => x"db",
          5763 => x"82",
          5764 => x"40",
          5765 => x"aa",
          5766 => x"ba",
          5767 => x"df",
          5768 => x"77",
          5769 => x"83",
          5770 => x"38",
          5771 => x"81",
          5772 => x"84",
          5773 => x"ff",
          5774 => x"78",
          5775 => x"9b",
          5776 => x"2b",
          5777 => x"56",
          5778 => x"76",
          5779 => x"51",
          5780 => x"08",
          5781 => x"38",
          5782 => x"3f",
          5783 => x"8c",
          5784 => x"9b",
          5785 => x"2b",
          5786 => x"5e",
          5787 => x"76",
          5788 => x"08",
          5789 => x"84",
          5790 => x"08",
          5791 => x"2e",
          5792 => x"80",
          5793 => x"51",
          5794 => x"05",
          5795 => x"38",
          5796 => x"70",
          5797 => x"81",
          5798 => x"38",
          5799 => x"82",
          5800 => x"08",
          5801 => x"56",
          5802 => x"38",
          5803 => x"5f",
          5804 => x"08",
          5805 => x"2e",
          5806 => x"e8",
          5807 => x"05",
          5808 => x"5e",
          5809 => x"1a",
          5810 => x"74",
          5811 => x"26",
          5812 => x"94",
          5813 => x"70",
          5814 => x"79",
          5815 => x"81",
          5816 => x"81",
          5817 => x"7c",
          5818 => x"e4",
          5819 => x"17",
          5820 => x"07",
          5821 => x"39",
          5822 => x"98",
          5823 => x"80",
          5824 => x"7a",
          5825 => x"8c",
          5826 => x"2e",
          5827 => x"54",
          5828 => x"53",
          5829 => x"fe",
          5830 => x"fc",
          5831 => x"17",
          5832 => x"31",
          5833 => x"a0",
          5834 => x"16",
          5835 => x"06",
          5836 => x"08",
          5837 => x"81",
          5838 => x"7c",
          5839 => x"e6",
          5840 => x"34",
          5841 => x"10",
          5842 => x"70",
          5843 => x"7a",
          5844 => x"fd",
          5845 => x"81",
          5846 => x"81",
          5847 => x"8e",
          5848 => x"19",
          5849 => x"05",
          5850 => x"fd",
          5851 => x"78",
          5852 => x"0d",
          5853 => x"55",
          5854 => x"74",
          5855 => x"73",
          5856 => x"86",
          5857 => x"78",
          5858 => x"72",
          5859 => x"91",
          5860 => x"8c",
          5861 => x"b9",
          5862 => x"76",
          5863 => x"11",
          5864 => x"73",
          5865 => x"ff",
          5866 => x"ba",
          5867 => x"53",
          5868 => x"ba",
          5869 => x"75",
          5870 => x"77",
          5871 => x"59",
          5872 => x"77",
          5873 => x"94",
          5874 => x"16",
          5875 => x"5a",
          5876 => x"73",
          5877 => x"84",
          5878 => x"08",
          5879 => x"2e",
          5880 => x"38",
          5881 => x"82",
          5882 => x"ae",
          5883 => x"53",
          5884 => x"0d",
          5885 => x"81",
          5886 => x"75",
          5887 => x"76",
          5888 => x"38",
          5889 => x"54",
          5890 => x"16",
          5891 => x"57",
          5892 => x"06",
          5893 => x"15",
          5894 => x"16",
          5895 => x"8b",
          5896 => x"0c",
          5897 => x"80",
          5898 => x"80",
          5899 => x"84",
          5900 => x"17",
          5901 => x"56",
          5902 => x"15",
          5903 => x"56",
          5904 => x"16",
          5905 => x"05",
          5906 => x"78",
          5907 => x"08",
          5908 => x"51",
          5909 => x"08",
          5910 => x"51",
          5911 => x"08",
          5912 => x"72",
          5913 => x"73",
          5914 => x"84",
          5915 => x"08",
          5916 => x"08",
          5917 => x"8c",
          5918 => x"0c",
          5919 => x"34",
          5920 => x"3d",
          5921 => x"89",
          5922 => x"53",
          5923 => x"84",
          5924 => x"8c",
          5925 => x"2e",
          5926 => x"73",
          5927 => x"04",
          5928 => x"ff",
          5929 => x"55",
          5930 => x"ab",
          5931 => x"80",
          5932 => x"70",
          5933 => x"80",
          5934 => x"9b",
          5935 => x"2b",
          5936 => x"55",
          5937 => x"88",
          5938 => x"84",
          5939 => x"99",
          5940 => x"74",
          5941 => x"ff",
          5942 => x"39",
          5943 => x"39",
          5944 => x"98",
          5945 => x"88",
          5946 => x"fa",
          5947 => x"80",
          5948 => x"80",
          5949 => x"80",
          5950 => x"16",
          5951 => x"38",
          5952 => x"73",
          5953 => x"88",
          5954 => x"fe",
          5955 => x"81",
          5956 => x"08",
          5957 => x"7a",
          5958 => x"2e",
          5959 => x"2e",
          5960 => x"2e",
          5961 => x"22",
          5962 => x"38",
          5963 => x"80",
          5964 => x"38",
          5965 => x"3f",
          5966 => x"8c",
          5967 => x"8c",
          5968 => x"ff",
          5969 => x"ff",
          5970 => x"84",
          5971 => x"2c",
          5972 => x"54",
          5973 => x"0d",
          5974 => x"ff",
          5975 => x"ff",
          5976 => x"84",
          5977 => x"2c",
          5978 => x"54",
          5979 => x"96",
          5980 => x"ba",
          5981 => x"14",
          5982 => x"ba",
          5983 => x"d8",
          5984 => x"d2",
          5985 => x"53",
          5986 => x"56",
          5987 => x"55",
          5988 => x"38",
          5989 => x"0d",
          5990 => x"a9",
          5991 => x"ba",
          5992 => x"05",
          5993 => x"74",
          5994 => x"38",
          5995 => x"3f",
          5996 => x"0d",
          5997 => x"95",
          5998 => x"68",
          5999 => x"05",
          6000 => x"84",
          6001 => x"08",
          6002 => x"9c",
          6003 => x"59",
          6004 => x"38",
          6005 => x"0c",
          6006 => x"08",
          6007 => x"82",
          6008 => x"ba",
          6009 => x"c1",
          6010 => x"56",
          6011 => x"38",
          6012 => x"81",
          6013 => x"17",
          6014 => x"b7",
          6015 => x"85",
          6016 => x"18",
          6017 => x"cc",
          6018 => x"82",
          6019 => x"11",
          6020 => x"71",
          6021 => x"72",
          6022 => x"ff",
          6023 => x"70",
          6024 => x"83",
          6025 => x"43",
          6026 => x"56",
          6027 => x"7a",
          6028 => x"07",
          6029 => x"ba",
          6030 => x"54",
          6031 => x"53",
          6032 => x"a6",
          6033 => x"fe",
          6034 => x"18",
          6035 => x"31",
          6036 => x"a0",
          6037 => x"17",
          6038 => x"06",
          6039 => x"08",
          6040 => x"81",
          6041 => x"77",
          6042 => x"92",
          6043 => x"ff",
          6044 => x"ff",
          6045 => x"08",
          6046 => x"8c",
          6047 => x"07",
          6048 => x"5a",
          6049 => x"26",
          6050 => x"18",
          6051 => x"77",
          6052 => x"17",
          6053 => x"71",
          6054 => x"25",
          6055 => x"1f",
          6056 => x"78",
          6057 => x"5a",
          6058 => x"7a",
          6059 => x"17",
          6060 => x"34",
          6061 => x"e7",
          6062 => x"56",
          6063 => x"55",
          6064 => x"54",
          6065 => x"22",
          6066 => x"2e",
          6067 => x"75",
          6068 => x"75",
          6069 => x"81",
          6070 => x"73",
          6071 => x"08",
          6072 => x"38",
          6073 => x"77",
          6074 => x"38",
          6075 => x"82",
          6076 => x"17",
          6077 => x"07",
          6078 => x"2e",
          6079 => x"55",
          6080 => x"0d",
          6081 => x"ff",
          6082 => x"ca",
          6083 => x"ba",
          6084 => x"84",
          6085 => x"38",
          6086 => x"e5",
          6087 => x"ff",
          6088 => x"82",
          6089 => x"94",
          6090 => x"27",
          6091 => x"0c",
          6092 => x"84",
          6093 => x"ff",
          6094 => x"51",
          6095 => x"08",
          6096 => x"73",
          6097 => x"80",
          6098 => x"56",
          6099 => x"39",
          6100 => x"fd",
          6101 => x"2e",
          6102 => x"81",
          6103 => x"38",
          6104 => x"19",
          6105 => x"8c",
          6106 => x"56",
          6107 => x"27",
          6108 => x"9c",
          6109 => x"80",
          6110 => x"75",
          6111 => x"8c",
          6112 => x"e3",
          6113 => x"d2",
          6114 => x"ba",
          6115 => x"84",
          6116 => x"38",
          6117 => x"fe",
          6118 => x"ff",
          6119 => x"80",
          6120 => x"94",
          6121 => x"27",
          6122 => x"84",
          6123 => x"17",
          6124 => x"a1",
          6125 => x"33",
          6126 => x"bb",
          6127 => x"56",
          6128 => x"82",
          6129 => x"86",
          6130 => x"33",
          6131 => x"90",
          6132 => x"84",
          6133 => x"56",
          6134 => x"53",
          6135 => x"3d",
          6136 => x"8c",
          6137 => x"2e",
          6138 => x"a7",
          6139 => x"08",
          6140 => x"ab",
          6141 => x"84",
          6142 => x"93",
          6143 => x"59",
          6144 => x"98",
          6145 => x"02",
          6146 => x"5d",
          6147 => x"7d",
          6148 => x"12",
          6149 => x"41",
          6150 => x"80",
          6151 => x"57",
          6152 => x"56",
          6153 => x"38",
          6154 => x"08",
          6155 => x"8b",
          6156 => x"84",
          6157 => x"ba",
          6158 => x"b4",
          6159 => x"ba",
          6160 => x"ba",
          6161 => x"16",
          6162 => x"71",
          6163 => x"5d",
          6164 => x"84",
          6165 => x"fe",
          6166 => x"08",
          6167 => x"d3",
          6168 => x"92",
          6169 => x"ba",
          6170 => x"30",
          6171 => x"7a",
          6172 => x"95",
          6173 => x"7b",
          6174 => x"26",
          6175 => x"d2",
          6176 => x"84",
          6177 => x"a7",
          6178 => x"19",
          6179 => x"76",
          6180 => x"7a",
          6181 => x"06",
          6182 => x"b8",
          6183 => x"f1",
          6184 => x"2e",
          6185 => x"b4",
          6186 => x"9c",
          6187 => x"0b",
          6188 => x"27",
          6189 => x"ff",
          6190 => x"56",
          6191 => x"96",
          6192 => x"fe",
          6193 => x"81",
          6194 => x"81",
          6195 => x"81",
          6196 => x"09",
          6197 => x"8c",
          6198 => x"a8",
          6199 => x"59",
          6200 => x"eb",
          6201 => x"2e",
          6202 => x"54",
          6203 => x"53",
          6204 => x"f1",
          6205 => x"79",
          6206 => x"74",
          6207 => x"84",
          6208 => x"08",
          6209 => x"8c",
          6210 => x"ba",
          6211 => x"80",
          6212 => x"9b",
          6213 => x"9c",
          6214 => x"58",
          6215 => x"38",
          6216 => x"33",
          6217 => x"79",
          6218 => x"80",
          6219 => x"f7",
          6220 => x"95",
          6221 => x"3d",
          6222 => x"05",
          6223 => x"3f",
          6224 => x"8c",
          6225 => x"ba",
          6226 => x"43",
          6227 => x"ff",
          6228 => x"56",
          6229 => x"0b",
          6230 => x"04",
          6231 => x"81",
          6232 => x"33",
          6233 => x"86",
          6234 => x"74",
          6235 => x"83",
          6236 => x"57",
          6237 => x"87",
          6238 => x"80",
          6239 => x"2e",
          6240 => x"7d",
          6241 => x"5d",
          6242 => x"19",
          6243 => x"80",
          6244 => x"17",
          6245 => x"05",
          6246 => x"17",
          6247 => x"76",
          6248 => x"55",
          6249 => x"22",
          6250 => x"81",
          6251 => x"17",
          6252 => x"ba",
          6253 => x"58",
          6254 => x"81",
          6255 => x"70",
          6256 => x"ee",
          6257 => x"08",
          6258 => x"18",
          6259 => x"31",
          6260 => x"ee",
          6261 => x"2e",
          6262 => x"54",
          6263 => x"53",
          6264 => x"ed",
          6265 => x"7b",
          6266 => x"fd",
          6267 => x"fd",
          6268 => x"f2",
          6269 => x"84",
          6270 => x"38",
          6271 => x"8d",
          6272 => x"fd",
          6273 => x"51",
          6274 => x"08",
          6275 => x"11",
          6276 => x"7b",
          6277 => x"0c",
          6278 => x"84",
          6279 => x"ff",
          6280 => x"9f",
          6281 => x"74",
          6282 => x"76",
          6283 => x"38",
          6284 => x"75",
          6285 => x"56",
          6286 => x"b8",
          6287 => x"c3",
          6288 => x"1a",
          6289 => x"0b",
          6290 => x"80",
          6291 => x"ff",
          6292 => x"34",
          6293 => x"17",
          6294 => x"81",
          6295 => x"d8",
          6296 => x"70",
          6297 => x"05",
          6298 => x"38",
          6299 => x"34",
          6300 => x"5b",
          6301 => x"78",
          6302 => x"34",
          6303 => x"f0",
          6304 => x"34",
          6305 => x"ba",
          6306 => x"fd",
          6307 => x"08",
          6308 => x"97",
          6309 => x"80",
          6310 => x"58",
          6311 => x"2a",
          6312 => x"5a",
          6313 => x"55",
          6314 => x"81",
          6315 => x"ed",
          6316 => x"75",
          6317 => x"04",
          6318 => x"17",
          6319 => x"ed",
          6320 => x"2a",
          6321 => x"88",
          6322 => x"7d",
          6323 => x"1b",
          6324 => x"90",
          6325 => x"88",
          6326 => x"55",
          6327 => x"81",
          6328 => x"ec",
          6329 => x"ff",
          6330 => x"b4",
          6331 => x"80",
          6332 => x"5b",
          6333 => x"ba",
          6334 => x"75",
          6335 => x"b1",
          6336 => x"51",
          6337 => x"08",
          6338 => x"8a",
          6339 => x"3d",
          6340 => x"3d",
          6341 => x"ff",
          6342 => x"56",
          6343 => x"81",
          6344 => x"86",
          6345 => x"3d",
          6346 => x"70",
          6347 => x"05",
          6348 => x"38",
          6349 => x"58",
          6350 => x"77",
          6351 => x"55",
          6352 => x"77",
          6353 => x"8c",
          6354 => x"d8",
          6355 => x"cb",
          6356 => x"b1",
          6357 => x"70",
          6358 => x"89",
          6359 => x"ff",
          6360 => x"2e",
          6361 => x"e5",
          6362 => x"5f",
          6363 => x"79",
          6364 => x"12",
          6365 => x"38",
          6366 => x"55",
          6367 => x"89",
          6368 => x"58",
          6369 => x"55",
          6370 => x"38",
          6371 => x"70",
          6372 => x"07",
          6373 => x"38",
          6374 => x"83",
          6375 => x"5a",
          6376 => x"fd",
          6377 => x"b1",
          6378 => x"51",
          6379 => x"08",
          6380 => x"38",
          6381 => x"2e",
          6382 => x"51",
          6383 => x"08",
          6384 => x"38",
          6385 => x"88",
          6386 => x"75",
          6387 => x"81",
          6388 => x"ef",
          6389 => x"19",
          6390 => x"81",
          6391 => x"a0",
          6392 => x"5d",
          6393 => x"33",
          6394 => x"75",
          6395 => x"08",
          6396 => x"19",
          6397 => x"07",
          6398 => x"83",
          6399 => x"18",
          6400 => x"27",
          6401 => x"71",
          6402 => x"75",
          6403 => x"5d",
          6404 => x"38",
          6405 => x"38",
          6406 => x"81",
          6407 => x"84",
          6408 => x"ff",
          6409 => x"7f",
          6410 => x"7b",
          6411 => x"79",
          6412 => x"6a",
          6413 => x"7b",
          6414 => x"58",
          6415 => x"5b",
          6416 => x"38",
          6417 => x"18",
          6418 => x"ed",
          6419 => x"18",
          6420 => x"3d",
          6421 => x"95",
          6422 => x"a2",
          6423 => x"ba",
          6424 => x"5c",
          6425 => x"16",
          6426 => x"33",
          6427 => x"81",
          6428 => x"53",
          6429 => x"fe",
          6430 => x"80",
          6431 => x"76",
          6432 => x"38",
          6433 => x"81",
          6434 => x"7b",
          6435 => x"fe",
          6436 => x"55",
          6437 => x"98",
          6438 => x"e1",
          6439 => x"7f",
          6440 => x"8c",
          6441 => x"0d",
          6442 => x"b1",
          6443 => x"19",
          6444 => x"07",
          6445 => x"39",
          6446 => x"fe",
          6447 => x"fe",
          6448 => x"b1",
          6449 => x"08",
          6450 => x"fe",
          6451 => x"8c",
          6452 => x"db",
          6453 => x"34",
          6454 => x"84",
          6455 => x"17",
          6456 => x"33",
          6457 => x"fe",
          6458 => x"a0",
          6459 => x"16",
          6460 => x"58",
          6461 => x"08",
          6462 => x"33",
          6463 => x"5c",
          6464 => x"84",
          6465 => x"17",
          6466 => x"8c",
          6467 => x"27",
          6468 => x"7c",
          6469 => x"38",
          6470 => x"08",
          6471 => x"51",
          6472 => x"e8",
          6473 => x"05",
          6474 => x"33",
          6475 => x"05",
          6476 => x"3f",
          6477 => x"8c",
          6478 => x"ba",
          6479 => x"5a",
          6480 => x"ff",
          6481 => x"56",
          6482 => x"80",
          6483 => x"86",
          6484 => x"61",
          6485 => x"7a",
          6486 => x"73",
          6487 => x"83",
          6488 => x"3f",
          6489 => x"0c",
          6490 => x"67",
          6491 => x"52",
          6492 => x"84",
          6493 => x"08",
          6494 => x"8c",
          6495 => x"66",
          6496 => x"95",
          6497 => x"84",
          6498 => x"cf",
          6499 => x"55",
          6500 => x"86",
          6501 => x"59",
          6502 => x"2a",
          6503 => x"2a",
          6504 => x"2a",
          6505 => x"81",
          6506 => x"e1",
          6507 => x"ba",
          6508 => x"3d",
          6509 => x"9a",
          6510 => x"ff",
          6511 => x"84",
          6512 => x"8c",
          6513 => x"7a",
          6514 => x"06",
          6515 => x"30",
          6516 => x"7b",
          6517 => x"76",
          6518 => x"80",
          6519 => x"80",
          6520 => x"f6",
          6521 => x"74",
          6522 => x"38",
          6523 => x"81",
          6524 => x"84",
          6525 => x"ff",
          6526 => x"78",
          6527 => x"56",
          6528 => x"8b",
          6529 => x"83",
          6530 => x"83",
          6531 => x"2b",
          6532 => x"70",
          6533 => x"07",
          6534 => x"56",
          6535 => x"0d",
          6536 => x"8e",
          6537 => x"3f",
          6538 => x"8c",
          6539 => x"84",
          6540 => x"80",
          6541 => x"77",
          6542 => x"70",
          6543 => x"dc",
          6544 => x"08",
          6545 => x"38",
          6546 => x"b4",
          6547 => x"ba",
          6548 => x"08",
          6549 => x"55",
          6550 => x"a0",
          6551 => x"17",
          6552 => x"33",
          6553 => x"81",
          6554 => x"16",
          6555 => x"ba",
          6556 => x"fe",
          6557 => x"f8",
          6558 => x"84",
          6559 => x"ba",
          6560 => x"5c",
          6561 => x"1b",
          6562 => x"81",
          6563 => x"8b",
          6564 => x"77",
          6565 => x"7b",
          6566 => x"a0",
          6567 => x"57",
          6568 => x"53",
          6569 => x"3d",
          6570 => x"8c",
          6571 => x"a6",
          6572 => x"55",
          6573 => x"ff",
          6574 => x"3d",
          6575 => x"5b",
          6576 => x"b7",
          6577 => x"75",
          6578 => x"74",
          6579 => x"83",
          6580 => x"51",
          6581 => x"ba",
          6582 => x"ba",
          6583 => x"76",
          6584 => x"9c",
          6585 => x"ff",
          6586 => x"81",
          6587 => x"99",
          6588 => x"ff",
          6589 => x"89",
          6590 => x"e9",
          6591 => x"81",
          6592 => x"f8",
          6593 => x"81",
          6594 => x"2a",
          6595 => x"34",
          6596 => x"05",
          6597 => x"70",
          6598 => x"58",
          6599 => x"8f",
          6600 => x"e5",
          6601 => x"38",
          6602 => x"33",
          6603 => x"06",
          6604 => x"38",
          6605 => x"3d",
          6606 => x"84",
          6607 => x"08",
          6608 => x"84",
          6609 => x"83",
          6610 => x"84",
          6611 => x"55",
          6612 => x"84",
          6613 => x"83",
          6614 => x"81",
          6615 => x"84",
          6616 => x"08",
          6617 => x"c4",
          6618 => x"76",
          6619 => x"81",
          6620 => x"ef",
          6621 => x"34",
          6622 => x"ba",
          6623 => x"39",
          6624 => x"56",
          6625 => x"84",
          6626 => x"80",
          6627 => x"75",
          6628 => x"ee",
          6629 => x"84",
          6630 => x"06",
          6631 => x"b8",
          6632 => x"80",
          6633 => x"38",
          6634 => x"09",
          6635 => x"76",
          6636 => x"51",
          6637 => x"08",
          6638 => x"59",
          6639 => x"be",
          6640 => x"57",
          6641 => x"9e",
          6642 => x"07",
          6643 => x"38",
          6644 => x"38",
          6645 => x"3f",
          6646 => x"8c",
          6647 => x"55",
          6648 => x"55",
          6649 => x"55",
          6650 => x"ff",
          6651 => x"88",
          6652 => x"59",
          6653 => x"33",
          6654 => x"15",
          6655 => x"76",
          6656 => x"81",
          6657 => x"da",
          6658 => x"7a",
          6659 => x"34",
          6660 => x"ba",
          6661 => x"57",
          6662 => x"08",
          6663 => x"fe",
          6664 => x"79",
          6665 => x"84",
          6666 => x"18",
          6667 => x"a0",
          6668 => x"33",
          6669 => x"ba",
          6670 => x"5a",
          6671 => x"3f",
          6672 => x"8c",
          6673 => x"ae",
          6674 => x"2e",
          6675 => x"54",
          6676 => x"53",
          6677 => x"d3",
          6678 => x"0d",
          6679 => x"05",
          6680 => x"80",
          6681 => x"80",
          6682 => x"80",
          6683 => x"18",
          6684 => x"c2",
          6685 => x"a5",
          6686 => x"9d",
          6687 => x"8c",
          6688 => x"33",
          6689 => x"74",
          6690 => x"11",
          6691 => x"54",
          6692 => x"ff",
          6693 => x"07",
          6694 => x"90",
          6695 => x"58",
          6696 => x"08",
          6697 => x"78",
          6698 => x"51",
          6699 => x"55",
          6700 => x"38",
          6701 => x"2e",
          6702 => x"ff",
          6703 => x"08",
          6704 => x"7d",
          6705 => x"81",
          6706 => x"73",
          6707 => x"04",
          6708 => x"3d",
          6709 => x"d0",
          6710 => x"06",
          6711 => x"08",
          6712 => x"2e",
          6713 => x"7c",
          6714 => x"74",
          6715 => x"77",
          6716 => x"84",
          6717 => x"08",
          6718 => x"17",
          6719 => x"7e",
          6720 => x"ff",
          6721 => x"8c",
          6722 => x"07",
          6723 => x"08",
          6724 => x"76",
          6725 => x"31",
          6726 => x"07",
          6727 => x"fe",
          6728 => x"74",
          6729 => x"54",
          6730 => x"39",
          6731 => x"ba",
          6732 => x"08",
          6733 => x"87",
          6734 => x"a2",
          6735 => x"80",
          6736 => x"05",
          6737 => x"75",
          6738 => x"38",
          6739 => x"d1",
          6740 => x"e5",
          6741 => x"05",
          6742 => x"84",
          6743 => x"ba",
          6744 => x"33",
          6745 => x"fe",
          6746 => x"81",
          6747 => x"83",
          6748 => x"2a",
          6749 => x"9f",
          6750 => x"52",
          6751 => x"ba",
          6752 => x"74",
          6753 => x"80",
          6754 => x"75",
          6755 => x"80",
          6756 => x"83",
          6757 => x"83",
          6758 => x"74",
          6759 => x"3d",
          6760 => x"59",
          6761 => x"ab",
          6762 => x"07",
          6763 => x"38",
          6764 => x"54",
          6765 => x"cd",
          6766 => x"08",
          6767 => x"33",
          6768 => x"2b",
          6769 => x"d4",
          6770 => x"38",
          6771 => x"11",
          6772 => x"e7",
          6773 => x"82",
          6774 => x"2b",
          6775 => x"88",
          6776 => x"1f",
          6777 => x"90",
          6778 => x"33",
          6779 => x"71",
          6780 => x"3d",
          6781 => x"45",
          6782 => x"8e",
          6783 => x"38",
          6784 => x"87",
          6785 => x"45",
          6786 => x"61",
          6787 => x"38",
          6788 => x"38",
          6789 => x"7a",
          6790 => x"7a",
          6791 => x"0b",
          6792 => x"80",
          6793 => x"38",
          6794 => x"17",
          6795 => x"2e",
          6796 => x"77",
          6797 => x"84",
          6798 => x"84",
          6799 => x"38",
          6800 => x"84",
          6801 => x"2a",
          6802 => x"15",
          6803 => x"7b",
          6804 => x"ff",
          6805 => x"4e",
          6806 => x"38",
          6807 => x"70",
          6808 => x"82",
          6809 => x"78",
          6810 => x"ff",
          6811 => x"62",
          6812 => x"2e",
          6813 => x"ff",
          6814 => x"82",
          6815 => x"18",
          6816 => x"38",
          6817 => x"76",
          6818 => x"84",
          6819 => x"fe",
          6820 => x"9f",
          6821 => x"7c",
          6822 => x"57",
          6823 => x"82",
          6824 => x"5d",
          6825 => x"80",
          6826 => x"08",
          6827 => x"5c",
          6828 => x"ff",
          6829 => x"26",
          6830 => x"06",
          6831 => x"99",
          6832 => x"ff",
          6833 => x"2a",
          6834 => x"06",
          6835 => x"7a",
          6836 => x"2a",
          6837 => x"2e",
          6838 => x"5f",
          6839 => x"7f",
          6840 => x"05",
          6841 => x"dd",
          6842 => x"fe",
          6843 => x"84",
          6844 => x"38",
          6845 => x"75",
          6846 => x"59",
          6847 => x"39",
          6848 => x"7a",
          6849 => x"61",
          6850 => x"2e",
          6851 => x"4a",
          6852 => x"8c",
          6853 => x"8b",
          6854 => x"27",
          6855 => x"ba",
          6856 => x"98",
          6857 => x"86",
          6858 => x"38",
          6859 => x"fd",
          6860 => x"80",
          6861 => x"15",
          6862 => x"e5",
          6863 => x"05",
          6864 => x"34",
          6865 => x"8b",
          6866 => x"8c",
          6867 => x"7b",
          6868 => x"8e",
          6869 => x"61",
          6870 => x"34",
          6871 => x"80",
          6872 => x"82",
          6873 => x"6c",
          6874 => x"ad",
          6875 => x"74",
          6876 => x"4c",
          6877 => x"95",
          6878 => x"80",
          6879 => x"05",
          6880 => x"61",
          6881 => x"67",
          6882 => x"4c",
          6883 => x"2a",
          6884 => x"08",
          6885 => x"85",
          6886 => x"80",
          6887 => x"05",
          6888 => x"7c",
          6889 => x"96",
          6890 => x"61",
          6891 => x"05",
          6892 => x"61",
          6893 => x"55",
          6894 => x"70",
          6895 => x"74",
          6896 => x"80",
          6897 => x"4b",
          6898 => x"53",
          6899 => x"3f",
          6900 => x"e7",
          6901 => x"87",
          6902 => x"76",
          6903 => x"55",
          6904 => x"62",
          6905 => x"ff",
          6906 => x"f8",
          6907 => x"7c",
          6908 => x"46",
          6909 => x"70",
          6910 => x"56",
          6911 => x"76",
          6912 => x"54",
          6913 => x"c5",
          6914 => x"e6",
          6915 => x"76",
          6916 => x"55",
          6917 => x"31",
          6918 => x"05",
          6919 => x"77",
          6920 => x"56",
          6921 => x"75",
          6922 => x"79",
          6923 => x"8c",
          6924 => x"76",
          6925 => x"58",
          6926 => x"6c",
          6927 => x"58",
          6928 => x"7d",
          6929 => x"06",
          6930 => x"61",
          6931 => x"57",
          6932 => x"80",
          6933 => x"60",
          6934 => x"81",
          6935 => x"05",
          6936 => x"67",
          6937 => x"c1",
          6938 => x"3f",
          6939 => x"8c",
          6940 => x"67",
          6941 => x"67",
          6942 => x"05",
          6943 => x"6b",
          6944 => x"98",
          6945 => x"61",
          6946 => x"45",
          6947 => x"90",
          6948 => x"34",
          6949 => x"cd",
          6950 => x"52",
          6951 => x"57",
          6952 => x"80",
          6953 => x"dd",
          6954 => x"f7",
          6955 => x"ba",
          6956 => x"98",
          6957 => x"74",
          6958 => x"39",
          6959 => x"81",
          6960 => x"74",
          6961 => x"98",
          6962 => x"82",
          6963 => x"80",
          6964 => x"38",
          6965 => x"3f",
          6966 => x"87",
          6967 => x"5c",
          6968 => x"80",
          6969 => x"0a",
          6970 => x"f8",
          6971 => x"ff",
          6972 => x"d3",
          6973 => x"bf",
          6974 => x"81",
          6975 => x"38",
          6976 => x"a0",
          6977 => x"61",
          6978 => x"7a",
          6979 => x"57",
          6980 => x"39",
          6981 => x"61",
          6982 => x"c5",
          6983 => x"05",
          6984 => x"88",
          6985 => x"7c",
          6986 => x"34",
          6987 => x"05",
          6988 => x"61",
          6989 => x"34",
          6990 => x"b0",
          6991 => x"86",
          6992 => x"05",
          6993 => x"34",
          6994 => x"61",
          6995 => x"57",
          6996 => x"76",
          6997 => x"55",
          6998 => x"70",
          6999 => x"05",
          7000 => x"38",
          7001 => x"60",
          7002 => x"81",
          7003 => x"38",
          7004 => x"62",
          7005 => x"ba",
          7006 => x"fe",
          7007 => x"0b",
          7008 => x"84",
          7009 => x"7b",
          7010 => x"34",
          7011 => x"ff",
          7012 => x"ff",
          7013 => x"05",
          7014 => x"61",
          7015 => x"34",
          7016 => x"34",
          7017 => x"86",
          7018 => x"be",
          7019 => x"80",
          7020 => x"17",
          7021 => x"d2",
          7022 => x"55",
          7023 => x"34",
          7024 => x"34",
          7025 => x"83",
          7026 => x"e5",
          7027 => x"05",
          7028 => x"34",
          7029 => x"e8",
          7030 => x"61",
          7031 => x"56",
          7032 => x"98",
          7033 => x"34",
          7034 => x"61",
          7035 => x"ee",
          7036 => x"34",
          7037 => x"34",
          7038 => x"79",
          7039 => x"81",
          7040 => x"bd",
          7041 => x"a6",
          7042 => x"5b",
          7043 => x"57",
          7044 => x"59",
          7045 => x"78",
          7046 => x"7b",
          7047 => x"8d",
          7048 => x"38",
          7049 => x"81",
          7050 => x"77",
          7051 => x"7a",
          7052 => x"84",
          7053 => x"f7",
          7054 => x"05",
          7055 => x"d5",
          7056 => x"24",
          7057 => x"8c",
          7058 => x"16",
          7059 => x"84",
          7060 => x"8b",
          7061 => x"54",
          7062 => x"51",
          7063 => x"70",
          7064 => x"30",
          7065 => x"0c",
          7066 => x"76",
          7067 => x"e3",
          7068 => x"8d",
          7069 => x"55",
          7070 => x"ff",
          7071 => x"08",
          7072 => x"38",
          7073 => x"38",
          7074 => x"77",
          7075 => x"24",
          7076 => x"19",
          7077 => x"24",
          7078 => x"55",
          7079 => x"51",
          7080 => x"08",
          7081 => x"ff",
          7082 => x"0d",
          7083 => x"75",
          7084 => x"ff",
          7085 => x"30",
          7086 => x"52",
          7087 => x"52",
          7088 => x"39",
          7089 => x"0d",
          7090 => x"05",
          7091 => x"72",
          7092 => x"ff",
          7093 => x"0c",
          7094 => x"73",
          7095 => x"81",
          7096 => x"38",
          7097 => x"2e",
          7098 => x"ff",
          7099 => x"8d",
          7100 => x"70",
          7101 => x"12",
          7102 => x"0c",
          7103 => x"0d",
          7104 => x"96",
          7105 => x"80",
          7106 => x"84",
          7107 => x"71",
          7108 => x"38",
          7109 => x"10",
          7110 => x"ba",
          7111 => x"fb",
          7112 => x"ff",
          7113 => x"ff",
          7114 => x"9f",
          7115 => x"82",
          7116 => x"80",
          7117 => x"53",
          7118 => x"05",
          7119 => x"56",
          7120 => x"70",
          7121 => x"73",
          7122 => x"22",
          7123 => x"79",
          7124 => x"2e",
          7125 => x"8c",
          7126 => x"c4",
          7127 => x"ea",
          7128 => x"05",
          7129 => x"70",
          7130 => x"51",
          7131 => x"ff",
          7132 => x"16",
          7133 => x"e6",
          7134 => x"06",
          7135 => x"83",
          7136 => x"e0",
          7137 => x"51",
          7138 => x"ff",
          7139 => x"73",
          7140 => x"83",
          7141 => x"a6",
          7142 => x"70",
          7143 => x"00",
          7144 => x"ff",
          7145 => x"00",
          7146 => x"00",
          7147 => x"00",
          7148 => x"00",
          7149 => x"00",
          7150 => x"00",
          7151 => x"00",
          7152 => x"00",
          7153 => x"00",
          7154 => x"00",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"00",
          7372 => x"00",
          7373 => x"00",
          7374 => x"00",
          7375 => x"00",
          7376 => x"00",
          7377 => x"00",
          7378 => x"00",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"74",
          7383 => x"74",
          7384 => x"74",
          7385 => x"64",
          7386 => x"63",
          7387 => x"61",
          7388 => x"79",
          7389 => x"66",
          7390 => x"70",
          7391 => x"6d",
          7392 => x"68",
          7393 => x"68",
          7394 => x"63",
          7395 => x"6a",
          7396 => x"61",
          7397 => x"74",
          7398 => x"00",
          7399 => x"00",
          7400 => x"7a",
          7401 => x"69",
          7402 => x"69",
          7403 => x"00",
          7404 => x"55",
          7405 => x"65",
          7406 => x"50",
          7407 => x"72",
          7408 => x"72",
          7409 => x"54",
          7410 => x"20",
          7411 => x"6c",
          7412 => x"49",
          7413 => x"69",
          7414 => x"6f",
          7415 => x"46",
          7416 => x"6c",
          7417 => x"54",
          7418 => x"20",
          7419 => x"6f",
          7420 => x"6c",
          7421 => x"46",
          7422 => x"62",
          7423 => x"4e",
          7424 => x"74",
          7425 => x"6c",
          7426 => x"20",
          7427 => x"6e",
          7428 => x"44",
          7429 => x"20",
          7430 => x"2e",
          7431 => x"65",
          7432 => x"20",
          7433 => x"6c",
          7434 => x"53",
          7435 => x"69",
          7436 => x"65",
          7437 => x"46",
          7438 => x"64",
          7439 => x"6c",
          7440 => x"46",
          7441 => x"65",
          7442 => x"73",
          7443 => x"41",
          7444 => x"65",
          7445 => x"49",
          7446 => x"66",
          7447 => x"2e",
          7448 => x"61",
          7449 => x"64",
          7450 => x"69",
          7451 => x"64",
          7452 => x"20",
          7453 => x"64",
          7454 => x"72",
          7455 => x"6f",
          7456 => x"20",
          7457 => x"53",
          7458 => x"00",
          7459 => x"20",
          7460 => x"73",
          7461 => x"20",
          7462 => x"65",
          7463 => x"72",
          7464 => x"25",
          7465 => x"3a",
          7466 => x"00",
          7467 => x"7c",
          7468 => x"25",
          7469 => x"20",
          7470 => x"00",
          7471 => x"2a",
          7472 => x"31",
          7473 => x"32",
          7474 => x"64",
          7475 => x"2c",
          7476 => x"32",
          7477 => x"73",
          7478 => x"5a",
          7479 => x"72",
          7480 => x"6e",
          7481 => x"55",
          7482 => x"20",
          7483 => x"70",
          7484 => x"31",
          7485 => x"65",
          7486 => x"55",
          7487 => x"20",
          7488 => x"70",
          7489 => x"30",
          7490 => x"65",
          7491 => x"49",
          7492 => x"20",
          7493 => x"70",
          7494 => x"4c",
          7495 => x"65",
          7496 => x"50",
          7497 => x"72",
          7498 => x"54",
          7499 => x"74",
          7500 => x"53",
          7501 => x"75",
          7502 => x"2e",
          7503 => x"6c",
          7504 => x"65",
          7505 => x"61",
          7506 => x"2e",
          7507 => x"7a",
          7508 => x"68",
          7509 => x"65",
          7510 => x"69",
          7511 => x"20",
          7512 => x"20",
          7513 => x"73",
          7514 => x"6d",
          7515 => x"2e",
          7516 => x"25",
          7517 => x"44",
          7518 => x"74",
          7519 => x"00",
          7520 => x"42",
          7521 => x"61",
          7522 => x"5a",
          7523 => x"25",
          7524 => x"73",
          7525 => x"43",
          7526 => x"6f",
          7527 => x"2e",
          7528 => x"61",
          7529 => x"70",
          7530 => x"6f",
          7531 => x"43",
          7532 => x"63",
          7533 => x"30",
          7534 => x"0a",
          7535 => x"20",
          7536 => x"64",
          7537 => x"25",
          7538 => x"45",
          7539 => x"67",
          7540 => x"20",
          7541 => x"2e",
          7542 => x"58",
          7543 => x"00",
          7544 => x"58",
          7545 => x"43",
          7546 => x"67",
          7547 => x"25",
          7548 => x"38",
          7549 => x"6c",
          7550 => x"0a",
          7551 => x"69",
          7552 => x"25",
          7553 => x"32",
          7554 => x"72",
          7555 => x"00",
          7556 => x"20",
          7557 => x"0a",
          7558 => x"65",
          7559 => x"25",
          7560 => x"4d",
          7561 => x"78",
          7562 => x"2c",
          7563 => x"20",
          7564 => x"20",
          7565 => x"2e",
          7566 => x"25",
          7567 => x"20",
          7568 => x"64",
          7569 => x"53",
          7570 => x"69",
          7571 => x"6e",
          7572 => x"76",
          7573 => x"70",
          7574 => x"64",
          7575 => x"65",
          7576 => x"20",
          7577 => x"52",
          7578 => x"63",
          7579 => x"72",
          7580 => x"30",
          7581 => x"20",
          7582 => x"4d",
          7583 => x"74",
          7584 => x"72",
          7585 => x"30",
          7586 => x"20",
          7587 => x"6b",
          7588 => x"41",
          7589 => x"20",
          7590 => x"30",
          7591 => x"4d",
          7592 => x"20",
          7593 => x"49",
          7594 => x"20",
          7595 => x"20",
          7596 => x"30",
          7597 => x"20",
          7598 => x"65",
          7599 => x"20",
          7600 => x"20",
          7601 => x"64",
          7602 => x"7a",
          7603 => x"57",
          7604 => x"20",
          7605 => x"6c",
          7606 => x"71",
          7607 => x"34",
          7608 => x"20",
          7609 => x"4d",
          7610 => x"46",
          7611 => x"20",
          7612 => x"64",
          7613 => x"7a",
          7614 => x"53",
          7615 => x"50",
          7616 => x"49",
          7617 => x"20",
          7618 => x"32",
          7619 => x"57",
          7620 => x"20",
          7621 => x"20",
          7622 => x"20",
          7623 => x"68",
          7624 => x"25",
          7625 => x"20",
          7626 => x"52",
          7627 => x"69",
          7628 => x"25",
          7629 => x"20",
          7630 => x"41",
          7631 => x"65",
          7632 => x"25",
          7633 => x"20",
          7634 => x"20",
          7635 => x"30",
          7636 => x"29",
          7637 => x"42",
          7638 => x"20",
          7639 => x"25",
          7640 => x"20",
          7641 => x"20",
          7642 => x"30",
          7643 => x"29",
          7644 => x"53",
          7645 => x"20",
          7646 => x"25",
          7647 => x"20",
          7648 => x"44",
          7649 => x"30",
          7650 => x"29",
          7651 => x"6f",
          7652 => x"6f",
          7653 => x"55",
          7654 => x"45",
          7655 => x"53",
          7656 => x"4d",
          7657 => x"46",
          7658 => x"45",
          7659 => x"01",
          7660 => x"00",
          7661 => x"00",
          7662 => x"01",
          7663 => x"00",
          7664 => x"00",
          7665 => x"01",
          7666 => x"00",
          7667 => x"00",
          7668 => x"01",
          7669 => x"00",
          7670 => x"00",
          7671 => x"01",
          7672 => x"00",
          7673 => x"00",
          7674 => x"01",
          7675 => x"00",
          7676 => x"00",
          7677 => x"04",
          7678 => x"00",
          7679 => x"00",
          7680 => x"03",
          7681 => x"00",
          7682 => x"00",
          7683 => x"04",
          7684 => x"00",
          7685 => x"00",
          7686 => x"03",
          7687 => x"00",
          7688 => x"00",
          7689 => x"03",
          7690 => x"00",
          7691 => x"00",
          7692 => x"1b",
          7693 => x"1b",
          7694 => x"1b",
          7695 => x"1b",
          7696 => x"1b",
          7697 => x"10",
          7698 => x"0d",
          7699 => x"08",
          7700 => x"05",
          7701 => x"03",
          7702 => x"01",
          7703 => x"6f",
          7704 => x"63",
          7705 => x"69",
          7706 => x"69",
          7707 => x"61",
          7708 => x"68",
          7709 => x"68",
          7710 => x"21",
          7711 => x"75",
          7712 => x"46",
          7713 => x"6f",
          7714 => x"74",
          7715 => x"6f",
          7716 => x"20",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"1b",
          7721 => x"1b",
          7722 => x"7e",
          7723 => x"7e",
          7724 => x"7e",
          7725 => x"7e",
          7726 => x"7e",
          7727 => x"7e",
          7728 => x"7e",
          7729 => x"7e",
          7730 => x"7e",
          7731 => x"7e",
          7732 => x"00",
          7733 => x"00",
          7734 => x"1b",
          7735 => x"1b",
          7736 => x"58",
          7737 => x"25",
          7738 => x"2c",
          7739 => x"00",
          7740 => x"2d",
          7741 => x"63",
          7742 => x"25",
          7743 => x"4b",
          7744 => x"25",
          7745 => x"25",
          7746 => x"52",
          7747 => x"72",
          7748 => x"72",
          7749 => x"30",
          7750 => x"00",
          7751 => x"30",
          7752 => x"00",
          7753 => x"30",
          7754 => x"42",
          7755 => x"2c",
          7756 => x"74",
          7757 => x"65",
          7758 => x"20",
          7759 => x"42",
          7760 => x"2c",
          7761 => x"74",
          7762 => x"65",
          7763 => x"6e",
          7764 => x"53",
          7765 => x"3e",
          7766 => x"2b",
          7767 => x"46",
          7768 => x"32",
          7769 => x"53",
          7770 => x"4e",
          7771 => x"20",
          7772 => x"20",
          7773 => x"41",
          7774 => x"41",
          7775 => x"00",
          7776 => x"00",
          7777 => x"01",
          7778 => x"14",
          7779 => x"80",
          7780 => x"45",
          7781 => x"90",
          7782 => x"59",
          7783 => x"41",
          7784 => x"a8",
          7785 => x"b0",
          7786 => x"b8",
          7787 => x"c0",
          7788 => x"c8",
          7789 => x"d0",
          7790 => x"d8",
          7791 => x"e0",
          7792 => x"e8",
          7793 => x"f0",
          7794 => x"f8",
          7795 => x"2b",
          7796 => x"5c",
          7797 => x"7f",
          7798 => x"00",
          7799 => x"00",
          7800 => x"00",
          7801 => x"00",
          7802 => x"00",
          7803 => x"00",
          7804 => x"00",
          7805 => x"00",
          7806 => x"00",
          7807 => x"00",
          7808 => x"00",
          7809 => x"20",
          7810 => x"00",
          7811 => x"00",
          7812 => x"00",
          7813 => x"00",
          7814 => x"25",
          7815 => x"25",
          7816 => x"25",
          7817 => x"25",
          7818 => x"25",
          7819 => x"25",
          7820 => x"25",
          7821 => x"25",
          7822 => x"25",
          7823 => x"25",
          7824 => x"25",
          7825 => x"25",
          7826 => x"03",
          7827 => x"00",
          7828 => x"03",
          7829 => x"03",
          7830 => x"22",
          7831 => x"00",
          7832 => x"00",
          7833 => x"25",
          7834 => x"00",
          7835 => x"00",
          7836 => x"01",
          7837 => x"01",
          7838 => x"01",
          7839 => x"01",
          7840 => x"01",
          7841 => x"01",
          7842 => x"01",
          7843 => x"01",
          7844 => x"01",
          7845 => x"01",
          7846 => x"01",
          7847 => x"01",
          7848 => x"01",
          7849 => x"01",
          7850 => x"01",
          7851 => x"01",
          7852 => x"01",
          7853 => x"01",
          7854 => x"01",
          7855 => x"01",
          7856 => x"01",
          7857 => x"01",
          7858 => x"01",
          7859 => x"01",
          7860 => x"00",
          7861 => x"01",
          7862 => x"02",
          7863 => x"02",
          7864 => x"02",
          7865 => x"01",
          7866 => x"01",
          7867 => x"02",
          7868 => x"02",
          7869 => x"01",
          7870 => x"02",
          7871 => x"01",
          7872 => x"02",
          7873 => x"02",
          7874 => x"02",
          7875 => x"02",
          7876 => x"02",
          7877 => x"01",
          7878 => x"02",
          7879 => x"01",
          7880 => x"02",
          7881 => x"02",
          7882 => x"00",
          7883 => x"03",
          7884 => x"03",
          7885 => x"03",
          7886 => x"03",
          7887 => x"03",
          7888 => x"01",
          7889 => x"03",
          7890 => x"03",
          7891 => x"03",
          7892 => x"07",
          7893 => x"01",
          7894 => x"00",
          7895 => x"05",
          7896 => x"1d",
          7897 => x"01",
          7898 => x"06",
          7899 => x"06",
          7900 => x"06",
          7901 => x"1f",
          7902 => x"1f",
          7903 => x"1f",
          7904 => x"1f",
          7905 => x"1f",
          7906 => x"1f",
          7907 => x"1f",
          7908 => x"1f",
          7909 => x"1f",
          7910 => x"1f",
          7911 => x"06",
          7912 => x"00",
          7913 => x"1f",
          7914 => x"21",
          7915 => x"21",
          7916 => x"04",
          7917 => x"01",
          7918 => x"01",
          7919 => x"03",
          7920 => x"00",
          7921 => x"00",
          7922 => x"00",
          7923 => x"00",
          7924 => x"00",
          7925 => x"00",
          7926 => x"00",
          7927 => x"00",
          7928 => x"00",
          7929 => x"00",
          7930 => x"00",
          7931 => x"00",
          7932 => x"00",
          7933 => x"00",
          7934 => x"00",
          7935 => x"00",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"00",
          7940 => x"00",
          7941 => x"00",
          7942 => x"00",
          7943 => x"00",
          7944 => x"00",
          7945 => x"00",
          7946 => x"00",
          7947 => x"00",
          7948 => x"00",
          7949 => x"00",
          7950 => x"00",
          7951 => x"00",
          7952 => x"00",
          7953 => x"00",
          7954 => x"00",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"00",
          7959 => x"00",
          7960 => x"00",
          7961 => x"00",
          7962 => x"00",
          7963 => x"00",
          7964 => x"00",
          7965 => x"00",
          7966 => x"00",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"00",
          7980 => x"00",
          7981 => x"01",
          7982 => x"00",
          7983 => x"00",
          7984 => x"05",
          7985 => x"00",
          7986 => x"01",
          7987 => x"01",
          7988 => x"00",
          7989 => x"00",
          7990 => x"00",
          7991 => x"00",
          7992 => x"00",
          7993 => x"00",
          7994 => x"00",
          7995 => x"00",
          7996 => x"00",
          7997 => x"00",
          7998 => x"00",
          7999 => x"00",
          8000 => x"01",
          8001 => x"01",
          8002 => x"02",
          8003 => x"1b",
          8004 => x"79",
          8005 => x"71",
          8006 => x"69",
          8007 => x"61",
          8008 => x"31",
          8009 => x"5c",
          8010 => x"f6",
          8011 => x"08",
          8012 => x"80",
          8013 => x"1b",
          8014 => x"59",
          8015 => x"51",
          8016 => x"49",
          8017 => x"41",
          8018 => x"31",
          8019 => x"5c",
          8020 => x"f6",
          8021 => x"08",
          8022 => x"80",
          8023 => x"1b",
          8024 => x"59",
          8025 => x"51",
          8026 => x"49",
          8027 => x"41",
          8028 => x"21",
          8029 => x"7c",
          8030 => x"f7",
          8031 => x"fb",
          8032 => x"85",
          8033 => x"1b",
          8034 => x"19",
          8035 => x"11",
          8036 => x"09",
          8037 => x"01",
          8038 => x"f0",
          8039 => x"f0",
          8040 => x"f0",
          8041 => x"f0",
          8042 => x"80",
          8043 => x"bf",
          8044 => x"35",
          8045 => x"7c",
          8046 => x"3d",
          8047 => x"46",
          8048 => x"3f",
          8049 => x"d3",
          8050 => x"c6",
          8051 => x"f0",
          8052 => x"80",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"00",
          9069 => x"00",
          9070 => x"00",
          9071 => x"00",
          9072 => x"00",
          9073 => x"00",
          9074 => x"00",
          9075 => x"00",
          9076 => x"00",
          9077 => x"00",
          9078 => x"00",
          9079 => x"00",
          9080 => x"00",
          9081 => x"00",
          9082 => x"00",
          9083 => x"00",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"ce",
          9090 => x"fc",
          9091 => x"c4",
          9092 => x"eb",
          9093 => x"64",
          9094 => x"2f",
          9095 => x"24",
          9096 => x"51",
          9097 => x"04",
          9098 => x"0c",
          9099 => x"14",
          9100 => x"59",
          9101 => x"84",
          9102 => x"8c",
          9103 => x"94",
          9104 => x"80",
          9105 => x"00",
          9106 => x"00",
          9107 => x"00",
          9108 => x"00",
          9109 => x"00",
          9110 => x"00",
          9111 => x"00",
          9112 => x"00",
          9113 => x"00",
          9114 => x"00",
          9115 => x"00",
          9116 => x"00",
          9117 => x"00",
          9118 => x"00",
          9119 => x"00",
          9120 => x"00",
          9121 => x"00",
        others => X"00"
    );

    signal RAM0_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM1_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM2_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM3_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM4_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM5_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM6_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM7_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM0_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM1_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM2_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM3_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM4_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM5_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM6_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM7_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal lowDataA          :     std_logic_vector(WORD_32BIT_RANGE);   -- Low word in 64 bit output from RAM matrix.
    signal highDataA         :     std_logic_vector(WORD_32BIT_RANGE);   -- High word in 64 bit output from RAM matrix.
    signal lowDataB          :     std_logic_vector(WORD_32BIT_RANGE);   -- Low word in 64 bit output from RAM matrix.
    signal highDataB         :     std_logic_vector(WORD_32BIT_RANGE);   -- High word in 64 bit output from RAM matrix.

begin

    -- Correctly assign the Little Endian value to the correct array, byte writes the data is in '7 downto 0', h-word writes
    -- the data is in '15 downto 0', word writes the data is in '31 downto 0'. Long words (64bits) are treated as two words for Endianness,
    -- and not as one continuous long word, this is because the ZPU is 32bit even when accessing a 64bit chunk.
    --
    RAM0_DATA <= memAWrite(7 downto 0)   when memAAddr(2) = '0'
                 else (others => '0');
    RAM1_DATA <= memAWrite(15 downto 8)  when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(15 downto 8)  when memAAddr(2) = '0' and (memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM4_DATA <= memAWrite(7 downto 0)   when memAAddr(2) = '1'
                 else (others => '0');
    RAM5_DATA <= memAWrite(15 downto 8)  when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM6_DATA <= memAWrite(23 downto 16) when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(7 downto 0);
    RAM7_DATA <= memAWrite(31 downto 24) when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(15 downto 8)  when memAAddr(2) = '1' and (memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "011") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "01"))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "010") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "01"))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "001") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "00"))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "000") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "00"))
                 else '0';
    RAM4_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "111") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "11"))
                 else '0';
    RAM5_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "110") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "11"))
                 else '0';
    RAM6_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "101") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "10"))
                 else '0';
    RAM7_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "100") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "10"))
                 else '0';

    memARead  <= lowDataA  when memAAddr(2) = '0'
                 else
                 highDataA;
    memBRead  <= lowDataB & highDataB;

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM0_DATA;
            else
                lowDataA(7 downto 0)    <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM1_DATA;
            else
                lowDataA(15 downto 8)   <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM2_DATA;
            else
                lowDataA(23 downto 16)  <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM3_DATA;
            else
                lowDataA(31 downto 24)  <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 4 - Port A - bits 39 to 32 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM4_WREN = '1' then
                RAM4(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM4_DATA;
            else
                highDataA(7 downto 0)   <= RAM4(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 5 - Port A - bits 47 to 40 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM5_WREN = '1' then
                RAM5(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM5_DATA;
            else
                highDataA(15 downto 8)  <= RAM5(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 6 - Port A - bits 56 to 48
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM6_WREN = '1' then
                RAM6(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM6_DATA;
            else
                highDataA(23 downto 16) <= RAM6(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 7 - Port A - bits 63 to 57 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM7_WREN = '1' then
                RAM7(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM7_DATA;
            else
                highDataA(31 downto 24) <= RAM7(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;


    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(7 downto 0);
                lowDataB(7 downto 0)    <= memBWrite(7 downto 0);
            else
                lowDataB(7 downto 0)    <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(15 downto 8);
                lowDataB(15 downto 8)    <= memBWrite(15 downto 8);
            else
                lowDataB(15 downto 8)    <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(23 downto 16);
                lowDataB(23 downto 16)  <= memBWrite(23 downto 16);
            else
                lowDataB(23 downto 16)  <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(31 downto 24);
                lowDataB(31 downto 24)  <= memBWrite(31 downto 24);
            else
                lowDataB(31 downto 24)  <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 4 - Port B - bits 39 downto 32
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM4(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(39 downto 32);
                highDataB(7 downto 0)   <= memBWrite(39 downto 32);
            else
                highDataB(7 downto 0)   <= RAM4(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 5 - Port B - bits 47 downto 40
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM5(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(47 downto 40);
                highDataB(15 downto 8)  <= memBWrite(47 downto 40);
            else
                highDataB(15 downto 8)  <= RAM5(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 6 - Port B - bits 55 downto 48
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM6(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(55 downto 48);
                highDataB(23 downto 16)  <= memBWrite(55 downto 48);
            else
                highDataB(23 downto 16)  <= RAM6(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 7 - Port B - bits 63 downto 56 
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM7(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(63 downto 56);
                highDataB(31 downto 24)  <= memBWrite(63 downto 56);
            else
                highDataB(31 downto 24)  <= RAM7(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

end arch;
