-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b87fa",
          2049 => x"f80d0b0b",
          2050 => x"0b93e904",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b93",
          2121 => x"cd040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b93b0",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b83be",
          2210 => x"bc738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"93b50400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b0bac",
          2219 => x"cc2d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b0bab",
          2227 => x"ab2d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"96040b0b",
          2317 => x"0b8ca604",
          2318 => x"0b0b0b8c",
          2319 => x"b6040b0b",
          2320 => x"0b8cc604",
          2321 => x"0b0b0b8c",
          2322 => x"d6040b0b",
          2323 => x"0b8ce604",
          2324 => x"0b0b0b8c",
          2325 => x"f6040b0b",
          2326 => x"0b8d8604",
          2327 => x"0b0b0b8d",
          2328 => x"96040b0b",
          2329 => x"0b8da604",
          2330 => x"0b0b0b8d",
          2331 => x"b6040b0b",
          2332 => x"0b8dc604",
          2333 => x"0b0b0b8d",
          2334 => x"d7040b0b",
          2335 => x"0b8de804",
          2336 => x"0b0b0b8d",
          2337 => x"f9040b0b",
          2338 => x"0b8e8a04",
          2339 => x"0b0b0b8e",
          2340 => x"9b040b0b",
          2341 => x"0b8eac04",
          2342 => x"0b0b0b8e",
          2343 => x"bd040b0b",
          2344 => x"0b8ece04",
          2345 => x"0b0b0b8e",
          2346 => x"df040b0b",
          2347 => x"0b8ef004",
          2348 => x"0b0b0b8f",
          2349 => x"81040b0b",
          2350 => x"0b8f9204",
          2351 => x"0b0b0b8f",
          2352 => x"a3040b0b",
          2353 => x"0b8fb404",
          2354 => x"0b0b0b8f",
          2355 => x"c5040b0b",
          2356 => x"0b8fd604",
          2357 => x"0b0b0b8f",
          2358 => x"e7040b0b",
          2359 => x"0b8ff804",
          2360 => x"0b0b0b90",
          2361 => x"89040b0b",
          2362 => x"0b909a04",
          2363 => x"0b0b0b90",
          2364 => x"ab040b0b",
          2365 => x"0b90bc04",
          2366 => x"0b0b0b90",
          2367 => x"cd040b0b",
          2368 => x"0b90de04",
          2369 => x"0b0b0b90",
          2370 => x"ef040b0b",
          2371 => x"0b918004",
          2372 => x"0b0b0b91",
          2373 => x"91040b0b",
          2374 => x"0b91a204",
          2375 => x"0b0b0b91",
          2376 => x"b3040b0b",
          2377 => x"0b91c404",
          2378 => x"0b0b0b91",
          2379 => x"d5040b0b",
          2380 => x"0b91e604",
          2381 => x"0b0b0b91",
          2382 => x"f7040b0b",
          2383 => x"0b928804",
          2384 => x"0b0b0b92",
          2385 => x"99040b0b",
          2386 => x"0b92aa04",
          2387 => x"0b0b0b92",
          2388 => x"bb040b0b",
          2389 => x"0b92cb04",
          2390 => x"0b0b0b92",
          2391 => x"dc040b0b",
          2392 => x"0b92ed04",
          2393 => x"0b0b0b92",
          2394 => x"fe04ffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0484ba98",
          2434 => x"0c80d5f6",
          2435 => x"2d84ba98",
          2436 => x"0880c080",
          2437 => x"900484ba",
          2438 => x"980ca2ee",
          2439 => x"2d84ba98",
          2440 => x"0880c080",
          2441 => x"900484ba",
          2442 => x"980ca0f3",
          2443 => x"2d84ba98",
          2444 => x"0880c080",
          2445 => x"900484ba",
          2446 => x"980ca0e0",
          2447 => x"2d84ba98",
          2448 => x"0880c080",
          2449 => x"900484ba",
          2450 => x"980c94a3",
          2451 => x"2d84ba98",
          2452 => x"0880c080",
          2453 => x"900484ba",
          2454 => x"980ca1f6",
          2455 => x"2d84ba98",
          2456 => x"0880c080",
          2457 => x"900484ba",
          2458 => x"980caf86",
          2459 => x"2d84ba98",
          2460 => x"0880c080",
          2461 => x"900484ba",
          2462 => x"980cad82",
          2463 => x"2d84ba98",
          2464 => x"0880c080",
          2465 => x"900484ba",
          2466 => x"980c9488",
          2467 => x"2d84ba98",
          2468 => x"0880c080",
          2469 => x"900484ba",
          2470 => x"980c95a8",
          2471 => x"2d84ba98",
          2472 => x"0880c080",
          2473 => x"900484ba",
          2474 => x"980c95d1",
          2475 => x"2d84ba98",
          2476 => x"0880c080",
          2477 => x"900484ba",
          2478 => x"980cb18a",
          2479 => x"2d84ba98",
          2480 => x"0880c080",
          2481 => x"900484ba",
          2482 => x"980c80d4",
          2483 => x"db2d84ba",
          2484 => x"980880c0",
          2485 => x"80900484",
          2486 => x"ba980c80",
          2487 => x"d5c02d84",
          2488 => x"ba980880",
          2489 => x"c0809004",
          2490 => x"84ba980c",
          2491 => x"80d2972d",
          2492 => x"84ba9808",
          2493 => x"80c08090",
          2494 => x"0484ba98",
          2495 => x"0c80d3ca",
          2496 => x"2d84ba98",
          2497 => x"0880c080",
          2498 => x"900484ba",
          2499 => x"980c82c9",
          2500 => x"f72d84ba",
          2501 => x"980880c0",
          2502 => x"80900484",
          2503 => x"ba980c82",
          2504 => x"e3c92d84",
          2505 => x"ba980880",
          2506 => x"c0809004",
          2507 => x"84ba980c",
          2508 => x"82d2e72d",
          2509 => x"84ba9808",
          2510 => x"80c08090",
          2511 => x"0484ba98",
          2512 => x"0c82d889",
          2513 => x"2d84ba98",
          2514 => x"0880c080",
          2515 => x"900484ba",
          2516 => x"980c82ed",
          2517 => x"e62d84ba",
          2518 => x"980880c0",
          2519 => x"80900484",
          2520 => x"ba980c82",
          2521 => x"faee2d84",
          2522 => x"ba980880",
          2523 => x"c0809004",
          2524 => x"84ba980c",
          2525 => x"82dfd02d",
          2526 => x"84ba9808",
          2527 => x"80c08090",
          2528 => x"0484ba98",
          2529 => x"0c82f287",
          2530 => x"2d84ba98",
          2531 => x"0880c080",
          2532 => x"900484ba",
          2533 => x"980c82f3",
          2534 => x"d42d84ba",
          2535 => x"980880c0",
          2536 => x"80900484",
          2537 => x"ba980c82",
          2538 => x"f4a92d84",
          2539 => x"ba980880",
          2540 => x"c0809004",
          2541 => x"84ba980c",
          2542 => x"8384eb2d",
          2543 => x"84ba9808",
          2544 => x"80c08090",
          2545 => x"0484ba98",
          2546 => x"0c82ffb0",
          2547 => x"2d84ba98",
          2548 => x"0880c080",
          2549 => x"900484ba",
          2550 => x"980c838b",
          2551 => x"cf2d84ba",
          2552 => x"980880c0",
          2553 => x"80900484",
          2554 => x"ba980c82",
          2555 => x"f6862d84",
          2556 => x"ba980880",
          2557 => x"c0809004",
          2558 => x"84ba980c",
          2559 => x"8394c62d",
          2560 => x"84ba9808",
          2561 => x"80c08090",
          2562 => x"0484ba98",
          2563 => x"0c8395d1",
          2564 => x"2d84ba98",
          2565 => x"0880c080",
          2566 => x"900484ba",
          2567 => x"980c82e6",
          2568 => x"992d84ba",
          2569 => x"980880c0",
          2570 => x"80900484",
          2571 => x"ba980c82",
          2572 => x"e4b02d84",
          2573 => x"ba980880",
          2574 => x"c0809004",
          2575 => x"84ba980c",
          2576 => x"82e7d72d",
          2577 => x"84ba9808",
          2578 => x"80c08090",
          2579 => x"0484ba98",
          2580 => x"0c82f6f0",
          2581 => x"2d84ba98",
          2582 => x"0880c080",
          2583 => x"900484ba",
          2584 => x"980c8396",
          2585 => x"e32d84ba",
          2586 => x"980880c0",
          2587 => x"80900484",
          2588 => x"ba980c83",
          2589 => x"9ac02d84",
          2590 => x"ba980880",
          2591 => x"c0809004",
          2592 => x"84ba980c",
          2593 => x"83a1b22d",
          2594 => x"84ba9808",
          2595 => x"80c08090",
          2596 => x"0484ba98",
          2597 => x"0c82c7c8",
          2598 => x"2d84ba98",
          2599 => x"0880c080",
          2600 => x"900484ba",
          2601 => x"980c83a4",
          2602 => x"db2d84ba",
          2603 => x"980880c0",
          2604 => x"80900484",
          2605 => x"ba980c83",
          2606 => x"b9dc2d84",
          2607 => x"ba980880",
          2608 => x"c0809004",
          2609 => x"84ba980c",
          2610 => x"83b88e2d",
          2611 => x"84ba9808",
          2612 => x"80c08090",
          2613 => x"0484ba98",
          2614 => x"0c81f4ac",
          2615 => x"2d84ba98",
          2616 => x"0880c080",
          2617 => x"900484ba",
          2618 => x"980c81f5",
          2619 => x"ab2d84ba",
          2620 => x"980880c0",
          2621 => x"80900484",
          2622 => x"ba980c81",
          2623 => x"f6aa2d84",
          2624 => x"ba980880",
          2625 => x"c0809004",
          2626 => x"84ba980c",
          2627 => x"80d0992d",
          2628 => x"84ba9808",
          2629 => x"80c08090",
          2630 => x"0484ba98",
          2631 => x"0c80d1e9",
          2632 => x"2d84ba98",
          2633 => x"0880c080",
          2634 => x"900484ba",
          2635 => x"980c80d7",
          2636 => x"942d84ba",
          2637 => x"980880c0",
          2638 => x"80900484",
          2639 => x"ba980cb1",
          2640 => x"9a2d84ba",
          2641 => x"980880c0",
          2642 => x"80900484",
          2643 => x"ba980c81",
          2644 => x"dbca2d84",
          2645 => x"ba980880",
          2646 => x"c0809004",
          2647 => x"84ba980c",
          2648 => x"81dd852d",
          2649 => x"84ba9808",
          2650 => x"80c08090",
          2651 => x"0484ba98",
          2652 => x"0c81f286",
          2653 => x"2d84ba98",
          2654 => x"0880c080",
          2655 => x"900484ba",
          2656 => x"980c81d5",
          2657 => x"da2d84ba",
          2658 => x"980880c0",
          2659 => x"8090043c",
          2660 => x"04101010",
          2661 => x"10101010",
          2662 => x"10101010",
          2663 => x"10101010",
          2664 => x"10101010",
          2665 => x"10101010",
          2666 => x"10101010",
          2667 => x"10101010",
          2668 => x"53510400",
          2669 => x"007381ff",
          2670 => x"06738306",
          2671 => x"09810583",
          2672 => x"05101010",
          2673 => x"2b0772fc",
          2674 => x"060c5151",
          2675 => x"04727280",
          2676 => x"728106ff",
          2677 => x"05097206",
          2678 => x"05711052",
          2679 => x"720a100a",
          2680 => x"5372ed38",
          2681 => x"51515351",
          2682 => x"0484ba8c",
          2683 => x"7084d5f8",
          2684 => x"278e3880",
          2685 => x"71708405",
          2686 => x"530c0b0b",
          2687 => x"0b93ec04",
          2688 => x"8c815180",
          2689 => x"cec40400",
          2690 => x"fc3d0d87",
          2691 => x"3d707084",
          2692 => x"05520856",
          2693 => x"53745284",
          2694 => x"d5f00851",
          2695 => x"81c53f86",
          2696 => x"3d0d04fa",
          2697 => x"3d0d787a",
          2698 => x"7c851133",
          2699 => x"81328106",
          2700 => x"80732507",
          2701 => x"56585557",
          2702 => x"80527272",
          2703 => x"2e098106",
          2704 => x"80d338ff",
          2705 => x"1477748a",
          2706 => x"32703070",
          2707 => x"72079f2a",
          2708 => x"51555556",
          2709 => x"54807425",
          2710 => x"b7387180",
          2711 => x"2eb23875",
          2712 => x"518efa3f",
          2713 => x"84ba8c08",
          2714 => x"5384ba8c",
          2715 => x"08ff2eae",
          2716 => x"3884ba8c",
          2717 => x"08757081",
          2718 => x"055734ff",
          2719 => x"14738a32",
          2720 => x"70307072",
          2721 => x"079f2a51",
          2722 => x"54545473",
          2723 => x"8024cb38",
          2724 => x"80753476",
          2725 => x"527184ba",
          2726 => x"8c0c883d",
          2727 => x"0d04800b",
          2728 => x"84ba8c0c",
          2729 => x"883d0d04",
          2730 => x"f53d0d7d",
          2731 => x"54860284",
          2732 => x"05990534",
          2733 => x"7356fe0a",
          2734 => x"588e3d88",
          2735 => x"05537e52",
          2736 => x"8d3de405",
          2737 => x"519d3f73",
          2738 => x"19548074",
          2739 => x"348d3d0d",
          2740 => x"04fd3d0d",
          2741 => x"863d8805",
          2742 => x"53765275",
          2743 => x"51853f85",
          2744 => x"3d0d04f1",
          2745 => x"3d0d6163",
          2746 => x"65425d5d",
          2747 => x"80708c1f",
          2748 => x"0c851e33",
          2749 => x"70812a81",
          2750 => x"32810655",
          2751 => x"555bff54",
          2752 => x"727b2e09",
          2753 => x"810680d2",
          2754 => x"387b3357",
          2755 => x"767b2e80",
          2756 => x"c538811c",
          2757 => x"7b810654",
          2758 => x"5c72802e",
          2759 => x"818138d0",
          2760 => x"175f7e89",
          2761 => x"2681a338",
          2762 => x"76b03270",
          2763 => x"30708025",
          2764 => x"51545578",
          2765 => x"ae387280",
          2766 => x"2ea9387a",
          2767 => x"832a7081",
          2768 => x"32810640",
          2769 => x"547e802e",
          2770 => x"9e387a82",
          2771 => x"80075b7b",
          2772 => x"335776ff",
          2773 => x"bd388c1d",
          2774 => x"08547384",
          2775 => x"ba8c0c91",
          2776 => x"3d0d047a",
          2777 => x"832a5478",
          2778 => x"10101079",
          2779 => x"10057098",
          2780 => x"2b70982c",
          2781 => x"19708180",
          2782 => x"0a298b0a",
          2783 => x"0570982c",
          2784 => x"525a5b56",
          2785 => x"5f807924",
          2786 => x"81863873",
          2787 => x"81065372",
          2788 => x"ffbd3878",
          2789 => x"7c335858",
          2790 => x"76fef738",
          2791 => x"ffb83976",
          2792 => x"a52e0981",
          2793 => x"06933881",
          2794 => x"73745a5a",
          2795 => x"5b8a7c33",
          2796 => x"585a76fe",
          2797 => x"dd38ff9e",
          2798 => x"397c5276",
          2799 => x"518baf3f",
          2800 => x"7b335776",
          2801 => x"fecc38ff",
          2802 => x"8d397a83",
          2803 => x"2a708106",
          2804 => x"5455788a",
          2805 => x"38817074",
          2806 => x"0640547e",
          2807 => x"9538e017",
          2808 => x"537280d8",
          2809 => x"26973872",
          2810 => x"101083ca",
          2811 => x"cc055473",
          2812 => x"080473e0",
          2813 => x"18545980",
          2814 => x"d87327eb",
          2815 => x"387c5276",
          2816 => x"518aeb3f",
          2817 => x"807c3358",
          2818 => x"5b76fe86",
          2819 => x"38fec739",
          2820 => x"80ff59fe",
          2821 => x"f639885a",
          2822 => x"7f608405",
          2823 => x"71087d83",
          2824 => x"ffcf065e",
          2825 => x"58415484",
          2826 => x"ba9c5e79",
          2827 => x"52755193",
          2828 => x"9a3f84ba",
          2829 => x"8c0881ff",
          2830 => x"0684ba8c",
          2831 => x"0818df05",
          2832 => x"56537289",
          2833 => x"26883884",
          2834 => x"ba8c08b0",
          2835 => x"0555747e",
          2836 => x"70810540",
          2837 => x"34795275",
          2838 => x"5190ca3f",
          2839 => x"84ba8c08",
          2840 => x"5684ba8c",
          2841 => x"08c5387d",
          2842 => x"84ba9c31",
          2843 => x"982b7bb2",
          2844 => x"0640567e",
          2845 => x"802e8f38",
          2846 => x"77848080",
          2847 => x"29fc8080",
          2848 => x"0570902c",
          2849 => x"59557a86",
          2850 => x"2a708106",
          2851 => x"555f7380",
          2852 => x"2e9e3877",
          2853 => x"84808029",
          2854 => x"f8808005",
          2855 => x"5379902e",
          2856 => x"8b387784",
          2857 => x"808029fc",
          2858 => x"80800553",
          2859 => x"72902c58",
          2860 => x"7a832a70",
          2861 => x"81065455",
          2862 => x"72802e9e",
          2863 => x"3875982c",
          2864 => x"7081ff06",
          2865 => x"54547873",
          2866 => x"2486cc38",
          2867 => x"7a83fff7",
          2868 => x"0670832a",
          2869 => x"71862a41",
          2870 => x"565b7481",
          2871 => x"06547380",
          2872 => x"2e85f038",
          2873 => x"77793190",
          2874 => x"2b70902c",
          2875 => x"7c838006",
          2876 => x"56595373",
          2877 => x"802e8596",
          2878 => x"387a812a",
          2879 => x"81065473",
          2880 => x"85eb387a",
          2881 => x"842a8106",
          2882 => x"54738698",
          2883 => x"387a852a",
          2884 => x"81065473",
          2885 => x"8697387e",
          2886 => x"81065473",
          2887 => x"858f387a",
          2888 => x"882a8106",
          2889 => x"5f7e802e",
          2890 => x"b2387778",
          2891 => x"84808029",
          2892 => x"fc808005",
          2893 => x"70902c5a",
          2894 => x"40548074",
          2895 => x"259d387c",
          2896 => x"52b05188",
          2897 => x"a93f7778",
          2898 => x"84808029",
          2899 => x"fc808005",
          2900 => x"70902c5a",
          2901 => x"40547380",
          2902 => x"24e53874",
          2903 => x"81065372",
          2904 => x"802eb238",
          2905 => x"78798180",
          2906 => x"0a2981ff",
          2907 => x"0a057098",
          2908 => x"2c5b5555",
          2909 => x"8075259d",
          2910 => x"387c52b0",
          2911 => x"5187ef3f",
          2912 => x"78798180",
          2913 => x"0a2981ff",
          2914 => x"0a057098",
          2915 => x"2c5b5555",
          2916 => x"748024e5",
          2917 => x"387a872a",
          2918 => x"7081065c",
          2919 => x"557a802e",
          2920 => x"81b93876",
          2921 => x"80e32e84",
          2922 => x"d8387680",
          2923 => x"f32e81ca",
          2924 => x"387680d3",
          2925 => x"2e81e238",
          2926 => x"7d84ba9c",
          2927 => x"2e96387c",
          2928 => x"52ff1e70",
          2929 => x"33525e87",
          2930 => x"a53f7d84",
          2931 => x"ba9c2e09",
          2932 => x"8106ec38",
          2933 => x"7481065b",
          2934 => x"7a802efc",
          2935 => x"a7387778",
          2936 => x"84808029",
          2937 => x"fc808005",
          2938 => x"70902c5a",
          2939 => x"40558075",
          2940 => x"25fc9138",
          2941 => x"7c52a051",
          2942 => x"86f43fe2",
          2943 => x"397a9007",
          2944 => x"5b7aa007",
          2945 => x"7c33585b",
          2946 => x"76fa8738",
          2947 => x"fac8397a",
          2948 => x"80c0075b",
          2949 => x"80f85790",
          2950 => x"60618405",
          2951 => x"71087e83",
          2952 => x"ffcf065f",
          2953 => x"5942555a",
          2954 => x"fbfd397f",
          2955 => x"60840577",
          2956 => x"fe800a06",
          2957 => x"83133370",
          2958 => x"982b7207",
          2959 => x"7c848080",
          2960 => x"29fc8080",
          2961 => x"0570902c",
          2962 => x"5e525a56",
          2963 => x"57415f7a",
          2964 => x"872a7081",
          2965 => x"065c557a",
          2966 => x"fec93877",
          2967 => x"78848080",
          2968 => x"29fc8080",
          2969 => x"0570902c",
          2970 => x"5a545f80",
          2971 => x"7f25feb3",
          2972 => x"387c52a0",
          2973 => x"5185f73f",
          2974 => x"e239ff1a",
          2975 => x"7083ffff",
          2976 => x"065b5779",
          2977 => x"83ffff2e",
          2978 => x"feca387c",
          2979 => x"52757081",
          2980 => x"05573351",
          2981 => x"85d83fe2",
          2982 => x"39ff1a70",
          2983 => x"83ffff06",
          2984 => x"5b547983",
          2985 => x"ffff2efe",
          2986 => x"ab387c52",
          2987 => x"75708105",
          2988 => x"57335185",
          2989 => x"b93fe239",
          2990 => x"75fc0a06",
          2991 => x"81fc0a07",
          2992 => x"78848080",
          2993 => x"29fc8080",
          2994 => x"0570902c",
          2995 => x"5a585680",
          2996 => x"e37b872a",
          2997 => x"7081065d",
          2998 => x"56577afd",
          2999 => x"c638fefb",
          3000 => x"397f6084",
          3001 => x"05710870",
          3002 => x"53404156",
          3003 => x"807e2482",
          3004 => x"df387a83",
          3005 => x"ffbf065b",
          3006 => x"84ba9c5e",
          3007 => x"faad397a",
          3008 => x"84077c33",
          3009 => x"585b76f8",
          3010 => x"8938f8ca",
          3011 => x"397a8807",
          3012 => x"5b807c33",
          3013 => x"585976f7",
          3014 => x"f938f8ba",
          3015 => x"397f6084",
          3016 => x"05710877",
          3017 => x"81065658",
          3018 => x"415f7282",
          3019 => x"8a387551",
          3020 => x"87f63f84",
          3021 => x"ba8c0883",
          3022 => x"ffff0678",
          3023 => x"7131902b",
          3024 => x"545a7290",
          3025 => x"2c58fe87",
          3026 => x"397a80c0",
          3027 => x"077c3358",
          3028 => x"5b76f7be",
          3029 => x"38f7ff39",
          3030 => x"7f608405",
          3031 => x"71087781",
          3032 => x"065d5841",
          3033 => x"547981cf",
          3034 => x"38755187",
          3035 => x"bb3f84ba",
          3036 => x"8c0883ff",
          3037 => x"ff067871",
          3038 => x"31902b54",
          3039 => x"5ac4397a",
          3040 => x"8180077c",
          3041 => x"33585b76",
          3042 => x"f78838f7",
          3043 => x"c9397778",
          3044 => x"84808029",
          3045 => x"fc808005",
          3046 => x"70902c5a",
          3047 => x"54548074",
          3048 => x"25fad638",
          3049 => x"7c52a051",
          3050 => x"83c43fe2",
          3051 => x"397c52b0",
          3052 => x"5183bb3f",
          3053 => x"79902e09",
          3054 => x"8106fae3",
          3055 => x"387c5276",
          3056 => x"5183ab3f",
          3057 => x"7a882a81",
          3058 => x"065f7e80",
          3059 => x"2efb8c38",
          3060 => x"fad83975",
          3061 => x"982c7871",
          3062 => x"31902b70",
          3063 => x"902c7d83",
          3064 => x"8006575a",
          3065 => x"515373fa",
          3066 => x"9038ffa2",
          3067 => x"397c52ad",
          3068 => x"5182fb3f",
          3069 => x"7e810654",
          3070 => x"73802efa",
          3071 => x"a238ffad",
          3072 => x"397c5275",
          3073 => x"982a5182",
          3074 => x"e53f7481",
          3075 => x"065b7a80",
          3076 => x"2ef7f138",
          3077 => x"fbc83978",
          3078 => x"7431982b",
          3079 => x"70982c5a",
          3080 => x"53f9b739",
          3081 => x"7c52ab51",
          3082 => x"82c43fc8",
          3083 => x"397c52a0",
          3084 => x"5182bb3f",
          3085 => x"ffbe3978",
          3086 => x"52755188",
          3087 => x"8b3f84ba",
          3088 => x"8c0883ff",
          3089 => x"ff067871",
          3090 => x"31902b54",
          3091 => x"5afdf339",
          3092 => x"7a82077e",
          3093 => x"307183ff",
          3094 => x"bf065257",
          3095 => x"5bfd9939",
          3096 => x"fe3d0d84",
          3097 => x"d5ec0853",
          3098 => x"75527451",
          3099 => x"f3b53f84",
          3100 => x"3d0d04fa",
          3101 => x"3d0d7855",
          3102 => x"800b84d5",
          3103 => x"f0088511",
          3104 => x"3370812a",
          3105 => x"81327081",
          3106 => x"06515658",
          3107 => x"5557ff56",
          3108 => x"72772e09",
          3109 => x"810680d5",
          3110 => x"38747081",
          3111 => x"05563353",
          3112 => x"72772eb0",
          3113 => x"3884d5f0",
          3114 => x"08527251",
          3115 => x"90140853",
          3116 => x"722d84ba",
          3117 => x"8c08802e",
          3118 => x"8338ff57",
          3119 => x"74708105",
          3120 => x"56335372",
          3121 => x"802e8838",
          3122 => x"84d5f008",
          3123 => x"54d73984",
          3124 => x"d5f00854",
          3125 => x"84d5f008",
          3126 => x"528a5190",
          3127 => x"14085574",
          3128 => x"2d84ba8c",
          3129 => x"08802e83",
          3130 => x"38ff5776",
          3131 => x"567584ba",
          3132 => x"8c0c883d",
          3133 => x"0d04fa3d",
          3134 => x"0d787a56",
          3135 => x"54800b85",
          3136 => x"16337081",
          3137 => x"2a813270",
          3138 => x"81065155",
          3139 => x"5757ff56",
          3140 => x"72772e09",
          3141 => x"81069238",
          3142 => x"73708105",
          3143 => x"55335372",
          3144 => x"772e0981",
          3145 => x"06983876",
          3146 => x"567584ba",
          3147 => x"8c0c883d",
          3148 => x"0d047370",
          3149 => x"81055533",
          3150 => x"5372802e",
          3151 => x"ea387452",
          3152 => x"72519015",
          3153 => x"0853722d",
          3154 => x"84ba8c08",
          3155 => x"802ee338",
          3156 => x"ff747081",
          3157 => x"05563354",
          3158 => x"5772e338",
          3159 => x"ca39ff3d",
          3160 => x"0d84d5f0",
          3161 => x"08527351",
          3162 => x"853f833d",
          3163 => x"0d04fa3d",
          3164 => x"0d787a85",
          3165 => x"11337081",
          3166 => x"2a813281",
          3167 => x"06565656",
          3168 => x"57ff5672",
          3169 => x"ae387382",
          3170 => x"2a810654",
          3171 => x"73802eac",
          3172 => x"388c1508",
          3173 => x"53728816",
          3174 => x"08259138",
          3175 => x"74085676",
          3176 => x"76347408",
          3177 => x"8105750c",
          3178 => x"8c150853",
          3179 => x"81138c16",
          3180 => x"0c765675",
          3181 => x"84ba8c0c",
          3182 => x"883d0d04",
          3183 => x"74527681",
          3184 => x"ff065190",
          3185 => x"15085473",
          3186 => x"2dff5684",
          3187 => x"ba8c08e3",
          3188 => x"388c1508",
          3189 => x"81058c16",
          3190 => x"0c7656d7",
          3191 => x"39fb3d0d",
          3192 => x"77851133",
          3193 => x"7081ff06",
          3194 => x"70813281",
          3195 => x"06555556",
          3196 => x"56ff5471",
          3197 => x"b3387286",
          3198 => x"2a810652",
          3199 => x"71b33872",
          3200 => x"822a8106",
          3201 => x"5271802e",
          3202 => x"80c33875",
          3203 => x"08703353",
          3204 => x"5371802e",
          3205 => x"80f03881",
          3206 => x"13760c8c",
          3207 => x"16088105",
          3208 => x"8c170c71",
          3209 => x"81ff0654",
          3210 => x"7384ba8c",
          3211 => x"0c873d0d",
          3212 => x"0474ffbf",
          3213 => x"06537285",
          3214 => x"17348c16",
          3215 => x"0881058c",
          3216 => x"170c8416",
          3217 => x"3384ba8c",
          3218 => x"0c873d0d",
          3219 => x"04755194",
          3220 => x"16085574",
          3221 => x"2d84ba8c",
          3222 => x"085284ba",
          3223 => x"8c088025",
          3224 => x"ffb93885",
          3225 => x"16337090",
          3226 => x"07545284",
          3227 => x"ba8c08ff",
          3228 => x"2e853871",
          3229 => x"a0075372",
          3230 => x"851734ff",
          3231 => x"547384ba",
          3232 => x"8c0c873d",
          3233 => x"0d0474a0",
          3234 => x"07537285",
          3235 => x"1734ff54",
          3236 => x"ec39fd3d",
          3237 => x"0d757771",
          3238 => x"54545471",
          3239 => x"70810553",
          3240 => x"335170f7",
          3241 => x"38ff1252",
          3242 => x"72708105",
          3243 => x"54335170",
          3244 => x"72708105",
          3245 => x"543470f0",
          3246 => x"387384ba",
          3247 => x"8c0c853d",
          3248 => x"0d04fc3d",
          3249 => x"0d767971",
          3250 => x"7a555552",
          3251 => x"5470802e",
          3252 => x"9d387372",
          3253 => x"27a13870",
          3254 => x"802e9338",
          3255 => x"71708105",
          3256 => x"53337370",
          3257 => x"81055534",
          3258 => x"ff115170",
          3259 => x"ef387384",
          3260 => x"ba8c0c86",
          3261 => x"3d0d0470",
          3262 => x"12557375",
          3263 => x"27d93870",
          3264 => x"14755353",
          3265 => x"ff13ff13",
          3266 => x"53537133",
          3267 => x"7334ff11",
          3268 => x"5170802e",
          3269 => x"d938ff13",
          3270 => x"ff135353",
          3271 => x"71337334",
          3272 => x"ff115170",
          3273 => x"df38c739",
          3274 => x"fe3d0d74",
          3275 => x"70535371",
          3276 => x"70810553",
          3277 => x"335170f7",
          3278 => x"38ff1270",
          3279 => x"743184ba",
          3280 => x"8c0c5184",
          3281 => x"3d0d04fd",
          3282 => x"3d0d7577",
          3283 => x"71545454",
          3284 => x"72708105",
          3285 => x"54335170",
          3286 => x"72708105",
          3287 => x"543470f0",
          3288 => x"387384ba",
          3289 => x"8c0c853d",
          3290 => x"0d04fd3d",
          3291 => x"0d757871",
          3292 => x"79555552",
          3293 => x"5470802e",
          3294 => x"93387170",
          3295 => x"81055333",
          3296 => x"73708105",
          3297 => x"5534ff11",
          3298 => x"5170ef38",
          3299 => x"7384ba8c",
          3300 => x"0c853d0d",
          3301 => x"04fc3d0d",
          3302 => x"76787a55",
          3303 => x"56547280",
          3304 => x"2ea13873",
          3305 => x"33757081",
          3306 => x"05573352",
          3307 => x"5271712e",
          3308 => x"0981069a",
          3309 => x"38811454",
          3310 => x"71802eb7",
          3311 => x"38ff1353",
          3312 => x"72e13880",
          3313 => x"517084ba",
          3314 => x"8c0c863d",
          3315 => x"0d047280",
          3316 => x"2ef13873",
          3317 => x"3353ff51",
          3318 => x"72802ee9",
          3319 => x"38ff1533",
          3320 => x"52815171",
          3321 => x"802ede38",
          3322 => x"72723184",
          3323 => x"ba8c0c86",
          3324 => x"3d0d0471",
          3325 => x"84ba8c0c",
          3326 => x"863d0d04",
          3327 => x"fb3d0d77",
          3328 => x"79537052",
          3329 => x"5680c13f",
          3330 => x"84ba8c08",
          3331 => x"84ba8c08",
          3332 => x"81055255",
          3333 => x"81b3b33f",
          3334 => x"84ba8c08",
          3335 => x"5484ba8c",
          3336 => x"08802e9b",
          3337 => x"3884ba8c",
          3338 => x"08155480",
          3339 => x"74347453",
          3340 => x"755284ba",
          3341 => x"8c0851fe",
          3342 => x"b13f84ba",
          3343 => x"8c085473",
          3344 => x"84ba8c0c",
          3345 => x"873d0d04",
          3346 => x"fd3d0d75",
          3347 => x"77717154",
          3348 => x"55535471",
          3349 => x"802e9f38",
          3350 => x"72708105",
          3351 => x"54335170",
          3352 => x"802e8c38",
          3353 => x"ff125271",
          3354 => x"ff2e0981",
          3355 => x"06ea38ff",
          3356 => x"13707531",
          3357 => x"52527084",
          3358 => x"ba8c0c85",
          3359 => x"3d0d04fd",
          3360 => x"3d0d7577",
          3361 => x"79725553",
          3362 => x"54547080",
          3363 => x"2e8e3872",
          3364 => x"72708105",
          3365 => x"5434ff11",
          3366 => x"5170f438",
          3367 => x"7384ba8c",
          3368 => x"0c853d0d",
          3369 => x"04fa3d0d",
          3370 => x"787a5854",
          3371 => x"a0527680",
          3372 => x"2e8b3876",
          3373 => x"5180f53f",
          3374 => x"84ba8c08",
          3375 => x"52e01253",
          3376 => x"73802e8d",
          3377 => x"38735180",
          3378 => x"e33f7184",
          3379 => x"ba8c0831",
          3380 => x"53805272",
          3381 => x"9f2680cb",
          3382 => x"38735272",
          3383 => x"9f2e80c3",
          3384 => x"38811374",
          3385 => x"712aa072",
          3386 => x"3176712b",
          3387 => x"57545455",
          3388 => x"80567476",
          3389 => x"2ea83872",
          3390 => x"10749f2a",
          3391 => x"07741077",
          3392 => x"07787231",
          3393 => x"ff119f2c",
          3394 => x"7081067b",
          3395 => x"72067571",
          3396 => x"31ff1c5c",
          3397 => x"56525255",
          3398 => x"58555374",
          3399 => x"da387310",
          3400 => x"76075271",
          3401 => x"84ba8c0c",
          3402 => x"883d0d04",
          3403 => x"fc3d0d76",
          3404 => x"70fc8080",
          3405 => x"06703070",
          3406 => x"72078025",
          3407 => x"70842b90",
          3408 => x"71317571",
          3409 => x"2a7083fe",
          3410 => x"80067030",
          3411 => x"70802583",
          3412 => x"2b887131",
          3413 => x"74712a70",
          3414 => x"81f00670",
          3415 => x"30708025",
          3416 => x"822b8471",
          3417 => x"3174712a",
          3418 => x"5553751b",
          3419 => x"05738c06",
          3420 => x"70307080",
          3421 => x"25108271",
          3422 => x"3177712a",
          3423 => x"70812a81",
          3424 => x"32708106",
          3425 => x"70308274",
          3426 => x"31067519",
          3427 => x"0584ba8c",
          3428 => x"0c515254",
          3429 => x"55515456",
          3430 => x"5a535555",
          3431 => x"55515656",
          3432 => x"56565158",
          3433 => x"56545286",
          3434 => x"3d0d04fd",
          3435 => x"3d0d7577",
          3436 => x"70547153",
          3437 => x"54548194",
          3438 => x"3f84ba8c",
          3439 => x"08732974",
          3440 => x"713184ba",
          3441 => x"8c0c5385",
          3442 => x"3d0d04fa",
          3443 => x"3d0d787a",
          3444 => x"5854a053",
          3445 => x"76802e8b",
          3446 => x"387651fe",
          3447 => x"cf3f84ba",
          3448 => x"8c0853e0",
          3449 => x"13527380",
          3450 => x"2e8d3873",
          3451 => x"51febd3f",
          3452 => x"7284ba8c",
          3453 => x"08315273",
          3454 => x"53719f26",
          3455 => x"80c53880",
          3456 => x"53719f2e",
          3457 => x"be388112",
          3458 => x"74712aa0",
          3459 => x"72317671",
          3460 => x"2b575454",
          3461 => x"55805674",
          3462 => x"762ea838",
          3463 => x"7210749f",
          3464 => x"2a077410",
          3465 => x"77077872",
          3466 => x"31ff119f",
          3467 => x"2c708106",
          3468 => x"7b720675",
          3469 => x"7131ff1c",
          3470 => x"5c565252",
          3471 => x"55585553",
          3472 => x"74da3872",
          3473 => x"84ba8c0c",
          3474 => x"883d0d04",
          3475 => x"fa3d0d78",
          3476 => x"9f2c7a9f",
          3477 => x"2c7a9f2c",
          3478 => x"7b327c9f",
          3479 => x"2c7d3273",
          3480 => x"73327174",
          3481 => x"31577275",
          3482 => x"31565956",
          3483 => x"595556fc",
          3484 => x"b43f84ba",
          3485 => x"8c087532",
          3486 => x"753184ba",
          3487 => x"8c0c883d",
          3488 => x"0d04f73d",
          3489 => x"0d7b7d5b",
          3490 => x"5780707b",
          3491 => x"0c770870",
          3492 => x"33565659",
          3493 => x"73a02e09",
          3494 => x"81068f38",
          3495 => x"81157078",
          3496 => x"0c703355",
          3497 => x"5573a02e",
          3498 => x"f33873ad",
          3499 => x"2e80f538",
          3500 => x"73b02e81",
          3501 => x"8338d014",
          3502 => x"58805677",
          3503 => x"892680db",
          3504 => x"388a5880",
          3505 => x"56a07427",
          3506 => x"80c43880",
          3507 => x"e0742789",
          3508 => x"38e01470",
          3509 => x"81ff0655",
          3510 => x"53d01470",
          3511 => x"81ff0651",
          3512 => x"53907327",
          3513 => x"8f38f913",
          3514 => x"7081ff06",
          3515 => x"54548973",
          3516 => x"27818938",
          3517 => x"72782781",
          3518 => x"83387776",
          3519 => x"29138116",
          3520 => x"70790c70",
          3521 => x"33565656",
          3522 => x"73a026ff",
          3523 => x"be387880",
          3524 => x"2e843875",
          3525 => x"3056757a",
          3526 => x"0c815675",
          3527 => x"84ba8c0c",
          3528 => x"8b3d0d04",
          3529 => x"81701670",
          3530 => x"790c7033",
          3531 => x"56565973",
          3532 => x"b02e0981",
          3533 => x"06feff38",
          3534 => x"81157078",
          3535 => x"0c703355",
          3536 => x"557380e2",
          3537 => x"2ea63890",
          3538 => x"587380f8",
          3539 => x"2ea03881",
          3540 => x"56a07427",
          3541 => x"c638d014",
          3542 => x"53805688",
          3543 => x"58897327",
          3544 => x"fee13875",
          3545 => x"84ba8c0c",
          3546 => x"8b3d0d04",
          3547 => x"82588115",
          3548 => x"70780c70",
          3549 => x"33555580",
          3550 => x"56feca39",
          3551 => x"800b84ba",
          3552 => x"8c0c8b3d",
          3553 => x"0d04f73d",
          3554 => x"0d7b7d5b",
          3555 => x"5780707b",
          3556 => x"0c770870",
          3557 => x"33565659",
          3558 => x"73a02e09",
          3559 => x"81068f38",
          3560 => x"81157078",
          3561 => x"0c703355",
          3562 => x"5573a02e",
          3563 => x"f33873ad",
          3564 => x"2e80f538",
          3565 => x"73b02e81",
          3566 => x"8338d014",
          3567 => x"58805677",
          3568 => x"892680db",
          3569 => x"388a5880",
          3570 => x"56a07427",
          3571 => x"80c43880",
          3572 => x"e0742789",
          3573 => x"38e01470",
          3574 => x"81ff0655",
          3575 => x"53d01470",
          3576 => x"81ff0651",
          3577 => x"53907327",
          3578 => x"8f38f913",
          3579 => x"7081ff06",
          3580 => x"54548973",
          3581 => x"27818938",
          3582 => x"72782781",
          3583 => x"83387776",
          3584 => x"29138116",
          3585 => x"70790c70",
          3586 => x"33565656",
          3587 => x"73a026ff",
          3588 => x"be387880",
          3589 => x"2e843875",
          3590 => x"3056757a",
          3591 => x"0c815675",
          3592 => x"84ba8c0c",
          3593 => x"8b3d0d04",
          3594 => x"81701670",
          3595 => x"790c7033",
          3596 => x"56565973",
          3597 => x"b02e0981",
          3598 => x"06feff38",
          3599 => x"81157078",
          3600 => x"0c703355",
          3601 => x"557380e2",
          3602 => x"2ea63890",
          3603 => x"587380f8",
          3604 => x"2ea03881",
          3605 => x"56a07427",
          3606 => x"c638d014",
          3607 => x"53805688",
          3608 => x"58897327",
          3609 => x"fee13875",
          3610 => x"84ba8c0c",
          3611 => x"8b3d0d04",
          3612 => x"82588115",
          3613 => x"70780c70",
          3614 => x"33555580",
          3615 => x"56feca39",
          3616 => x"800b84ba",
          3617 => x"8c0c8b3d",
          3618 => x"0d0480d6",
          3619 => x"dc3f84ba",
          3620 => x"8c0881ff",
          3621 => x"0684ba8c",
          3622 => x"0c04ff3d",
          3623 => x"0d735271",
          3624 => x"93268c38",
          3625 => x"71101083",
          3626 => x"becc0552",
          3627 => x"71080483",
          3628 => x"cee451ef",
          3629 => x"be3f833d",
          3630 => x"0d0483ce",
          3631 => x"f451efb3",
          3632 => x"3f833d0d",
          3633 => x"0483cf8c",
          3634 => x"51efa83f",
          3635 => x"833d0d04",
          3636 => x"83cfa451",
          3637 => x"ef9d3f83",
          3638 => x"3d0d0483",
          3639 => x"cfbc51ef",
          3640 => x"923f833d",
          3641 => x"0d0483cf",
          3642 => x"cc51ef87",
          3643 => x"3f833d0d",
          3644 => x"0483cfec",
          3645 => x"51eefc3f",
          3646 => x"833d0d04",
          3647 => x"83cffc51",
          3648 => x"eef13f83",
          3649 => x"3d0d0483",
          3650 => x"d0a451ee",
          3651 => x"e63f833d",
          3652 => x"0d0483d0",
          3653 => x"b851eedb",
          3654 => x"3f833d0d",
          3655 => x"0483d0d4",
          3656 => x"51eed03f",
          3657 => x"833d0d04",
          3658 => x"83d0ec51",
          3659 => x"eec53f83",
          3660 => x"3d0d0483",
          3661 => x"d18451ee",
          3662 => x"ba3f833d",
          3663 => x"0d0483d1",
          3664 => x"9c51eeaf",
          3665 => x"3f833d0d",
          3666 => x"0483d1ac",
          3667 => x"51eea43f",
          3668 => x"833d0d04",
          3669 => x"83d1c051",
          3670 => x"ee993f83",
          3671 => x"3d0d0483",
          3672 => x"d1d051ee",
          3673 => x"8e3f833d",
          3674 => x"0d0483d1",
          3675 => x"e051ee83",
          3676 => x"3f833d0d",
          3677 => x"0483d1f0",
          3678 => x"51edf83f",
          3679 => x"833d0d04",
          3680 => x"83d28051",
          3681 => x"eded3f83",
          3682 => x"3d0d0483",
          3683 => x"d28c51ed",
          3684 => x"e23f833d",
          3685 => x"0d04ec3d",
          3686 => x"0d660284",
          3687 => x"0580e305",
          3688 => x"335b5880",
          3689 => x"68793070",
          3690 => x"7b077325",
          3691 => x"51575759",
          3692 => x"78577587",
          3693 => x"ff268338",
          3694 => x"81577477",
          3695 => x"077081ff",
          3696 => x"06515593",
          3697 => x"577480e2",
          3698 => x"38815377",
          3699 => x"528c3d70",
          3700 => x"52588296",
          3701 => x"a23f84ba",
          3702 => x"8c085784",
          3703 => x"ba8c0880",
          3704 => x"2e80d038",
          3705 => x"775182af",
          3706 => x"e03f7630",
          3707 => x"70780780",
          3708 => x"257b3070",
          3709 => x"9f2a7206",
          3710 => x"53575758",
          3711 => x"77802eaa",
          3712 => x"3887c098",
          3713 => x"88085574",
          3714 => x"87e72680",
          3715 => x"e0387452",
          3716 => x"7887e829",
          3717 => x"51f58e3f",
          3718 => x"84ba8c08",
          3719 => x"5483d2bc",
          3720 => x"53785283",
          3721 => x"d29851df",
          3722 => x"df3f7684",
          3723 => x"ba8c0c96",
          3724 => x"3d0d0484",
          3725 => x"ba8c0887",
          3726 => x"c098880c",
          3727 => x"84ba8c08",
          3728 => x"59963dd4",
          3729 => x"05548480",
          3730 => x"53755277",
          3731 => x"51829e97",
          3732 => x"3f84ba8c",
          3733 => x"085784ba",
          3734 => x"8c08ff88",
          3735 => x"387a5574",
          3736 => x"802eff80",
          3737 => x"38741975",
          3738 => x"175759d5",
          3739 => x"3987e852",
          3740 => x"7451f4b1",
          3741 => x"3f84ba8c",
          3742 => x"08527851",
          3743 => x"f4a73f84",
          3744 => x"ba8c0854",
          3745 => x"83d2bc53",
          3746 => x"785283d2",
          3747 => x"9851def8",
          3748 => x"3fff9739",
          3749 => x"f83d0d7c",
          3750 => x"028405b7",
          3751 => x"05335859",
          3752 => x"ff588053",
          3753 => x"7b527a51",
          3754 => x"fdec3f84",
          3755 => x"ba8c088b",
          3756 => x"3876802e",
          3757 => x"91387681",
          3758 => x"2e8a3877",
          3759 => x"84ba8c0c",
          3760 => x"8a3d0d04",
          3761 => x"780484d5",
          3762 => x"ec566155",
          3763 => x"605484ba",
          3764 => x"8c537f52",
          3765 => x"7e51782d",
          3766 => x"84ba8c08",
          3767 => x"84ba8c0c",
          3768 => x"8a3d0d04",
          3769 => x"f33d0d7f",
          3770 => x"6163028c",
          3771 => x"0580cf05",
          3772 => x"33737315",
          3773 => x"68415f5c",
          3774 => x"5c5f5d5e",
          3775 => x"78802e83",
          3776 => x"82387a52",
          3777 => x"83d2c451",
          3778 => x"ddfe3f83",
          3779 => x"d2cc51dd",
          3780 => x"f73f8054",
          3781 => x"737927b2",
          3782 => x"387c902e",
          3783 => x"81ed387c",
          3784 => x"a02e82a8",
          3785 => x"38731853",
          3786 => x"727a2781",
          3787 => x"a7387233",
          3788 => x"5283d2d0",
          3789 => x"51ddd13f",
          3790 => x"811484d5",
          3791 => x"f0085354",
          3792 => x"a051ecaa",
          3793 => x"3f787426",
          3794 => x"dc3883d2",
          3795 => x"d851ddb8",
          3796 => x"3f805675",
          3797 => x"792780c0",
          3798 => x"38751870",
          3799 => x"33555380",
          3800 => x"55727a27",
          3801 => x"83388155",
          3802 => x"80539f74",
          3803 => x"27833881",
          3804 => x"53747306",
          3805 => x"7081ff06",
          3806 => x"56577480",
          3807 => x"2e883880",
          3808 => x"fe742781",
          3809 => x"ee3884d5",
          3810 => x"f00852a0",
          3811 => x"51ebdf3f",
          3812 => x"81165678",
          3813 => x"7626c238",
          3814 => x"83d2dc51",
          3815 => x"e9d53f78",
          3816 => x"18791c5c",
          3817 => x"5880519d",
          3818 => x"b23f84ba",
          3819 => x"8c08982b",
          3820 => x"70982c58",
          3821 => x"5476a02e",
          3822 => x"81ee3876",
          3823 => x"9b2e82c3",
          3824 => x"387b1e57",
          3825 => x"767826fe",
          3826 => x"b938ff0b",
          3827 => x"84ba8c0c",
          3828 => x"8f3d0d04",
          3829 => x"83d2e051",
          3830 => x"dcae3f81",
          3831 => x"1484d5f0",
          3832 => x"085354a0",
          3833 => x"51eb873f",
          3834 => x"787426fe",
          3835 => x"b838feda",
          3836 => x"3983d2f0",
          3837 => x"51dc913f",
          3838 => x"821484d5",
          3839 => x"f0085354",
          3840 => x"a051eaea",
          3841 => x"3f737927",
          3842 => x"fec03873",
          3843 => x"1853727a",
          3844 => x"27df3872",
          3845 => x"225283d2",
          3846 => x"e451dbec",
          3847 => x"3f821484",
          3848 => x"d5f00853",
          3849 => x"54a051ea",
          3850 => x"c53f7874",
          3851 => x"26dd38fe",
          3852 => x"993983d2",
          3853 => x"ec51dbd0",
          3854 => x"3f841484",
          3855 => x"d5f00853",
          3856 => x"54a051ea",
          3857 => x"a93f7379",
          3858 => x"27fdff38",
          3859 => x"73185372",
          3860 => x"7a27df38",
          3861 => x"72085283",
          3862 => x"d2c451db",
          3863 => x"ab3f8414",
          3864 => x"84d5f008",
          3865 => x"5354a051",
          3866 => x"ea843f78",
          3867 => x"7426dd38",
          3868 => x"fdd83984",
          3869 => x"d5f00852",
          3870 => x"7351e9f2",
          3871 => x"3f811656",
          3872 => x"fe913980",
          3873 => x"cee33f84",
          3874 => x"ba8c0881",
          3875 => x"ff065388",
          3876 => x"5972a82e",
          3877 => x"fcec38a0",
          3878 => x"597280d0",
          3879 => x"2e098106",
          3880 => x"fce03890",
          3881 => x"59fcdb39",
          3882 => x"80519baf",
          3883 => x"3f84ba8c",
          3884 => x"08982b70",
          3885 => x"982c70a0",
          3886 => x"32703072",
          3887 => x"9b327030",
          3888 => x"70720773",
          3889 => x"75070651",
          3890 => x"55585957",
          3891 => x"58537280",
          3892 => x"25fde838",
          3893 => x"80519b83",
          3894 => x"3f84ba8c",
          3895 => x"08982b70",
          3896 => x"982c70a0",
          3897 => x"32703072",
          3898 => x"9b327030",
          3899 => x"70720773",
          3900 => x"75070651",
          3901 => x"55585957",
          3902 => x"58538073",
          3903 => x"24ffa938",
          3904 => x"fdb93980",
          3905 => x"0b84ba8c",
          3906 => x"0c8f3d0d",
          3907 => x"04fe3d0d",
          3908 => x"87c09680",
          3909 => x"0853aad1",
          3910 => x"3f81519c",
          3911 => x"f73f83d3",
          3912 => x"b4519d88",
          3913 => x"3f80519c",
          3914 => x"eb3f7281",
          3915 => x"2a708106",
          3916 => x"51527182",
          3917 => x"b7387282",
          3918 => x"2a708106",
          3919 => x"51527182",
          3920 => x"89387283",
          3921 => x"2a708106",
          3922 => x"51527181",
          3923 => x"db387284",
          3924 => x"2a708106",
          3925 => x"51527181",
          3926 => x"ad387285",
          3927 => x"2a708106",
          3928 => x"51527180",
          3929 => x"ff387286",
          3930 => x"2a708106",
          3931 => x"51527180",
          3932 => x"d2387287",
          3933 => x"2a708106",
          3934 => x"515271a9",
          3935 => x"3872882a",
          3936 => x"81065372",
          3937 => x"8838a9e9",
          3938 => x"3f843d0d",
          3939 => x"0481519c",
          3940 => x"833f83d3",
          3941 => x"cc519c94",
          3942 => x"3f80519b",
          3943 => x"f73fa9d1",
          3944 => x"3f843d0d",
          3945 => x"0481519b",
          3946 => x"eb3f83d3",
          3947 => x"e0519bfc",
          3948 => x"3f80519b",
          3949 => x"df3f7288",
          3950 => x"2a810653",
          3951 => x"72802ec6",
          3952 => x"38cb3981",
          3953 => x"519bcd3f",
          3954 => x"83d3f451",
          3955 => x"9bde3f80",
          3956 => x"519bc13f",
          3957 => x"72872a70",
          3958 => x"81065152",
          3959 => x"71802eff",
          3960 => x"9c38c239",
          3961 => x"81519bac",
          3962 => x"3f83d488",
          3963 => x"519bbd3f",
          3964 => x"80519ba0",
          3965 => x"3f72862a",
          3966 => x"70810651",
          3967 => x"5271802e",
          3968 => x"fef038ff",
          3969 => x"be398151",
          3970 => x"9b8a3f83",
          3971 => x"d49c519b",
          3972 => x"9b3f8051",
          3973 => x"9afe3f72",
          3974 => x"852a7081",
          3975 => x"06515271",
          3976 => x"802efec2",
          3977 => x"38ffbd39",
          3978 => x"81519ae8",
          3979 => x"3f83d4b0",
          3980 => x"519af93f",
          3981 => x"80519adc",
          3982 => x"3f72842a",
          3983 => x"70810651",
          3984 => x"5271802e",
          3985 => x"fe9438ff",
          3986 => x"bd398151",
          3987 => x"9ac63f83",
          3988 => x"d4c4519a",
          3989 => x"d73f8051",
          3990 => x"9aba3f72",
          3991 => x"832a7081",
          3992 => x"06515271",
          3993 => x"802efde6",
          3994 => x"38ffbd39",
          3995 => x"81519aa4",
          3996 => x"3f83d4d4",
          3997 => x"519ab53f",
          3998 => x"80519a98",
          3999 => x"3f72822a",
          4000 => x"70810651",
          4001 => x"5271802e",
          4002 => x"fdb838ff",
          4003 => x"bd39ca3d",
          4004 => x"0d807041",
          4005 => x"41ff6184",
          4006 => x"d1980c42",
          4007 => x"81526051",
          4008 => x"81b6d53f",
          4009 => x"84ba8c08",
          4010 => x"81ff069b",
          4011 => x"3d405978",
          4012 => x"612e84b1",
          4013 => x"3883d5a8",
          4014 => x"51e3b83f",
          4015 => x"983d4383",
          4016 => x"d5e051d6",
          4017 => x"c33f7e48",
          4018 => x"80f85380",
          4019 => x"527e51eb",
          4020 => x"ae3f0b0b",
          4021 => x"83ef8033",
          4022 => x"7081ff06",
          4023 => x"5b597980",
          4024 => x"2e82f138",
          4025 => x"79812e83",
          4026 => x"88387881",
          4027 => x"ff065e7d",
          4028 => x"822e83c1",
          4029 => x"3867705a",
          4030 => x"5a79802e",
          4031 => x"83dc3879",
          4032 => x"335c7ba0",
          4033 => x"2e098106",
          4034 => x"8c38811a",
          4035 => x"70335d5a",
          4036 => x"7ba02ef6",
          4037 => x"38805c7b",
          4038 => x"9b26be38",
          4039 => x"7b902983",
          4040 => x"ef840570",
          4041 => x"08525be7",
          4042 => x"ff3f84ba",
          4043 => x"8c0884ba",
          4044 => x"8c08547a",
          4045 => x"537b0852",
          4046 => x"5de8da3f",
          4047 => x"84ba8c08",
          4048 => x"8b38841b",
          4049 => x"335e7d81",
          4050 => x"2e838038",
          4051 => x"811c7081",
          4052 => x"ff065d5b",
          4053 => x"9b7c27c4",
          4054 => x"389a3d33",
          4055 => x"5c7b802e",
          4056 => x"fedd3880",
          4057 => x"f8527e51",
          4058 => x"e9923f84",
          4059 => x"ba8c085e",
          4060 => x"84ba8c08",
          4061 => x"802e8dd3",
          4062 => x"3884ba8c",
          4063 => x"0848b83d",
          4064 => x"ff800551",
          4065 => x"91933f84",
          4066 => x"ba8c0860",
          4067 => x"62065c5c",
          4068 => x"7a802e81",
          4069 => x"843884ba",
          4070 => x"8c0851e7",
          4071 => x"8b3f84ba",
          4072 => x"8c088f26",
          4073 => x"80f33881",
          4074 => x"0ba53d5e",
          4075 => x"5b7a822e",
          4076 => x"8d8f387a",
          4077 => x"82248cec",
          4078 => x"387a812e",
          4079 => x"82ee387b",
          4080 => x"54805383",
          4081 => x"d5e4527c",
          4082 => x"51d5dd3f",
          4083 => x"83f2c858",
          4084 => x"84babc57",
          4085 => x"7d566755",
          4086 => x"80549080",
          4087 => x"0a539080",
          4088 => x"0a527c51",
          4089 => x"f5ae3f84",
          4090 => x"ba8c0884",
          4091 => x"ba8c0809",
          4092 => x"70307072",
          4093 => x"07802551",
          4094 => x"5b5b4280",
          4095 => x"5a7a8326",
          4096 => x"8338815a",
          4097 => x"787a0659",
          4098 => x"78802e8d",
          4099 => x"38811b70",
          4100 => x"81ff065c",
          4101 => x"5a7aff95",
          4102 => x"387f8132",
          4103 => x"61813207",
          4104 => x"5d7c81f8",
          4105 => x"3861ff2e",
          4106 => x"81f2387d",
          4107 => x"518195aa",
          4108 => x"3f83d5e0",
          4109 => x"51d3d13f",
          4110 => x"7e4880f8",
          4111 => x"5380527e",
          4112 => x"51e8bc3f",
          4113 => x"0b0b83ef",
          4114 => x"80337081",
          4115 => x"ff065b59",
          4116 => x"79fd9138",
          4117 => x"815383d5",
          4118 => x"8c5284d1",
          4119 => x"9c518289",
          4120 => x"963f84ba",
          4121 => x"8c0880c5",
          4122 => x"38810b0b",
          4123 => x"0b83ef80",
          4124 => x"3484d19c",
          4125 => x"5380f852",
          4126 => x"7e5182f7",
          4127 => x"913f84ba",
          4128 => x"8c08802e",
          4129 => x"a03884ba",
          4130 => x"8c0851df",
          4131 => x"e63f0b0b",
          4132 => x"83ef8033",
          4133 => x"7081ff06",
          4134 => x"5f597d82",
          4135 => x"2e098106",
          4136 => x"fcd33891",
          4137 => x"3984d19c",
          4138 => x"5182a29d",
          4139 => x"3f820b0b",
          4140 => x"0b83ef80",
          4141 => x"3483d59c",
          4142 => x"5380f852",
          4143 => x"7e51a7ce",
          4144 => x"3f67705a",
          4145 => x"5a79fcb7",
          4146 => x"3890397c",
          4147 => x"1a630c85",
          4148 => x"1b335978",
          4149 => x"818926fd",
          4150 => x"80387810",
          4151 => x"1083bf9c",
          4152 => x"055a7908",
          4153 => x"0483d5ec",
          4154 => x"51df883f",
          4155 => x"9a3d5f83",
          4156 => x"5383d680",
          4157 => x"527e51e4",
          4158 => x"f13f6053",
          4159 => x"7e5284bb",
          4160 => x"b8518285",
          4161 => x"c33f84ba",
          4162 => x"8c08612e",
          4163 => x"098106fb",
          4164 => x"a4388170",
          4165 => x"9a3d4541",
          4166 => x"41fba439",
          4167 => x"83d68451",
          4168 => x"ded13f7d",
          4169 => x"518193b2",
          4170 => x"3ffe8639",
          4171 => x"83d69456",
          4172 => x"7b5583d6",
          4173 => x"98548053",
          4174 => x"83d69c52",
          4175 => x"7c51d2e8",
          4176 => x"3ffd8939",
          4177 => x"818ce33f",
          4178 => x"faf5399a",
          4179 => x"dd3ffaef",
          4180 => x"39815283",
          4181 => x"51bf943f",
          4182 => x"fae53981",
          4183 => x"8e953ffa",
          4184 => x"de3983d6",
          4185 => x"ac51de8b",
          4186 => x"3f805978",
          4187 => x"0483d6c0",
          4188 => x"51de803f",
          4189 => x"d0f33ffa",
          4190 => x"c639b83d",
          4191 => x"ff841153",
          4192 => x"ff800551",
          4193 => x"ec803f84",
          4194 => x"ba8c0880",
          4195 => x"2efab038",
          4196 => x"685283d6",
          4197 => x"dc51d0f0",
          4198 => x"3f685a79",
          4199 => x"2d84ba8c",
          4200 => x"08802efa",
          4201 => x"9a3884ba",
          4202 => x"8c085283",
          4203 => x"d6f851d0",
          4204 => x"d73ffa8b",
          4205 => x"39b83dff",
          4206 => x"841153ff",
          4207 => x"800551eb",
          4208 => x"c53f84ba",
          4209 => x"8c08802e",
          4210 => x"f9f53868",
          4211 => x"5283d794",
          4212 => x"51d0b53f",
          4213 => x"68597804",
          4214 => x"b83dfef4",
          4215 => x"1153ff80",
          4216 => x"0551e99e",
          4217 => x"3f84ba8c",
          4218 => x"08802ef9",
          4219 => x"d238b83d",
          4220 => x"fef01153",
          4221 => x"ff800551",
          4222 => x"e9883f84",
          4223 => x"ba8c0886",
          4224 => x"d0386459",
          4225 => x"78085378",
          4226 => x"5283d7b0",
          4227 => x"51cff93f",
          4228 => x"84d5ec08",
          4229 => x"5380f852",
          4230 => x"7e51d087",
          4231 => x"3f7e487e",
          4232 => x"335978ae",
          4233 => x"2ef99838",
          4234 => x"789f2687",
          4235 => x"d3386484",
          4236 => x"05704659",
          4237 => x"cf39b83d",
          4238 => x"fef41153",
          4239 => x"ff800551",
          4240 => x"e8c03f84",
          4241 => x"ba8c0880",
          4242 => x"2ef8f438",
          4243 => x"b83dfef0",
          4244 => x"1153ff80",
          4245 => x"0551e8aa",
          4246 => x"3f84ba8c",
          4247 => x"0886b038",
          4248 => x"64597822",
          4249 => x"53785283",
          4250 => x"d7c051cf",
          4251 => x"9b3f84d5",
          4252 => x"ec085380",
          4253 => x"f8527e51",
          4254 => x"cfa93f7e",
          4255 => x"487e3359",
          4256 => x"78ae2ef8",
          4257 => x"ba38789f",
          4258 => x"2687ca38",
          4259 => x"64820570",
          4260 => x"4659cf39",
          4261 => x"b83dff84",
          4262 => x"1153ff80",
          4263 => x"0551e9e6",
          4264 => x"3f84ba8c",
          4265 => x"08802ef8",
          4266 => x"9638b83d",
          4267 => x"fefc1153",
          4268 => x"ff800551",
          4269 => x"e9d03f84",
          4270 => x"ba8c0880",
          4271 => x"2ef88038",
          4272 => x"b83dfef8",
          4273 => x"1153ff80",
          4274 => x"0551e9ba",
          4275 => x"3f84ba8c",
          4276 => x"08802ef7",
          4277 => x"ea3883d7",
          4278 => x"cc51ceac",
          4279 => x"3f68675d",
          4280 => x"59787c27",
          4281 => x"838d3865",
          4282 => x"70337a33",
          4283 => x"5f5c5a7a",
          4284 => x"7d2e9538",
          4285 => x"7a557954",
          4286 => x"78335378",
          4287 => x"5283d7dc",
          4288 => x"51ce853f",
          4289 => x"66665b5c",
          4290 => x"8119811b",
          4291 => x"4759d239",
          4292 => x"b83dff84",
          4293 => x"1153ff80",
          4294 => x"0551e8ea",
          4295 => x"3f84ba8c",
          4296 => x"08802ef7",
          4297 => x"9a38b83d",
          4298 => x"fefc1153",
          4299 => x"ff800551",
          4300 => x"e8d43f84",
          4301 => x"ba8c0880",
          4302 => x"2ef78438",
          4303 => x"b83dfef8",
          4304 => x"1153ff80",
          4305 => x"0551e8be",
          4306 => x"3f84ba8c",
          4307 => x"08802ef6",
          4308 => x"ee3883d7",
          4309 => x"f851cdb0",
          4310 => x"3f685a79",
          4311 => x"67278293",
          4312 => x"38655c79",
          4313 => x"7081055b",
          4314 => x"337c3465",
          4315 => x"810546eb",
          4316 => x"39b83dff",
          4317 => x"841153ff",
          4318 => x"800551e8",
          4319 => x"893f84ba",
          4320 => x"8c08802e",
          4321 => x"f6b938b8",
          4322 => x"3dfefc11",
          4323 => x"53ff8005",
          4324 => x"51e7f33f",
          4325 => x"84ba8c08",
          4326 => x"b1386870",
          4327 => x"33545283",
          4328 => x"d88451cc",
          4329 => x"e33f84d5",
          4330 => x"ec085380",
          4331 => x"f8527e51",
          4332 => x"ccf13f7e",
          4333 => x"487e3359",
          4334 => x"78ae2ef6",
          4335 => x"8238789f",
          4336 => x"26849738",
          4337 => x"68810549",
          4338 => x"d1396859",
          4339 => x"0280db05",
          4340 => x"33793468",
          4341 => x"810549b8",
          4342 => x"3dfefc11",
          4343 => x"53ff8005",
          4344 => x"51e7a33f",
          4345 => x"84ba8c08",
          4346 => x"802ef5d3",
          4347 => x"38685902",
          4348 => x"80db0533",
          4349 => x"79346881",
          4350 => x"0549b83d",
          4351 => x"fefc1153",
          4352 => x"ff800551",
          4353 => x"e7803f84",
          4354 => x"ba8c08ff",
          4355 => x"bd38f5af",
          4356 => x"39b83dff",
          4357 => x"841153ff",
          4358 => x"800551e6",
          4359 => x"e93f84ba",
          4360 => x"8c08802e",
          4361 => x"f59938b8",
          4362 => x"3dfefc11",
          4363 => x"53ff8005",
          4364 => x"51e6d33f",
          4365 => x"84ba8c08",
          4366 => x"802ef583",
          4367 => x"38b83dfe",
          4368 => x"f81153ff",
          4369 => x"800551e6",
          4370 => x"bd3f84ba",
          4371 => x"8c088638",
          4372 => x"84ba8c08",
          4373 => x"4683d890",
          4374 => x"51cbad3f",
          4375 => x"68675b59",
          4376 => x"787a278f",
          4377 => x"38655b7a",
          4378 => x"79708405",
          4379 => x"5b0c7979",
          4380 => x"26f5388a",
          4381 => x"51d9e73f",
          4382 => x"f4c539b8",
          4383 => x"3dff8005",
          4384 => x"5187963f",
          4385 => x"84ba8c08",
          4386 => x"b93dff80",
          4387 => x"05525988",
          4388 => x"d83f8153",
          4389 => x"84ba8c08",
          4390 => x"527851e9",
          4391 => x"f93f84ba",
          4392 => x"8c08802e",
          4393 => x"f4993884",
          4394 => x"ba8c0851",
          4395 => x"e7ec3ff4",
          4396 => x"8e39b83d",
          4397 => x"ff841153",
          4398 => x"ff800551",
          4399 => x"e5c83f84",
          4400 => x"ba8c0891",
          4401 => x"3883f390",
          4402 => x"335a7980",
          4403 => x"2e83c038",
          4404 => x"83f2c808",
          4405 => x"49b83dfe",
          4406 => x"fc1153ff",
          4407 => x"800551e5",
          4408 => x"a53f84ba",
          4409 => x"8c089138",
          4410 => x"83f39033",
          4411 => x"5a79802e",
          4412 => x"838a3883",
          4413 => x"f2cc0847",
          4414 => x"b83dfef8",
          4415 => x"1153ff80",
          4416 => x"0551e582",
          4417 => x"3f84ba8c",
          4418 => x"08802ea5",
          4419 => x"3880665c",
          4420 => x"5c7a882e",
          4421 => x"8338815c",
          4422 => x"7a903270",
          4423 => x"30707207",
          4424 => x"9f2a7e06",
          4425 => x"5c5f5d79",
          4426 => x"802e8838",
          4427 => x"7aa02e83",
          4428 => x"38884683",
          4429 => x"d8a051d6",
          4430 => x"ba3f8055",
          4431 => x"68546553",
          4432 => x"66526851",
          4433 => x"eb9e3f83",
          4434 => x"d8ac51d6",
          4435 => x"a63ff2ef",
          4436 => x"39646471",
          4437 => x"0c596484",
          4438 => x"0545b83d",
          4439 => x"fef01153",
          4440 => x"ff800551",
          4441 => x"e29c3f84",
          4442 => x"ba8c0880",
          4443 => x"2ef2d038",
          4444 => x"6464710c",
          4445 => x"59648405",
          4446 => x"45b83dfe",
          4447 => x"f01153ff",
          4448 => x"800551e1",
          4449 => x"fd3f84ba",
          4450 => x"8c08c638",
          4451 => x"f2b13964",
          4452 => x"5e0280ce",
          4453 => x"05227e70",
          4454 => x"82054023",
          4455 => x"7d45b83d",
          4456 => x"fef01153",
          4457 => x"ff800551",
          4458 => x"e1d83f84",
          4459 => x"ba8c0880",
          4460 => x"2ef28c38",
          4461 => x"645e0280",
          4462 => x"ce05227e",
          4463 => x"70820540",
          4464 => x"237d45b8",
          4465 => x"3dfef011",
          4466 => x"53ff8005",
          4467 => x"51e1b33f",
          4468 => x"84ba8c08",
          4469 => x"ffb938f1",
          4470 => x"e639b83d",
          4471 => x"fefc1153",
          4472 => x"ff800551",
          4473 => x"e3a03f84",
          4474 => x"ba8c0880",
          4475 => x"2e81dc38",
          4476 => x"685c0280",
          4477 => x"db05337c",
          4478 => x"34688105",
          4479 => x"49fb9b39",
          4480 => x"b83dfef0",
          4481 => x"1153ff80",
          4482 => x"0551e0f6",
          4483 => x"3f84ba8c",
          4484 => x"08802e81",
          4485 => x"98386464",
          4486 => x"710c5d64",
          4487 => x"84057046",
          4488 => x"59f7e139",
          4489 => x"7a832e09",
          4490 => x"8106f393",
          4491 => x"387b5583",
          4492 => x"d6985480",
          4493 => x"5383d8b8",
          4494 => x"527c51c8",
          4495 => x"eb3ff38c",
          4496 => x"397b527c",
          4497 => x"51da803f",
          4498 => x"f3823983",
          4499 => x"d8c451d4",
          4500 => x"a23ff0eb",
          4501 => x"39b83dfe",
          4502 => x"f01153ff",
          4503 => x"800551e0",
          4504 => x"a13f84ba",
          4505 => x"8c08802e",
          4506 => x"b8386459",
          4507 => x"0280ce05",
          4508 => x"22797082",
          4509 => x"055b2378",
          4510 => x"45f7e739",
          4511 => x"83f39133",
          4512 => x"5c7b802e",
          4513 => x"80cf3883",
          4514 => x"f2d40847",
          4515 => x"fcea3983",
          4516 => x"f391335c",
          4517 => x"7b802ea1",
          4518 => x"3883f2d0",
          4519 => x"0849fcb5",
          4520 => x"3983d8f0",
          4521 => x"51d3cc3f",
          4522 => x"6459f7b6",
          4523 => x"3983d8f0",
          4524 => x"51d3c03f",
          4525 => x"6459f6cc",
          4526 => x"3983f392",
          4527 => x"33597880",
          4528 => x"2ea53883",
          4529 => x"f2d80849",
          4530 => x"fc8b3983",
          4531 => x"d8f051d3",
          4532 => x"a23ff9c6",
          4533 => x"3983f392",
          4534 => x"33597880",
          4535 => x"2e9b3883",
          4536 => x"f2dc0847",
          4537 => x"fc923983",
          4538 => x"f393335e",
          4539 => x"7d802e9b",
          4540 => x"3883f2e0",
          4541 => x"0849fbdd",
          4542 => x"3983f393",
          4543 => x"335e7d80",
          4544 => x"2e9b3883",
          4545 => x"f2e40847",
          4546 => x"fbee3983",
          4547 => x"f38e335d",
          4548 => x"7c802e9b",
          4549 => x"3883f2e8",
          4550 => x"0849fbb9",
          4551 => x"3983f38e",
          4552 => x"335d7c80",
          4553 => x"2e943883",
          4554 => x"f2ec0847",
          4555 => x"fbca3983",
          4556 => x"f2f808fc",
          4557 => x"800549fb",
          4558 => x"9c3983f2",
          4559 => x"f8088805",
          4560 => x"47fbb539",
          4561 => x"f33d0d80",
          4562 => x"0b84babc",
          4563 => x"3487c094",
          4564 => x"8c700856",
          4565 => x"57878480",
          4566 => x"527451da",
          4567 => x"c83f84ba",
          4568 => x"8c08902b",
          4569 => x"77085755",
          4570 => x"87848052",
          4571 => x"7551dab5",
          4572 => x"3f7484ba",
          4573 => x"8c080777",
          4574 => x"0c87c094",
          4575 => x"9c700856",
          4576 => x"57878480",
          4577 => x"527451da",
          4578 => x"9c3f84ba",
          4579 => x"8c08902b",
          4580 => x"77085755",
          4581 => x"87848052",
          4582 => x"7551da89",
          4583 => x"3f7484ba",
          4584 => x"8c080777",
          4585 => x"0c8c8083",
          4586 => x"0b87c094",
          4587 => x"840c8c80",
          4588 => x"830b87c0",
          4589 => x"94940c81",
          4590 => x"bcec5c81",
          4591 => x"c7eb5d83",
          4592 => x"028405a1",
          4593 => x"0534805e",
          4594 => x"84d5ec0b",
          4595 => x"893d7088",
          4596 => x"130c7072",
          4597 => x"0c84d5f0",
          4598 => x"0c56b6f5",
          4599 => x"3f89833f",
          4600 => x"95873fba",
          4601 => x"8d5194fc",
          4602 => x"3f83d2f8",
          4603 => x"5283d2fc",
          4604 => x"51c4953f",
          4605 => x"83f2fc70",
          4606 => x"22525594",
          4607 => x"873f83d3",
          4608 => x"845483d3",
          4609 => x"90538115",
          4610 => x"335283d3",
          4611 => x"9851c3f8",
          4612 => x"3f8d973f",
          4613 => x"ecf83f80",
          4614 => x"04fb3d0d",
          4615 => x"77700856",
          4616 => x"56807552",
          4617 => x"5374732e",
          4618 => x"81833874",
          4619 => x"337081ff",
          4620 => x"06525270",
          4621 => x"a02e0981",
          4622 => x"06913881",
          4623 => x"15703370",
          4624 => x"81ff0653",
          4625 => x"535570a0",
          4626 => x"2ef13871",
          4627 => x"81ff0654",
          4628 => x"73a22e81",
          4629 => x"82387452",
          4630 => x"72812e80",
          4631 => x"e7388072",
          4632 => x"337081ff",
          4633 => x"06535454",
          4634 => x"70a02e83",
          4635 => x"38815470",
          4636 => x"802e8b38",
          4637 => x"73802e86",
          4638 => x"38811252",
          4639 => x"e1398073",
          4640 => x"81ff0652",
          4641 => x"5470a02e",
          4642 => x"09810683",
          4643 => x"38815470",
          4644 => x"a2327030",
          4645 => x"70802576",
          4646 => x"07525253",
          4647 => x"72802e88",
          4648 => x"38807270",
          4649 => x"81055434",
          4650 => x"71760c74",
          4651 => x"517084ba",
          4652 => x"8c0c873d",
          4653 => x"0d047080",
          4654 => x"2ec43873",
          4655 => x"802effbe",
          4656 => x"38811252",
          4657 => x"80723370",
          4658 => x"81ff0653",
          4659 => x"545470a2",
          4660 => x"2ee43881",
          4661 => x"54e03981",
          4662 => x"15558175",
          4663 => x"53537281",
          4664 => x"2e098106",
          4665 => x"fef838dc",
          4666 => x"39fc3d0d",
          4667 => x"76537208",
          4668 => x"8b38800b",
          4669 => x"84ba8c0c",
          4670 => x"863d0d04",
          4671 => x"863dfc05",
          4672 => x"527251da",
          4673 => x"fd3f84ba",
          4674 => x"8c08802e",
          4675 => x"e5387484",
          4676 => x"ba8c0c86",
          4677 => x"3d0d04fc",
          4678 => x"3d0d7682",
          4679 => x"1133ff05",
          4680 => x"52538152",
          4681 => x"708b2681",
          4682 => x"98388313",
          4683 => x"33ff0554",
          4684 => x"8252739e",
          4685 => x"26818a38",
          4686 => x"84133351",
          4687 => x"83527097",
          4688 => x"2680fe38",
          4689 => x"85133354",
          4690 => x"845273bb",
          4691 => x"2680f238",
          4692 => x"86133355",
          4693 => x"855274bb",
          4694 => x"2680e638",
          4695 => x"88132255",
          4696 => x"86527487",
          4697 => x"e72680d9",
          4698 => x"388a1322",
          4699 => x"54875273",
          4700 => x"87e72680",
          4701 => x"cc38810b",
          4702 => x"87c0989c",
          4703 => x"0c722287",
          4704 => x"c098bc0c",
          4705 => x"82133387",
          4706 => x"c098b80c",
          4707 => x"83133387",
          4708 => x"c098b40c",
          4709 => x"84133387",
          4710 => x"c098b00c",
          4711 => x"85133387",
          4712 => x"c098ac0c",
          4713 => x"86133387",
          4714 => x"c098a80c",
          4715 => x"7487c098",
          4716 => x"a40c7387",
          4717 => x"c098a00c",
          4718 => x"800b87c0",
          4719 => x"989c0c80",
          4720 => x"527184ba",
          4721 => x"8c0c863d",
          4722 => x"0d04f33d",
          4723 => x"0d7f5b87",
          4724 => x"c0989c5d",
          4725 => x"817d0c87",
          4726 => x"c098bc08",
          4727 => x"5e7d7b23",
          4728 => x"87c098b8",
          4729 => x"085c7b82",
          4730 => x"1c3487c0",
          4731 => x"98b4085a",
          4732 => x"79831c34",
          4733 => x"87c098b0",
          4734 => x"085c7b84",
          4735 => x"1c3487c0",
          4736 => x"98ac085a",
          4737 => x"79851c34",
          4738 => x"87c098a8",
          4739 => x"085c7b86",
          4740 => x"1c3487c0",
          4741 => x"98a4085c",
          4742 => x"7b881c23",
          4743 => x"87c098a0",
          4744 => x"085a798a",
          4745 => x"1c23807d",
          4746 => x"0c7983ff",
          4747 => x"ff06597b",
          4748 => x"83ffff06",
          4749 => x"58861b33",
          4750 => x"57851b33",
          4751 => x"56841b33",
          4752 => x"55831b33",
          4753 => x"54821b33",
          4754 => x"537d83ff",
          4755 => x"ff065283",
          4756 => x"d8f451ff",
          4757 => x"bfb23f8f",
          4758 => x"3d0d04fe",
          4759 => x"3d0d0293",
          4760 => x"05335372",
          4761 => x"812ea838",
          4762 => x"725180e8",
          4763 => x"b13f84ba",
          4764 => x"8c08982b",
          4765 => x"70982c51",
          4766 => x"5271ff2e",
          4767 => x"09810686",
          4768 => x"3872832e",
          4769 => x"e3387184",
          4770 => x"ba8c0c84",
          4771 => x"3d0d0472",
          4772 => x"5180e88a",
          4773 => x"3f84ba8c",
          4774 => x"08982b70",
          4775 => x"982c5152",
          4776 => x"71ff2e09",
          4777 => x"8106df38",
          4778 => x"725180e7",
          4779 => x"f13f84ba",
          4780 => x"8c08982b",
          4781 => x"70982c51",
          4782 => x"5271ff2e",
          4783 => x"d238c739",
          4784 => x"fd3d0d80",
          4785 => x"70545271",
          4786 => x"882b5481",
          4787 => x"5180e7ce",
          4788 => x"3f84ba8c",
          4789 => x"08982b70",
          4790 => x"982c5152",
          4791 => x"71ff2eeb",
          4792 => x"38737207",
          4793 => x"81145452",
          4794 => x"837325db",
          4795 => x"387184ba",
          4796 => x"8c0c853d",
          4797 => x"0d04fc3d",
          4798 => x"0d029b05",
          4799 => x"3383f2c4",
          4800 => x"337081ff",
          4801 => x"06535555",
          4802 => x"70802e80",
          4803 => x"f43887c0",
          4804 => x"94940870",
          4805 => x"962a7081",
          4806 => x"06535452",
          4807 => x"70802e8c",
          4808 => x"3871912a",
          4809 => x"70810651",
          4810 => x"5170e338",
          4811 => x"72813281",
          4812 => x"06537280",
          4813 => x"2e8a3871",
          4814 => x"932a8106",
          4815 => x"5271cf38",
          4816 => x"7381ff06",
          4817 => x"5187c094",
          4818 => x"80527080",
          4819 => x"2e863887",
          4820 => x"c0949052",
          4821 => x"74720c74",
          4822 => x"84ba8c0c",
          4823 => x"863d0d04",
          4824 => x"71912a70",
          4825 => x"81065151",
          4826 => x"70973872",
          4827 => x"81328106",
          4828 => x"5372802e",
          4829 => x"cb387193",
          4830 => x"2a810652",
          4831 => x"71802ec0",
          4832 => x"3887c094",
          4833 => x"84087096",
          4834 => x"2a708106",
          4835 => x"53545270",
          4836 => x"cf38d839",
          4837 => x"ff3d0d02",
          4838 => x"8f053370",
          4839 => x"30709f2a",
          4840 => x"51525270",
          4841 => x"83f2c434",
          4842 => x"833d0d04",
          4843 => x"fa3d0d78",
          4844 => x"55807533",
          4845 => x"70565257",
          4846 => x"70772e80",
          4847 => x"e7388115",
          4848 => x"83f2c433",
          4849 => x"7081ff06",
          4850 => x"54575571",
          4851 => x"802e80ff",
          4852 => x"3887c094",
          4853 => x"94087096",
          4854 => x"2a708106",
          4855 => x"53545270",
          4856 => x"802e8c38",
          4857 => x"71912a70",
          4858 => x"81065151",
          4859 => x"70e33872",
          4860 => x"81328106",
          4861 => x"5372802e",
          4862 => x"8a387193",
          4863 => x"2a810652",
          4864 => x"71cf3875",
          4865 => x"81ff0651",
          4866 => x"87c09480",
          4867 => x"5270802e",
          4868 => x"863887c0",
          4869 => x"94905273",
          4870 => x"720c8117",
          4871 => x"75335557",
          4872 => x"73ff9b38",
          4873 => x"7684ba8c",
          4874 => x"0c883d0d",
          4875 => x"0471912a",
          4876 => x"70810651",
          4877 => x"51709838",
          4878 => x"72813281",
          4879 => x"06537280",
          4880 => x"2ec13871",
          4881 => x"932a8106",
          4882 => x"5271802e",
          4883 => x"ffb53887",
          4884 => x"c0948408",
          4885 => x"70962a70",
          4886 => x"81065354",
          4887 => x"5270ce38",
          4888 => x"d739ff3d",
          4889 => x"0d87c09e",
          4890 => x"8008709c",
          4891 => x"2a8a0652",
          4892 => x"5270802e",
          4893 => x"84ab3887",
          4894 => x"c09ea408",
          4895 => x"83f2c80c",
          4896 => x"87c09ea8",
          4897 => x"0883f2cc",
          4898 => x"0c87c09e",
          4899 => x"940883f2",
          4900 => x"d00c87c0",
          4901 => x"9e980883",
          4902 => x"f2d40c87",
          4903 => x"c09e9c08",
          4904 => x"83f2d80c",
          4905 => x"87c09ea0",
          4906 => x"0883f2dc",
          4907 => x"0c87c09e",
          4908 => x"ac0883f2",
          4909 => x"e00c87c0",
          4910 => x"9eb00883",
          4911 => x"f2e40c87",
          4912 => x"c09eb408",
          4913 => x"83f2e80c",
          4914 => x"87c09eb8",
          4915 => x"0883f2ec",
          4916 => x"0c87c09e",
          4917 => x"bc0883f2",
          4918 => x"f00c87c0",
          4919 => x"9ec00883",
          4920 => x"f2f40c87",
          4921 => x"c09ec408",
          4922 => x"83f2f80c",
          4923 => x"87c09e80",
          4924 => x"08527183",
          4925 => x"f2fc2387",
          4926 => x"c09e8408",
          4927 => x"83f3800c",
          4928 => x"87c09e88",
          4929 => x"0883f384",
          4930 => x"0c87c09e",
          4931 => x"8c0883f3",
          4932 => x"880c810b",
          4933 => x"83f38c34",
          4934 => x"800b87c0",
          4935 => x"9e900870",
          4936 => x"84800a06",
          4937 => x"51525270",
          4938 => x"82fb3871",
          4939 => x"83f38d34",
          4940 => x"800b87c0",
          4941 => x"9e900870",
          4942 => x"88800a06",
          4943 => x"51525270",
          4944 => x"802e8338",
          4945 => x"81527183",
          4946 => x"f38e3480",
          4947 => x"0b87c09e",
          4948 => x"90087090",
          4949 => x"800a0651",
          4950 => x"52527080",
          4951 => x"2e833881",
          4952 => x"527183f3",
          4953 => x"8f34800b",
          4954 => x"87c09e90",
          4955 => x"08708880",
          4956 => x"80065152",
          4957 => x"5270802e",
          4958 => x"83388152",
          4959 => x"7183f390",
          4960 => x"34800b87",
          4961 => x"c09e9008",
          4962 => x"70a08080",
          4963 => x"06515252",
          4964 => x"70802e83",
          4965 => x"38815271",
          4966 => x"83f39134",
          4967 => x"800b87c0",
          4968 => x"9e900870",
          4969 => x"90808006",
          4970 => x"51525270",
          4971 => x"802e8338",
          4972 => x"81527183",
          4973 => x"f3923480",
          4974 => x"0b87c09e",
          4975 => x"90087084",
          4976 => x"80800651",
          4977 => x"52527080",
          4978 => x"2e833881",
          4979 => x"527183f3",
          4980 => x"9334800b",
          4981 => x"87c09e90",
          4982 => x"08708280",
          4983 => x"80065152",
          4984 => x"5270802e",
          4985 => x"83388152",
          4986 => x"7183f394",
          4987 => x"34800b87",
          4988 => x"c09e9008",
          4989 => x"70818080",
          4990 => x"06515252",
          4991 => x"70802e83",
          4992 => x"38815271",
          4993 => x"83f39534",
          4994 => x"800b87c0",
          4995 => x"9e900870",
          4996 => x"80c08006",
          4997 => x"51525270",
          4998 => x"802e8338",
          4999 => x"81527183",
          5000 => x"f3963480",
          5001 => x"0b87c09e",
          5002 => x"900870a0",
          5003 => x"80065152",
          5004 => x"5270802e",
          5005 => x"83388152",
          5006 => x"7183f397",
          5007 => x"3487c09e",
          5008 => x"90089880",
          5009 => x"06708a2a",
          5010 => x"53517183",
          5011 => x"f3983480",
          5012 => x"0b87c09e",
          5013 => x"90087084",
          5014 => x"80065152",
          5015 => x"5270802e",
          5016 => x"83388152",
          5017 => x"7183f399",
          5018 => x"3487c09e",
          5019 => x"900883f0",
          5020 => x"0670842a",
          5021 => x"53517183",
          5022 => x"f39a3480",
          5023 => x"0b87c09e",
          5024 => x"90087088",
          5025 => x"06515252",
          5026 => x"70802e83",
          5027 => x"38815271",
          5028 => x"83f39b34",
          5029 => x"87c09e90",
          5030 => x"08870651",
          5031 => x"7083f39c",
          5032 => x"34833d0d",
          5033 => x"048152fd",
          5034 => x"8239fb3d",
          5035 => x"0d83d98c",
          5036 => x"51ffb6d4",
          5037 => x"3f83f38c",
          5038 => x"33547386",
          5039 => x"aa3883d9",
          5040 => x"a051c3af",
          5041 => x"3f83f38e",
          5042 => x"33557485",
          5043 => x"fa3883f3",
          5044 => x"93335473",
          5045 => x"85d13883",
          5046 => x"f3903356",
          5047 => x"7585a838",
          5048 => x"83f39133",
          5049 => x"557484ff",
          5050 => x"3883f392",
          5051 => x"33547384",
          5052 => x"d63883f3",
          5053 => x"97335675",
          5054 => x"84b33883",
          5055 => x"f39b3354",
          5056 => x"73849038",
          5057 => x"83f39933",
          5058 => x"557483ed",
          5059 => x"3883f38d",
          5060 => x"33567583",
          5061 => x"cf3883f3",
          5062 => x"8f335473",
          5063 => x"83b13883",
          5064 => x"f3943355",
          5065 => x"74839338",
          5066 => x"83f39533",
          5067 => x"567582f4",
          5068 => x"3883f396",
          5069 => x"33547381",
          5070 => x"ec3883d9",
          5071 => x"b851c2b3",
          5072 => x"3f83f2f0",
          5073 => x"085283d9",
          5074 => x"c451ffb5",
          5075 => x"bb3f83f2",
          5076 => x"f4085283",
          5077 => x"d9ec51ff",
          5078 => x"b5ae3f83",
          5079 => x"f2f80852",
          5080 => x"83da9451",
          5081 => x"ffb5a13f",
          5082 => x"83dabc51",
          5083 => x"c2853f83",
          5084 => x"f2fc2252",
          5085 => x"83dac451",
          5086 => x"ffb58d3f",
          5087 => x"83f38008",
          5088 => x"56bd84c0",
          5089 => x"527551ca",
          5090 => x"9c3f84ba",
          5091 => x"8c08bd84",
          5092 => x"c0297671",
          5093 => x"31545484",
          5094 => x"ba8c0852",
          5095 => x"83daec51",
          5096 => x"ffb4e53f",
          5097 => x"83f39333",
          5098 => x"557480c3",
          5099 => x"3883f38e",
          5100 => x"3355748a",
          5101 => x"388a51c3",
          5102 => x"a53f873d",
          5103 => x"0d0483f3",
          5104 => x"880856bd",
          5105 => x"84c05275",
          5106 => x"51c9da3f",
          5107 => x"84ba8c08",
          5108 => x"bd84c029",
          5109 => x"76713154",
          5110 => x"5484ba8c",
          5111 => x"085283db",
          5112 => x"9851ffb4",
          5113 => x"a33f8a51",
          5114 => x"c2f43f87",
          5115 => x"3d0d0483",
          5116 => x"f3840856",
          5117 => x"bd84c052",
          5118 => x"7551c9a9",
          5119 => x"3f84ba8c",
          5120 => x"08bd84c0",
          5121 => x"29767131",
          5122 => x"545484ba",
          5123 => x"8c085283",
          5124 => x"dbc451ff",
          5125 => x"b3f23f83",
          5126 => x"f38e3355",
          5127 => x"74802eff",
          5128 => x"9438ff9a",
          5129 => x"3983dbf0",
          5130 => x"51c0c83f",
          5131 => x"83d9b851",
          5132 => x"c0c13f83",
          5133 => x"f2f00852",
          5134 => x"83d9c451",
          5135 => x"ffb3c93f",
          5136 => x"83f2f408",
          5137 => x"5283d9ec",
          5138 => x"51ffb3bc",
          5139 => x"3f83f2f8",
          5140 => x"085283da",
          5141 => x"9451ffb3",
          5142 => x"af3f83da",
          5143 => x"bc51c093",
          5144 => x"3f83f2fc",
          5145 => x"225283da",
          5146 => x"c451ffb3",
          5147 => x"9b3f83f3",
          5148 => x"800856bd",
          5149 => x"84c05275",
          5150 => x"51c8aa3f",
          5151 => x"84ba8c08",
          5152 => x"bd84c029",
          5153 => x"76713154",
          5154 => x"5484ba8c",
          5155 => x"085283da",
          5156 => x"ec51ffb2",
          5157 => x"f33f83f3",
          5158 => x"93335574",
          5159 => x"802efe8d",
          5160 => x"38fecc39",
          5161 => x"83dbf851",
          5162 => x"ffbfc83f",
          5163 => x"83f39633",
          5164 => x"5473802e",
          5165 => x"fd8438fe",
          5166 => x"ec3983dc",
          5167 => x"8051ffbf",
          5168 => x"b23f83f3",
          5169 => x"95335675",
          5170 => x"802efce5",
          5171 => x"38d63983",
          5172 => x"dc8c51ff",
          5173 => x"bf9d3f83",
          5174 => x"f3943355",
          5175 => x"74802efc",
          5176 => x"c738d739",
          5177 => x"83dc9851",
          5178 => x"ffbf883f",
          5179 => x"83f38f33",
          5180 => x"5473802e",
          5181 => x"fca938d7",
          5182 => x"3983f39a",
          5183 => x"335283dc",
          5184 => x"ac51ffb2",
          5185 => x"833f83f3",
          5186 => x"8d335675",
          5187 => x"802efc86",
          5188 => x"38d23983",
          5189 => x"f39c3352",
          5190 => x"83dccc51",
          5191 => x"ffb1e93f",
          5192 => x"83f39933",
          5193 => x"5574802e",
          5194 => x"fbe338cd",
          5195 => x"3983f398",
          5196 => x"335283dc",
          5197 => x"ec51ffb1",
          5198 => x"cf3f83f3",
          5199 => x"9b335473",
          5200 => x"802efbc0",
          5201 => x"38cd3983",
          5202 => x"f2d80883",
          5203 => x"f2dc0811",
          5204 => x"545283dd",
          5205 => x"8c51ffb1",
          5206 => x"af3f83f3",
          5207 => x"97335675",
          5208 => x"802efb97",
          5209 => x"38c73983",
          5210 => x"f2d00883",
          5211 => x"f2d40811",
          5212 => x"545283dd",
          5213 => x"a851ffb1",
          5214 => x"8f3f83f3",
          5215 => x"92335473",
          5216 => x"802efaee",
          5217 => x"38c13983",
          5218 => x"f2c80883",
          5219 => x"f2cc0811",
          5220 => x"545283dd",
          5221 => x"c451ffb0",
          5222 => x"ef3f83f3",
          5223 => x"91335574",
          5224 => x"802efac5",
          5225 => x"38c13983",
          5226 => x"f2e00883",
          5227 => x"f2e40811",
          5228 => x"545283dd",
          5229 => x"e051ffb0",
          5230 => x"cf3f83f3",
          5231 => x"90335675",
          5232 => x"802efa9c",
          5233 => x"38c13983",
          5234 => x"f2e80883",
          5235 => x"f2ec0811",
          5236 => x"545283dd",
          5237 => x"fc51ffb0",
          5238 => x"af3f83f3",
          5239 => x"93335473",
          5240 => x"802ef9f3",
          5241 => x"38c13983",
          5242 => x"de9851ff",
          5243 => x"b09a3f83",
          5244 => x"d9a051ff",
          5245 => x"bcfd3f83",
          5246 => x"f38e3355",
          5247 => x"74802ef9",
          5248 => x"cd38c439",
          5249 => x"ff3d0d02",
          5250 => x"8e053352",
          5251 => x"7185268c",
          5252 => x"38711010",
          5253 => x"83c3c405",
          5254 => x"52710804",
          5255 => x"83deac51",
          5256 => x"ffafe53f",
          5257 => x"833d0d04",
          5258 => x"83deb451",
          5259 => x"ffafd93f",
          5260 => x"833d0d04",
          5261 => x"83debc51",
          5262 => x"ffafcd3f",
          5263 => x"833d0d04",
          5264 => x"83dec451",
          5265 => x"ffafc13f",
          5266 => x"833d0d04",
          5267 => x"83decc51",
          5268 => x"ffafb53f",
          5269 => x"833d0d04",
          5270 => x"83ded451",
          5271 => x"ffafa93f",
          5272 => x"833d0d04",
          5273 => x"7188800c",
          5274 => x"04800b87",
          5275 => x"c096840c",
          5276 => x"0483f3a0",
          5277 => x"0887c096",
          5278 => x"840c04d9",
          5279 => x"3d0daa3d",
          5280 => x"08ad3d08",
          5281 => x"5a5a8170",
          5282 => x"57588052",
          5283 => x"83f3f808",
          5284 => x"518288d2",
          5285 => x"3f84ba8c",
          5286 => x"0880ed38",
          5287 => x"8b3d57ff",
          5288 => x"0b83f3f8",
          5289 => x"08545580",
          5290 => x"f8527651",
          5291 => x"82d2df3f",
          5292 => x"84ba8c08",
          5293 => x"802ea438",
          5294 => x"7651c0ec",
          5295 => x"3f84ba8c",
          5296 => x"08811757",
          5297 => x"55800b84",
          5298 => x"ba8c0825",
          5299 => x"8e3884ba",
          5300 => x"8c08ff05",
          5301 => x"70185555",
          5302 => x"80743474",
          5303 => x"09703070",
          5304 => x"72079f2a",
          5305 => x"51555578",
          5306 => x"762e8538",
          5307 => x"73ffb038",
          5308 => x"83f3f808",
          5309 => x"8c110853",
          5310 => x"518287ea",
          5311 => x"3f84ba8c",
          5312 => x"088f3878",
          5313 => x"762e9a38",
          5314 => x"7784ba8c",
          5315 => x"0ca93d0d",
          5316 => x"0483e284",
          5317 => x"51ffadf0",
          5318 => x"3f78762e",
          5319 => x"098106e8",
          5320 => x"38765279",
          5321 => x"51c0a03f",
          5322 => x"7951ffbf",
          5323 => x"fb3fab3d",
          5324 => x"085684ba",
          5325 => x"8c087634",
          5326 => x"765283e2",
          5327 => x"b051ffad",
          5328 => x"c73f800b",
          5329 => x"84ba8c0c",
          5330 => x"a93d0d04",
          5331 => x"d83d0dab",
          5332 => x"3d08ad3d",
          5333 => x"0871725d",
          5334 => x"72335757",
          5335 => x"5a5773a0",
          5336 => x"2e819138",
          5337 => x"800b8d3d",
          5338 => x"59567510",
          5339 => x"101083f4",
          5340 => x"80057008",
          5341 => x"5254ffbf",
          5342 => x"af3f84ba",
          5343 => x"8c085379",
          5344 => x"52730851",
          5345 => x"c08f3f84",
          5346 => x"ba8c0890",
          5347 => x"38841433",
          5348 => x"5473812e",
          5349 => x"81883873",
          5350 => x"822e9938",
          5351 => x"81167081",
          5352 => x"ff065754",
          5353 => x"827627c2",
          5354 => x"38805473",
          5355 => x"84ba8c0c",
          5356 => x"aa3d0d04",
          5357 => x"811a5aaa",
          5358 => x"3dff8411",
          5359 => x"53ff8005",
          5360 => x"51c7c33f",
          5361 => x"84ba8c08",
          5362 => x"802ed138",
          5363 => x"ff1b5378",
          5364 => x"527651fd",
          5365 => x"a63f84ba",
          5366 => x"8c0881ff",
          5367 => x"06547380",
          5368 => x"2ec93881",
          5369 => x"167081ff",
          5370 => x"06575482",
          5371 => x"7627fefa",
          5372 => x"38ffb639",
          5373 => x"78337705",
          5374 => x"56767627",
          5375 => x"fee63881",
          5376 => x"15705b70",
          5377 => x"33555573",
          5378 => x"a02e0981",
          5379 => x"06fed538",
          5380 => x"757526eb",
          5381 => x"38800b8d",
          5382 => x"3d5956fe",
          5383 => x"cd397384",
          5384 => x"ba8c0853",
          5385 => x"83f3f808",
          5386 => x"52568285",
          5387 => x"b93f84ba",
          5388 => x"8c0880d0",
          5389 => x"3883f3f8",
          5390 => x"085380f8",
          5391 => x"52775182",
          5392 => x"cfcc3f84",
          5393 => x"ba8c0880",
          5394 => x"2eba3877",
          5395 => x"51ffbdd8",
          5396 => x"3f84ba8c",
          5397 => x"0855800b",
          5398 => x"84ba8c08",
          5399 => x"259d3884",
          5400 => x"ba8c08ff",
          5401 => x"05701958",
          5402 => x"55807734",
          5403 => x"77537552",
          5404 => x"811683e1",
          5405 => x"f85256ff",
          5406 => x"ab8e3f74",
          5407 => x"ff2e0981",
          5408 => x"06ffb238",
          5409 => x"810b84ba",
          5410 => x"8c0caa3d",
          5411 => x"0d04ce3d",
          5412 => x"0db53d08",
          5413 => x"b73d08b9",
          5414 => x"3d085a41",
          5415 => x"5c800bb4",
          5416 => x"3d3483f3",
          5417 => x"fc3383f3",
          5418 => x"f808565d",
          5419 => x"749e3874",
          5420 => x"83f3f433",
          5421 => x"56567480",
          5422 => x"2e82cb38",
          5423 => x"77802e91",
          5424 => x"8d388170",
          5425 => x"77065a57",
          5426 => x"7890a038",
          5427 => x"77802e90",
          5428 => x"fd38933d",
          5429 => x"b43d5f5f",
          5430 => x"8051eaff",
          5431 => x"3f84ba8c",
          5432 => x"08982b70",
          5433 => x"982c5b56",
          5434 => x"79ff2eec",
          5435 => x"387981ff",
          5436 => x"0684d1c8",
          5437 => x"3370982b",
          5438 => x"70982c84",
          5439 => x"d1c43370",
          5440 => x"982b7097",
          5441 => x"2c71982c",
          5442 => x"05701010",
          5443 => x"83ded805",
          5444 => x"70081570",
          5445 => x"3352535c",
          5446 => x"5d46525b",
          5447 => x"585c5981",
          5448 => x"5774792e",
          5449 => x"80cd3878",
          5450 => x"75278187",
          5451 => x"38758180",
          5452 => x"0a2981ff",
          5453 => x"0a057098",
          5454 => x"2c575580",
          5455 => x"762481cb",
          5456 => x"38751016",
          5457 => x"70822b56",
          5458 => x"57800b83",
          5459 => x"dedc1633",
          5460 => x"42577761",
          5461 => x"25913883",
          5462 => x"ded81508",
          5463 => x"18703356",
          5464 => x"4178752e",
          5465 => x"81953876",
          5466 => x"802ec238",
          5467 => x"7584d1c4",
          5468 => x"34815776",
          5469 => x"802e8199",
          5470 => x"38811b70",
          5471 => x"982b7098",
          5472 => x"2c84d1c4",
          5473 => x"3370982b",
          5474 => x"70972c71",
          5475 => x"982c0570",
          5476 => x"822b83de",
          5477 => x"dc11335f",
          5478 => x"535f5d58",
          5479 => x"5d57577a",
          5480 => x"782e8190",
          5481 => x"387684d1",
          5482 => x"c834feac",
          5483 => x"39815776",
          5484 => x"ffba3875",
          5485 => x"81800a29",
          5486 => x"81800a05",
          5487 => x"70982c70",
          5488 => x"81ff0659",
          5489 => x"57417695",
          5490 => x"2680c038",
          5491 => x"75101670",
          5492 => x"822b5155",
          5493 => x"800b83de",
          5494 => x"dc163342",
          5495 => x"57776125",
          5496 => x"ce3883de",
          5497 => x"d8150818",
          5498 => x"70334255",
          5499 => x"78612eff",
          5500 => x"bc387680",
          5501 => x"2effbc38",
          5502 => x"fef23981",
          5503 => x"5776802e",
          5504 => x"feab38fe",
          5505 => x"e7398156",
          5506 => x"fdb23980",
          5507 => x"5776fee9",
          5508 => x"387684d1",
          5509 => x"c8347684",
          5510 => x"d1c43479",
          5511 => x"7e34767f",
          5512 => x"0c625574",
          5513 => x"9526fdb0",
          5514 => x"38741010",
          5515 => x"83c3dc05",
          5516 => x"57760804",
          5517 => x"83dee015",
          5518 => x"087f0c80",
          5519 => x"0b84d1c8",
          5520 => x"34800b84",
          5521 => x"d1c434d9",
          5522 => x"3984d1d0",
          5523 => x"33567580",
          5524 => x"2efd8538",
          5525 => x"84d5f008",
          5526 => x"528851ff",
          5527 => x"b6903f84",
          5528 => x"d1d033ff",
          5529 => x"05577684",
          5530 => x"d1d034fc",
          5531 => x"eb3984d1",
          5532 => x"d0337081",
          5533 => x"ff0684d1",
          5534 => x"cc335b57",
          5535 => x"55757927",
          5536 => x"fcd63884",
          5537 => x"d5f00852",
          5538 => x"81155877",
          5539 => x"84d1d034",
          5540 => x"7b167033",
          5541 => x"5255ffb5",
          5542 => x"d53ffcbc",
          5543 => x"397c932e",
          5544 => x"8bda387c",
          5545 => x"101083f3",
          5546 => x"a8057008",
          5547 => x"5759758f",
          5548 => x"83387584",
          5549 => x"d1cc3475",
          5550 => x"7c3484d1",
          5551 => x"cc3384d1",
          5552 => x"d0335656",
          5553 => x"74802eb6",
          5554 => x"3884d5f0",
          5555 => x"08528851",
          5556 => x"ffb59b3f",
          5557 => x"84d5f008",
          5558 => x"52a051ff",
          5559 => x"b5903f84",
          5560 => x"d5f00852",
          5561 => x"8851ffb5",
          5562 => x"853f84d1",
          5563 => x"d033ff05",
          5564 => x"5b7a84d1",
          5565 => x"d0347a81",
          5566 => x"ff065574",
          5567 => x"cc387b51",
          5568 => x"ffa6853f",
          5569 => x"7584d1d0",
          5570 => x"34fbcd39",
          5571 => x"7c8a3883",
          5572 => x"f3f00856",
          5573 => x"758d9e38",
          5574 => x"7c101083",
          5575 => x"f3a405fc",
          5576 => x"11085755",
          5577 => x"758ef938",
          5578 => x"74085675",
          5579 => x"802efba8",
          5580 => x"387551ff",
          5581 => x"b7f23f84",
          5582 => x"ba8c0884",
          5583 => x"d1cc3484",
          5584 => x"ba8c0881",
          5585 => x"ff068105",
          5586 => x"5375527b",
          5587 => x"51ffb89a",
          5588 => x"3f84d1cc",
          5589 => x"3384d1d0",
          5590 => x"33565674",
          5591 => x"802eff9e",
          5592 => x"3884d5f0",
          5593 => x"08528851",
          5594 => x"ffb4833f",
          5595 => x"84d5f008",
          5596 => x"52a051ff",
          5597 => x"b3f83f84",
          5598 => x"d5f00852",
          5599 => x"8851ffb3",
          5600 => x"ed3f84d1",
          5601 => x"d033ff05",
          5602 => x"557484d1",
          5603 => x"d0347481",
          5604 => x"ff0655c7",
          5605 => x"3984d1d0",
          5606 => x"337081ff",
          5607 => x"0684d1cc",
          5608 => x"335b5755",
          5609 => x"757927fa",
          5610 => x"af3884d5",
          5611 => x"f0085281",
          5612 => x"15577684",
          5613 => x"d1d0347b",
          5614 => x"16703352",
          5615 => x"55ffb3ae",
          5616 => x"3f84d1d0",
          5617 => x"337081ff",
          5618 => x"0684d1cc",
          5619 => x"335a5755",
          5620 => x"757827fa",
          5621 => x"833884d5",
          5622 => x"f0085281",
          5623 => x"15577684",
          5624 => x"d1d0347b",
          5625 => x"16703352",
          5626 => x"55ffb382",
          5627 => x"3f84d1d0",
          5628 => x"337081ff",
          5629 => x"0684d1cc",
          5630 => x"335a5755",
          5631 => x"777626ff",
          5632 => x"a938f9d4",
          5633 => x"3984d1d0",
          5634 => x"3384d1cc",
          5635 => x"33565674",
          5636 => x"762ef9c4",
          5637 => x"38ff155b",
          5638 => x"7a84d1cc",
          5639 => x"3475982b",
          5640 => x"70982c7c",
          5641 => x"81ff0643",
          5642 => x"575a6076",
          5643 => x"2480ef38",
          5644 => x"84d5f008",
          5645 => x"52a051ff",
          5646 => x"b2b43f84",
          5647 => x"d1d03370",
          5648 => x"982b7098",
          5649 => x"2c84d1cc",
          5650 => x"335a5757",
          5651 => x"41747724",
          5652 => x"f9863884",
          5653 => x"d5f00852",
          5654 => x"8851ffb2",
          5655 => x"913f7481",
          5656 => x"800a2981",
          5657 => x"800a0570",
          5658 => x"982c84d1",
          5659 => x"cc335d56",
          5660 => x"5a747b24",
          5661 => x"f8e23884",
          5662 => x"d5f00852",
          5663 => x"8851ffb1",
          5664 => x"ed3f7481",
          5665 => x"800a2981",
          5666 => x"800a0570",
          5667 => x"982c84d1",
          5668 => x"cc335d56",
          5669 => x"5a7a7525",
          5670 => x"ffb938f8",
          5671 => x"bb397b16",
          5672 => x"58811833",
          5673 => x"783484d5",
          5674 => x"f0085277",
          5675 => x"3351ffb1",
          5676 => x"bd3f7581",
          5677 => x"800a2981",
          5678 => x"800a0570",
          5679 => x"982c84d1",
          5680 => x"cc335b57",
          5681 => x"55757925",
          5682 => x"fee6387b",
          5683 => x"16588118",
          5684 => x"33783484",
          5685 => x"d5f00852",
          5686 => x"773351ff",
          5687 => x"b1903f75",
          5688 => x"81800a29",
          5689 => x"81800a05",
          5690 => x"70982c84",
          5691 => x"d1cc335b",
          5692 => x"57557876",
          5693 => x"24ffa738",
          5694 => x"feb63984",
          5695 => x"d1d03355",
          5696 => x"74802ef7",
          5697 => x"d33884d5",
          5698 => x"f0085288",
          5699 => x"51ffb0de",
          5700 => x"3f84d1d0",
          5701 => x"33ff0557",
          5702 => x"7684d1d0",
          5703 => x"347681ff",
          5704 => x"0655dd39",
          5705 => x"84d1cc33",
          5706 => x"7c055f80",
          5707 => x"7f3484d5",
          5708 => x"f008528a",
          5709 => x"51ffb0b6",
          5710 => x"3f84d1cc",
          5711 => x"527b51f4",
          5712 => x"8b3f84ba",
          5713 => x"8c0881ff",
          5714 => x"06587789",
          5715 => x"cf3884d1",
          5716 => x"cc335776",
          5717 => x"802e80d8",
          5718 => x"3883f3fc",
          5719 => x"33701010",
          5720 => x"83f3a405",
          5721 => x"7008575e",
          5722 => x"56748ba0",
          5723 => x"3875822b",
          5724 => x"87fc0683",
          5725 => x"f3a40581",
          5726 => x"18705357",
          5727 => x"5b80e8ca",
          5728 => x"3f84ba8c",
          5729 => x"087b0c83",
          5730 => x"f3fc3370",
          5731 => x"101083f3",
          5732 => x"a4057008",
          5733 => x"57414174",
          5734 => x"8bad3883",
          5735 => x"f3f80856",
          5736 => x"75802e8c",
          5737 => x"3883f3f4",
          5738 => x"33587780",
          5739 => x"2e8bbc38",
          5740 => x"800b84d1",
          5741 => x"d034800b",
          5742 => x"84d1cc34",
          5743 => x"7b84ba8c",
          5744 => x"0cb43d0d",
          5745 => x"0484d1d0",
          5746 => x"33557480",
          5747 => x"2eb63884",
          5748 => x"d5f00852",
          5749 => x"8851ffaf",
          5750 => x"953f84d5",
          5751 => x"f00852a0",
          5752 => x"51ffaf8a",
          5753 => x"3f84d5f0",
          5754 => x"08528851",
          5755 => x"ffaeff3f",
          5756 => x"84d1d033",
          5757 => x"ff055675",
          5758 => x"84d1d034",
          5759 => x"7581ff06",
          5760 => x"5574cc38",
          5761 => x"83d2b851",
          5762 => x"ff9ffd3f",
          5763 => x"800b84d1",
          5764 => x"d034800b",
          5765 => x"84d1cc34",
          5766 => x"f5be3983",
          5767 => x"7c34800b",
          5768 => x"811d3484",
          5769 => x"d1d03355",
          5770 => x"74802eb6",
          5771 => x"3884d5f0",
          5772 => x"08528851",
          5773 => x"ffaeb73f",
          5774 => x"84d5f008",
          5775 => x"52a051ff",
          5776 => x"aeac3f84",
          5777 => x"d5f00852",
          5778 => x"8851ffae",
          5779 => x"a13f84d1",
          5780 => x"d033ff05",
          5781 => x"5d7c84d1",
          5782 => x"d0347c81",
          5783 => x"ff065574",
          5784 => x"cc3883d2",
          5785 => x"b851ff9f",
          5786 => x"9f3f800b",
          5787 => x"84d1d034",
          5788 => x"800b84d1",
          5789 => x"cc347b84",
          5790 => x"ba8c0cb4",
          5791 => x"3d0d0484",
          5792 => x"d1d03370",
          5793 => x"81ff065c",
          5794 => x"567a802e",
          5795 => x"f4ca3884",
          5796 => x"d1cc33ff",
          5797 => x"05597884",
          5798 => x"d1cc34ff",
          5799 => x"16587784",
          5800 => x"d1d03484",
          5801 => x"d5f00852",
          5802 => x"8851ffad",
          5803 => x"c13f84d1",
          5804 => x"d0337098",
          5805 => x"2b70982c",
          5806 => x"84d1cc33",
          5807 => x"5a525b56",
          5808 => x"76762480",
          5809 => x"ef3884d5",
          5810 => x"f00852a0",
          5811 => x"51ffad9e",
          5812 => x"3f84d1d0",
          5813 => x"3370982b",
          5814 => x"70982c84",
          5815 => x"d1cc335d",
          5816 => x"57595674",
          5817 => x"7a24f3f0",
          5818 => x"3884d5f0",
          5819 => x"08528851",
          5820 => x"ffacfb3f",
          5821 => x"7481800a",
          5822 => x"2981800a",
          5823 => x"0570982c",
          5824 => x"84d1cc33",
          5825 => x"5b515574",
          5826 => x"7924f3cc",
          5827 => x"3884d5f0",
          5828 => x"08528851",
          5829 => x"ffacd73f",
          5830 => x"7481800a",
          5831 => x"2981800a",
          5832 => x"0570982c",
          5833 => x"84d1cc33",
          5834 => x"5b515578",
          5835 => x"7525ffb9",
          5836 => x"38f3a539",
          5837 => x"7b165781",
          5838 => x"17337734",
          5839 => x"84d5f008",
          5840 => x"52763351",
          5841 => x"ffaca73f",
          5842 => x"7581800a",
          5843 => x"2981800a",
          5844 => x"0570982c",
          5845 => x"84d1cc33",
          5846 => x"43575b75",
          5847 => x"6125fee6",
          5848 => x"387b1657",
          5849 => x"81173377",
          5850 => x"3484d5f0",
          5851 => x"08527633",
          5852 => x"51ffabfa",
          5853 => x"3f758180",
          5854 => x"0a298180",
          5855 => x"0a057098",
          5856 => x"2c84d1cc",
          5857 => x"3343575b",
          5858 => x"607624ff",
          5859 => x"a738feb6",
          5860 => x"3984d1d0",
          5861 => x"337081ff",
          5862 => x"06585876",
          5863 => x"602ef2b8",
          5864 => x"3884d1cc",
          5865 => x"33557675",
          5866 => x"27ae3874",
          5867 => x"982b7098",
          5868 => x"2c574176",
          5869 => x"7624a138",
          5870 => x"7b165b7a",
          5871 => x"33811c34",
          5872 => x"7581800a",
          5873 => x"2981ff0a",
          5874 => x"0570982c",
          5875 => x"84d1d033",
          5876 => x"52575875",
          5877 => x"7825e138",
          5878 => x"81185574",
          5879 => x"84d1d034",
          5880 => x"7781ff06",
          5881 => x"7c055ab3",
          5882 => x"3d337a34",
          5883 => x"84d1cc33",
          5884 => x"57766025",
          5885 => x"8b388117",
          5886 => x"567584d1",
          5887 => x"cc347557",
          5888 => x"84d1d033",
          5889 => x"7081800a",
          5890 => x"2981ff0a",
          5891 => x"0570982c",
          5892 => x"7981ff06",
          5893 => x"44585c58",
          5894 => x"60762481",
          5895 => x"ef387798",
          5896 => x"2b70982c",
          5897 => x"7881ff06",
          5898 => x"5c575975",
          5899 => x"7a25f1a8",
          5900 => x"3884d5f0",
          5901 => x"08528851",
          5902 => x"ffaab33f",
          5903 => x"7581800a",
          5904 => x"2981800a",
          5905 => x"0570982c",
          5906 => x"84d1cc33",
          5907 => x"57574175",
          5908 => x"7525f184",
          5909 => x"3884d5f0",
          5910 => x"08528851",
          5911 => x"ffaa8f3f",
          5912 => x"7581800a",
          5913 => x"2981800a",
          5914 => x"0570982c",
          5915 => x"84d1cc33",
          5916 => x"57574174",
          5917 => x"7624ffb9",
          5918 => x"38f0dd39",
          5919 => x"83f3a408",
          5920 => x"5675802e",
          5921 => x"f49d3875",
          5922 => x"51ffad9c",
          5923 => x"3f84ba8c",
          5924 => x"0884d1cc",
          5925 => x"3484ba8c",
          5926 => x"0881ff06",
          5927 => x"81055375",
          5928 => x"527b51ff",
          5929 => x"adc43f84",
          5930 => x"d1cc3384",
          5931 => x"d1d03356",
          5932 => x"5674802e",
          5933 => x"f4c83884",
          5934 => x"d5f00852",
          5935 => x"8851ffa9",
          5936 => x"ad3f84d5",
          5937 => x"f00852a0",
          5938 => x"51ffa9a2",
          5939 => x"3f84d5f0",
          5940 => x"08528851",
          5941 => x"ffa9973f",
          5942 => x"84d1d033",
          5943 => x"ff055b7a",
          5944 => x"84d1d034",
          5945 => x"7a81ff06",
          5946 => x"55c739a8",
          5947 => x"5180e1da",
          5948 => x"3f84ba8c",
          5949 => x"0883f3f8",
          5950 => x"0c84ba8c",
          5951 => x"0885a538",
          5952 => x"7683f3f4",
          5953 => x"3477efca",
          5954 => x"3880c339",
          5955 => x"84d5f008",
          5956 => x"527b1670",
          5957 => x"335258ff",
          5958 => x"a8d43f75",
          5959 => x"81800a29",
          5960 => x"81800a05",
          5961 => x"70982c84",
          5962 => x"d1cc3352",
          5963 => x"57577676",
          5964 => x"24da3884",
          5965 => x"d1d03370",
          5966 => x"982b7098",
          5967 => x"2c7981ff",
          5968 => x"065d585a",
          5969 => x"58757a25",
          5970 => x"ef8e38fd",
          5971 => x"e43983f3",
          5972 => x"f808802e",
          5973 => x"eefc3883",
          5974 => x"f3a45793",
          5975 => x"56760855",
          5976 => x"74bb38ff",
          5977 => x"16841858",
          5978 => x"56758025",
          5979 => x"f038800b",
          5980 => x"83f3fc34",
          5981 => x"83f3f808",
          5982 => x"5574802e",
          5983 => x"eed43874",
          5984 => x"5181e8c5",
          5985 => x"3f83f3f8",
          5986 => x"085180da",
          5987 => x"cd3f800b",
          5988 => x"83f3f80c",
          5989 => x"933db43d",
          5990 => x"5f5feebc",
          5991 => x"39745180",
          5992 => x"dab83f80",
          5993 => x"770cff16",
          5994 => x"84185856",
          5995 => x"758025ff",
          5996 => x"ac38ffba",
          5997 => x"397551ff",
          5998 => x"aaee3f84",
          5999 => x"ba8c0884",
          6000 => x"d1cc3484",
          6001 => x"ba8c0881",
          6002 => x"ff068105",
          6003 => x"5375527b",
          6004 => x"51ffab96",
          6005 => x"3f930b84",
          6006 => x"d1cc3384",
          6007 => x"d1d03357",
          6008 => x"575d7480",
          6009 => x"2ef29738",
          6010 => x"84d5f008",
          6011 => x"528851ff",
          6012 => x"a6fc3f84",
          6013 => x"d5f00852",
          6014 => x"a051ffa6",
          6015 => x"f13f84d5",
          6016 => x"f0085288",
          6017 => x"51ffa6e6",
          6018 => x"3f84d1d0",
          6019 => x"33ff055a",
          6020 => x"7984d1d0",
          6021 => x"347981ff",
          6022 => x"0655c739",
          6023 => x"807c3480",
          6024 => x"0b84d1d0",
          6025 => x"34800b84",
          6026 => x"d1cc347b",
          6027 => x"84ba8c0c",
          6028 => x"b43d0d04",
          6029 => x"7551ffa9",
          6030 => x"ef3f84ba",
          6031 => x"8c0884d1",
          6032 => x"cc3484ba",
          6033 => x"8c0881ff",
          6034 => x"06810553",
          6035 => x"75527b51",
          6036 => x"ffaa973f",
          6037 => x"811d7081",
          6038 => x"ff0684d1",
          6039 => x"cc3384d1",
          6040 => x"d0335852",
          6041 => x"5e567480",
          6042 => x"2ef19338",
          6043 => x"84d5f008",
          6044 => x"528851ff",
          6045 => x"a5f83f84",
          6046 => x"d5f00852",
          6047 => x"a051ffa5",
          6048 => x"ed3f84d5",
          6049 => x"f0085288",
          6050 => x"51ffa5e2",
          6051 => x"3f84d1d0",
          6052 => x"33ff0557",
          6053 => x"7684d1d0",
          6054 => x"347681ff",
          6055 => x"0655c739",
          6056 => x"7551ffa9",
          6057 => x"833f84ba",
          6058 => x"8c0884d1",
          6059 => x"cc3484ba",
          6060 => x"8c0881ff",
          6061 => x"06810553",
          6062 => x"75527b51",
          6063 => x"ffa9ab3f",
          6064 => x"ff1d7081",
          6065 => x"ff0684d1",
          6066 => x"cc3384d1",
          6067 => x"d0335858",
          6068 => x"5e587480",
          6069 => x"2ef0a738",
          6070 => x"84d5f008",
          6071 => x"528851ff",
          6072 => x"a58c3f84",
          6073 => x"d5f00852",
          6074 => x"a051ffa5",
          6075 => x"813f84d5",
          6076 => x"f0085288",
          6077 => x"51ffa4f6",
          6078 => x"3f84d1d0",
          6079 => x"33ff0541",
          6080 => x"6084d1d0",
          6081 => x"346081ff",
          6082 => x"0655c739",
          6083 => x"745180d7",
          6084 => x"c93f83f3",
          6085 => x"fc337082",
          6086 => x"2b87fc06",
          6087 => x"83f3a405",
          6088 => x"81197054",
          6089 => x"525c5680",
          6090 => x"dda03f84",
          6091 => x"ba8c087b",
          6092 => x"0c83f3fc",
          6093 => x"33701010",
          6094 => x"83f3a405",
          6095 => x"70085741",
          6096 => x"4174802e",
          6097 => x"f4d53875",
          6098 => x"537b5274",
          6099 => x"51ffa89a",
          6100 => x"3f83f3fc",
          6101 => x"33810570",
          6102 => x"81ff065a",
          6103 => x"56937927",
          6104 => x"82f23877",
          6105 => x"83f3fc34",
          6106 => x"f4b139b4",
          6107 => x"3dfef805",
          6108 => x"5476537b",
          6109 => x"52755181",
          6110 => x"d98f3f83",
          6111 => x"f3f80852",
          6112 => x"8a5182ba",
          6113 => x"d73f83f3",
          6114 => x"f8085181",
          6115 => x"e0c23f80",
          6116 => x"0b84d1d0",
          6117 => x"34800b84",
          6118 => x"d1cc347b",
          6119 => x"84ba8c0c",
          6120 => x"b43d0d04",
          6121 => x"93537752",
          6122 => x"84ba8c08",
          6123 => x"5181cac7",
          6124 => x"3f84ba8c",
          6125 => x"0882a538",
          6126 => x"84ba8c08",
          6127 => x"963d5c5d",
          6128 => x"83f3f808",
          6129 => x"5380f852",
          6130 => x"7a5182b8",
          6131 => x"c13f84ba",
          6132 => x"8c085a84",
          6133 => x"ba8c087b",
          6134 => x"2e098106",
          6135 => x"e9ee3884",
          6136 => x"ba8c0851",
          6137 => x"ffa6c13f",
          6138 => x"84ba8c08",
          6139 => x"56800b84",
          6140 => x"ba8c0825",
          6141 => x"80e33884",
          6142 => x"ba8c08ff",
          6143 => x"05701b58",
          6144 => x"56807734",
          6145 => x"7581ff06",
          6146 => x"83f3fc33",
          6147 => x"70101083",
          6148 => x"f3a40570",
          6149 => x"08584058",
          6150 => x"597480f2",
          6151 => x"3876822b",
          6152 => x"87fc0683",
          6153 => x"f3a40581",
          6154 => x"1a705358",
          6155 => x"5580db9a",
          6156 => x"3f84ba8c",
          6157 => x"08750c83",
          6158 => x"f3fc3370",
          6159 => x"101083f3",
          6160 => x"a4057008",
          6161 => x"57404174",
          6162 => x"a038811d",
          6163 => x"7081ff06",
          6164 => x"5e57937d",
          6165 => x"27833880",
          6166 => x"5d75ff2e",
          6167 => x"098106fe",
          6168 => x"df3877e8",
          6169 => x"ed38f9e6",
          6170 => x"39765379",
          6171 => x"527451ff",
          6172 => x"a5f83f83",
          6173 => x"f3fc3381",
          6174 => x"057081ff",
          6175 => x"065b5793",
          6176 => x"7a2780c8",
          6177 => x"38800b83",
          6178 => x"f3fc34ff",
          6179 => x"bd397451",
          6180 => x"80d4c73f",
          6181 => x"83f3fc33",
          6182 => x"70822b87",
          6183 => x"fc0683f3",
          6184 => x"a405811b",
          6185 => x"70545256",
          6186 => x"5780da9e",
          6187 => x"3f84ba8c",
          6188 => x"08750c83",
          6189 => x"f3fc3370",
          6190 => x"101083f3",
          6191 => x"a4057008",
          6192 => x"57404174",
          6193 => x"802eff82",
          6194 => x"38ff9e39",
          6195 => x"7683f3fc",
          6196 => x"34fef739",
          6197 => x"7583f3fc",
          6198 => x"34f1c039",
          6199 => x"83e1b851",
          6200 => x"ff9f903f",
          6201 => x"77e7eb38",
          6202 => x"f8e439f2",
          6203 => x"3d0d0280",
          6204 => x"c3053302",
          6205 => x"840580c7",
          6206 => x"05335b53",
          6207 => x"72832681",
          6208 => x"8d387281",
          6209 => x"2e818b38",
          6210 => x"81732583",
          6211 => x"9e387282",
          6212 => x"2e82a838",
          6213 => x"87a3a080",
          6214 => x"5987a3b0",
          6215 => x"80705e57",
          6216 => x"80569fa0",
          6217 => x"5879762e",
          6218 => x"90387583",
          6219 => x"f9bc3475",
          6220 => x"83f9bd34",
          6221 => x"7583f9ba",
          6222 => x"2383f9b8",
          6223 => x"3370982b",
          6224 => x"71902b07",
          6225 => x"71882b07",
          6226 => x"71077a7f",
          6227 => x"5656565b",
          6228 => x"78772794",
          6229 => x"38807470",
          6230 => x"8405560c",
          6231 => x"74737084",
          6232 => x"05550c76",
          6233 => x"7426ee38",
          6234 => x"757827a2",
          6235 => x"3883f9b8",
          6236 => x"338498de",
          6237 => x"17797831",
          6238 => x"555555a0",
          6239 => x"0be0e015",
          6240 => x"34747470",
          6241 => x"81055634",
          6242 => x"ff135372",
          6243 => x"ee38903d",
          6244 => x"0d0487a3",
          6245 => x"a0800b83",
          6246 => x"f9bc3370",
          6247 => x"10101183",
          6248 => x"f9bd3371",
          6249 => x"90291174",
          6250 => x"055b4158",
          6251 => x"405987a3",
          6252 => x"b0800b84",
          6253 => x"b8803370",
          6254 => x"81ff0684",
          6255 => x"b7ff3370",
          6256 => x"81ff0683",
          6257 => x"f9ba2270",
          6258 => x"83ffff06",
          6259 => x"7075295d",
          6260 => x"595d585e",
          6261 => x"575b5d73",
          6262 => x"73268738",
          6263 => x"72743175",
          6264 => x"29567981",
          6265 => x"ff067e81",
          6266 => x"ff067c81",
          6267 => x"ff067a83",
          6268 => x"ffff0662",
          6269 => x"81ff0670",
          6270 => x"7529145d",
          6271 => x"4257575b",
          6272 => x"5c747426",
          6273 => x"8f3883f9",
          6274 => x"bc337476",
          6275 => x"3105707d",
          6276 => x"291b595f",
          6277 => x"7683065c",
          6278 => x"7b802efe",
          6279 => x"9c38787d",
          6280 => x"55537277",
          6281 => x"26fec138",
          6282 => x"80737081",
          6283 => x"05553483",
          6284 => x"f9b83374",
          6285 => x"70810556",
          6286 => x"34e83987",
          6287 => x"a3a08059",
          6288 => x"87a3b080",
          6289 => x"7084b880",
          6290 => x"337081ff",
          6291 => x"0684b7ff",
          6292 => x"337081ff",
          6293 => x"0683f9ba",
          6294 => x"22707429",
          6295 => x"5d5b5d57",
          6296 => x"5e565e57",
          6297 => x"74782781",
          6298 => x"df387381",
          6299 => x"ff067381",
          6300 => x"ff067171",
          6301 => x"29185a54",
          6302 => x"5479802e",
          6303 => x"fdbb3880",
          6304 => x"0b83f9bc",
          6305 => x"34800b83",
          6306 => x"f9bd3483",
          6307 => x"f9b83370",
          6308 => x"982b7190",
          6309 => x"2b077188",
          6310 => x"2b077107",
          6311 => x"7a7f5656",
          6312 => x"565b7679",
          6313 => x"26fdae38",
          6314 => x"fdbe3972",
          6315 => x"fce63883",
          6316 => x"f9bc3370",
          6317 => x"81ff0670",
          6318 => x"10101183",
          6319 => x"f9bd3371",
          6320 => x"90291187",
          6321 => x"a3a08011",
          6322 => x"5e575b56",
          6323 => x"565f87a3",
          6324 => x"b0807014",
          6325 => x"84b88033",
          6326 => x"7081ff06",
          6327 => x"84b7ff33",
          6328 => x"7081ff06",
          6329 => x"83f9ba22",
          6330 => x"7083ffff",
          6331 => x"067c7529",
          6332 => x"60055e5a",
          6333 => x"415f585f",
          6334 => x"405e5779",
          6335 => x"73268b38",
          6336 => x"727a3115",
          6337 => x"707d2919",
          6338 => x"57537d81",
          6339 => x"ff067481",
          6340 => x"ff067171",
          6341 => x"297d83ff",
          6342 => x"ff066281",
          6343 => x"ff067075",
          6344 => x"29585f5b",
          6345 => x"5c5d557b",
          6346 => x"78268538",
          6347 => x"77752953",
          6348 => x"79733116",
          6349 => x"7983065b",
          6350 => x"5879fde2",
          6351 => x"38768306",
          6352 => x"5c7bfdda",
          6353 => x"38fbf239",
          6354 => x"7478317b",
          6355 => x"2956fe9a",
          6356 => x"39fb3d0d",
          6357 => x"86ee809c",
          6358 => x"5480f474",
          6359 => x"34ffb074",
          6360 => x"3486ee80",
          6361 => x"98538073",
          6362 => x"34807334",
          6363 => x"86ee8094",
          6364 => x"568a7634",
          6365 => x"807634ff",
          6366 => x"80743486",
          6367 => x"ee808c55",
          6368 => x"ff8a7534",
          6369 => x"87753485",
          6370 => x"75348175",
          6371 => x"34815283",
          6372 => x"51fad83f",
          6373 => x"879087e0",
          6374 => x"70085454",
          6375 => x"81f85687",
          6376 => x"8c81f873",
          6377 => x"77068407",
          6378 => x"54557275",
          6379 => x"34730870",
          6380 => x"80ff0680",
          6381 => x"c0075153",
          6382 => x"72753487",
          6383 => x"9087cc08",
          6384 => x"70770681",
          6385 => x"07515372",
          6386 => x"878c81f3",
          6387 => x"34730881",
          6388 => x"f7068807",
          6389 => x"53727534",
          6390 => x"80d00b84",
          6391 => x"b8803480",
          6392 => x"0b84ba8c",
          6393 => x"0c873d0d",
          6394 => x"0484b880",
          6395 => x"3384ba8c",
          6396 => x"0c04f73d",
          6397 => x"0d02af05",
          6398 => x"33028405",
          6399 => x"b3053384",
          6400 => x"b7ff335b",
          6401 => x"59568153",
          6402 => x"75792682",
          6403 => x"da3884b8",
          6404 => x"803383f9",
          6405 => x"bd3383f9",
          6406 => x"bc337271",
          6407 => x"291287a3",
          6408 => x"a0801183",
          6409 => x"f9ba225f",
          6410 => x"51575971",
          6411 => x"7c290570",
          6412 => x"83ffff06",
          6413 => x"83f89233",
          6414 => x"53575853",
          6415 => x"72812e83",
          6416 => x"c43883f9",
          6417 => x"ba227605",
          6418 => x"557483f9",
          6419 => x"ba2383f9",
          6420 => x"bc337605",
          6421 => x"7081ff06",
          6422 => x"7a81ff06",
          6423 => x"555b5572",
          6424 => x"7a26828c",
          6425 => x"38ff1953",
          6426 => x"7283f9bc",
          6427 => x"3483f9ba",
          6428 => x"227083ff",
          6429 => x"ff0684b7",
          6430 => x"fe335c55",
          6431 => x"57797426",
          6432 => x"82893884",
          6433 => x"b8803376",
          6434 => x"71295458",
          6435 => x"8054729f",
          6436 => x"9f26ac38",
          6437 => x"8498de70",
          6438 => x"145455e0",
          6439 => x"e01333e0",
          6440 => x"e0163472",
          6441 => x"70810554",
          6442 => x"33757081",
          6443 => x"05573481",
          6444 => x"145484b7",
          6445 => x"fd7327e3",
          6446 => x"38739f9f",
          6447 => x"26a13883",
          6448 => x"f9b83384",
          6449 => x"98de1554",
          6450 => x"55a00be0",
          6451 => x"e0143474",
          6452 => x"73708105",
          6453 => x"55348114",
          6454 => x"549f9f74",
          6455 => x"27eb3884",
          6456 => x"b7fe33ff",
          6457 => x"05567583",
          6458 => x"f9ba2375",
          6459 => x"577881ff",
          6460 => x"067783ff",
          6461 => x"ff065454",
          6462 => x"73732681",
          6463 => x"fd387274",
          6464 => x"31810584",
          6465 => x"b8803371",
          6466 => x"71295855",
          6467 => x"57755587",
          6468 => x"a3a08058",
          6469 => x"87a3b080",
          6470 => x"7981ff06",
          6471 => x"7581ff06",
          6472 => x"71712919",
          6473 => x"5c5c5457",
          6474 => x"757927b9",
          6475 => x"388498de",
          6476 => x"1654e0e0",
          6477 => x"14335384",
          6478 => x"b8881333",
          6479 => x"78708105",
          6480 => x"5a347370",
          6481 => x"81055533",
          6482 => x"77708105",
          6483 => x"59348115",
          6484 => x"84b88033",
          6485 => x"84b7ff33",
          6486 => x"71712919",
          6487 => x"565c5a55",
          6488 => x"727526ce",
          6489 => x"38805372",
          6490 => x"84ba8c0c",
          6491 => x"8b3d0d04",
          6492 => x"7483f9bc",
          6493 => x"3483f9ba",
          6494 => x"227083ff",
          6495 => x"ff0684b7",
          6496 => x"fe335c55",
          6497 => x"57737a27",
          6498 => x"fdf93877",
          6499 => x"802efedd",
          6500 => x"387881ff",
          6501 => x"06ff0583",
          6502 => x"f9bc3356",
          6503 => x"5372752e",
          6504 => x"098106fe",
          6505 => x"c8387376",
          6506 => x"31810584",
          6507 => x"b8803371",
          6508 => x"71297872",
          6509 => x"29115652",
          6510 => x"59547373",
          6511 => x"27feae38",
          6512 => x"83f9b833",
          6513 => x"8498de15",
          6514 => x"74763155",
          6515 => x"5656a00b",
          6516 => x"e0e01634",
          6517 => x"75757081",
          6518 => x"055734ff",
          6519 => x"13537280",
          6520 => x"2efe8a38",
          6521 => x"a00be0e0",
          6522 => x"16347575",
          6523 => x"70810557",
          6524 => x"34ff1353",
          6525 => x"72d838fd",
          6526 => x"f439800b",
          6527 => x"84b88033",
          6528 => x"5556fe89",
          6529 => x"3983f9be",
          6530 => x"15335984",
          6531 => x"b8881933",
          6532 => x"743484b7",
          6533 => x"ff3359fc",
          6534 => x"a939fc3d",
          6535 => x"0d760284",
          6536 => x"059f0533",
          6537 => x"53517086",
          6538 => x"269b3870",
          6539 => x"101083c4",
          6540 => x"b4055170",
          6541 => x"080484b8",
          6542 => x"80335171",
          6543 => x"71278638",
          6544 => x"7183f9bd",
          6545 => x"34800b84",
          6546 => x"ba8c0c86",
          6547 => x"3d0d0480",
          6548 => x"0b83f9bd",
          6549 => x"3483f9bc",
          6550 => x"337081ff",
          6551 => x"06545272",
          6552 => x"802ee238",
          6553 => x"ff125170",
          6554 => x"83f9bc34",
          6555 => x"800b84ba",
          6556 => x"8c0c863d",
          6557 => x"0d0483f9",
          6558 => x"bc337073",
          6559 => x"31700970",
          6560 => x"9f2c7206",
          6561 => x"54555354",
          6562 => x"7083f9bc",
          6563 => x"34de3983",
          6564 => x"f9bc3372",
          6565 => x"0584b7ff",
          6566 => x"33ff1155",
          6567 => x"56517075",
          6568 => x"25833870",
          6569 => x"537283f9",
          6570 => x"bc34800b",
          6571 => x"84ba8c0c",
          6572 => x"863d0d04",
          6573 => x"83f9bd33",
          6574 => x"70733170",
          6575 => x"09709f2c",
          6576 => x"72065456",
          6577 => x"53557083",
          6578 => x"f9bd3480",
          6579 => x"0b84ba8c",
          6580 => x"0c863d0d",
          6581 => x"0483f9bd",
          6582 => x"33720584",
          6583 => x"b88033ff",
          6584 => x"11555551",
          6585 => x"70742583",
          6586 => x"38705372",
          6587 => x"83f9bd34",
          6588 => x"800b84ba",
          6589 => x"8c0c863d",
          6590 => x"0d04800b",
          6591 => x"83f9bd34",
          6592 => x"83f9bc33",
          6593 => x"84b7ff33",
          6594 => x"ff055652",
          6595 => x"717525fe",
          6596 => x"b4388112",
          6597 => x"517083f9",
          6598 => x"bc34fed0",
          6599 => x"39ff3d0d",
          6600 => x"028f0533",
          6601 => x"5170b126",
          6602 => x"b3387010",
          6603 => x"1083c4d0",
          6604 => x"05517008",
          6605 => x"0483f9b8",
          6606 => x"337080f0",
          6607 => x"0671842b",
          6608 => x"80f00670",
          6609 => x"72842a07",
          6610 => x"51525351",
          6611 => x"7180f02e",
          6612 => x"0981069c",
          6613 => x"3880f20b",
          6614 => x"83f9b834",
          6615 => x"800b84ba",
          6616 => x"8c0c833d",
          6617 => x"0d0483f9",
          6618 => x"b833819f",
          6619 => x"06900751",
          6620 => x"7083f9b8",
          6621 => x"34800b84",
          6622 => x"ba8c0c83",
          6623 => x"3d0d0483",
          6624 => x"f9b83380",
          6625 => x"f0075170",
          6626 => x"83f9b834",
          6627 => x"e83983f9",
          6628 => x"b83381fe",
          6629 => x"06860751",
          6630 => x"7083f9b8",
          6631 => x"34d73980",
          6632 => x"f10b83f9",
          6633 => x"b834800b",
          6634 => x"84ba8c0c",
          6635 => x"833d0d04",
          6636 => x"83f9b833",
          6637 => x"81fc0684",
          6638 => x"07517083",
          6639 => x"f9b834ff",
          6640 => x"b43983f9",
          6641 => x"b8338707",
          6642 => x"517083f9",
          6643 => x"b834ffa5",
          6644 => x"3983f9b8",
          6645 => x"3381fd06",
          6646 => x"85075170",
          6647 => x"83f9b834",
          6648 => x"ff933983",
          6649 => x"f9b83381",
          6650 => x"fb068307",
          6651 => x"517083f9",
          6652 => x"b834ff81",
          6653 => x"3983f9b8",
          6654 => x"3381f906",
          6655 => x"81075170",
          6656 => x"83f9b834",
          6657 => x"feef3983",
          6658 => x"f9b83381",
          6659 => x"f8065170",
          6660 => x"83f9b834",
          6661 => x"fedf3983",
          6662 => x"f9b83381",
          6663 => x"df0680d0",
          6664 => x"07517083",
          6665 => x"f9b834fe",
          6666 => x"cc3983f9",
          6667 => x"b83381bf",
          6668 => x"06b00751",
          6669 => x"7083f9b8",
          6670 => x"34feba39",
          6671 => x"83f9b833",
          6672 => x"81ef0680",
          6673 => x"e0075170",
          6674 => x"83f9b834",
          6675 => x"fea73983",
          6676 => x"f9b83381",
          6677 => x"cf0680c0",
          6678 => x"07517083",
          6679 => x"f9b834fe",
          6680 => x"943983f9",
          6681 => x"b83381af",
          6682 => x"06a00751",
          6683 => x"7083f9b8",
          6684 => x"34fe8239",
          6685 => x"83f9b833",
          6686 => x"818f0651",
          6687 => x"7083f9b8",
          6688 => x"34fdf239",
          6689 => x"83f9b833",
          6690 => x"81fa0682",
          6691 => x"07517083",
          6692 => x"f9b834fd",
          6693 => x"e039f33d",
          6694 => x"0d02bf05",
          6695 => x"33028405",
          6696 => x"80c30533",
          6697 => x"83f9bc33",
          6698 => x"83f9bb33",
          6699 => x"83f9bd33",
          6700 => x"84b88233",
          6701 => x"43415f5d",
          6702 => x"5b597882",
          6703 => x"2e82a138",
          6704 => x"788224a5",
          6705 => x"3878812e",
          6706 => x"8182387d",
          6707 => x"84b88234",
          6708 => x"800b84b8",
          6709 => x"84347a83",
          6710 => x"f9bc347b",
          6711 => x"83f9ba23",
          6712 => x"7c83f9bd",
          6713 => x"348f3d0d",
          6714 => x"0478832e",
          6715 => x"098106db",
          6716 => x"38800b84",
          6717 => x"b8823481",
          6718 => x"0b84b884",
          6719 => x"34820b83",
          6720 => x"f9bc34a8",
          6721 => x"0b83f9bd",
          6722 => x"34820b83",
          6723 => x"f9ba2379",
          6724 => x"5884b880",
          6725 => x"335784b7",
          6726 => x"ff335684",
          6727 => x"b7fe3355",
          6728 => x"7b547c53",
          6729 => x"7a5283e3",
          6730 => x"c451ff81",
          6731 => x"db3f7d84",
          6732 => x"b8823480",
          6733 => x"0b84b884",
          6734 => x"347a83f9",
          6735 => x"bc347b83",
          6736 => x"f9ba237c",
          6737 => x"83f9bd34",
          6738 => x"8f3d0d04",
          6739 => x"800b84b8",
          6740 => x"8234810b",
          6741 => x"84b88434",
          6742 => x"800b83f9",
          6743 => x"bc34a80b",
          6744 => x"83f9bd34",
          6745 => x"800b83f9",
          6746 => x"ba2384b9",
          6747 => x"8f335884",
          6748 => x"b98e3357",
          6749 => x"84b98d33",
          6750 => x"5679557b",
          6751 => x"547c537a",
          6752 => x"5283e3e0",
          6753 => x"51ff8180",
          6754 => x"3f800b84",
          6755 => x"b98d335a",
          6756 => x"5a797927",
          6757 => x"a5387910",
          6758 => x"84b9e005",
          6759 => x"70225359",
          6760 => x"83e3f851",
          6761 => x"ff80e13f",
          6762 => x"811a7081",
          6763 => x"ff0684b9",
          6764 => x"8d33525b",
          6765 => x"59787a26",
          6766 => x"dd3883d2",
          6767 => x"ec51ff80",
          6768 => x"c73f7d84",
          6769 => x"b8823480",
          6770 => x"0b84b884",
          6771 => x"347a83f9",
          6772 => x"bc347b83",
          6773 => x"f9ba237c",
          6774 => x"83f9bd34",
          6775 => x"8f3d0d04",
          6776 => x"800b84b8",
          6777 => x"8234810b",
          6778 => x"84b88434",
          6779 => x"810b83f9",
          6780 => x"bc34a80b",
          6781 => x"83f9bd34",
          6782 => x"810b83f9",
          6783 => x"ba2383f7",
          6784 => x"f051ff92",
          6785 => x"a33f84ba",
          6786 => x"8c085283",
          6787 => x"e3fc51fe",
          6788 => x"fff63f80",
          6789 => x"5983f7f0",
          6790 => x"51ff928c",
          6791 => x"3f7884ba",
          6792 => x"8c0827fd",
          6793 => x"a63883f7",
          6794 => x"f0193352",
          6795 => x"83e48451",
          6796 => x"feffd53f",
          6797 => x"81197081",
          6798 => x"ff065a5a",
          6799 => x"d839f93d",
          6800 => x"0d7a0284",
          6801 => x"05a70533",
          6802 => x"84b88033",
          6803 => x"83f9bd33",
          6804 => x"83f9bc33",
          6805 => x"72712912",
          6806 => x"87a3a080",
          6807 => x"1183f9ba",
          6808 => x"22535159",
          6809 => x"5c717c29",
          6810 => x"057083ff",
          6811 => x"ff0683f8",
          6812 => x"92335259",
          6813 => x"51555757",
          6814 => x"72812e81",
          6815 => x"e9387589",
          6816 => x"2e81f938",
          6817 => x"75892481",
          6818 => x"b9387581",
          6819 => x"2e838538",
          6820 => x"75882e82",
          6821 => x"d53884b8",
          6822 => x"803383f9",
          6823 => x"bc3383f9",
          6824 => x"bd337272",
          6825 => x"29055556",
          6826 => x"5484b888",
          6827 => x"163387a3",
          6828 => x"a0801434",
          6829 => x"84b88033",
          6830 => x"83f9bd33",
          6831 => x"83f9ba22",
          6832 => x"72712912",
          6833 => x"5a5a5653",
          6834 => x"7583f9be",
          6835 => x"183483f9",
          6836 => x"bc337371",
          6837 => x"29165854",
          6838 => x"83f9b833",
          6839 => x"87a3b080",
          6840 => x"183484b8",
          6841 => x"80337081",
          6842 => x"ff0683f9",
          6843 => x"ba2283f9",
          6844 => x"bd337272",
          6845 => x"2911575b",
          6846 => x"57555783",
          6847 => x"f9b83384",
          6848 => x"98de1434",
          6849 => x"81187081",
          6850 => x"ff065955",
          6851 => x"73782681",
          6852 => x"993884b8",
          6853 => x"81335877",
          6854 => x"81ea38ff",
          6855 => x"17537283",
          6856 => x"f9bd3484",
          6857 => x"b8833353",
          6858 => x"72802e8c",
          6859 => x"3884b884",
          6860 => x"33577680",
          6861 => x"2e80fb38",
          6862 => x"800b84ba",
          6863 => x"8c0c893d",
          6864 => x"0d04758d",
          6865 => x"2e973875",
          6866 => x"8d2480f7",
          6867 => x"38758a2e",
          6868 => x"098106fe",
          6869 => x"c1388152",
          6870 => x"8151f196",
          6871 => x"3f800b83",
          6872 => x"f9bd34ff",
          6873 => x"be3983f9",
          6874 => x"be153353",
          6875 => x"84b88813",
          6876 => x"33743475",
          6877 => x"892e0981",
          6878 => x"06fe8938",
          6879 => x"80537652",
          6880 => x"a051fdba",
          6881 => x"3f811370",
          6882 => x"81ff0654",
          6883 => x"54728326",
          6884 => x"ff913876",
          6885 => x"52a051fd",
          6886 => x"a53f8113",
          6887 => x"7081ff06",
          6888 => x"54548373",
          6889 => x"27d838fe",
          6890 => x"fa397483",
          6891 => x"f9bd34fe",
          6892 => x"f2397552",
          6893 => x"8351f9de",
          6894 => x"3f800b84",
          6895 => x"ba8c0c89",
          6896 => x"3d0d0475",
          6897 => x"80ff2e09",
          6898 => x"8106fdca",
          6899 => x"3883f9bd",
          6900 => x"337081ff",
          6901 => x"0655ff05",
          6902 => x"53738338",
          6903 => x"73537283",
          6904 => x"f9bd3476",
          6905 => x"52a051fc",
          6906 => x"d53f83f9",
          6907 => x"bd337081",
          6908 => x"ff0655ff",
          6909 => x"055373fe",
          6910 => x"a5387353",
          6911 => x"7283f9bd",
          6912 => x"34fea039",
          6913 => x"800b83f9",
          6914 => x"bd348152",
          6915 => x"8151efe2",
          6916 => x"3ffe9039",
          6917 => x"80527551",
          6918 => x"efd83ffe",
          6919 => x"8639e63d",
          6920 => x"0d0280f3",
          6921 => x"053384b9",
          6922 => x"88085759",
          6923 => x"75812e81",
          6924 => x"b8387582",
          6925 => x"2e838238",
          6926 => x"788a2e84",
          6927 => x"b538788a",
          6928 => x"2482d138",
          6929 => x"78882e84",
          6930 => x"b9387889",
          6931 => x"2e888f38",
          6932 => x"84b88033",
          6933 => x"83f9bc33",
          6934 => x"83f9bd33",
          6935 => x"72722905",
          6936 => x"585e5c84",
          6937 => x"b8881933",
          6938 => x"87a3a080",
          6939 => x"173484b8",
          6940 => x"803383f9",
          6941 => x"bd3383f9",
          6942 => x"ba227271",
          6943 => x"29125a5a",
          6944 => x"42407883",
          6945 => x"f9be1834",
          6946 => x"83f9bc33",
          6947 => x"60712962",
          6948 => x"05405a83",
          6949 => x"f9b8337f",
          6950 => x"87a3b080",
          6951 => x"053484b8",
          6952 => x"80337081",
          6953 => x"ff0683f9",
          6954 => x"ba2283f9",
          6955 => x"bd337272",
          6956 => x"29114240",
          6957 => x"5d585983",
          6958 => x"f9b83384",
          6959 => x"98de1f34",
          6960 => x"811d7081",
          6961 => x"ff064258",
          6962 => x"76612681",
          6963 => x"b83884b8",
          6964 => x"81335a79",
          6965 => x"86f138ff",
          6966 => x"19567583",
          6967 => x"f9bd3480",
          6968 => x"0b84ba8c",
          6969 => x"0c9c3d0d",
          6970 => x"0478b72e",
          6971 => x"848a38b7",
          6972 => x"792581fd",
          6973 => x"3878b82e",
          6974 => x"9bb33878",
          6975 => x"80db2e89",
          6976 => x"cc38800b",
          6977 => x"84b9880c",
          6978 => x"84b88033",
          6979 => x"83f9bc33",
          6980 => x"83f9bd33",
          6981 => x"72722905",
          6982 => x"5e404084",
          6983 => x"b8881933",
          6984 => x"87a3a080",
          6985 => x"1d3484b8",
          6986 => x"803383f9",
          6987 => x"bd3383f9",
          6988 => x"ba227271",
          6989 => x"2912415f",
          6990 => x"59567883",
          6991 => x"f9be1f34",
          6992 => x"83f9bc33",
          6993 => x"76712919",
          6994 => x"5b5783f9",
          6995 => x"b83387a3",
          6996 => x"b0801b34",
          6997 => x"84b88033",
          6998 => x"7081ff06",
          6999 => x"83f9ba22",
          7000 => x"83f9bd33",
          7001 => x"72722911",
          7002 => x"44424358",
          7003 => x"5983f9b8",
          7004 => x"33608498",
          7005 => x"de053481",
          7006 => x"1f587781",
          7007 => x"ff064160",
          7008 => x"7727feca",
          7009 => x"387783f9",
          7010 => x"bd34800b",
          7011 => x"84ba8c0c",
          7012 => x"9c3d0d04",
          7013 => x"789b2e82",
          7014 => x"b738789b",
          7015 => x"24838138",
          7016 => x"788d2e09",
          7017 => x"8106fda8",
          7018 => x"38800b83",
          7019 => x"f9bd3480",
          7020 => x"0b84ba8c",
          7021 => x"0c9c3d0d",
          7022 => x"04789b2e",
          7023 => x"82aa38d0",
          7024 => x"19567589",
          7025 => x"2684d038",
          7026 => x"84b98c33",
          7027 => x"81115957",
          7028 => x"7784b98c",
          7029 => x"347884b9",
          7030 => x"90183477",
          7031 => x"81ff0659",
          7032 => x"800b84b9",
          7033 => x"901a3480",
          7034 => x"0b84ba8c",
          7035 => x"0c9c3d0d",
          7036 => x"04789b2e",
          7037 => x"fde93880",
          7038 => x"0b84b988",
          7039 => x"0c84b880",
          7040 => x"3383f9bc",
          7041 => x"3383f9bd",
          7042 => x"33727229",
          7043 => x"055e4040",
          7044 => x"84b88819",
          7045 => x"3387a3a0",
          7046 => x"801d3484",
          7047 => x"b8803383",
          7048 => x"f9bd3383",
          7049 => x"f9ba2272",
          7050 => x"71291241",
          7051 => x"5f595678",
          7052 => x"83f9be1f",
          7053 => x"3483f9bc",
          7054 => x"33767129",
          7055 => x"195b5783",
          7056 => x"f9b83387",
          7057 => x"a3b0801b",
          7058 => x"3484b880",
          7059 => x"337081ff",
          7060 => x"0683f9ba",
          7061 => x"2283f9bd",
          7062 => x"33727229",
          7063 => x"11444243",
          7064 => x"585983f9",
          7065 => x"b8336084",
          7066 => x"98de0534",
          7067 => x"811f58fe",
          7068 => x"89398152",
          7069 => x"8151eafa",
          7070 => x"3f800b83",
          7071 => x"f9bd34fe",
          7072 => x"ae3984b8",
          7073 => x"803383f9",
          7074 => x"bd337081",
          7075 => x"ff0683f9",
          7076 => x"bc337371",
          7077 => x"291287a3",
          7078 => x"a0800583",
          7079 => x"f9ba2240",
          7080 => x"515d727e",
          7081 => x"29057083",
          7082 => x"ffff0683",
          7083 => x"f892335a",
          7084 => x"51595a5c",
          7085 => x"75812e86",
          7086 => x"a4387881",
          7087 => x"ff06ff1a",
          7088 => x"575776fc",
          7089 => x"95387656",
          7090 => x"7583f9bd",
          7091 => x"34fc9039",
          7092 => x"800b84b9",
          7093 => x"8c34800b",
          7094 => x"84b98d34",
          7095 => x"800b84b9",
          7096 => x"8e34800b",
          7097 => x"84b98f34",
          7098 => x"810b84b9",
          7099 => x"880c800b",
          7100 => x"84ba8c0c",
          7101 => x"9c3d0d04",
          7102 => x"83f9bc33",
          7103 => x"84b9f434",
          7104 => x"83f9bd33",
          7105 => x"84b9f534",
          7106 => x"83f9bb33",
          7107 => x"84b9f634",
          7108 => x"800b84b9",
          7109 => x"880c800b",
          7110 => x"84ba8c0c",
          7111 => x"9c3d0d04",
          7112 => x"7880ff2e",
          7113 => x"098106fa",
          7114 => x"a73883f9",
          7115 => x"bc3384b8",
          7116 => x"80337081",
          7117 => x"ff0683f9",
          7118 => x"bd337081",
          7119 => x"ff067275",
          7120 => x"291187a3",
          7121 => x"a0800583",
          7122 => x"f9ba225c",
          7123 => x"40727b29",
          7124 => x"057083ff",
          7125 => x"ff0683f8",
          7126 => x"9233445c",
          7127 => x"435c425b",
          7128 => x"5c7d812e",
          7129 => x"85fe3878",
          7130 => x"81ff06ff",
          7131 => x"1a585675",
          7132 => x"83387557",
          7133 => x"7683f9bd",
          7134 => x"347b81ff",
          7135 => x"067a81ff",
          7136 => x"067881ff",
          7137 => x"06727229",
          7138 => x"055f405b",
          7139 => x"84b8a833",
          7140 => x"87a3a080",
          7141 => x"1e3484b8",
          7142 => x"803383f9",
          7143 => x"bd3383f9",
          7144 => x"ba227271",
          7145 => x"29125a5e",
          7146 => x"4240a00b",
          7147 => x"83f9be18",
          7148 => x"3483f9bc",
          7149 => x"33607129",
          7150 => x"62055a56",
          7151 => x"83f9b833",
          7152 => x"87a3b080",
          7153 => x"1a3484b8",
          7154 => x"80337081",
          7155 => x"ff0683f9",
          7156 => x"ba2283f9",
          7157 => x"bd337272",
          7158 => x"2911435d",
          7159 => x"5a5e5983",
          7160 => x"f9b8337f",
          7161 => x"8498de05",
          7162 => x"34811a70",
          7163 => x"81ff065c",
          7164 => x"587c7b26",
          7165 => x"95ea3884",
          7166 => x"b881335a",
          7167 => x"7996d038",
          7168 => x"ff195877",
          7169 => x"83f9bd34",
          7170 => x"83f9bd33",
          7171 => x"7081ff06",
          7172 => x"58ff0556",
          7173 => x"fdac3978",
          7174 => x"bb2e95d8",
          7175 => x"3878bd2e",
          7176 => x"83d73878",
          7177 => x"bf2e95a8",
          7178 => x"3884b98c",
          7179 => x"335f7e83",
          7180 => x"f938ffbf",
          7181 => x"195675b4",
          7182 => x"2684c838",
          7183 => x"75101083",
          7184 => x"c6980558",
          7185 => x"77080480",
          7186 => x"0b83f9bd",
          7187 => x"34805281",
          7188 => x"51e79f3f",
          7189 => x"800b84ba",
          7190 => x"8c0c9c3d",
          7191 => x"0d0483f9",
          7192 => x"bc3384b8",
          7193 => x"80337081",
          7194 => x"ff0683f9",
          7195 => x"bd337081",
          7196 => x"ff067275",
          7197 => x"291187a3",
          7198 => x"a0800583",
          7199 => x"f9ba225c",
          7200 => x"41727b29",
          7201 => x"057083ff",
          7202 => x"ff0683f8",
          7203 => x"92334653",
          7204 => x"455c595b",
          7205 => x"5b7f812e",
          7206 => x"82ef3880",
          7207 => x"5c7a81ff",
          7208 => x"067a81ff",
          7209 => x"067a81ff",
          7210 => x"06727229",
          7211 => x"055c5840",
          7212 => x"84b8a833",
          7213 => x"87a3a080",
          7214 => x"1b3484b8",
          7215 => x"803383f9",
          7216 => x"bd3383f9",
          7217 => x"ba227271",
          7218 => x"29125e41",
          7219 => x"5e56a00b",
          7220 => x"83f9be1c",
          7221 => x"3483f9bc",
          7222 => x"33767129",
          7223 => x"1e5a5e83",
          7224 => x"f9b83387",
          7225 => x"a3b0801a",
          7226 => x"3484b880",
          7227 => x"337081ff",
          7228 => x"0683f9ba",
          7229 => x"2283f9bd",
          7230 => x"33727229",
          7231 => x"115b445a",
          7232 => x"405983f9",
          7233 => x"b8338498",
          7234 => x"de183460",
          7235 => x"81057081",
          7236 => x"ff065b58",
          7237 => x"7e7a2681",
          7238 => x"ac3884b8",
          7239 => x"81335877",
          7240 => x"92fb38ff",
          7241 => x"19567583",
          7242 => x"f9bd3481",
          7243 => x"1c7081ff",
          7244 => x"065d597b",
          7245 => x"8326f7a7",
          7246 => x"3883f9bc",
          7247 => x"3384b880",
          7248 => x"3383f9bd",
          7249 => x"337281ff",
          7250 => x"067281ff",
          7251 => x"067281ff",
          7252 => x"06727229",
          7253 => x"05545b43",
          7254 => x"5b5b5b84",
          7255 => x"b8a83387",
          7256 => x"a3a0801b",
          7257 => x"3484b880",
          7258 => x"3383f9bd",
          7259 => x"3383f9ba",
          7260 => x"22727129",
          7261 => x"125e415e",
          7262 => x"56a00b83",
          7263 => x"f9be1c34",
          7264 => x"83f9bc33",
          7265 => x"7671291e",
          7266 => x"5a5e83f9",
          7267 => x"b83387a3",
          7268 => x"b0801a34",
          7269 => x"84b88033",
          7270 => x"7081ff06",
          7271 => x"83f9ba22",
          7272 => x"83f9bd33",
          7273 => x"72722911",
          7274 => x"5b445a40",
          7275 => x"5983f9b8",
          7276 => x"338498de",
          7277 => x"18346081",
          7278 => x"057081ff",
          7279 => x"065b5879",
          7280 => x"7f27fed6",
          7281 => x"387783f9",
          7282 => x"bd34fedf",
          7283 => x"39820b84",
          7284 => x"b9880c80",
          7285 => x"0b84ba8c",
          7286 => x"0c9c3d0d",
          7287 => x"0483f9be",
          7288 => x"17335984",
          7289 => x"b8881933",
          7290 => x"7a3483f9",
          7291 => x"bd337081",
          7292 => x"ff0658ff",
          7293 => x"0556f9ca",
          7294 => x"39810b84",
          7295 => x"b98e3480",
          7296 => x"0b84ba8c",
          7297 => x"0c9c3d0d",
          7298 => x"0483f9be",
          7299 => x"17335b84",
          7300 => x"b8881b33",
          7301 => x"7c3483f9",
          7302 => x"bc3384b8",
          7303 => x"803383f9",
          7304 => x"bd335b5b",
          7305 => x"5b805cfc",
          7306 => x"f43984b9",
          7307 => x"90429c3d",
          7308 => x"dc1153d8",
          7309 => x"0551ff8a",
          7310 => x"cd3f84ba",
          7311 => x"8c08802e",
          7312 => x"fbf03884",
          7313 => x"b98d3381",
          7314 => x"11575a75",
          7315 => x"84b98d34",
          7316 => x"791083fe",
          7317 => x"06410280",
          7318 => x"ca052261",
          7319 => x"84b9e005",
          7320 => x"23fbcf39",
          7321 => x"83f9be17",
          7322 => x"335c84b8",
          7323 => x"881c337b",
          7324 => x"3483f9bc",
          7325 => x"3384b880",
          7326 => x"3383f9bd",
          7327 => x"335b5b5c",
          7328 => x"f9e53984",
          7329 => x"b8803383",
          7330 => x"f9bc3383",
          7331 => x"f9bd3372",
          7332 => x"72290541",
          7333 => x"5d5b84b8",
          7334 => x"8819337f",
          7335 => x"87a3a080",
          7336 => x"053484b8",
          7337 => x"803383f9",
          7338 => x"bd3383f9",
          7339 => x"ba227271",
          7340 => x"29125a43",
          7341 => x"5b567883",
          7342 => x"f9be1834",
          7343 => x"83f9bc33",
          7344 => x"7671291b",
          7345 => x"415e83f9",
          7346 => x"b8336087",
          7347 => x"a3b08005",
          7348 => x"3484b880",
          7349 => x"337081ff",
          7350 => x"0683f9ba",
          7351 => x"2283f9bd",
          7352 => x"33727229",
          7353 => x"11415f5a",
          7354 => x"425a83f9",
          7355 => x"b8338498",
          7356 => x"de1e3481",
          7357 => x"1c7081ff",
          7358 => x"065c5860",
          7359 => x"7b2690a2",
          7360 => x"3884b881",
          7361 => x"33587790",
          7362 => x"e238ff1a",
          7363 => x"567583f9",
          7364 => x"bd34800b",
          7365 => x"84b9880c",
          7366 => x"84b88333",
          7367 => x"407f802e",
          7368 => x"f3bd3884",
          7369 => x"b8843356",
          7370 => x"75f3b438",
          7371 => x"78528151",
          7372 => x"eae43f80",
          7373 => x"0b84ba8c",
          7374 => x"0c9c3d0d",
          7375 => x"0484b9f4",
          7376 => x"3383f9bc",
          7377 => x"3484b9f5",
          7378 => x"3383f9bd",
          7379 => x"3484b9f6",
          7380 => x"33577683",
          7381 => x"f9ba23ff",
          7382 => x"b93983f9",
          7383 => x"bc3384b9",
          7384 => x"f43483f9",
          7385 => x"bd3384b9",
          7386 => x"f53483f9",
          7387 => x"bb3384b9",
          7388 => x"f634ff9e",
          7389 => x"3984b98d",
          7390 => x"335b7a80",
          7391 => x"2eff9338",
          7392 => x"84b9e022",
          7393 => x"5d7c862e",
          7394 => x"098106ff",
          7395 => x"853883f9",
          7396 => x"bd338105",
          7397 => x"5583f9bc",
          7398 => x"33810554",
          7399 => x"9b5383e4",
          7400 => x"8c52943d",
          7401 => x"705257fe",
          7402 => x"edfe3f76",
          7403 => x"51fefef8",
          7404 => x"3f84ba8c",
          7405 => x"0881ff06",
          7406 => x"83f89033",
          7407 => x"57760541",
          7408 => x"60a024fe",
          7409 => x"cd387652",
          7410 => x"83f7f051",
          7411 => x"fefdc33f",
          7412 => x"fec03980",
          7413 => x"0b84b98d",
          7414 => x"335b5879",
          7415 => x"81ff065b",
          7416 => x"777b27fe",
          7417 => x"ad387710",
          7418 => x"84b9e005",
          7419 => x"81113357",
          7420 => x"4175b126",
          7421 => x"8aa53875",
          7422 => x"101083c7",
          7423 => x"ec055f7e",
          7424 => x"080484b9",
          7425 => x"8d335e7d",
          7426 => x"802e8fa4",
          7427 => x"3883f9bc",
          7428 => x"3384b9e1",
          7429 => x"33717131",
          7430 => x"7009709f",
          7431 => x"2c72065a",
          7432 => x"42595e5c",
          7433 => x"7583f9bc",
          7434 => x"34fde739",
          7435 => x"84b98d33",
          7436 => x"5675802e",
          7437 => x"8ee73884",
          7438 => x"b9e133ff",
          7439 => x"057081ff",
          7440 => x"0684b880",
          7441 => x"335d575f",
          7442 => x"757b27fd",
          7443 => x"c5387583",
          7444 => x"f9bd34fd",
          7445 => x"bd39800b",
          7446 => x"83f9bd34",
          7447 => x"83f9bc33",
          7448 => x"7081ff06",
          7449 => x"5d577b80",
          7450 => x"2efda738",
          7451 => x"ff175675",
          7452 => x"83f9bc34",
          7453 => x"fd9c3980",
          7454 => x"0b83f9bd",
          7455 => x"3483f9bc",
          7456 => x"3384b7ff",
          7457 => x"33ff0557",
          7458 => x"57767625",
          7459 => x"fd843881",
          7460 => x"17567583",
          7461 => x"f9bc34fc",
          7462 => x"f93984b9",
          7463 => x"8d33407f",
          7464 => x"802e8de0",
          7465 => x"3883f9bd",
          7466 => x"3384b9e1",
          7467 => x"33717131",
          7468 => x"7009709f",
          7469 => x"2c72065a",
          7470 => x"4159425a",
          7471 => x"7583f9bd",
          7472 => x"34fccf39",
          7473 => x"84b98d33",
          7474 => x"5b7a802e",
          7475 => x"fcc43884",
          7476 => x"b9e02241",
          7477 => x"60992e09",
          7478 => x"8106fcb6",
          7479 => x"3884b880",
          7480 => x"3383f9bd",
          7481 => x"3383f9bc",
          7482 => x"33727129",
          7483 => x"1287a3a0",
          7484 => x"801183f9",
          7485 => x"ba224351",
          7486 => x"5a587160",
          7487 => x"29057083",
          7488 => x"ffff0683",
          7489 => x"f8900887",
          7490 => x"fffe8006",
          7491 => x"425a5d5d",
          7492 => x"7e848280",
          7493 => x"2e92bf38",
          7494 => x"800b83f8",
          7495 => x"9134fbf2",
          7496 => x"3984b98d",
          7497 => x"335a7980",
          7498 => x"2efbe738",
          7499 => x"84b9e022",
          7500 => x"5877992e",
          7501 => x"098106fb",
          7502 => x"d938810b",
          7503 => x"83f89134",
          7504 => x"fbd03984",
          7505 => x"b98d3356",
          7506 => x"75802e90",
          7507 => x"be3884b9",
          7508 => x"e13383f9",
          7509 => x"bd335d7c",
          7510 => x"0584b880",
          7511 => x"33ff1159",
          7512 => x"5e56757d",
          7513 => x"25833875",
          7514 => x"577683f9",
          7515 => x"bd34fba2",
          7516 => x"3984b98d",
          7517 => x"33577680",
          7518 => x"2e8cc838",
          7519 => x"84b9e133",
          7520 => x"83f9bc33",
          7521 => x"42610584",
          7522 => x"b7ff33ff",
          7523 => x"11594156",
          7524 => x"75602583",
          7525 => x"38755776",
          7526 => x"83f9bc34",
          7527 => x"faf43983",
          7528 => x"e49851fe",
          7529 => x"e8e23f80",
          7530 => x"0b84b98d",
          7531 => x"33575776",
          7532 => x"76278bc7",
          7533 => x"38761084",
          7534 => x"b9e00570",
          7535 => x"22535a83",
          7536 => x"e3f851fe",
          7537 => x"e8c23f81",
          7538 => x"177081ff",
          7539 => x"0684b98d",
          7540 => x"33585858",
          7541 => x"da39820b",
          7542 => x"84b98d33",
          7543 => x"5f577d80",
          7544 => x"2e8d3884",
          7545 => x"b9e02256",
          7546 => x"75832683",
          7547 => x"38755781",
          7548 => x"527681ff",
          7549 => x"0651d5f3",
          7550 => x"3ffa9739",
          7551 => x"84b98d33",
          7552 => x"57817727",
          7553 => x"8eb73884",
          7554 => x"b9e333ff",
          7555 => x"057081ff",
          7556 => x"0684b9e1",
          7557 => x"33ff0570",
          7558 => x"81ff0684",
          7559 => x"b7ff3370",
          7560 => x"81ff06ff",
          7561 => x"11404352",
          7562 => x"5b595c5c",
          7563 => x"777e2783",
          7564 => x"38775a79",
          7565 => x"83f9ba23",
          7566 => x"7681ff06",
          7567 => x"ff18585f",
          7568 => x"777f2783",
          7569 => x"38775776",
          7570 => x"83f9bc34",
          7571 => x"84b88033",
          7572 => x"ff115740",
          7573 => x"7a6027f9",
          7574 => x"b4387a56",
          7575 => x"7583f9bd",
          7576 => x"34f9af39",
          7577 => x"84b98d33",
          7578 => x"5f7e802e",
          7579 => x"8aef3884",
          7580 => x"b9e13384",
          7581 => x"b7ff3340",
          7582 => x"5b7a7f26",
          7583 => x"f9943883",
          7584 => x"f9bc3384",
          7585 => x"b8803370",
          7586 => x"81ff0683",
          7587 => x"f9bd3371",
          7588 => x"74291187",
          7589 => x"a3a08005",
          7590 => x"83f9ba22",
          7591 => x"5f40717e",
          7592 => x"29057083",
          7593 => x"ffff0683",
          7594 => x"f8923346",
          7595 => x"5259595f",
          7596 => x"5d60812e",
          7597 => x"84f03879",
          7598 => x"83ffff06",
          7599 => x"707c315d",
          7600 => x"57807c24",
          7601 => x"8efe3884",
          7602 => x"b7ff3356",
          7603 => x"7676278e",
          7604 => x"d638ff16",
          7605 => x"567583f9",
          7606 => x"ba237c81",
          7607 => x"ff06707c",
          7608 => x"31415780",
          7609 => x"60248ee5",
          7610 => x"3884b7ff",
          7611 => x"33567676",
          7612 => x"278dee38",
          7613 => x"ff165675",
          7614 => x"83f9bc34",
          7615 => x"7e81ff06",
          7616 => x"83f9ba22",
          7617 => x"5757805a",
          7618 => x"76762690",
          7619 => x"38757731",
          7620 => x"81057e81",
          7621 => x"ff067171",
          7622 => x"295c5e5b",
          7623 => x"795887a3",
          7624 => x"a0805b87",
          7625 => x"a3b0807f",
          7626 => x"81ff067f",
          7627 => x"81ff0671",
          7628 => x"71291d42",
          7629 => x"58425c79",
          7630 => x"7f27f7d6",
          7631 => x"388498de",
          7632 => x"1a57e0e0",
          7633 => x"17335f84",
          7634 => x"b8881f33",
          7635 => x"7b708105",
          7636 => x"5d347670",
          7637 => x"81055833",
          7638 => x"7c708105",
          7639 => x"5e348118",
          7640 => x"84b88033",
          7641 => x"84b7ff33",
          7642 => x"7171291d",
          7643 => x"43405e58",
          7644 => x"776027f7",
          7645 => x"9d38e0e0",
          7646 => x"17335f84",
          7647 => x"b8881f33",
          7648 => x"7b708105",
          7649 => x"5d347670",
          7650 => x"81055833",
          7651 => x"7c708105",
          7652 => x"5e348118",
          7653 => x"84b88033",
          7654 => x"84b7ff33",
          7655 => x"7171291d",
          7656 => x"43405e58",
          7657 => x"7f7826ff",
          7658 => x"9938f6e6",
          7659 => x"3984b98d",
          7660 => x"33567580",
          7661 => x"2e87e038",
          7662 => x"805284b9",
          7663 => x"e13351d8",
          7664 => x"b13ff6ce",
          7665 => x"39800b84",
          7666 => x"b88033ff",
          7667 => x"1184b98d",
          7668 => x"335d5940",
          7669 => x"5879782e",
          7670 => x"943884b9",
          7671 => x"e0225675",
          7672 => x"782e0981",
          7673 => x"068bbe38",
          7674 => x"83f9bd33",
          7675 => x"587681ff",
          7676 => x"0683f9bc",
          7677 => x"3379435c",
          7678 => x"5c76ff2e",
          7679 => x"81ed3884",
          7680 => x"b7ff3340",
          7681 => x"7a6026f6",
          7682 => x"89387e81",
          7683 => x"ff065660",
          7684 => x"7626f5fe",
          7685 => x"387b7626",
          7686 => x"617d2707",
          7687 => x"5776f5f2",
          7688 => x"387a1010",
          7689 => x"1b709029",
          7690 => x"620587a3",
          7691 => x"a0801170",
          7692 => x"1f5d5a87",
          7693 => x"a3b08005",
          7694 => x"79830658",
          7695 => x"515d758b",
          7696 => x"ac387983",
          7697 => x"0657768b",
          7698 => x"a43883f9",
          7699 => x"b8337098",
          7700 => x"2b71902b",
          7701 => x"0771882b",
          7702 => x"07710779",
          7703 => x"7f59525f",
          7704 => x"57777a27",
          7705 => x"9e388077",
          7706 => x"70840559",
          7707 => x"0c7d7670",
          7708 => x"8405580c",
          7709 => x"797726ee",
          7710 => x"3884b880",
          7711 => x"3384b7ff",
          7712 => x"33415f7e",
          7713 => x"81ff0660",
          7714 => x"81ff0683",
          7715 => x"f9ba227d",
          7716 => x"73296405",
          7717 => x"5959595a",
          7718 => x"7777268c",
          7719 => x"38767831",
          7720 => x"1b707b29",
          7721 => x"62055740",
          7722 => x"75761d57",
          7723 => x"57767626",
          7724 => x"f4e03883",
          7725 => x"f9b83384",
          7726 => x"98de1859",
          7727 => x"5aa00be0",
          7728 => x"e0193479",
          7729 => x"78708105",
          7730 => x"5a348117",
          7731 => x"57767626",
          7732 => x"f4c038a0",
          7733 => x"0be0e019",
          7734 => x"34797870",
          7735 => x"81055a34",
          7736 => x"81175775",
          7737 => x"7727d638",
          7738 => x"f4a839ff",
          7739 => x"1f7081ff",
          7740 => x"065d58fe",
          7741 => x"8a3983f9",
          7742 => x"b8337080",
          7743 => x"f0067184",
          7744 => x"2b80f006",
          7745 => x"71842a07",
          7746 => x"585d577b",
          7747 => x"80f02e09",
          7748 => x"8106be38",
          7749 => x"80f20b83",
          7750 => x"f9b83481",
          7751 => x"187081ff",
          7752 => x"065956f5",
          7753 => x"b63983f9",
          7754 => x"be17335e",
          7755 => x"84b8881e",
          7756 => x"337c3483",
          7757 => x"f9bc3384",
          7758 => x"b8803383",
          7759 => x"f9ba2284",
          7760 => x"b7ff3342",
          7761 => x"5c5f5dfa",
          7762 => x"ee3983f9",
          7763 => x"b8338707",
          7764 => x"567583f9",
          7765 => x"b8348118",
          7766 => x"7081ff06",
          7767 => x"5956f4fb",
          7768 => x"3983f9b8",
          7769 => x"3381fd06",
          7770 => x"85075675",
          7771 => x"83f9b834",
          7772 => x"e53983f9",
          7773 => x"b83381fb",
          7774 => x"06830756",
          7775 => x"7583f9b8",
          7776 => x"34d43983",
          7777 => x"f9b83381",
          7778 => x"f9068107",
          7779 => x"567583f9",
          7780 => x"b834c339",
          7781 => x"83f9b833",
          7782 => x"819f0690",
          7783 => x"07567583",
          7784 => x"f9b834ff",
          7785 => x"b13980f1",
          7786 => x"0b83f9b8",
          7787 => x"34811870",
          7788 => x"81ff0659",
          7789 => x"56f4a439",
          7790 => x"83f9b833",
          7791 => x"818f0656",
          7792 => x"7583f9b8",
          7793 => x"34ff8f39",
          7794 => x"83f9b833",
          7795 => x"819f0690",
          7796 => x"07567583",
          7797 => x"f9b834fe",
          7798 => x"fd3983f9",
          7799 => x"b83381ef",
          7800 => x"0680e007",
          7801 => x"567583f9",
          7802 => x"b834feea",
          7803 => x"3983f9b8",
          7804 => x"3381cf06",
          7805 => x"80c00756",
          7806 => x"7583f9b8",
          7807 => x"34fed739",
          7808 => x"83f9b833",
          7809 => x"81af06a0",
          7810 => x"07567583",
          7811 => x"f9b834fe",
          7812 => x"c53983f9",
          7813 => x"b83381fe",
          7814 => x"06860756",
          7815 => x"7583f9b8",
          7816 => x"34feb339",
          7817 => x"83f9b833",
          7818 => x"81fc0684",
          7819 => x"07567583",
          7820 => x"f9b834fe",
          7821 => x"a13983f9",
          7822 => x"b83381fa",
          7823 => x"06820756",
          7824 => x"7583f9b8",
          7825 => x"34fe8f39",
          7826 => x"83f9b833",
          7827 => x"81f80656",
          7828 => x"7583f9b8",
          7829 => x"34fdff39",
          7830 => x"83f9b833",
          7831 => x"80f00756",
          7832 => x"7583f9b8",
          7833 => x"34fdef39",
          7834 => x"83f9b833",
          7835 => x"80f00756",
          7836 => x"7583f9b8",
          7837 => x"34fddf39",
          7838 => x"83f9b833",
          7839 => x"81df0680",
          7840 => x"d0075675",
          7841 => x"83f9b834",
          7842 => x"fdcc3983",
          7843 => x"f9b83381",
          7844 => x"bf06b007",
          7845 => x"567583f9",
          7846 => x"b834fdba",
          7847 => x"39800b83",
          7848 => x"f9bd3480",
          7849 => x"528151d2",
          7850 => x"c93fecff",
          7851 => x"3984b9f4",
          7852 => x"3383f9bc",
          7853 => x"3484b9f5",
          7854 => x"3383f9bd",
          7855 => x"3484b9f6",
          7856 => x"33597883",
          7857 => x"f9ba2380",
          7858 => x"0b84b988",
          7859 => x"0ce8c739",
          7860 => x"810b84b9",
          7861 => x"8f34800b",
          7862 => x"84ba8c0c",
          7863 => x"9c3d0d04",
          7864 => x"7783f9bd",
          7865 => x"3483f9bd",
          7866 => x"337081ff",
          7867 => x"0658ff05",
          7868 => x"56e7cf39",
          7869 => x"84b99042",
          7870 => x"9c3ddc11",
          7871 => x"53d80551",
          7872 => x"fef9833f",
          7873 => x"84ba8c08",
          7874 => x"a13884ba",
          7875 => x"8c0884b9",
          7876 => x"880c800b",
          7877 => x"84b98c34",
          7878 => x"800b84ba",
          7879 => x"8c0c9c3d",
          7880 => x"0d047783",
          7881 => x"f9bd34ef",
          7882 => x"e93984b9",
          7883 => x"8d338111",
          7884 => x"5c5c7a84",
          7885 => x"b98d347b",
          7886 => x"1083fe06",
          7887 => x"5d0280ca",
          7888 => x"052284b9",
          7889 => x"e01e2380",
          7890 => x"0b84b98c",
          7891 => x"34ca3980",
          7892 => x"0b83f9bd",
          7893 => x"34805281",
          7894 => x"51d1973f",
          7895 => x"83f9bd33",
          7896 => x"7081ff06",
          7897 => x"58ff0556",
          7898 => x"e6d83980",
          7899 => x"0b83f9bd",
          7900 => x"34805281",
          7901 => x"51d0fb3f",
          7902 => x"ef98398a",
          7903 => x"51feebde",
          7904 => x"3fef8f39",
          7905 => x"83f9bd33",
          7906 => x"ff057009",
          7907 => x"709f2c72",
          7908 => x"06585f57",
          7909 => x"f2a63975",
          7910 => x"528151d9",
          7911 => x"3984b880",
          7912 => x"33407560",
          7913 => x"27eeeb38",
          7914 => x"7583f9bd",
          7915 => x"34eee339",
          7916 => x"83f9bc33",
          7917 => x"ff057009",
          7918 => x"709f2c72",
          7919 => x"06584057",
          7920 => x"f0e23983",
          7921 => x"f9bc3381",
          7922 => x"0584b7ff",
          7923 => x"33ff1159",
          7924 => x"59567578",
          7925 => x"25f3c038",
          7926 => x"7557f3bb",
          7927 => x"3984b7ff",
          7928 => x"337081ff",
          7929 => x"06585c81",
          7930 => x"7726eea6",
          7931 => x"3883f9bc",
          7932 => x"3384b880",
          7933 => x"337081ff",
          7934 => x"0683f9bd",
          7935 => x"33717429",
          7936 => x"1187a3a0",
          7937 => x"800583f9",
          7938 => x"ba225f5f",
          7939 => x"717e2905",
          7940 => x"7083ffff",
          7941 => x"0683f892",
          7942 => x"335d5b44",
          7943 => x"425f5d77",
          7944 => x"812e81f5",
          7945 => x"387983ff",
          7946 => x"ff06ff11",
          7947 => x"5c57807b",
          7948 => x"24848938",
          7949 => x"84b7ff33",
          7950 => x"56767627",
          7951 => x"839838ff",
          7952 => x"16567583",
          7953 => x"f9ba237c",
          7954 => x"81ff06ff",
          7955 => x"11575780",
          7956 => x"762483df",
          7957 => x"3884b7ff",
          7958 => x"33567676",
          7959 => x"2782ec38",
          7960 => x"ff165675",
          7961 => x"83f9bc34",
          7962 => x"7b81ff06",
          7963 => x"83f9ba22",
          7964 => x"5757805a",
          7965 => x"76762690",
          7966 => x"38757731",
          7967 => x"81057e81",
          7968 => x"ff067171",
          7969 => x"295c5e5f",
          7970 => x"795887a3",
          7971 => x"a0805b87",
          7972 => x"a3b0807c",
          7973 => x"81ff067f",
          7974 => x"81ff0671",
          7975 => x"71291d41",
          7976 => x"42425d79",
          7977 => x"7e27ecea",
          7978 => x"388498de",
          7979 => x"1a57e0e0",
          7980 => x"17335e84",
          7981 => x"b8881e33",
          7982 => x"7b708105",
          7983 => x"5d347670",
          7984 => x"81055833",
          7985 => x"7d708105",
          7986 => x"5f348118",
          7987 => x"84b88033",
          7988 => x"84b7ff33",
          7989 => x"7171291d",
          7990 => x"59415d58",
          7991 => x"777627ec",
          7992 => x"b138e0e0",
          7993 => x"17335e84",
          7994 => x"b8881e33",
          7995 => x"7b708105",
          7996 => x"5d347670",
          7997 => x"81055833",
          7998 => x"7d708105",
          7999 => x"5f348118",
          8000 => x"84b88033",
          8001 => x"84b7ff33",
          8002 => x"7171291d",
          8003 => x"59415d58",
          8004 => x"757826ff",
          8005 => x"9938ebfa",
          8006 => x"3983f9be",
          8007 => x"17335c84",
          8008 => x"b8881c33",
          8009 => x"7b3483f9",
          8010 => x"bc3384b8",
          8011 => x"803383f9",
          8012 => x"ba2284b7",
          8013 => x"ff335f5c",
          8014 => x"5f5dfde9",
          8015 => x"3976ebd2",
          8016 => x"3884b7ff",
          8017 => x"337081ff",
          8018 => x"06ff115c",
          8019 => x"42587661",
          8020 => x"27833876",
          8021 => x"5a7983f9",
          8022 => x"ba237781",
          8023 => x"ff06ff19",
          8024 => x"585a807a",
          8025 => x"27833880",
          8026 => x"577683f9",
          8027 => x"bc3484b8",
          8028 => x"80337081",
          8029 => x"ff06ff12",
          8030 => x"52595680",
          8031 => x"7827eb8d",
          8032 => x"38805675",
          8033 => x"83f9bd34",
          8034 => x"eb883983",
          8035 => x"f9bd3381",
          8036 => x"0584b880",
          8037 => x"33ff1159",
          8038 => x"4056757f",
          8039 => x"25efca38",
          8040 => x"7557efc5",
          8041 => x"3975812e",
          8042 => x"098106f4",
          8043 => x"c03883f9",
          8044 => x"bd337081",
          8045 => x"ff0683f9",
          8046 => x"bc337a44",
          8047 => x"5d5d5776",
          8048 => x"ff2e0981",
          8049 => x"06f4b838",
          8050 => x"f6a139ff",
          8051 => x"1d567583",
          8052 => x"f9bc34fd",
          8053 => x"9339ff1a",
          8054 => x"567583f9",
          8055 => x"ba23fce7",
          8056 => x"397c7b31",
          8057 => x"567583f9",
          8058 => x"bc34f290",
          8059 => x"39777d58",
          8060 => x"56777a26",
          8061 => x"f58d3880",
          8062 => x"76708105",
          8063 => x"583483f9",
          8064 => x"b8337770",
          8065 => x"81055934",
          8066 => x"757a26f4",
          8067 => x"ec388076",
          8068 => x"70810558",
          8069 => x"3483f9b8",
          8070 => x"33777081",
          8071 => x"05593479",
          8072 => x"7627d438",
          8073 => x"f4d33979",
          8074 => x"7b315675",
          8075 => x"83f9ba23",
          8076 => x"f1a83980",
          8077 => x"0b83f9bc",
          8078 => x"34fcad39",
          8079 => x"7e83f9ba",
          8080 => x"23fc8439",
          8081 => x"800b83f9",
          8082 => x"ba23f18e",
          8083 => x"39800b83",
          8084 => x"f9bc34f1",
          8085 => x"a73983f9",
          8086 => x"be18335a",
          8087 => x"84b8881a",
          8088 => x"33773480",
          8089 => x"0b83f891",
          8090 => x"34e9a739",
          8091 => x"fd3d0d02",
          8092 => x"97053384",
          8093 => x"b8823354",
          8094 => x"5472802e",
          8095 => x"90387351",
          8096 => x"db9c3f80",
          8097 => x"0b84ba8c",
          8098 => x"0c853d0d",
          8099 => x"04765273",
          8100 => x"51d7ab3f",
          8101 => x"800b84ba",
          8102 => x"8c0c853d",
          8103 => x"0d04f33d",
          8104 => x"0d02bf05",
          8105 => x"335cff0b",
          8106 => x"83f89033",
          8107 => x"7081ff06",
          8108 => x"83f7f011",
          8109 => x"33585555",
          8110 => x"5974802e",
          8111 => x"80d63881",
          8112 => x"14567583",
          8113 => x"f8903474",
          8114 => x"597884ba",
          8115 => x"8c0c8f3d",
          8116 => x"0d0483f7",
          8117 => x"ec085482",
          8118 => x"5373802e",
          8119 => x"91387373",
          8120 => x"32703071",
          8121 => x"07700970",
          8122 => x"9f2a565d",
          8123 => x"5e587283",
          8124 => x"f7ec0cff",
          8125 => x"5980547b",
          8126 => x"812e0981",
          8127 => x"0683387b",
          8128 => x"547b8332",
          8129 => x"70307080",
          8130 => x"2576075c",
          8131 => x"5c5d7980",
          8132 => x"2e85c438",
          8133 => x"84b88033",
          8134 => x"83f9bd33",
          8135 => x"83f9bc33",
          8136 => x"72712912",
          8137 => x"87a3a080",
          8138 => x"0583f9ba",
          8139 => x"225b595d",
          8140 => x"71792905",
          8141 => x"7083ffff",
          8142 => x"0683f891",
          8143 => x"33585955",
          8144 => x"5874812e",
          8145 => x"838c3881",
          8146 => x"f0547386",
          8147 => x"ee808034",
          8148 => x"800b87c0",
          8149 => x"98880c87",
          8150 => x"c0988808",
          8151 => x"5675802e",
          8152 => x"f63886ee",
          8153 => x"80840857",
          8154 => x"7683f5bc",
          8155 => x"15348114",
          8156 => x"7081ff06",
          8157 => x"555581f9",
          8158 => x"7427cf38",
          8159 => x"805483f7",
          8160 => x"ac143370",
          8161 => x"81ff0683",
          8162 => x"f7b61633",
          8163 => x"58545572",
          8164 => x"762e85c1",
          8165 => x"387281ff",
          8166 => x"2e86b438",
          8167 => x"7483f7c0",
          8168 => x"15347581",
          8169 => x"ff065a79",
          8170 => x"81ff2e85",
          8171 => x"cd387583",
          8172 => x"f7ca1534",
          8173 => x"83f7ac14",
          8174 => x"3383f7b6",
          8175 => x"15348114",
          8176 => x"7081ff06",
          8177 => x"555e8974",
          8178 => x"27ffb338",
          8179 => x"83f7b433",
          8180 => x"70982b70",
          8181 => x"80255856",
          8182 => x"547583f7",
          8183 => x"e4347381",
          8184 => x"ff067086",
          8185 => x"2a813270",
          8186 => x"81065154",
          8187 => x"5872802e",
          8188 => x"85e73881",
          8189 => x"0b83f7e5",
          8190 => x"34730981",
          8191 => x"06537280",
          8192 => x"2e85e438",
          8193 => x"810b83f7",
          8194 => x"e634800b",
          8195 => x"83f7e533",
          8196 => x"83f7ec08",
          8197 => x"83f7e633",
          8198 => x"7083f7e8",
          8199 => x"3383f7e7",
          8200 => x"335d5d42",
          8201 => x"5e5c5e56",
          8202 => x"83f7c016",
          8203 => x"33557481",
          8204 => x"ff2e8d38",
          8205 => x"83f7d416",
          8206 => x"33547380",
          8207 => x"2e828238",
          8208 => x"83f7ca16",
          8209 => x"33537281",
          8210 => x"ff2e8b38",
          8211 => x"83f7d416",
          8212 => x"33547381",
          8213 => x"ec387481",
          8214 => x"ff065473",
          8215 => x"81ff2e8d",
          8216 => x"3883f7d4",
          8217 => x"16335372",
          8218 => x"812e81da",
          8219 => x"387481ff",
          8220 => x"06537281",
          8221 => x"ff2e848c",
          8222 => x"3883f7d4",
          8223 => x"16335481",
          8224 => x"74278480",
          8225 => x"3883f7e0",
          8226 => x"0887e805",
          8227 => x"87c0989c",
          8228 => x"08545473",
          8229 => x"732783ec",
          8230 => x"38810b87",
          8231 => x"c0989c08",
          8232 => x"83f7e00c",
          8233 => x"58811670",
          8234 => x"81ff0657",
          8235 => x"54897627",
          8236 => x"fef63876",
          8237 => x"83f7e734",
          8238 => x"7783f7e8",
          8239 => x"34fe9e19",
          8240 => x"53729c26",
          8241 => x"828b3872",
          8242 => x"101083c9",
          8243 => x"b4055a79",
          8244 => x"080483f8",
          8245 => x"94085473",
          8246 => x"802e9138",
          8247 => x"83f41487",
          8248 => x"c0989c08",
          8249 => x"5e5e7d7d",
          8250 => x"27fcdc38",
          8251 => x"800b83f8",
          8252 => x"92335454",
          8253 => x"72812e83",
          8254 => x"38745473",
          8255 => x"83f89234",
          8256 => x"87c0989c",
          8257 => x"0883f894",
          8258 => x"0c7381ff",
          8259 => x"06587781",
          8260 => x"2e943883",
          8261 => x"f9be1733",
          8262 => x"5484b888",
          8263 => x"14337634",
          8264 => x"81f054fc",
          8265 => x"a53983f7",
          8266 => x"ec085372",
          8267 => x"802e829c",
          8268 => x"3872812e",
          8269 => x"83f43880",
          8270 => x"c3763481",
          8271 => x"f054fc8a",
          8272 => x"398058fe",
          8273 => x"e0398074",
          8274 => x"56578359",
          8275 => x"7c812e9b",
          8276 => x"3879772e",
          8277 => x"09810683",
          8278 => x"b4387d81",
          8279 => x"2e80ed38",
          8280 => x"79812e80",
          8281 => x"d7387981",
          8282 => x"ff065987",
          8283 => x"77277598",
          8284 => x"2b545472",
          8285 => x"8025a138",
          8286 => x"73802e9c",
          8287 => x"38811770",
          8288 => x"81ff0676",
          8289 => x"1081fe06",
          8290 => x"87722771",
          8291 => x"982b5753",
          8292 => x"57585480",
          8293 => x"7324e138",
          8294 => x"78101010",
          8295 => x"79100576",
          8296 => x"11832b78",
          8297 => x"0583f49c",
          8298 => x"0570335b",
          8299 => x"56547887",
          8300 => x"c0989c08",
          8301 => x"83f7e00c",
          8302 => x"57fdea39",
          8303 => x"80597d81",
          8304 => x"2effa838",
          8305 => x"7981ff06",
          8306 => x"59ffa039",
          8307 => x"8259ff9b",
          8308 => x"3978ff2e",
          8309 => x"fa9f3880",
          8310 => x"0b84b882",
          8311 => x"33545472",
          8312 => x"812e83e8",
          8313 => x"387b8232",
          8314 => x"70307080",
          8315 => x"25760740",
          8316 => x"59567d8a",
          8317 => x"387b832e",
          8318 => x"098106f9",
          8319 => x"cc3878ff",
          8320 => x"2ef9c638",
          8321 => x"80537210",
          8322 => x"101083f8",
          8323 => x"98057033",
          8324 => x"5d54787c",
          8325 => x"2e83ba38",
          8326 => x"81137081",
          8327 => x"ff065457",
          8328 => x"937327e2",
          8329 => x"3884b883",
          8330 => x"33537280",
          8331 => x"2ef99a38",
          8332 => x"84b88433",
          8333 => x"5574f991",
          8334 => x"387881ff",
          8335 => x"06528251",
          8336 => x"ccd43f78",
          8337 => x"84ba8c0c",
          8338 => x"8f3d0d04",
          8339 => x"be763481",
          8340 => x"f054f9f6",
          8341 => x"397281ff",
          8342 => x"2e923883",
          8343 => x"f7d41433",
          8344 => x"81055b7a",
          8345 => x"83f7d415",
          8346 => x"34fac939",
          8347 => x"800b83f7",
          8348 => x"d41534ff",
          8349 => x"0b83f7c0",
          8350 => x"1534ff0b",
          8351 => x"83f7ca15",
          8352 => x"34fab139",
          8353 => x"7481ff06",
          8354 => x"537281ff",
          8355 => x"2efc9638",
          8356 => x"83f7d416",
          8357 => x"33558175",
          8358 => x"27fc8a38",
          8359 => x"7781ff06",
          8360 => x"5473812e",
          8361 => x"098106fb",
          8362 => x"fc3883f7",
          8363 => x"e00881fa",
          8364 => x"0587c098",
          8365 => x"9c085455",
          8366 => x"747327fb",
          8367 => x"e83887c0",
          8368 => x"989c0883",
          8369 => x"f7e00c76",
          8370 => x"81ff0659",
          8371 => x"fbd739ff",
          8372 => x"0b83f7c0",
          8373 => x"1534f9ca",
          8374 => x"397283f7",
          8375 => x"e5347309",
          8376 => x"81065372",
          8377 => x"fa9e3872",
          8378 => x"83f7e634",
          8379 => x"800b83f7",
          8380 => x"e53383f7",
          8381 => x"ec0883f7",
          8382 => x"e6337083",
          8383 => x"f7e83383",
          8384 => x"f7e7335d",
          8385 => x"5d425e5c",
          8386 => x"5e56fa9c",
          8387 => x"3979822e",
          8388 => x"098106fc",
          8389 => x"cb387a59",
          8390 => x"7a812efc",
          8391 => x"ce387981",
          8392 => x"2e098106",
          8393 => x"fcc038fd",
          8394 => x"9339ef76",
          8395 => x"3481f054",
          8396 => x"f8983980",
          8397 => x"0b84b883",
          8398 => x"33575475",
          8399 => x"83388154",
          8400 => x"7384b883",
          8401 => x"34ff59f7",
          8402 => x"ac39800b",
          8403 => x"84b88233",
          8404 => x"58547683",
          8405 => x"38815473",
          8406 => x"84b88234",
          8407 => x"ff59f795",
          8408 => x"39815383",
          8409 => x"f7ec0884",
          8410 => x"2ef78338",
          8411 => x"840b83f7",
          8412 => x"ec0cf6ff",
          8413 => x"3984b7ff",
          8414 => x"337081ff",
          8415 => x"06ff1157",
          8416 => x"5a548079",
          8417 => x"27833880",
          8418 => x"557483f9",
          8419 => x"ba237381",
          8420 => x"ff06ff15",
          8421 => x"55538073",
          8422 => x"27833880",
          8423 => x"547383f9",
          8424 => x"bc3484b8",
          8425 => x"80337081",
          8426 => x"ff0656ff",
          8427 => x"05538075",
          8428 => x"27833880",
          8429 => x"537283f9",
          8430 => x"bd34ff59",
          8431 => x"f6b73981",
          8432 => x"528351ff",
          8433 => x"baa53fff",
          8434 => x"59f6aa39",
          8435 => x"7254fc95",
          8436 => x"39841408",
          8437 => x"5283f7f0",
          8438 => x"51fedeeb",
          8439 => x"3f810b83",
          8440 => x"f8903483",
          8441 => x"f7f03359",
          8442 => x"fcbb3980",
          8443 => x"3d0d8151",
          8444 => x"f5ac3f82",
          8445 => x"3d0d04f9",
          8446 => x"3d0d800b",
          8447 => x"83f49808",
          8448 => x"545802a7",
          8449 => x"05338214",
          8450 => x"3483f498",
          8451 => x"085280e0",
          8452 => x"7234850b",
          8453 => x"83f49808",
          8454 => x"5657fe0b",
          8455 => x"81163480",
          8456 => x"0b86f080",
          8457 => x"e83487c0",
          8458 => x"989c0883",
          8459 => x"f4980856",
          8460 => x"80ce9005",
          8461 => x"5487c098",
          8462 => x"9c085387",
          8463 => x"c0989c08",
          8464 => x"5271732e",
          8465 => x"f6388115",
          8466 => x"3387c098",
          8467 => x"9c085753",
          8468 => x"75742787",
          8469 => x"387281fe",
          8470 => x"2edb3887",
          8471 => x"c098a408",
          8472 => x"52ff5671",
          8473 => x"742780cd",
          8474 => x"38725672",
          8475 => x"ff2e80c5",
          8476 => x"3887c098",
          8477 => x"9c0880ce",
          8478 => x"90055487",
          8479 => x"c0989c08",
          8480 => x"5387c098",
          8481 => x"9c085675",
          8482 => x"732ef638",
          8483 => x"81153387",
          8484 => x"c0989c08",
          8485 => x"53537174",
          8486 => x"27873872",
          8487 => x"81ff2edb",
          8488 => x"3887c098",
          8489 => x"a40852ff",
          8490 => x"56717427",
          8491 => x"a4387256",
          8492 => x"72ff2e9d",
          8493 => x"3876802e",
          8494 => x"a3387581",
          8495 => x"ff065372",
          8496 => x"fed83875",
          8497 => x"ff2e9538",
          8498 => x"7784ba8c",
          8499 => x"0c893d0d",
          8500 => x"04ff1770",
          8501 => x"81ff0658",
          8502 => x"5476df38",
          8503 => x"810b83e4",
          8504 => x"d45258fe",
          8505 => x"d78d3f77",
          8506 => x"84ba8c0c",
          8507 => x"893d0d04",
          8508 => x"f93d0d7a",
          8509 => x"028405a7",
          8510 => x"05335753",
          8511 => x"800b83f4",
          8512 => x"98087488",
          8513 => x"2b87fc80",
          8514 => x"80067076",
          8515 => x"982a0751",
          8516 => x"56565872",
          8517 => x"83163473",
          8518 => x"902a5271",
          8519 => x"84163472",
          8520 => x"902a5776",
          8521 => x"85163473",
          8522 => x"86163483",
          8523 => x"f4980853",
          8524 => x"75821434",
          8525 => x"83f49808",
          8526 => x"5280e172",
          8527 => x"34850b83",
          8528 => x"f4980856",
          8529 => x"57fe0b81",
          8530 => x"1634800b",
          8531 => x"86f080e8",
          8532 => x"3487c098",
          8533 => x"9c0883f4",
          8534 => x"98085680",
          8535 => x"ce900554",
          8536 => x"87c0989c",
          8537 => x"085387c0",
          8538 => x"989c0852",
          8539 => x"71732ef6",
          8540 => x"38811533",
          8541 => x"87c0989c",
          8542 => x"08575375",
          8543 => x"74278738",
          8544 => x"7281fe2e",
          8545 => x"db3887c0",
          8546 => x"98a40852",
          8547 => x"ff567174",
          8548 => x"2780cf38",
          8549 => x"725672ff",
          8550 => x"2e80c738",
          8551 => x"87c0989c",
          8552 => x"0880ce90",
          8553 => x"055487c0",
          8554 => x"989c0853",
          8555 => x"87c0989c",
          8556 => x"08567573",
          8557 => x"2ef63881",
          8558 => x"153387c0",
          8559 => x"989c0853",
          8560 => x"53717427",
          8561 => x"87387281",
          8562 => x"ff2edb38",
          8563 => x"87c098a4",
          8564 => x"0852ff56",
          8565 => x"71742780",
          8566 => x"df387256",
          8567 => x"72ff2e80",
          8568 => x"d7387680",
          8569 => x"2e80dd38",
          8570 => x"7581ff06",
          8571 => x"5372fed5",
          8572 => x"38755271",
          8573 => x"81ff0657",
          8574 => x"76aa3880",
          8575 => x"c6157c84",
          8576 => x"80115653",
          8577 => x"53717427",
          8578 => x"92387270",
          8579 => x"81055433",
          8580 => x"72708105",
          8581 => x"54347372",
          8582 => x"26f03877",
          8583 => x"84ba8c0c",
          8584 => x"893d0d04",
          8585 => x"810b83e4",
          8586 => x"e85258fe",
          8587 => x"d4c53f77",
          8588 => x"84ba8c0c",
          8589 => x"893d0d04",
          8590 => x"ff177081",
          8591 => x"ff065854",
          8592 => x"76ffa538",
          8593 => x"ff52ffab",
          8594 => x"39f93d0d",
          8595 => x"7a028405",
          8596 => x"a7053357",
          8597 => x"57800b83",
          8598 => x"f4980878",
          8599 => x"882b87fc",
          8600 => x"80800670",
          8601 => x"7a982a07",
          8602 => x"51565658",
          8603 => x"76831634",
          8604 => x"73902a52",
          8605 => x"71841634",
          8606 => x"76902a53",
          8607 => x"72851634",
          8608 => x"73861634",
          8609 => x"7b83f498",
          8610 => x"0880c611",
          8611 => x"84801357",
          8612 => x"55565271",
          8613 => x"74279738",
          8614 => x"71708105",
          8615 => x"53337370",
          8616 => x"81055534",
          8617 => x"737226f0",
          8618 => x"3883f498",
          8619 => x"08557582",
          8620 => x"163483f4",
          8621 => x"98085680",
          8622 => x"e2763485",
          8623 => x"0b83f498",
          8624 => x"085657fe",
          8625 => x"0b811634",
          8626 => x"800b86f0",
          8627 => x"80e83487",
          8628 => x"c0989c08",
          8629 => x"83f49808",
          8630 => x"5680ce90",
          8631 => x"055487c0",
          8632 => x"989c0853",
          8633 => x"87c0989c",
          8634 => x"08527173",
          8635 => x"2ef63881",
          8636 => x"153387c0",
          8637 => x"989c0857",
          8638 => x"53757427",
          8639 => x"87387281",
          8640 => x"fe2edb38",
          8641 => x"87c098a4",
          8642 => x"0852ff56",
          8643 => x"71742780",
          8644 => x"cd387256",
          8645 => x"72ff2e80",
          8646 => x"c53887c0",
          8647 => x"989c0880",
          8648 => x"ce900554",
          8649 => x"87c0989c",
          8650 => x"085387c0",
          8651 => x"989c0856",
          8652 => x"75732ef6",
          8653 => x"38811533",
          8654 => x"87c0989c",
          8655 => x"08535371",
          8656 => x"74278738",
          8657 => x"7281ff2e",
          8658 => x"db3887c0",
          8659 => x"98a40852",
          8660 => x"ff567174",
          8661 => x"27a93872",
          8662 => x"5672ff2e",
          8663 => x"a2387680",
          8664 => x"2ea83875",
          8665 => x"81ff0653",
          8666 => x"72fed838",
          8667 => x"757081ff",
          8668 => x"06565274",
          8669 => x"a1387784",
          8670 => x"ba8c0c89",
          8671 => x"3d0d04ff",
          8672 => x"177081ff",
          8673 => x"06585476",
          8674 => x"da38ff70",
          8675 => x"81ff0656",
          8676 => x"5274802e",
          8677 => x"e138810b",
          8678 => x"83e4fc52",
          8679 => x"58fed1d3",
          8680 => x"3f7784ba",
          8681 => x"8c0c893d",
          8682 => x"0d04fb3d",
          8683 => x"0d83f498",
          8684 => x"085180d0",
          8685 => x"7134850b",
          8686 => x"83f49808",
          8687 => x"5656fe0b",
          8688 => x"81163480",
          8689 => x"0b86f080",
          8690 => x"e83487c0",
          8691 => x"989c0883",
          8692 => x"f4980856",
          8693 => x"80ce9005",
          8694 => x"5487c098",
          8695 => x"9c085287",
          8696 => x"c0989c08",
          8697 => x"5372722e",
          8698 => x"f6388115",
          8699 => x"3387c098",
          8700 => x"9c085252",
          8701 => x"70742787",
          8702 => x"387181fe",
          8703 => x"2edb3887",
          8704 => x"c098a408",
          8705 => x"51ff5370",
          8706 => x"742780cd",
          8707 => x"38715371",
          8708 => x"ff2e80c5",
          8709 => x"3887c098",
          8710 => x"9c0880ce",
          8711 => x"90055487",
          8712 => x"c0989c08",
          8713 => x"5287c098",
          8714 => x"9c085372",
          8715 => x"722ef638",
          8716 => x"81153387",
          8717 => x"c0989c08",
          8718 => x"52527074",
          8719 => x"27873871",
          8720 => x"81ff2edb",
          8721 => x"3887c098",
          8722 => x"a40851ff",
          8723 => x"53707427",
          8724 => x"98387153",
          8725 => x"71ff2e91",
          8726 => x"3875802e",
          8727 => x"8a387281",
          8728 => x"ff065271",
          8729 => x"fed838ff",
          8730 => x"39ff1670",
          8731 => x"81ff0657",
          8732 => x"54e73980",
          8733 => x"3d0d83e5",
          8734 => x"9051fecf",
          8735 => x"f63f823d",
          8736 => x"0d04f93d",
          8737 => x"0d84b9fc",
          8738 => x"087a7131",
          8739 => x"832a7083",
          8740 => x"ffff0670",
          8741 => x"832b7311",
          8742 => x"70338112",
          8743 => x"33718b2b",
          8744 => x"71832b07",
          8745 => x"77117033",
          8746 => x"81123371",
          8747 => x"982b7190",
          8748 => x"2b075c54",
          8749 => x"4153535d",
          8750 => x"57595256",
          8751 => x"57538071",
          8752 => x"2481af38",
          8753 => x"72168211",
          8754 => x"33831233",
          8755 => x"718b2b71",
          8756 => x"832b0776",
          8757 => x"05703381",
          8758 => x"12337198",
          8759 => x"2b71902b",
          8760 => x"0757535c",
          8761 => x"52595652",
          8762 => x"80712483",
          8763 => x"9e388413",
          8764 => x"33851433",
          8765 => x"718b2b71",
          8766 => x"832b0775",
          8767 => x"0576882a",
          8768 => x"52545657",
          8769 => x"74861334",
          8770 => x"7381ff06",
          8771 => x"54738713",
          8772 => x"3484b9fc",
          8773 => x"08701784",
          8774 => x"12338513",
          8775 => x"3371882b",
          8776 => x"0770882a",
          8777 => x"5c555954",
          8778 => x"51778414",
          8779 => x"34718514",
          8780 => x"3484b9fc",
          8781 => x"08165280",
          8782 => x"0b861334",
          8783 => x"800b8713",
          8784 => x"3484b9fc",
          8785 => x"08537484",
          8786 => x"14347385",
          8787 => x"143484b9",
          8788 => x"fc081670",
          8789 => x"33811233",
          8790 => x"71882b07",
          8791 => x"82808007",
          8792 => x"70882a58",
          8793 => x"58525274",
          8794 => x"72347581",
          8795 => x"1334893d",
          8796 => x"0d048612",
          8797 => x"33871333",
          8798 => x"718b2b71",
          8799 => x"832b0775",
          8800 => x"11841633",
          8801 => x"85173371",
          8802 => x"882b0770",
          8803 => x"882a5858",
          8804 => x"54515358",
          8805 => x"58718412",
          8806 => x"34728512",
          8807 => x"3484b9fc",
          8808 => x"08701684",
          8809 => x"11338512",
          8810 => x"33718b2b",
          8811 => x"71832b07",
          8812 => x"565a5a52",
          8813 => x"72058612",
          8814 => x"33871333",
          8815 => x"71882b07",
          8816 => x"70882a52",
          8817 => x"55595277",
          8818 => x"86133472",
          8819 => x"87133484",
          8820 => x"b9fc0815",
          8821 => x"70338112",
          8822 => x"3371882b",
          8823 => x"0781ffff",
          8824 => x"0670882a",
          8825 => x"5a5a5452",
          8826 => x"76723477",
          8827 => x"81133484",
          8828 => x"b9fc0870",
          8829 => x"17703381",
          8830 => x"1233718b",
          8831 => x"2b71832b",
          8832 => x"07740570",
          8833 => x"33811233",
          8834 => x"71882b07",
          8835 => x"70832b8f",
          8836 => x"fff80677",
          8837 => x"057b882a",
          8838 => x"54525354",
          8839 => x"5c5a5754",
          8840 => x"52778214",
          8841 => x"34738314",
          8842 => x"3484b9fc",
          8843 => x"08701770",
          8844 => x"33811233",
          8845 => x"718b2b71",
          8846 => x"832b0774",
          8847 => x"05703381",
          8848 => x"12337188",
          8849 => x"2b0781ff",
          8850 => x"ff067088",
          8851 => x"2a5f5253",
          8852 => x"555a5754",
          8853 => x"52777334",
          8854 => x"70811434",
          8855 => x"84b9fc08",
          8856 => x"70178211",
          8857 => x"33831233",
          8858 => x"718b2b71",
          8859 => x"832b0774",
          8860 => x"05703381",
          8861 => x"12337198",
          8862 => x"2b71902b",
          8863 => x"0758535d",
          8864 => x"525a5753",
          8865 => x"53708025",
          8866 => x"fce43871",
          8867 => x"33811333",
          8868 => x"71882b07",
          8869 => x"82808007",
          8870 => x"70882a59",
          8871 => x"59547675",
          8872 => x"34778116",
          8873 => x"3484b9fc",
          8874 => x"08701770",
          8875 => x"33811233",
          8876 => x"718b2b71",
          8877 => x"832b0774",
          8878 => x"05821433",
          8879 => x"83153371",
          8880 => x"882b0770",
          8881 => x"882a575c",
          8882 => x"5c525856",
          8883 => x"52537282",
          8884 => x"15347583",
          8885 => x"1534893d",
          8886 => x"0d04f93d",
          8887 => x"0d7984b9",
          8888 => x"fc085858",
          8889 => x"76802e8f",
          8890 => x"3877802e",
          8891 => x"86387751",
          8892 => x"fb903f89",
          8893 => x"3d0d0484",
          8894 => x"fff40b84",
          8895 => x"b9fc0ca0",
          8896 => x"800b84b9",
          8897 => x"f8238280",
          8898 => x"80537652",
          8899 => x"84fff451",
          8900 => x"fed2ec3f",
          8901 => x"84b9fc08",
          8902 => x"55767534",
          8903 => x"810b8116",
          8904 => x"3484b9fc",
          8905 => x"08547684",
          8906 => x"1534810b",
          8907 => x"85153484",
          8908 => x"b9fc0856",
          8909 => x"76861734",
          8910 => x"810b8717",
          8911 => x"3484b9fc",
          8912 => x"0884b9f8",
          8913 => x"22ff05fe",
          8914 => x"80800770",
          8915 => x"83ffff06",
          8916 => x"70882a58",
          8917 => x"51555674",
          8918 => x"88173473",
          8919 => x"89173484",
          8920 => x"b9f82270",
          8921 => x"10101084",
          8922 => x"b9fc0805",
          8923 => x"f8055555",
          8924 => x"76821534",
          8925 => x"810b8315",
          8926 => x"34feee39",
          8927 => x"f73d0d7b",
          8928 => x"52805381",
          8929 => x"51847227",
          8930 => x"8e38fb12",
          8931 => x"832a8205",
          8932 => x"7083ffff",
          8933 => x"06515170",
          8934 => x"83ffff06",
          8935 => x"84b9fc08",
          8936 => x"84113385",
          8937 => x"12337188",
          8938 => x"2b077052",
          8939 => x"595a5855",
          8940 => x"81ffff54",
          8941 => x"75802e80",
          8942 => x"cc387510",
          8943 => x"10101770",
          8944 => x"33811233",
          8945 => x"71882b07",
          8946 => x"7081ffff",
          8947 => x"06793170",
          8948 => x"83ffff06",
          8949 => x"707a2756",
          8950 => x"535c5c54",
          8951 => x"52727427",
          8952 => x"8a387080",
          8953 => x"2e853875",
          8954 => x"73555884",
          8955 => x"12338513",
          8956 => x"3371882b",
          8957 => x"07575a75",
          8958 => x"c1387381",
          8959 => x"ffff2e85",
          8960 => x"38777454",
          8961 => x"56807683",
          8962 => x"2b781170",
          8963 => x"33811233",
          8964 => x"71882b07",
          8965 => x"7081ffff",
          8966 => x"0656565d",
          8967 => x"56595970",
          8968 => x"792e8338",
          8969 => x"81598051",
          8970 => x"74732682",
          8971 => x"8d387851",
          8972 => x"78802e82",
          8973 => x"85387275",
          8974 => x"2e828838",
          8975 => x"74167083",
          8976 => x"2b781174",
          8977 => x"82808007",
          8978 => x"70882a5b",
          8979 => x"5c56565a",
          8980 => x"76743478",
          8981 => x"81153484",
          8982 => x"b9fc0815",
          8983 => x"76882a53",
          8984 => x"53718214",
          8985 => x"34758314",
          8986 => x"3484b9fc",
          8987 => x"08701970",
          8988 => x"33811233",
          8989 => x"71882b07",
          8990 => x"70832b8f",
          8991 => x"fff80674",
          8992 => x"057e83ff",
          8993 => x"ff067088",
          8994 => x"2a5c5853",
          8995 => x"57595252",
          8996 => x"75821234",
          8997 => x"7281ff06",
          8998 => x"53728312",
          8999 => x"3484b9fc",
          9000 => x"08185475",
          9001 => x"74347281",
          9002 => x"153484b9",
          9003 => x"fc087019",
          9004 => x"86113387",
          9005 => x"1233718b",
          9006 => x"2b71832b",
          9007 => x"07740558",
          9008 => x"5c5c5357",
          9009 => x"75841534",
          9010 => x"72851534",
          9011 => x"84b9fc08",
          9012 => x"70165578",
          9013 => x"05861133",
          9014 => x"87123371",
          9015 => x"882b0770",
          9016 => x"882a5454",
          9017 => x"58597086",
          9018 => x"15347187",
          9019 => x"153484b9",
          9020 => x"fc087019",
          9021 => x"84113385",
          9022 => x"1233718b",
          9023 => x"2b71832b",
          9024 => x"07740558",
          9025 => x"5a5c5a52",
          9026 => x"75861534",
          9027 => x"72871534",
          9028 => x"84b9fc08",
          9029 => x"70165578",
          9030 => x"05841133",
          9031 => x"85123371",
          9032 => x"882b0770",
          9033 => x"882a545c",
          9034 => x"57597084",
          9035 => x"15347985",
          9036 => x"153484b9",
          9037 => x"fc081884",
          9038 => x"05517084",
          9039 => x"ba8c0c8b",
          9040 => x"3d0d0486",
          9041 => x"14338715",
          9042 => x"33718b2b",
          9043 => x"71832b07",
          9044 => x"79058417",
          9045 => x"33851833",
          9046 => x"71882b07",
          9047 => x"70882a5a",
          9048 => x"5b595354",
          9049 => x"52748412",
          9050 => x"34768512",
          9051 => x"3484b9fc",
          9052 => x"08701984",
          9053 => x"11338512",
          9054 => x"33718b2b",
          9055 => x"71832b07",
          9056 => x"74058614",
          9057 => x"33871533",
          9058 => x"71882b07",
          9059 => x"70882a58",
          9060 => x"5d5f5256",
          9061 => x"5b575270",
          9062 => x"861a3476",
          9063 => x"871a3484",
          9064 => x"b9fc0818",
          9065 => x"70338112",
          9066 => x"3371882b",
          9067 => x"0781ffff",
          9068 => x"0670882a",
          9069 => x"59575457",
          9070 => x"75773474",
          9071 => x"81183484",
          9072 => x"b9fc0818",
          9073 => x"840551fe",
          9074 => x"f139f93d",
          9075 => x"0d7984b9",
          9076 => x"fc085858",
          9077 => x"76802ea0",
          9078 => x"38775477",
          9079 => x"8a387384",
          9080 => x"ba8c0c89",
          9081 => x"3d0d0477",
          9082 => x"51fb913f",
          9083 => x"84ba8c08",
          9084 => x"84ba8c0c",
          9085 => x"893d0d04",
          9086 => x"84fff40b",
          9087 => x"84b9fc0c",
          9088 => x"a0800b84",
          9089 => x"b9f82382",
          9090 => x"80805376",
          9091 => x"5284fff4",
          9092 => x"51fecceb",
          9093 => x"3f84b9fc",
          9094 => x"08557675",
          9095 => x"34810b81",
          9096 => x"163484b9",
          9097 => x"fc085476",
          9098 => x"84153481",
          9099 => x"0b851534",
          9100 => x"84b9fc08",
          9101 => x"56768617",
          9102 => x"34810b87",
          9103 => x"173484b9",
          9104 => x"fc0884b9",
          9105 => x"f822ff05",
          9106 => x"fe808007",
          9107 => x"7083ffff",
          9108 => x"0670882a",
          9109 => x"58515556",
          9110 => x"74881734",
          9111 => x"73891734",
          9112 => x"84b9f822",
          9113 => x"70101010",
          9114 => x"84b9fc08",
          9115 => x"05f80555",
          9116 => x"55768215",
          9117 => x"34810b83",
          9118 => x"15347754",
          9119 => x"77802efe",
          9120 => x"dd38fee3",
          9121 => x"39ed3d0d",
          9122 => x"6567415f",
          9123 => x"807084b9",
          9124 => x"fc085945",
          9125 => x"4176612e",
          9126 => x"84aa387e",
          9127 => x"802e85af",
          9128 => x"387f802e",
          9129 => x"88d73881",
          9130 => x"54846027",
          9131 => x"8f387ffb",
          9132 => x"05832a82",
          9133 => x"057083ff",
          9134 => x"ff065558",
          9135 => x"7383ffff",
          9136 => x"067f7831",
          9137 => x"832a7083",
          9138 => x"ffff0670",
          9139 => x"832b7a11",
          9140 => x"70338112",
          9141 => x"3371882b",
          9142 => x"07707531",
          9143 => x"7083ffff",
          9144 => x"06701010",
          9145 => x"10fc0573",
          9146 => x"832b6111",
          9147 => x"70338112",
          9148 => x"3371882b",
          9149 => x"0770902b",
          9150 => x"70902c53",
          9151 => x"42454644",
          9152 => x"53544344",
          9153 => x"5c485952",
          9154 => x"5e5f4280",
          9155 => x"7a2485fd",
          9156 => x"38821533",
          9157 => x"83163371",
          9158 => x"882b0770",
          9159 => x"10101019",
          9160 => x"70338112",
          9161 => x"3371982b",
          9162 => x"71902b07",
          9163 => x"535c5356",
          9164 => x"56568074",
          9165 => x"2485c938",
          9166 => x"7a622782",
          9167 => x"f638631b",
          9168 => x"5877622e",
          9169 => x"87a23860",
          9170 => x"802e85f9",
          9171 => x"38601b58",
          9172 => x"77622587",
          9173 => x"be386318",
          9174 => x"59617924",
          9175 => x"92f73876",
          9176 => x"1e703381",
          9177 => x"1233718b",
          9178 => x"2b71832b",
          9179 => x"077a1170",
          9180 => x"33811233",
          9181 => x"71982b71",
          9182 => x"902b0747",
          9183 => x"43595253",
          9184 => x"575b5880",
          9185 => x"60248cba",
          9186 => x"38761e82",
          9187 => x"11338312",
          9188 => x"33718b2b",
          9189 => x"71832b07",
          9190 => x"7a118611",
          9191 => x"33871233",
          9192 => x"718b2b71",
          9193 => x"832b077e",
          9194 => x"05841433",
          9195 => x"85153371",
          9196 => x"882b0770",
          9197 => x"882a5957",
          9198 => x"48525b41",
          9199 => x"58535c59",
          9200 => x"5677841d",
          9201 => x"3479851d",
          9202 => x"3484b9fc",
          9203 => x"08701784",
          9204 => x"11338512",
          9205 => x"33718b2b",
          9206 => x"71832b07",
          9207 => x"74058614",
          9208 => x"33871533",
          9209 => x"71882b07",
          9210 => x"70882a5f",
          9211 => x"425e5240",
          9212 => x"57415777",
          9213 => x"8616347b",
          9214 => x"87163484",
          9215 => x"b9fc0816",
          9216 => x"70338112",
          9217 => x"3371882b",
          9218 => x"0781ffff",
          9219 => x"0670882a",
          9220 => x"5a5c5e59",
          9221 => x"76793479",
          9222 => x"811a3484",
          9223 => x"b9fc0870",
          9224 => x"1f821133",
          9225 => x"83123371",
          9226 => x"8b2b7183",
          9227 => x"2b077405",
          9228 => x"73338115",
          9229 => x"3371882b",
          9230 => x"0770882a",
          9231 => x"415c455d",
          9232 => x"5f5a5555",
          9233 => x"79793475",
          9234 => x"811a3484",
          9235 => x"b9fc0870",
          9236 => x"1f703381",
          9237 => x"1233718b",
          9238 => x"2b71832b",
          9239 => x"07740582",
          9240 => x"14338315",
          9241 => x"3371882b",
          9242 => x"0770882a",
          9243 => x"415c455d",
          9244 => x"5f5a5555",
          9245 => x"79821a34",
          9246 => x"75831a34",
          9247 => x"84b9fc08",
          9248 => x"701f8211",
          9249 => x"33831233",
          9250 => x"71882b07",
          9251 => x"66576256",
          9252 => x"70832b42",
          9253 => x"525a5d7e",
          9254 => x"05840551",
          9255 => x"fec4a33f",
          9256 => x"84b9fc08",
          9257 => x"1e840561",
          9258 => x"65051c70",
          9259 => x"83ffff06",
          9260 => x"5d445f7a",
          9261 => x"622681b6",
          9262 => x"387e5473",
          9263 => x"84ba8c0c",
          9264 => x"953d0d04",
          9265 => x"84fff40b",
          9266 => x"84b9fc0c",
          9267 => x"a0800b84",
          9268 => x"b9f82382",
          9269 => x"80805360",
          9270 => x"5284fff4",
          9271 => x"51fec79f",
          9272 => x"3f84b9fc",
          9273 => x"085e607e",
          9274 => x"34810b81",
          9275 => x"1f3484b9",
          9276 => x"fc085d60",
          9277 => x"841e3481",
          9278 => x"0b851e34",
          9279 => x"84b9fc08",
          9280 => x"5c60861d",
          9281 => x"34810b87",
          9282 => x"1d3484b9",
          9283 => x"fc0884b9",
          9284 => x"f822ff05",
          9285 => x"fe808007",
          9286 => x"7083ffff",
          9287 => x"0670882a",
          9288 => x"5c5a5b57",
          9289 => x"78881834",
          9290 => x"77891834",
          9291 => x"84b9f822",
          9292 => x"70101010",
          9293 => x"84b9fc08",
          9294 => x"05f80555",
          9295 => x"56608215",
          9296 => x"34810b83",
          9297 => x"153484b9",
          9298 => x"fc08577e",
          9299 => x"fad33876",
          9300 => x"802e828c",
          9301 => x"387e547f",
          9302 => x"802efedf",
          9303 => x"387f51f4",
          9304 => x"9b3f84ba",
          9305 => x"8c0884ba",
          9306 => x"8c0c953d",
          9307 => x"0d04611c",
          9308 => x"84b9fc08",
          9309 => x"71832b71",
          9310 => x"115e447f",
          9311 => x"05703381",
          9312 => x"12337188",
          9313 => x"2b0781ff",
          9314 => x"ff067088",
          9315 => x"2a48445b",
          9316 => x"5e40637b",
          9317 => x"3460811c",
          9318 => x"346184b9",
          9319 => x"fc08057c",
          9320 => x"882a5758",
          9321 => x"75821934",
          9322 => x"7b831934",
          9323 => x"84b9fc08",
          9324 => x"701f7033",
          9325 => x"81123371",
          9326 => x"882b0770",
          9327 => x"832b8fff",
          9328 => x"f8067405",
          9329 => x"6483ffff",
          9330 => x"0670882a",
          9331 => x"4a5c4757",
          9332 => x"5e5b5d63",
          9333 => x"63820534",
          9334 => x"7681ff06",
          9335 => x"41606383",
          9336 => x"053484b9",
          9337 => x"fc081e5b",
          9338 => x"637b3460",
          9339 => x"811c3461",
          9340 => x"84b9fc08",
          9341 => x"05840551",
          9342 => x"ed883f7e",
          9343 => x"54fdbc39",
          9344 => x"7b753170",
          9345 => x"83ffff06",
          9346 => x"4254faac",
          9347 => x"397781ff",
          9348 => x"ff067631",
          9349 => x"7083ffff",
          9350 => x"06821733",
          9351 => x"83183371",
          9352 => x"882b0770",
          9353 => x"1010101b",
          9354 => x"70338112",
          9355 => x"3371982b",
          9356 => x"71902b07",
          9357 => x"535e5354",
          9358 => x"58584554",
          9359 => x"738025f9",
          9360 => x"f738ffbc",
          9361 => x"39617824",
          9362 => x"fa833880",
          9363 => x"7a248b8f",
          9364 => x"387783ff",
          9365 => x"ff065b61",
          9366 => x"7b27fcdd",
          9367 => x"38fe8f39",
          9368 => x"84fff40b",
          9369 => x"84b9fc0c",
          9370 => x"a0800b84",
          9371 => x"b9f82382",
          9372 => x"8080537e",
          9373 => x"5284fff4",
          9374 => x"51fec483",
          9375 => x"3f84b9fc",
          9376 => x"085a7e7a",
          9377 => x"34810b81",
          9378 => x"1b3484b9",
          9379 => x"fc08597e",
          9380 => x"841a3481",
          9381 => x"0b851a34",
          9382 => x"84b9fc08",
          9383 => x"587e8619",
          9384 => x"34810b87",
          9385 => x"193484b9",
          9386 => x"fc0884b9",
          9387 => x"f822ff05",
          9388 => x"fe808007",
          9389 => x"7083ffff",
          9390 => x"0670882a",
          9391 => x"58565744",
          9392 => x"74648805",
          9393 => x"34736489",
          9394 => x"053484b9",
          9395 => x"f8227010",
          9396 => x"101084b9",
          9397 => x"fc0805f8",
          9398 => x"0542437e",
          9399 => x"61820534",
          9400 => x"81618305",
          9401 => x"34fcee39",
          9402 => x"807a2483",
          9403 => x"de386183",
          9404 => x"ffff065b",
          9405 => x"617b27fb",
          9406 => x"c038fcf2",
          9407 => x"3976802e",
          9408 => x"82bd387e",
          9409 => x"51eafb3f",
          9410 => x"7f547384",
          9411 => x"ba8c0c95",
          9412 => x"3d0d0476",
          9413 => x"1e821133",
          9414 => x"83123371",
          9415 => x"8b2b7183",
          9416 => x"2b077a11",
          9417 => x"86113387",
          9418 => x"1233718b",
          9419 => x"2b71832b",
          9420 => x"077e0584",
          9421 => x"14338515",
          9422 => x"3371882b",
          9423 => x"0770882a",
          9424 => x"43444556",
          9425 => x"5b465853",
          9426 => x"5c455678",
          9427 => x"64840534",
          9428 => x"7a648505",
          9429 => x"3484b9fc",
          9430 => x"08701784",
          9431 => x"11338512",
          9432 => x"33718b2b",
          9433 => x"71832b07",
          9434 => x"74058614",
          9435 => x"33871533",
          9436 => x"71882b07",
          9437 => x"70882a5b",
          9438 => x"4142485d",
          9439 => x"595d4173",
          9440 => x"64860534",
          9441 => x"7a648705",
          9442 => x"3484b9fc",
          9443 => x"08167033",
          9444 => x"81123371",
          9445 => x"882b0781",
          9446 => x"ffff0670",
          9447 => x"882a5f5c",
          9448 => x"5a5d7b7d",
          9449 => x"3479811e",
          9450 => x"3484b9fc",
          9451 => x"08701f82",
          9452 => x"11338312",
          9453 => x"33718b2b",
          9454 => x"71832b07",
          9455 => x"74057333",
          9456 => x"81153371",
          9457 => x"882b0770",
          9458 => x"882a5e5c",
          9459 => x"5e404357",
          9460 => x"4554767c",
          9461 => x"3475811d",
          9462 => x"3484b9fc",
          9463 => x"08701f70",
          9464 => x"33811233",
          9465 => x"718b2b71",
          9466 => x"832b0774",
          9467 => x"05821433",
          9468 => x"83153371",
          9469 => x"882b0770",
          9470 => x"882a4047",
          9471 => x"405b405c",
          9472 => x"55557882",
          9473 => x"18346083",
          9474 => x"183484b9",
          9475 => x"fc08701f",
          9476 => x"82113383",
          9477 => x"12337188",
          9478 => x"2b076657",
          9479 => x"62567083",
          9480 => x"2b425258",
          9481 => x"5d7e0584",
          9482 => x"0551febd",
          9483 => x"953f84b9",
          9484 => x"fc081e84",
          9485 => x"057883ff",
          9486 => x"ff065c5f",
          9487 => x"fc993984",
          9488 => x"fff40b84",
          9489 => x"b9fc0ca0",
          9490 => x"800b84b9",
          9491 => x"f8238280",
          9492 => x"80537f52",
          9493 => x"84fff451",
          9494 => x"fec0a43f",
          9495 => x"84b9fc08",
          9496 => x"567f7634",
          9497 => x"810b8117",
          9498 => x"3484b9fc",
          9499 => x"08557f84",
          9500 => x"1634810b",
          9501 => x"85163484",
          9502 => x"b9fc0854",
          9503 => x"7f861534",
          9504 => x"810b8715",
          9505 => x"3484b9fc",
          9506 => x"0884b9f8",
          9507 => x"22ff05fe",
          9508 => x"80800770",
          9509 => x"83ffff06",
          9510 => x"70882a45",
          9511 => x"43445e61",
          9512 => x"881f3460",
          9513 => x"891f3484",
          9514 => x"b9f82270",
          9515 => x"10101084",
          9516 => x"b9fc0805",
          9517 => x"f8055c5d",
          9518 => x"7f821c34",
          9519 => x"810b831c",
          9520 => x"347e51e7",
          9521 => x"bd3f7f54",
          9522 => x"fcc03986",
          9523 => x"1933871a",
          9524 => x"33718b2b",
          9525 => x"71832b07",
          9526 => x"7905841c",
          9527 => x"33851d33",
          9528 => x"71882b07",
          9529 => x"70882a5c",
          9530 => x"485e4359",
          9531 => x"55766184",
          9532 => x"05346361",
          9533 => x"85053484",
          9534 => x"b9fc0870",
          9535 => x"1e841133",
          9536 => x"85123371",
          9537 => x"8b2b7183",
          9538 => x"2b077405",
          9539 => x"86143387",
          9540 => x"15337188",
          9541 => x"2b077088",
          9542 => x"2a415f48",
          9543 => x"48595659",
          9544 => x"40796486",
          9545 => x"05347864",
          9546 => x"87053484",
          9547 => x"b9fc081d",
          9548 => x"70338112",
          9549 => x"3371882b",
          9550 => x"0781ffff",
          9551 => x"0670882a",
          9552 => x"59425858",
          9553 => x"7578347f",
          9554 => x"81193484",
          9555 => x"b9fc0870",
          9556 => x"1f703381",
          9557 => x"1233718b",
          9558 => x"2b71832b",
          9559 => x"07740570",
          9560 => x"33811233",
          9561 => x"71882b07",
          9562 => x"70832b8f",
          9563 => x"fff80677",
          9564 => x"0563882a",
          9565 => x"485d5d5a",
          9566 => x"5d405d44",
          9567 => x"417f8217",
          9568 => x"347b8317",
          9569 => x"3484b9fc",
          9570 => x"08701f70",
          9571 => x"33811233",
          9572 => x"718b2b71",
          9573 => x"832b0774",
          9574 => x"05703381",
          9575 => x"12337188",
          9576 => x"2b0781ff",
          9577 => x"ff067088",
          9578 => x"2a485d5e",
          9579 => x"5e465a41",
          9580 => x"5b606034",
          9581 => x"76608105",
          9582 => x"346183ff",
          9583 => x"ff065bfa",
          9584 => x"b3398615",
          9585 => x"33871633",
          9586 => x"718b2b71",
          9587 => x"832b0779",
          9588 => x"05841833",
          9589 => x"85193371",
          9590 => x"882b0770",
          9591 => x"882a5e5e",
          9592 => x"5a52415d",
          9593 => x"78841e34",
          9594 => x"79851e34",
          9595 => x"84b9fc08",
          9596 => x"70198411",
          9597 => x"33851233",
          9598 => x"718b2b71",
          9599 => x"832b0774",
          9600 => x"05861433",
          9601 => x"87153371",
          9602 => x"882b0770",
          9603 => x"882a4456",
          9604 => x"5e525a42",
          9605 => x"55567c60",
          9606 => x"86053475",
          9607 => x"60870534",
          9608 => x"84b9fc08",
          9609 => x"18703381",
          9610 => x"12337188",
          9611 => x"2b0781ff",
          9612 => x"ff067088",
          9613 => x"2a5b5b58",
          9614 => x"55777534",
          9615 => x"78811634",
          9616 => x"84b9fc08",
          9617 => x"701f7033",
          9618 => x"81123371",
          9619 => x"8b2b7183",
          9620 => x"2b077405",
          9621 => x"70338112",
          9622 => x"3371882b",
          9623 => x"0770832b",
          9624 => x"8ffff806",
          9625 => x"77056388",
          9626 => x"2a56545f",
          9627 => x"5f585942",
          9628 => x"5e557f82",
          9629 => x"17347b83",
          9630 => x"173484b9",
          9631 => x"fc08701f",
          9632 => x"70338112",
          9633 => x"33718b2b",
          9634 => x"71832b07",
          9635 => x"74057033",
          9636 => x"81123371",
          9637 => x"882b0781",
          9638 => x"ffff0670",
          9639 => x"882a5d54",
          9640 => x"5e585b59",
          9641 => x"5d55757c",
          9642 => x"3476811d",
          9643 => x"3484b9fc",
          9644 => x"08701f82",
          9645 => x"11338312",
          9646 => x"33718b2b",
          9647 => x"71832b07",
          9648 => x"74118611",
          9649 => x"33871233",
          9650 => x"718b2b71",
          9651 => x"832b0778",
          9652 => x"05841433",
          9653 => x"85153371",
          9654 => x"882b0770",
          9655 => x"882a5957",
          9656 => x"49525c42",
          9657 => x"59535d5a",
          9658 => x"57577784",
          9659 => x"1d347985",
          9660 => x"1d3484b9",
          9661 => x"fc087017",
          9662 => x"84113385",
          9663 => x"1233718b",
          9664 => x"2b71832b",
          9665 => x"07740586",
          9666 => x"14338715",
          9667 => x"3371882b",
          9668 => x"0770882a",
          9669 => x"5f425e52",
          9670 => x"40574157",
          9671 => x"77861634",
          9672 => x"7b871634",
          9673 => x"84b9fc08",
          9674 => x"16703381",
          9675 => x"12337188",
          9676 => x"2b0781ff",
          9677 => x"ff067088",
          9678 => x"2a5a5c5e",
          9679 => x"59767934",
          9680 => x"79811a34",
          9681 => x"84b9fc08",
          9682 => x"701f8211",
          9683 => x"33831233",
          9684 => x"718b2b71",
          9685 => x"832b0774",
          9686 => x"05733381",
          9687 => x"15337188",
          9688 => x"2b077088",
          9689 => x"2a415c45",
          9690 => x"5d5f5a55",
          9691 => x"55797934",
          9692 => x"75811a34",
          9693 => x"84b9fc08",
          9694 => x"701f7033",
          9695 => x"81123371",
          9696 => x"8b2b7183",
          9697 => x"2b077405",
          9698 => x"82143383",
          9699 => x"15337188",
          9700 => x"2b077088",
          9701 => x"2a415c45",
          9702 => x"5d5f5a55",
          9703 => x"5579821a",
          9704 => x"3475831a",
          9705 => x"3484b9fc",
          9706 => x"08701f82",
          9707 => x"11338312",
          9708 => x"3371882b",
          9709 => x"07665762",
          9710 => x"5670832b",
          9711 => x"42525a5d",
          9712 => x"7e058405",
          9713 => x"51feb5fa",
          9714 => x"3f84b9fc",
          9715 => x"081e8405",
          9716 => x"6165051c",
          9717 => x"7083ffff",
          9718 => x"065d445f",
          9719 => x"f1d53986",
          9720 => x"1933871a",
          9721 => x"33718b2b",
          9722 => x"71832b07",
          9723 => x"7905841c",
          9724 => x"33851d33",
          9725 => x"71882b07",
          9726 => x"70882a40",
          9727 => x"485d4341",
          9728 => x"557a6184",
          9729 => x"05346361",
          9730 => x"85053484",
          9731 => x"b9fc0870",
          9732 => x"1e841133",
          9733 => x"85123371",
          9734 => x"8b2b7183",
          9735 => x"2b077405",
          9736 => x"86143387",
          9737 => x"15337188",
          9738 => x"2b077088",
          9739 => x"2a5b415f",
          9740 => x"485c5941",
          9741 => x"56736486",
          9742 => x"05347a64",
          9743 => x"87053484",
          9744 => x"b9fc081d",
          9745 => x"70338112",
          9746 => x"3371882b",
          9747 => x"0781ffff",
          9748 => x"0670882a",
          9749 => x"5c5f4255",
          9750 => x"7875347c",
          9751 => x"81163484",
          9752 => x"b9fc0870",
          9753 => x"1f703381",
          9754 => x"1233718b",
          9755 => x"2b71832b",
          9756 => x"07740570",
          9757 => x"33811233",
          9758 => x"71882b07",
          9759 => x"70832b8f",
          9760 => x"fff80677",
          9761 => x"0563882a",
          9762 => x"5d445c49",
          9763 => x"585e4558",
          9764 => x"4074821e",
          9765 => x"347b831e",
          9766 => x"3484b9fc",
          9767 => x"08701f70",
          9768 => x"33811233",
          9769 => x"718b2b71",
          9770 => x"832b0774",
          9771 => x"05703381",
          9772 => x"12337188",
          9773 => x"2b0781ff",
          9774 => x"ff067088",
          9775 => x"2a475f49",
          9776 => x"5846595e",
          9777 => x"5b7f7d34",
          9778 => x"78811e34",
          9779 => x"7783ffff",
          9780 => x"065bf383",
          9781 => x"397e6052",
          9782 => x"54e5a13f",
          9783 => x"84ba8c08",
          9784 => x"5f84ba8c",
          9785 => x"08802e93",
          9786 => x"38625373",
          9787 => x"5284ba8c",
          9788 => x"0851feb4",
          9789 => x"f53f7351",
          9790 => x"df883f61",
          9791 => x"5b617b27",
          9792 => x"efb738f0",
          9793 => x"e939f93d",
          9794 => x"0d7a7a29",
          9795 => x"84b9fc08",
          9796 => x"58587680",
          9797 => x"2eb73877",
          9798 => x"54778a38",
          9799 => x"7384ba8c",
          9800 => x"0c893d0d",
          9801 => x"047751e4",
          9802 => x"d33f84ba",
          9803 => x"8c085484",
          9804 => x"ba8c0880",
          9805 => x"2ee63877",
          9806 => x"53805284",
          9807 => x"ba8c0851",
          9808 => x"feb6bc3f",
          9809 => x"7384ba8c",
          9810 => x"0c893d0d",
          9811 => x"0484fff4",
          9812 => x"0b84b9fc",
          9813 => x"0ca0800b",
          9814 => x"84b9f823",
          9815 => x"82808053",
          9816 => x"765284ff",
          9817 => x"f451feb6",
          9818 => x"963f84b9",
          9819 => x"fc085576",
          9820 => x"7534810b",
          9821 => x"81163484",
          9822 => x"b9fc0854",
          9823 => x"76841534",
          9824 => x"810b8515",
          9825 => x"3484b9fc",
          9826 => x"08567686",
          9827 => x"1734810b",
          9828 => x"87173484",
          9829 => x"b9fc0884",
          9830 => x"b9f822ff",
          9831 => x"05fe8080",
          9832 => x"077083ff",
          9833 => x"ff067088",
          9834 => x"2a585155",
          9835 => x"56748817",
          9836 => x"34738917",
          9837 => x"3484b9f8",
          9838 => x"22701010",
          9839 => x"1084b9fc",
          9840 => x"0805f805",
          9841 => x"55557682",
          9842 => x"1534810b",
          9843 => x"83153477",
          9844 => x"5477802e",
          9845 => x"fec638fe",
          9846 => x"cc39ff3d",
          9847 => x"0d028f05",
          9848 => x"33518152",
          9849 => x"70722687",
          9850 => x"3884ba88",
          9851 => x"11335271",
          9852 => x"84ba8c0c",
          9853 => x"833d0d04",
          9854 => x"fe3d0d02",
          9855 => x"93053352",
          9856 => x"83537181",
          9857 => x"269d3871",
          9858 => x"51d3ec3f",
          9859 => x"84ba8c08",
          9860 => x"81ff0653",
          9861 => x"72873872",
          9862 => x"84ba8813",
          9863 => x"3484ba88",
          9864 => x"12335372",
          9865 => x"84ba8c0c",
          9866 => x"843d0d04",
          9867 => x"f73d0d7c",
          9868 => x"7e60028c",
          9869 => x"05af0533",
          9870 => x"5a5c5759",
          9871 => x"81547674",
          9872 => x"26873884",
          9873 => x"ba881733",
          9874 => x"54738106",
          9875 => x"54835573",
          9876 => x"bd387358",
          9877 => x"850b87c0",
          9878 => x"988c0c78",
          9879 => x"53755276",
          9880 => x"51d58d3f",
          9881 => x"84ba8c08",
          9882 => x"81ff0655",
          9883 => x"74802ea7",
          9884 => x"3887c098",
          9885 => x"8c085473",
          9886 => x"e2387978",
          9887 => x"26d63874",
          9888 => x"fc808006",
          9889 => x"5473802e",
          9890 => x"83388154",
          9891 => x"73557484",
          9892 => x"ba8c0c8b",
          9893 => x"3d0d0484",
          9894 => x"80168119",
          9895 => x"7081ff06",
          9896 => x"5a555679",
          9897 => x"7826ffac",
          9898 => x"38d539f7",
          9899 => x"3d0d7c7e",
          9900 => x"60028c05",
          9901 => x"af05335a",
          9902 => x"5c575981",
          9903 => x"54767426",
          9904 => x"873884ba",
          9905 => x"88173354",
          9906 => x"73810654",
          9907 => x"835573bd",
          9908 => x"38735885",
          9909 => x"0b87c098",
          9910 => x"8c0c7853",
          9911 => x"75527651",
          9912 => x"d6e73f84",
          9913 => x"ba8c0881",
          9914 => x"ff065574",
          9915 => x"802ea738",
          9916 => x"87c0988c",
          9917 => x"085473e2",
          9918 => x"38797826",
          9919 => x"d63874fc",
          9920 => x"80800654",
          9921 => x"73802e83",
          9922 => x"38815473",
          9923 => x"557484ba",
          9924 => x"8c0c8b3d",
          9925 => x"0d048480",
          9926 => x"16811970",
          9927 => x"81ff065a",
          9928 => x"55567978",
          9929 => x"26ffac38",
          9930 => x"d539fc3d",
          9931 => x"0d780284",
          9932 => x"059b0533",
          9933 => x"0288059f",
          9934 => x"05335353",
          9935 => x"55815371",
          9936 => x"73268738",
          9937 => x"84ba8812",
          9938 => x"33537281",
          9939 => x"06548353",
          9940 => x"739b3885",
          9941 => x"0b87c098",
          9942 => x"8c0c8153",
          9943 => x"70732e96",
          9944 => x"38727125",
          9945 => x"ad387083",
          9946 => x"2e9a3884",
          9947 => x"537284ba",
          9948 => x"8c0c863d",
          9949 => x"0d048880",
          9950 => x"0a750c73",
          9951 => x"84ba8c0c",
          9952 => x"863d0d04",
          9953 => x"8180750c",
          9954 => x"800b84ba",
          9955 => x"8c0c863d",
          9956 => x"0d047184",
          9957 => x"2b87c092",
          9958 => x"8c115354",
          9959 => x"70cd3871",
          9960 => x"0870812a",
          9961 => x"81065151",
          9962 => x"70802e8a",
          9963 => x"3887c098",
          9964 => x"8c085574",
          9965 => x"ea3887c0",
          9966 => x"988c0851",
          9967 => x"70ca3881",
          9968 => x"720c87c0",
          9969 => x"928c1452",
          9970 => x"71088206",
          9971 => x"5473802e",
          9972 => x"ff9b3871",
          9973 => x"08820654",
          9974 => x"73ee38ff",
          9975 => x"9039f63d",
          9976 => x"0d7c5880",
          9977 => x"0b831933",
          9978 => x"715b5657",
          9979 => x"74772e09",
          9980 => x"8106a838",
          9981 => x"77335675",
          9982 => x"832e8187",
          9983 => x"38805380",
          9984 => x"52811833",
          9985 => x"51fea33f",
          9986 => x"84ba8c08",
          9987 => x"802e8338",
          9988 => x"81597884",
          9989 => x"ba8c0c8c",
          9990 => x"3d0d0481",
          9991 => x"54b41808",
          9992 => x"53b81870",
          9993 => x"53811933",
          9994 => x"525afcff",
          9995 => x"3f815984",
          9996 => x"ba8c0877",
          9997 => x"2e098106",
          9998 => x"d93884ba",
          9999 => x"8c088319",
         10000 => x"34b41808",
         10001 => x"70a81a08",
         10002 => x"31a01a08",
         10003 => x"84ba8c08",
         10004 => x"5c58565b",
         10005 => x"747627ff",
         10006 => x"9b388218",
         10007 => x"33557482",
         10008 => x"2e098106",
         10009 => x"ff8e3881",
         10010 => x"54751b53",
         10011 => x"79528118",
         10012 => x"3351fcb7",
         10013 => x"3f767833",
         10014 => x"57597583",
         10015 => x"2e098106",
         10016 => x"fefb3884",
         10017 => x"18335776",
         10018 => x"812e0981",
         10019 => x"06feee38",
         10020 => x"b8185a84",
         10021 => x"807a5657",
         10022 => x"80757081",
         10023 => x"055734ff",
         10024 => x"175776f4",
         10025 => x"3880d50b",
         10026 => x"84b61934",
         10027 => x"ffaa0b84",
         10028 => x"b7193480",
         10029 => x"d27a3480",
         10030 => x"d20bb919",
         10031 => x"3480e10b",
         10032 => x"ba193480",
         10033 => x"c10bbb19",
         10034 => x"3480f20b",
         10035 => x"849c1934",
         10036 => x"80f20b84",
         10037 => x"9d193480",
         10038 => x"c10b849e",
         10039 => x"193480e1",
         10040 => x"0b849f19",
         10041 => x"34941808",
         10042 => x"557484a0",
         10043 => x"19347488",
         10044 => x"2a5b7a84",
         10045 => x"a1193474",
         10046 => x"902a5675",
         10047 => x"84a21934",
         10048 => x"74982a5b",
         10049 => x"7a84a319",
         10050 => x"34901808",
         10051 => x"5b7a84a4",
         10052 => x"19347a88",
         10053 => x"2a557484",
         10054 => x"a519347a",
         10055 => x"902a5675",
         10056 => x"84a61934",
         10057 => x"7a982a55",
         10058 => x"7484a719",
         10059 => x"34a41808",
         10060 => x"810570b4",
         10061 => x"1a0c5b81",
         10062 => x"547a5379",
         10063 => x"52811833",
         10064 => x"51fae83f",
         10065 => x"76841934",
         10066 => x"80538052",
         10067 => x"81183351",
         10068 => x"fbd83f84",
         10069 => x"ba8c0880",
         10070 => x"2efdb738",
         10071 => x"fdb239f3",
         10072 => x"3d0d6060",
         10073 => x"70085956",
         10074 => x"56817627",
         10075 => x"88389c17",
         10076 => x"0876268c",
         10077 => x"38815877",
         10078 => x"84ba8c0c",
         10079 => x"8f3d0d04",
         10080 => x"ff773356",
         10081 => x"5874822e",
         10082 => x"81cc3874",
         10083 => x"822482a5",
         10084 => x"3874812e",
         10085 => x"098106dd",
         10086 => x"3875812a",
         10087 => x"1670892a",
         10088 => x"a8190805",
         10089 => x"5a5a805b",
         10090 => x"b4170879",
         10091 => x"2eb03883",
         10092 => x"17335c7b",
         10093 => x"7b2e0981",
         10094 => x"0683de38",
         10095 => x"81547853",
         10096 => x"b8175281",
         10097 => x"173351f8",
         10098 => x"e33f84ba",
         10099 => x"8c08802e",
         10100 => x"8538ff59",
         10101 => x"815b78b4",
         10102 => x"180c7aff",
         10103 => x"9a387983",
         10104 => x"ff0617b8",
         10105 => x"1133811c",
         10106 => x"70892aa8",
         10107 => x"1b080553",
         10108 => x"5d5d59b4",
         10109 => x"1708792e",
         10110 => x"b538800b",
         10111 => x"83183371",
         10112 => x"5c565d74",
         10113 => x"7d2e0981",
         10114 => x"0684b538",
         10115 => x"81547853",
         10116 => x"b8175281",
         10117 => x"173351f8",
         10118 => x"933f84ba",
         10119 => x"8c08802e",
         10120 => x"8538ff59",
         10121 => x"815a78b4",
         10122 => x"180c79fe",
         10123 => x"ca387a83",
         10124 => x"ff0617b8",
         10125 => x"11337088",
         10126 => x"2b7e0778",
         10127 => x"81067184",
         10128 => x"2a535d59",
         10129 => x"595d79fe",
         10130 => x"ae38769f",
         10131 => x"ff0684ba",
         10132 => x"8c0c8f3d",
         10133 => x"0d047588",
         10134 => x"2aa81808",
         10135 => x"0559b417",
         10136 => x"08792eb5",
         10137 => x"38800b83",
         10138 => x"1833715c",
         10139 => x"5d5b7b7b",
         10140 => x"2e098106",
         10141 => x"81c23881",
         10142 => x"547853b8",
         10143 => x"17528117",
         10144 => x"3351f7a8",
         10145 => x"3f84ba8c",
         10146 => x"08802e85",
         10147 => x"38ff5981",
         10148 => x"5a78b418",
         10149 => x"0c79fddf",
         10150 => x"38751083",
         10151 => x"fe067705",
         10152 => x"b8058111",
         10153 => x"33713371",
         10154 => x"882b0784",
         10155 => x"ba8c0c57",
         10156 => x"5b8f3d0d",
         10157 => x"0474832e",
         10158 => x"098106fd",
         10159 => x"b8387587",
         10160 => x"2aa81808",
         10161 => x"0559b417",
         10162 => x"08792eb5",
         10163 => x"38800b83",
         10164 => x"1833715c",
         10165 => x"5e5b7c7b",
         10166 => x"2e098106",
         10167 => x"82813881",
         10168 => x"547853b8",
         10169 => x"17528117",
         10170 => x"3351f6c0",
         10171 => x"3f84ba8c",
         10172 => x"08802e85",
         10173 => x"38ff5981",
         10174 => x"5a78b418",
         10175 => x"0c79fcf7",
         10176 => x"3875822b",
         10177 => x"83fc0677",
         10178 => x"05b80583",
         10179 => x"11338212",
         10180 => x"3371902b",
         10181 => x"71882b07",
         10182 => x"81143370",
         10183 => x"7207882b",
         10184 => x"75337180",
         10185 => x"fffffe80",
         10186 => x"060784ba",
         10187 => x"8c0c415c",
         10188 => x"5e595a56",
         10189 => x"8f3d0d04",
         10190 => x"8154b417",
         10191 => x"0853b817",
         10192 => x"70538118",
         10193 => x"33525cf6",
         10194 => x"e23f815a",
         10195 => x"84ba8c08",
         10196 => x"7b2e0981",
         10197 => x"06febe38",
         10198 => x"84ba8c08",
         10199 => x"831834b4",
         10200 => x"1708a818",
         10201 => x"083184ba",
         10202 => x"8c085b5e",
         10203 => x"7da01808",
         10204 => x"27fe8438",
         10205 => x"82173355",
         10206 => x"74822e09",
         10207 => x"8106fdf7",
         10208 => x"388154b4",
         10209 => x"1708a018",
         10210 => x"0805537b",
         10211 => x"52811733",
         10212 => x"51f6983f",
         10213 => x"7a5afddf",
         10214 => x"398154b4",
         10215 => x"170853b8",
         10216 => x"17705381",
         10217 => x"1833525c",
         10218 => x"f6813f84",
         10219 => x"ba8c087b",
         10220 => x"2e098106",
         10221 => x"82813884",
         10222 => x"ba8c0883",
         10223 => x"1834b417",
         10224 => x"08a81808",
         10225 => x"315d7ca0",
         10226 => x"1808278b",
         10227 => x"38821733",
         10228 => x"5e7d822e",
         10229 => x"81cb3884",
         10230 => x"ba8c085b",
         10231 => x"fbde3981",
         10232 => x"54b41708",
         10233 => x"53b81770",
         10234 => x"53811833",
         10235 => x"525cf5bb",
         10236 => x"3f815a84",
         10237 => x"ba8c087b",
         10238 => x"2e098106",
         10239 => x"fdff3884",
         10240 => x"ba8c0883",
         10241 => x"1834b417",
         10242 => x"08a81808",
         10243 => x"3184ba8c",
         10244 => x"085b5e7d",
         10245 => x"a0180827",
         10246 => x"fdc53882",
         10247 => x"17335574",
         10248 => x"822e0981",
         10249 => x"06fdb838",
         10250 => x"8154b417",
         10251 => x"08a01808",
         10252 => x"05537b52",
         10253 => x"81173351",
         10254 => x"f4f13f7a",
         10255 => x"5afda039",
         10256 => x"8154b417",
         10257 => x"0853b817",
         10258 => x"70538118",
         10259 => x"33525ef4",
         10260 => x"da3f815a",
         10261 => x"84ba8c08",
         10262 => x"7d2e0981",
         10263 => x"06fbcb38",
         10264 => x"84ba8c08",
         10265 => x"831834b4",
         10266 => x"1708a818",
         10267 => x"083184ba",
         10268 => x"8c085b55",
         10269 => x"74a01808",
         10270 => x"27fb9138",
         10271 => x"82173355",
         10272 => x"74822e09",
         10273 => x"8106fb84",
         10274 => x"388154b4",
         10275 => x"1708a018",
         10276 => x"0805537d",
         10277 => x"52811733",
         10278 => x"51f4903f",
         10279 => x"7c5afaec",
         10280 => x"398154b4",
         10281 => x"1708a018",
         10282 => x"0805537b",
         10283 => x"52811733",
         10284 => x"51f3f83f",
         10285 => x"fa863981",
         10286 => x"5b7af9bb",
         10287 => x"38fa9f39",
         10288 => x"f23d0d60",
         10289 => x"62645d57",
         10290 => x"59825881",
         10291 => x"76279c38",
         10292 => x"759c1a08",
         10293 => x"27953878",
         10294 => x"33557478",
         10295 => x"2e963874",
         10296 => x"78248180",
         10297 => x"3874812e",
         10298 => x"828a3877",
         10299 => x"84ba8c0c",
         10300 => x"903d0d04",
         10301 => x"75882aa8",
         10302 => x"1a080558",
         10303 => x"800bb41a",
         10304 => x"08585c76",
         10305 => x"782e86b6",
         10306 => x"38831933",
         10307 => x"7c5b5d7c",
         10308 => x"7c2e0981",
         10309 => x"0683fa38",
         10310 => x"81547753",
         10311 => x"b8195281",
         10312 => x"193351f2",
         10313 => x"873f84ba",
         10314 => x"8c08802e",
         10315 => x"8538ff58",
         10316 => x"815a77b4",
         10317 => x"1a0c7958",
         10318 => x"79ffb038",
         10319 => x"751083fe",
         10320 => x"0679057b",
         10321 => x"83ffff06",
         10322 => x"585e76b8",
         10323 => x"1f347688",
         10324 => x"2a5a79b9",
         10325 => x"1f34810b",
         10326 => x"831a3477",
         10327 => x"84ba8c0c",
         10328 => x"903d0d04",
         10329 => x"74832e09",
         10330 => x"8106feff",
         10331 => x"3875872a",
         10332 => x"a81a0805",
         10333 => x"58800bb4",
         10334 => x"1a08585c",
         10335 => x"76782e85",
         10336 => x"e1388319",
         10337 => x"337c5b5d",
         10338 => x"7c7c2e09",
         10339 => x"810684bd",
         10340 => x"38815477",
         10341 => x"53b81952",
         10342 => x"81193351",
         10343 => x"f18e3f84",
         10344 => x"ba8c0880",
         10345 => x"2e8538ff",
         10346 => x"58815a77",
         10347 => x"b41a0c79",
         10348 => x"5879feb7",
         10349 => x"3875822b",
         10350 => x"83fc0679",
         10351 => x"05b81183",
         10352 => x"11337098",
         10353 => x"2b8f0a06",
         10354 => x"7ef00a06",
         10355 => x"0741575e",
         10356 => x"5c7d7d34",
         10357 => x"7d882a56",
         10358 => x"75b91d34",
         10359 => x"7d902a5a",
         10360 => x"79ba1d34",
         10361 => x"7d982a5b",
         10362 => x"7abb1d34",
         10363 => x"810b831a",
         10364 => x"34fee839",
         10365 => x"75812a16",
         10366 => x"70892aa8",
         10367 => x"1b0805b4",
         10368 => x"1b085959",
         10369 => x"5a76782e",
         10370 => x"b738800b",
         10371 => x"831a3371",
         10372 => x"5e565d74",
         10373 => x"7d2e0981",
         10374 => x"0682d438",
         10375 => x"81547753",
         10376 => x"b8195281",
         10377 => x"193351f0",
         10378 => x"833f84ba",
         10379 => x"8c08802e",
         10380 => x"8538ff58",
         10381 => x"815c77b4",
         10382 => x"1a0c7b58",
         10383 => x"7bfdac38",
         10384 => x"7983ff06",
         10385 => x"19b80581",
         10386 => x"1b778106",
         10387 => x"5f5f577a",
         10388 => x"557c802e",
         10389 => x"8f387a84",
         10390 => x"2b9ff006",
         10391 => x"77338f06",
         10392 => x"7107565a",
         10393 => x"74773481",
         10394 => x"0b831a34",
         10395 => x"7d892aa8",
         10396 => x"1a080556",
         10397 => x"800bb41a",
         10398 => x"08565f74",
         10399 => x"762e83dd",
         10400 => x"38815474",
         10401 => x"53b81970",
         10402 => x"53811a33",
         10403 => x"5257f09b",
         10404 => x"3f815884",
         10405 => x"ba8c087f",
         10406 => x"2e098106",
         10407 => x"80c73884",
         10408 => x"ba8c0883",
         10409 => x"1a34b419",
         10410 => x"0870a81b",
         10411 => x"0831a01b",
         10412 => x"0884ba8c",
         10413 => x"085b5c56",
         10414 => x"5c747a27",
         10415 => x"8b388219",
         10416 => x"33557482",
         10417 => x"2e82e438",
         10418 => x"81547553",
         10419 => x"76528119",
         10420 => x"3351eed8",
         10421 => x"3f84ba8c",
         10422 => x"08802e85",
         10423 => x"38ff5681",
         10424 => x"5875b41a",
         10425 => x"0c77fc83",
         10426 => x"387d83ff",
         10427 => x"0619b805",
         10428 => x"7b842a56",
         10429 => x"567c8f38",
         10430 => x"7a882a76",
         10431 => x"3381f006",
         10432 => x"718f0607",
         10433 => x"565c7476",
         10434 => x"34810b83",
         10435 => x"1a34fccb",
         10436 => x"39815476",
         10437 => x"53b81970",
         10438 => x"53811a33",
         10439 => x"525def8b",
         10440 => x"3f815a84",
         10441 => x"ba8c087c",
         10442 => x"2e098106",
         10443 => x"fc883884",
         10444 => x"ba8c0883",
         10445 => x"1a34b419",
         10446 => x"0870a81b",
         10447 => x"0831a01b",
         10448 => x"0884ba8c",
         10449 => x"085d5940",
         10450 => x"5e7e7727",
         10451 => x"fbca3882",
         10452 => x"19335574",
         10453 => x"822e0981",
         10454 => x"06fbbd38",
         10455 => x"8154761e",
         10456 => x"537c5281",
         10457 => x"193351ee",
         10458 => x"c23f7b5a",
         10459 => x"fbaa3981",
         10460 => x"547653b8",
         10461 => x"19705381",
         10462 => x"1a335257",
         10463 => x"eead3f81",
         10464 => x"5c84ba8c",
         10465 => x"087d2e09",
         10466 => x"8106fdae",
         10467 => x"3884ba8c",
         10468 => x"08831a34",
         10469 => x"b4190870",
         10470 => x"a81b0831",
         10471 => x"a01b0884",
         10472 => x"ba8c085f",
         10473 => x"40565f74",
         10474 => x"7e27fcf0",
         10475 => x"38821933",
         10476 => x"5574822e",
         10477 => x"098106fc",
         10478 => x"e3388154",
         10479 => x"7d1f5376",
         10480 => x"52811933",
         10481 => x"51ede43f",
         10482 => x"7c5cfcd0",
         10483 => x"39815476",
         10484 => x"53b81970",
         10485 => x"53811a33",
         10486 => x"5257edcf",
         10487 => x"3f815a84",
         10488 => x"ba8c087c",
         10489 => x"2e098106",
         10490 => x"fbc53884",
         10491 => x"ba8c0883",
         10492 => x"1a34b419",
         10493 => x"0870a81b",
         10494 => x"0831a01b",
         10495 => x"0884ba8c",
         10496 => x"085d5f40",
         10497 => x"5e7e7d27",
         10498 => x"fb873882",
         10499 => x"19335574",
         10500 => x"822e0981",
         10501 => x"06fafa38",
         10502 => x"81547c1e",
         10503 => x"53765281",
         10504 => x"193351ed",
         10505 => x"863f7b5a",
         10506 => x"fae73981",
         10507 => x"54791c53",
         10508 => x"76528119",
         10509 => x"3351ecf3",
         10510 => x"3f7e58fd",
         10511 => x"8b397b76",
         10512 => x"1083fe06",
         10513 => x"7a057c83",
         10514 => x"ffff0659",
         10515 => x"5f5876b8",
         10516 => x"1f347688",
         10517 => x"2a5a79b9",
         10518 => x"1f34f9fa",
         10519 => x"397e58fd",
         10520 => x"88397b76",
         10521 => x"822b83fc",
         10522 => x"067a05b8",
         10523 => x"11831133",
         10524 => x"70982b8f",
         10525 => x"0a067ff0",
         10526 => x"0a060742",
         10527 => x"585f5d58",
         10528 => x"7d7d347d",
         10529 => x"882a5675",
         10530 => x"b91d347d",
         10531 => x"902a5a79",
         10532 => x"ba1d347d",
         10533 => x"982a5b7a",
         10534 => x"bb1d34fa",
         10535 => x"cf39f63d",
         10536 => x"0d7c7e71",
         10537 => x"085b5c5a",
         10538 => x"7a818a38",
         10539 => x"90190857",
         10540 => x"76802e80",
         10541 => x"f438769c",
         10542 => x"1a082780",
         10543 => x"ec389419",
         10544 => x"08705654",
         10545 => x"73802e80",
         10546 => x"d738767b",
         10547 => x"2e819338",
         10548 => x"76568116",
         10549 => x"569c1908",
         10550 => x"76268938",
         10551 => x"82567577",
         10552 => x"2682b238",
         10553 => x"75527951",
         10554 => x"f0f53f84",
         10555 => x"ba8c0880",
         10556 => x"2e81d038",
         10557 => x"805884ba",
         10558 => x"8c08812e",
         10559 => x"b13884ba",
         10560 => x"8c080970",
         10561 => x"30707207",
         10562 => x"8025707b",
         10563 => x"07515155",
         10564 => x"557382aa",
         10565 => x"3875772e",
         10566 => x"098106ff",
         10567 => x"b5387355",
         10568 => x"7484ba8c",
         10569 => x"0c8c3d0d",
         10570 => x"048157ff",
         10571 => x"913984ba",
         10572 => x"8c0858ca",
         10573 => x"397a5279",
         10574 => x"51f0a43f",
         10575 => x"81557484",
         10576 => x"ba8c0827",
         10577 => x"db3884ba",
         10578 => x"8c085584",
         10579 => x"ba8c08ff",
         10580 => x"2ece389c",
         10581 => x"190884ba",
         10582 => x"8c0826c4",
         10583 => x"387a57fe",
         10584 => x"dd39811b",
         10585 => x"569c1908",
         10586 => x"76268338",
         10587 => x"82567552",
         10588 => x"7951efeb",
         10589 => x"3f805884",
         10590 => x"ba8c0881",
         10591 => x"2e81a038",
         10592 => x"84ba8c08",
         10593 => x"09703070",
         10594 => x"72078025",
         10595 => x"707b0784",
         10596 => x"ba8c0854",
         10597 => x"51515555",
         10598 => x"73ff8538",
         10599 => x"84ba8c08",
         10600 => x"802e9a38",
         10601 => x"90190854",
         10602 => x"817427fe",
         10603 => x"a338739c",
         10604 => x"1a0827fe",
         10605 => x"9b387370",
         10606 => x"5757fe96",
         10607 => x"3975802e",
         10608 => x"fe8e38ff",
         10609 => x"53755278",
         10610 => x"51f5f53f",
         10611 => x"84ba8c08",
         10612 => x"84ba8c08",
         10613 => x"307084ba",
         10614 => x"8c080780",
         10615 => x"25565855",
         10616 => x"7a80c438",
         10617 => x"7480e338",
         10618 => x"75901a0c",
         10619 => x"9c1908fe",
         10620 => x"05941a08",
         10621 => x"56587478",
         10622 => x"268638ff",
         10623 => x"15941a0c",
         10624 => x"84193381",
         10625 => x"075a7984",
         10626 => x"1a347555",
         10627 => x"7484ba8c",
         10628 => x"0c8c3d0d",
         10629 => x"04800b84",
         10630 => x"ba8c0c8c",
         10631 => x"3d0d0484",
         10632 => x"ba8c0858",
         10633 => x"feda3973",
         10634 => x"802effb8",
         10635 => x"3875537a",
         10636 => x"527851f5",
         10637 => x"8b3f84ba",
         10638 => x"8c0855ff",
         10639 => x"a73984ba",
         10640 => x"8c0884ba",
         10641 => x"8c0c8c3d",
         10642 => x"0d04ff56",
         10643 => x"74812eff",
         10644 => x"b9388155",
         10645 => x"ffb639f8",
         10646 => x"3d0d7a7c",
         10647 => x"71085955",
         10648 => x"5873f080",
         10649 => x"0a2680df",
         10650 => x"38739f06",
         10651 => x"537280d7",
         10652 => x"38739019",
         10653 => x"0c881808",
         10654 => x"557480df",
         10655 => x"38763356",
         10656 => x"75822680",
         10657 => x"cc387385",
         10658 => x"2a53820b",
         10659 => x"8818225a",
         10660 => x"56727927",
         10661 => x"a938ac17",
         10662 => x"0898190c",
         10663 => x"7494190c",
         10664 => x"98180853",
         10665 => x"82567280",
         10666 => x"2e943873",
         10667 => x"892a1398",
         10668 => x"190c7383",
         10669 => x"ff0617b8",
         10670 => x"059c190c",
         10671 => x"80567584",
         10672 => x"ba8c0c8a",
         10673 => x"3d0d0482",
         10674 => x"0b84ba8c",
         10675 => x"0c8a3d0d",
         10676 => x"04ac1708",
         10677 => x"5574802e",
         10678 => x"ffac388a",
         10679 => x"17227089",
         10680 => x"2b575973",
         10681 => x"7627a538",
         10682 => x"9c170853",
         10683 => x"fe15fe14",
         10684 => x"54568059",
         10685 => x"7573278d",
         10686 => x"388a1722",
         10687 => x"767129b0",
         10688 => x"1908055a",
         10689 => x"53789819",
         10690 => x"0cff9139",
         10691 => x"74527751",
         10692 => x"eccd3f84",
         10693 => x"ba8c0855",
         10694 => x"84ba8c08",
         10695 => x"ff2ea438",
         10696 => x"810b84ba",
         10697 => x"8c0827ff",
         10698 => x"9e389c17",
         10699 => x"085384ba",
         10700 => x"8c087327",
         10701 => x"ff913873",
         10702 => x"76315473",
         10703 => x"7627cd38",
         10704 => x"ffaa3981",
         10705 => x"0b84ba8c",
         10706 => x"0c8a3d0d",
         10707 => x"04f33d0d",
         10708 => x"7f700890",
         10709 => x"1208a005",
         10710 => x"5c5a57f0",
         10711 => x"800a7a27",
         10712 => x"8638800b",
         10713 => x"98180c98",
         10714 => x"17085584",
         10715 => x"5674802e",
         10716 => x"b2387983",
         10717 => x"ff065b7a",
         10718 => x"9d388115",
         10719 => x"94180857",
         10720 => x"5875a938",
         10721 => x"79852a88",
         10722 => x"1a225755",
         10723 => x"74762781",
         10724 => x"f5387798",
         10725 => x"180c7990",
         10726 => x"180c781b",
         10727 => x"b8059c18",
         10728 => x"0c805675",
         10729 => x"84ba8c0c",
         10730 => x"8f3d0d04",
         10731 => x"7798180c",
         10732 => x"8a1922ff",
         10733 => x"057a892a",
         10734 => x"065c7bda",
         10735 => x"38755276",
         10736 => x"51eb9c3f",
         10737 => x"84ba8c08",
         10738 => x"5d825681",
         10739 => x"0b84ba8c",
         10740 => x"0827d038",
         10741 => x"815684ba",
         10742 => x"8c08ff2e",
         10743 => x"c6389c19",
         10744 => x"0884ba8c",
         10745 => x"08268291",
         10746 => x"3860802e",
         10747 => x"81983894",
         10748 => x"17085276",
         10749 => x"51f9a73f",
         10750 => x"84ba8c08",
         10751 => x"5d875684",
         10752 => x"ba8c0880",
         10753 => x"2eff9c38",
         10754 => x"825684ba",
         10755 => x"8c08812e",
         10756 => x"ff913881",
         10757 => x"5684ba8c",
         10758 => x"08ff2eff",
         10759 => x"863884ba",
         10760 => x"8c08831a",
         10761 => x"335f587d",
         10762 => x"80ea38fe",
         10763 => x"189c1a08",
         10764 => x"fe055956",
         10765 => x"805c7578",
         10766 => x"278d388a",
         10767 => x"19227671",
         10768 => x"29b01b08",
         10769 => x"055d5e7b",
         10770 => x"b41a0cb8",
         10771 => x"19588480",
         10772 => x"78575580",
         10773 => x"76708105",
         10774 => x"5834ff15",
         10775 => x"5574f438",
         10776 => x"74568a19",
         10777 => x"22557575",
         10778 => x"27818038",
         10779 => x"8154751c",
         10780 => x"53775281",
         10781 => x"193351e4",
         10782 => x"b23f84ba",
         10783 => x"8c0880e7",
         10784 => x"38811656",
         10785 => x"dd397a98",
         10786 => x"180c840b",
         10787 => x"84ba8c0c",
         10788 => x"8f3d0d04",
         10789 => x"7554b419",
         10790 => x"0853b819",
         10791 => x"7053811a",
         10792 => x"335256e4",
         10793 => x"863f84ba",
         10794 => x"8c0880f3",
         10795 => x"3884ba8c",
         10796 => x"08831a34",
         10797 => x"b41908a8",
         10798 => x"1a083155",
         10799 => x"74a01a08",
         10800 => x"27fee838",
         10801 => x"8219335c",
         10802 => x"7b822e09",
         10803 => x"8106fedb",
         10804 => x"388154b4",
         10805 => x"1908a01a",
         10806 => x"08055375",
         10807 => x"52811933",
         10808 => x"51e3c83f",
         10809 => x"fec5398a",
         10810 => x"19225574",
         10811 => x"83ffff06",
         10812 => x"5574762e",
         10813 => x"098106a7",
         10814 => x"387c9418",
         10815 => x"0cfe1d9c",
         10816 => x"1a08fe05",
         10817 => x"5e568058",
         10818 => x"757d27fd",
         10819 => x"85388a19",
         10820 => x"22767129",
         10821 => x"b01b0805",
         10822 => x"98190c5c",
         10823 => x"fcf83981",
         10824 => x"0b84ba8c",
         10825 => x"0c8f3d0d",
         10826 => x"04ee3d0d",
         10827 => x"6466415c",
         10828 => x"847c085a",
         10829 => x"5b81ff70",
         10830 => x"981e0858",
         10831 => x"5e5e7580",
         10832 => x"2e82d238",
         10833 => x"b8195f75",
         10834 => x"5a8058b4",
         10835 => x"1908762e",
         10836 => x"82d13883",
         10837 => x"19337858",
         10838 => x"5574782e",
         10839 => x"09810681",
         10840 => x"94388154",
         10841 => x"7553b819",
         10842 => x"52811933",
         10843 => x"51e1bd3f",
         10844 => x"84ba8c08",
         10845 => x"802e8538",
         10846 => x"ff5a8157",
         10847 => x"79b41a0c",
         10848 => x"765b7682",
         10849 => x"90389c1c",
         10850 => x"08703358",
         10851 => x"5876802e",
         10852 => x"8281388b",
         10853 => x"1833bf06",
         10854 => x"7081ff06",
         10855 => x"5b416086",
         10856 => x"1d347681",
         10857 => x"e5327030",
         10858 => x"78ae3270",
         10859 => x"30728025",
         10860 => x"71802507",
         10861 => x"54454557",
         10862 => x"55749338",
         10863 => x"747adf06",
         10864 => x"43566188",
         10865 => x"2e81bf38",
         10866 => x"75602e81",
         10867 => x"863881ff",
         10868 => x"5d80527b",
         10869 => x"51faf63f",
         10870 => x"84ba8c08",
         10871 => x"5b84ba8c",
         10872 => x"0881b238",
         10873 => x"981c0856",
         10874 => x"75fedc38",
         10875 => x"7a84ba8c",
         10876 => x"0c943d0d",
         10877 => x"048154b4",
         10878 => x"1908537e",
         10879 => x"52811933",
         10880 => x"51e1a83f",
         10881 => x"815784ba",
         10882 => x"8c08782e",
         10883 => x"098106fe",
         10884 => x"ef3884ba",
         10885 => x"8c08831a",
         10886 => x"34b41908",
         10887 => x"a81a0831",
         10888 => x"84ba8c08",
         10889 => x"585b7aa0",
         10890 => x"1a0827fe",
         10891 => x"b5388219",
         10892 => x"33416082",
         10893 => x"2e098106",
         10894 => x"fea83881",
         10895 => x"54b41908",
         10896 => x"a01a0805",
         10897 => x"537e5281",
         10898 => x"193351e0",
         10899 => x"de3f7757",
         10900 => x"fe903979",
         10901 => x"8f2e0981",
         10902 => x"0681e738",
         10903 => x"76862a81",
         10904 => x"065b7a80",
         10905 => x"2e93388d",
         10906 => x"18337781",
         10907 => x"bf067090",
         10908 => x"1f087fac",
         10909 => x"050c595e",
         10910 => x"5e767d2e",
         10911 => x"ab3881ff",
         10912 => x"55745dfe",
         10913 => x"cc398156",
         10914 => x"75602e09",
         10915 => x"8106febe",
         10916 => x"38c13984",
         10917 => x"5b800b98",
         10918 => x"1d0c7a84",
         10919 => x"ba8c0c94",
         10920 => x"3d0d0477",
         10921 => x"5bfddf39",
         10922 => x"8d183357",
         10923 => x"7d772e09",
         10924 => x"8106cb38",
         10925 => x"8c19089b",
         10926 => x"19339a1a",
         10927 => x"3371882b",
         10928 => x"07585641",
         10929 => x"75ffb738",
         10930 => x"77337081",
         10931 => x"bf068d29",
         10932 => x"f305515a",
         10933 => x"8176585b",
         10934 => x"83e68c17",
         10935 => x"33780581",
         10936 => x"11337133",
         10937 => x"71882b07",
         10938 => x"5244567a",
         10939 => x"802e80c5",
         10940 => x"387981fe",
         10941 => x"26ff8738",
         10942 => x"79106105",
         10943 => x"765c4275",
         10944 => x"6223811a",
         10945 => x"5a811757",
         10946 => x"8c7727cc",
         10947 => x"38773370",
         10948 => x"862a8106",
         10949 => x"59577780",
         10950 => x"2e903879",
         10951 => x"81fe26fe",
         10952 => x"dd387910",
         10953 => x"61054380",
         10954 => x"6323ff1d",
         10955 => x"7081ff06",
         10956 => x"5e41fd9d",
         10957 => x"397583ff",
         10958 => x"ff2eca38",
         10959 => x"81ff55fe",
         10960 => x"c0397ca8",
         10961 => x"387c558b",
         10962 => x"5774812a",
         10963 => x"75818029",
         10964 => x"05787081",
         10965 => x"055a3340",
         10966 => x"7f057081",
         10967 => x"ff06ff19",
         10968 => x"59565976",
         10969 => x"e438747e",
         10970 => x"2efd8138",
         10971 => x"ff0bac1d",
         10972 => x"0c7a84ba",
         10973 => x"8c0c943d",
         10974 => x"0d04ef3d",
         10975 => x"0d637008",
         10976 => x"5c5c8052",
         10977 => x"7b51f5cf",
         10978 => x"3f84ba8c",
         10979 => x"085a84ba",
         10980 => x"8c088280",
         10981 => x"3881ff70",
         10982 => x"405dff0b",
         10983 => x"ac1d0cb8",
         10984 => x"1b5e981c",
         10985 => x"08568058",
         10986 => x"b41b0876",
         10987 => x"2e82cc38",
         10988 => x"831b3378",
         10989 => x"58557478",
         10990 => x"2e098106",
         10991 => x"81df3881",
         10992 => x"547553b8",
         10993 => x"1b52811b",
         10994 => x"3351dce0",
         10995 => x"3f84ba8c",
         10996 => x"08802e85",
         10997 => x"38ff5681",
         10998 => x"5775b41c",
         10999 => x"0c765a76",
         11000 => x"81b2389c",
         11001 => x"1c087033",
         11002 => x"58597680",
         11003 => x"2e849938",
         11004 => x"8b1933bf",
         11005 => x"067081ff",
         11006 => x"06575877",
         11007 => x"861d3476",
         11008 => x"81e52e80",
         11009 => x"f2387583",
         11010 => x"2a810655",
         11011 => x"758f2e81",
         11012 => x"ef387480",
         11013 => x"e238758f",
         11014 => x"2e81e538",
         11015 => x"7caa3878",
         11016 => x"7d56588b",
         11017 => x"5774812a",
         11018 => x"75818029",
         11019 => x"05787081",
         11020 => x"055a3357",
         11021 => x"76057081",
         11022 => x"ff06ff19",
         11023 => x"59565d76",
         11024 => x"e438747f",
         11025 => x"2e80cd38",
         11026 => x"ab1c3381",
         11027 => x"065776a7",
         11028 => x"388b0ba0",
         11029 => x"1d595778",
         11030 => x"7081055a",
         11031 => x"33787081",
         11032 => x"055a3371",
         11033 => x"7131ff1a",
         11034 => x"5a584240",
         11035 => x"76802e81",
         11036 => x"dc387580",
         11037 => x"2ee13881",
         11038 => x"ff5dff0b",
         11039 => x"ac1d0c80",
         11040 => x"527b51f5",
         11041 => x"c83f84ba",
         11042 => x"8c085a84",
         11043 => x"ba8c0880",
         11044 => x"2efe8f38",
         11045 => x"7984ba8c",
         11046 => x"0c933d0d",
         11047 => x"048154b4",
         11048 => x"1b08537d",
         11049 => x"52811b33",
         11050 => x"51dc803f",
         11051 => x"815784ba",
         11052 => x"8c08782e",
         11053 => x"098106fe",
         11054 => x"a43884ba",
         11055 => x"8c08831c",
         11056 => x"34b41b08",
         11057 => x"a81c0831",
         11058 => x"84ba8c08",
         11059 => x"585978a0",
         11060 => x"1c0827fd",
         11061 => x"ea38821b",
         11062 => x"335a7982",
         11063 => x"2e098106",
         11064 => x"fddd3881",
         11065 => x"54b41b08",
         11066 => x"a01c0805",
         11067 => x"537d5281",
         11068 => x"1b3351db",
         11069 => x"b63f7757",
         11070 => x"fdc53977",
         11071 => x"5afde439",
         11072 => x"ab1c3370",
         11073 => x"862a8106",
         11074 => x"425560fe",
         11075 => x"f2387686",
         11076 => x"2a81065a",
         11077 => x"79802e93",
         11078 => x"388d1933",
         11079 => x"7781bf06",
         11080 => x"70901f08",
         11081 => x"7fac050c",
         11082 => x"595e5f76",
         11083 => x"7d2eaf38",
         11084 => x"81ff5574",
         11085 => x"5d80527b",
         11086 => x"51f4923f",
         11087 => x"84ba8c08",
         11088 => x"5a84ba8c",
         11089 => x"08802efc",
         11090 => x"d938fec8",
         11091 => x"3975802e",
         11092 => x"fec23881",
         11093 => x"ff5dff0b",
         11094 => x"ac1d0cfe",
         11095 => x"a2398d19",
         11096 => x"33577e77",
         11097 => x"2e098106",
         11098 => x"c7388c1b",
         11099 => x"089b1a33",
         11100 => x"9a1b3371",
         11101 => x"882b0759",
         11102 => x"424076ff",
         11103 => x"b3387833",
         11104 => x"70bf068d",
         11105 => x"29f3055b",
         11106 => x"55817759",
         11107 => x"5683e68c",
         11108 => x"18337905",
         11109 => x"81113371",
         11110 => x"3371882b",
         11111 => x"07524257",
         11112 => x"75802e80",
         11113 => x"ed387981",
         11114 => x"fe26ff84",
         11115 => x"38765181",
         11116 => x"a18a3f84",
         11117 => x"ba8c087a",
         11118 => x"10610570",
         11119 => x"22534381",
         11120 => x"1b5b5681",
         11121 => x"a0f63f75",
         11122 => x"84ba8c08",
         11123 => x"2e098106",
         11124 => x"fede3876",
         11125 => x"56811858",
         11126 => x"8c7827ff",
         11127 => x"b0387833",
         11128 => x"70862a81",
         11129 => x"06565975",
         11130 => x"802e9238",
         11131 => x"74802e8d",
         11132 => x"38791060",
         11133 => x"05702241",
         11134 => x"417ffeb4",
         11135 => x"38ff1d70",
         11136 => x"81ff065e",
         11137 => x"5afeae39",
         11138 => x"840b84ba",
         11139 => x"8c0c933d",
         11140 => x"0d047683",
         11141 => x"ffff2eff",
         11142 => x"bc3881ff",
         11143 => x"55fe9439",
         11144 => x"ea3d0d68",
         11145 => x"700870ab",
         11146 => x"133381a0",
         11147 => x"06585a5d",
         11148 => x"5e865674",
         11149 => x"85b53874",
         11150 => x"8c1d0870",
         11151 => x"2257575d",
         11152 => x"74802e8e",
         11153 => x"38811d70",
         11154 => x"10177022",
         11155 => x"51565d74",
         11156 => x"f438953d",
         11157 => x"a01f5b40",
         11158 => x"8c607b58",
         11159 => x"58557570",
         11160 => x"81055733",
         11161 => x"77708105",
         11162 => x"5934ff15",
         11163 => x"5574ef38",
         11164 => x"0280db05",
         11165 => x"33708106",
         11166 => x"58567680",
         11167 => x"2e82aa38",
         11168 => x"80c00bab",
         11169 => x"1f34810b",
         11170 => x"943d405b",
         11171 => x"8c1c087b",
         11172 => x"58598b7a",
         11173 => x"615a5755",
         11174 => x"77708105",
         11175 => x"59337670",
         11176 => x"81055834",
         11177 => x"ff155574",
         11178 => x"ef38857b",
         11179 => x"2780c238",
         11180 => x"7a792256",
         11181 => x"5774802e",
         11182 => x"b8387482",
         11183 => x"1a5a568f",
         11184 => x"58758106",
         11185 => x"77100776",
         11186 => x"812a7083",
         11187 => x"ffff0672",
         11188 => x"902a8106",
         11189 => x"44585657",
         11190 => x"60802e87",
         11191 => x"387684a0",
         11192 => x"a13257ff",
         11193 => x"18587780",
         11194 => x"25d73878",
         11195 => x"225574ca",
         11196 => x"38870284",
         11197 => x"0580cf05",
         11198 => x"575876b0",
         11199 => x"07bf0655",
         11200 => x"b9752784",
         11201 => x"38871555",
         11202 => x"747634ff",
         11203 => x"16ff1978",
         11204 => x"842a5959",
         11205 => x"5676e338",
         11206 => x"771f5980",
         11207 => x"fe793476",
         11208 => x"7a585680",
         11209 => x"7827a038",
         11210 => x"79335574",
         11211 => x"a02e9838",
         11212 => x"81165675",
         11213 => x"782788a2",
         11214 => x"38751a70",
         11215 => x"33565774",
         11216 => x"a02e0981",
         11217 => x"06ea3881",
         11218 => x"1656a055",
         11219 => x"7787268e",
         11220 => x"38983d78",
         11221 => x"05ec0581",
         11222 => x"19713357",
         11223 => x"59417477",
         11224 => x"34877627",
         11225 => x"87f4387d",
         11226 => x"51f88f3f",
         11227 => x"84ba8c08",
         11228 => x"8b38811b",
         11229 => x"5b80e37b",
         11230 => x"27fe9138",
         11231 => x"87567a80",
         11232 => x"e42e82e7",
         11233 => x"3884ba8c",
         11234 => x"085684ba",
         11235 => x"8c08842e",
         11236 => x"09810682",
         11237 => x"d6380280",
         11238 => x"db0533ab",
         11239 => x"1f347d08",
         11240 => x"02840580",
         11241 => x"db053357",
         11242 => x"5875812a",
         11243 => x"81065f81",
         11244 => x"5b7e802e",
         11245 => x"90388d52",
         11246 => x"8c1d51fe",
         11247 => x"89e73f84",
         11248 => x"ba8c081b",
         11249 => x"5b80527d",
         11250 => x"51ed8c3f",
         11251 => x"84ba8c08",
         11252 => x"5684ba8c",
         11253 => x"08818238",
         11254 => x"84ba8c08",
         11255 => x"b8195e59",
         11256 => x"981e0856",
         11257 => x"8057b418",
         11258 => x"08762e85",
         11259 => x"f3388318",
         11260 => x"33407f77",
         11261 => x"2e098106",
         11262 => x"82a33881",
         11263 => x"547553b8",
         11264 => x"18528118",
         11265 => x"3351d4a4",
         11266 => x"3f84ba8c",
         11267 => x"08802e85",
         11268 => x"38ff5681",
         11269 => x"5775b419",
         11270 => x"0c765676",
         11271 => x"bc389c1e",
         11272 => x"08703356",
         11273 => x"427481e5",
         11274 => x"2e81c938",
         11275 => x"74307080",
         11276 => x"25780756",
         11277 => x"5f74802e",
         11278 => x"81c93881",
         11279 => x"1959787b",
         11280 => x"2e868938",
         11281 => x"81527d51",
         11282 => x"ee833f84",
         11283 => x"ba8c0856",
         11284 => x"84ba8c08",
         11285 => x"802eff88",
         11286 => x"38875875",
         11287 => x"842e8189",
         11288 => x"38755875",
         11289 => x"818338ff",
         11290 => x"1b407f81",
         11291 => x"f338981e",
         11292 => x"0857b41c",
         11293 => x"08772eaf",
         11294 => x"38831c33",
         11295 => x"7857407f",
         11296 => x"84823881",
         11297 => x"547653b8",
         11298 => x"1c52811c",
         11299 => x"3351d39c",
         11300 => x"3f84ba8c",
         11301 => x"08802e85",
         11302 => x"38ff5781",
         11303 => x"5676b41d",
         11304 => x"0c755875",
         11305 => x"80c338a0",
         11306 => x"0b9c1f08",
         11307 => x"57558076",
         11308 => x"70810558",
         11309 => x"34ff1555",
         11310 => x"74f4388b",
         11311 => x"0b9c1f08",
         11312 => x"7b585855",
         11313 => x"75708105",
         11314 => x"57337770",
         11315 => x"81055934",
         11316 => x"ff155574",
         11317 => x"ef389c1e",
         11318 => x"08ab1f33",
         11319 => x"98065e5a",
         11320 => x"7c8c1b34",
         11321 => x"810b831d",
         11322 => x"34775675",
         11323 => x"84ba8c0c",
         11324 => x"983d0d04",
         11325 => x"81753070",
         11326 => x"80257207",
         11327 => x"57405774",
         11328 => x"feb93874",
         11329 => x"5981527d",
         11330 => x"51ecc23f",
         11331 => x"84ba8c08",
         11332 => x"5684ba8c",
         11333 => x"08802efd",
         11334 => x"c738febd",
         11335 => x"398154b4",
         11336 => x"1808537c",
         11337 => x"52811833",
         11338 => x"51d3803f",
         11339 => x"84ba8c08",
         11340 => x"772e0981",
         11341 => x"0683bf38",
         11342 => x"84ba8c08",
         11343 => x"831934b4",
         11344 => x"1808a819",
         11345 => x"08315574",
         11346 => x"a0190827",
         11347 => x"8b388218",
         11348 => x"33416082",
         11349 => x"2e84ac38",
         11350 => x"84ba8c08",
         11351 => x"57fd9c39",
         11352 => x"7f852b90",
         11353 => x"1f087131",
         11354 => x"53587d51",
         11355 => x"e9e93f84",
         11356 => x"ba8c0858",
         11357 => x"84ba8c08",
         11358 => x"feef3879",
         11359 => x"84ba8c08",
         11360 => x"56588b57",
         11361 => x"74812a75",
         11362 => x"81802905",
         11363 => x"78708105",
         11364 => x"5a335776",
         11365 => x"057081ff",
         11366 => x"06ff1959",
         11367 => x"565d76e4",
         11368 => x"387481ff",
         11369 => x"06b81d43",
         11370 => x"41981e08",
         11371 => x"578056b4",
         11372 => x"1c08772e",
         11373 => x"b238831c",
         11374 => x"335b7a76",
         11375 => x"2e098106",
         11376 => x"82c93881",
         11377 => x"547653b8",
         11378 => x"1c52811c",
         11379 => x"3351d0dc",
         11380 => x"3f84ba8c",
         11381 => x"08802e85",
         11382 => x"38ff5781",
         11383 => x"5676b41d",
         11384 => x"0c755875",
         11385 => x"fe83388c",
         11386 => x"1c089c1f",
         11387 => x"086181ff",
         11388 => x"065f5c5f",
         11389 => x"608d1c34",
         11390 => x"8f0b8b1c",
         11391 => x"34758c1c",
         11392 => x"34759a1c",
         11393 => x"34759b1c",
         11394 => x"347c8d29",
         11395 => x"f3057677",
         11396 => x"5a585976",
         11397 => x"83ffff2e",
         11398 => x"8b387810",
         11399 => x"1f702281",
         11400 => x"1b5b5856",
         11401 => x"83e68c18",
         11402 => x"337b0555",
         11403 => x"76757081",
         11404 => x"05573476",
         11405 => x"882a5675",
         11406 => x"75347685",
         11407 => x"3883ffff",
         11408 => x"57811858",
         11409 => x"8c7827cb",
         11410 => x"387683ff",
         11411 => x"ff2e81b3",
         11412 => x"3878101f",
         11413 => x"70225858",
         11414 => x"76802e81",
         11415 => x"a6387c7b",
         11416 => x"34810b83",
         11417 => x"1d348052",
         11418 => x"7d51e9e1",
         11419 => x"3f84ba8c",
         11420 => x"085884ba",
         11421 => x"8c08fcf1",
         11422 => x"387fff05",
         11423 => x"407ffea9",
         11424 => x"38fbeb39",
         11425 => x"8154b41c",
         11426 => x"0853b81c",
         11427 => x"7053811d",
         11428 => x"335259d0",
         11429 => x"963f8156",
         11430 => x"84ba8c08",
         11431 => x"fc833884",
         11432 => x"ba8c0883",
         11433 => x"1d34b41c",
         11434 => x"08a81d08",
         11435 => x"3184ba8c",
         11436 => x"08574160",
         11437 => x"a01d0827",
         11438 => x"fbc93882",
         11439 => x"1c334261",
         11440 => x"822e0981",
         11441 => x"06fbbc38",
         11442 => x"8154b41c",
         11443 => x"08a01d08",
         11444 => x"05537852",
         11445 => x"811c3351",
         11446 => x"cfd13f77",
         11447 => x"56fba439",
         11448 => x"769c1f08",
         11449 => x"70335743",
         11450 => x"567481e5",
         11451 => x"2e098106",
         11452 => x"faba38fb",
         11453 => x"ff398170",
         11454 => x"57577680",
         11455 => x"2efa9f38",
         11456 => x"fad7397c",
         11457 => x"80c0075d",
         11458 => x"fed43981",
         11459 => x"54b41c08",
         11460 => x"53615281",
         11461 => x"1c3351cf",
         11462 => x"923f84ba",
         11463 => x"8c08762e",
         11464 => x"098106bc",
         11465 => x"3884ba8c",
         11466 => x"08831d34",
         11467 => x"b41c08a8",
         11468 => x"1d083155",
         11469 => x"74a01d08",
         11470 => x"278a3882",
         11471 => x"1c335f7e",
         11472 => x"822eaa38",
         11473 => x"84ba8c08",
         11474 => x"56fcf839",
         11475 => x"75ff1c41",
         11476 => x"587f802e",
         11477 => x"fa9838fc",
         11478 => x"8739751a",
         11479 => x"57f7e839",
         11480 => x"81705956",
         11481 => x"75802efc",
         11482 => x"fe38fafd",
         11483 => x"398154b4",
         11484 => x"1c08a01d",
         11485 => x"08055361",
         11486 => x"52811c33",
         11487 => x"51ceac3f",
         11488 => x"fcc13981",
         11489 => x"54b41808",
         11490 => x"a0190805",
         11491 => x"537c5281",
         11492 => x"183351ce",
         11493 => x"963ff8e3",
         11494 => x"39f33d0d",
         11495 => x"7f617108",
         11496 => x"405e5c80",
         11497 => x"0b961e34",
         11498 => x"981c0880",
         11499 => x"2e82b538",
         11500 => x"ac1c08ff",
         11501 => x"2e80d938",
         11502 => x"80707160",
         11503 => x"8c050870",
         11504 => x"2257585b",
         11505 => x"5c587278",
         11506 => x"2ebc3877",
         11507 => x"54741470",
         11508 => x"22811b5b",
         11509 => x"55567a82",
         11510 => x"953880d0",
         11511 => x"80147083",
         11512 => x"ffff0658",
         11513 => x"5a768fff",
         11514 => x"26828338",
         11515 => x"73791a76",
         11516 => x"1170225d",
         11517 => x"58555b79",
         11518 => x"d4387a30",
         11519 => x"70802570",
         11520 => x"307a065a",
         11521 => x"5c5e7c18",
         11522 => x"94055780",
         11523 => x"0b821834",
         11524 => x"8070891f",
         11525 => x"5957589c",
         11526 => x"1c081670",
         11527 => x"33811858",
         11528 => x"565374a0",
         11529 => x"2eb23874",
         11530 => x"852e81bc",
         11531 => x"38758932",
         11532 => x"70307072",
         11533 => x"07802555",
         11534 => x"5b54778b",
         11535 => x"26903872",
         11536 => x"802e8b38",
         11537 => x"ae777081",
         11538 => x"05593481",
         11539 => x"18587477",
         11540 => x"70810559",
         11541 => x"34811858",
         11542 => x"8a7627ff",
         11543 => x"ba387c18",
         11544 => x"88055580",
         11545 => x"0b811634",
         11546 => x"961d3353",
         11547 => x"72a53877",
         11548 => x"81f338bf",
         11549 => x"0b961e34",
         11550 => x"81577c17",
         11551 => x"94055680",
         11552 => x"0b821734",
         11553 => x"9c1c088c",
         11554 => x"11335553",
         11555 => x"73893873",
         11556 => x"891e349c",
         11557 => x"1c08538b",
         11558 => x"1333881e",
         11559 => x"349c1c08",
         11560 => x"9c118311",
         11561 => x"33821233",
         11562 => x"71902b71",
         11563 => x"882b0781",
         11564 => x"14337072",
         11565 => x"07882b75",
         11566 => x"33710764",
         11567 => x"0c599716",
         11568 => x"33961733",
         11569 => x"71882b07",
         11570 => x"5f415b40",
         11571 => x"5a565b55",
         11572 => x"77861e23",
         11573 => x"99153398",
         11574 => x"16337188",
         11575 => x"2b075d54",
         11576 => x"7b841e23",
         11577 => x"8f3d0d04",
         11578 => x"81e555fe",
         11579 => x"c039771d",
         11580 => x"961181ff",
         11581 => x"7a31585b",
         11582 => x"5783b552",
         11583 => x"7a902b74",
         11584 => x"07518191",
         11585 => x"893f84ba",
         11586 => x"8c0883ff",
         11587 => x"ff065581",
         11588 => x"ff7527ad",
         11589 => x"38817627",
         11590 => x"81b33874",
         11591 => x"882a5473",
         11592 => x"7a347497",
         11593 => x"18348278",
         11594 => x"0558800b",
         11595 => x"8c1f0856",
         11596 => x"5b781975",
         11597 => x"1170225c",
         11598 => x"575479fd",
         11599 => x"9038fdba",
         11600 => x"39743076",
         11601 => x"30707807",
         11602 => x"80257280",
         11603 => x"25075855",
         11604 => x"577580f9",
         11605 => x"38747a34",
         11606 => x"81780558",
         11607 => x"800b8c1f",
         11608 => x"08565bcd",
         11609 => x"39727389",
         11610 => x"1f335a57",
         11611 => x"5777802e",
         11612 => x"fe88387c",
         11613 => x"961e7e57",
         11614 => x"59548914",
         11615 => x"33ffbf11",
         11616 => x"5a547899",
         11617 => x"26a4389c",
         11618 => x"1c088c11",
         11619 => x"33545b88",
         11620 => x"7627b438",
         11621 => x"72842a53",
         11622 => x"7281065e",
         11623 => x"7d802e8a",
         11624 => x"38a01470",
         11625 => x"83ffff06",
         11626 => x"55537378",
         11627 => x"7081055a",
         11628 => x"34811681",
         11629 => x"16811971",
         11630 => x"8913335e",
         11631 => x"57595656",
         11632 => x"79ffb738",
         11633 => x"fdb43972",
         11634 => x"832a53cc",
         11635 => x"39807b30",
         11636 => x"70802570",
         11637 => x"30730653",
         11638 => x"5d5f58fc",
         11639 => x"a939ef3d",
         11640 => x"0d637008",
         11641 => x"7042575c",
         11642 => x"80657033",
         11643 => x"57555374",
         11644 => x"af2e8338",
         11645 => x"81537480",
         11646 => x"dc2e81df",
         11647 => x"3872802e",
         11648 => x"81d93898",
         11649 => x"1608881d",
         11650 => x"0c733396",
         11651 => x"3d943d41",
         11652 => x"42559f75",
         11653 => x"2782a738",
         11654 => x"73428c16",
         11655 => x"08588057",
         11656 => x"61707081",
         11657 => x"05523355",
         11658 => x"537381df",
         11659 => x"38727f0c",
         11660 => x"73ff2e81",
         11661 => x"ec3883ff",
         11662 => x"ff74278b",
         11663 => x"38761018",
         11664 => x"56807623",
         11665 => x"81175773",
         11666 => x"83ffff06",
         11667 => x"70af3270",
         11668 => x"309f7327",
         11669 => x"71802507",
         11670 => x"575b5b55",
         11671 => x"73829038",
         11672 => x"7480dc2e",
         11673 => x"82893874",
         11674 => x"80ff26b2",
         11675 => x"3883e5a8",
         11676 => x"0b83e5a8",
         11677 => x"337081ff",
         11678 => x"06565456",
         11679 => x"73802e81",
         11680 => x"ab387375",
         11681 => x"2e8f3881",
         11682 => x"16703370",
         11683 => x"81ff0656",
         11684 => x"545673ee",
         11685 => x"387281ff",
         11686 => x"065b7a81",
         11687 => x"84387681",
         11688 => x"fe2680fd",
         11689 => x"38761018",
         11690 => x"5d747d23",
         11691 => x"81176270",
         11692 => x"70810552",
         11693 => x"33565457",
         11694 => x"73802efe",
         11695 => x"f03880cb",
         11696 => x"39817380",
         11697 => x"dc327030",
         11698 => x"70802573",
         11699 => x"07515558",
         11700 => x"5572802e",
         11701 => x"a1388114",
         11702 => x"70465480",
         11703 => x"74335455",
         11704 => x"72af2edd",
         11705 => x"387280dc",
         11706 => x"32703070",
         11707 => x"80257707",
         11708 => x"51545772",
         11709 => x"e1387288",
         11710 => x"1d0c7333",
         11711 => x"963d943d",
         11712 => x"41425574",
         11713 => x"9f26fe90",
         11714 => x"38b43983",
         11715 => x"b5527351",
         11716 => x"818de73f",
         11717 => x"84ba8c08",
         11718 => x"83ffff06",
         11719 => x"5473fe8d",
         11720 => x"38865473",
         11721 => x"84ba8c0c",
         11722 => x"933d0d04",
         11723 => x"83e5a833",
         11724 => x"7081ff06",
         11725 => x"5c537a80",
         11726 => x"2efee338",
         11727 => x"e439ff80",
         11728 => x"0bab1d34",
         11729 => x"80527b51",
         11730 => x"de8d3f84",
         11731 => x"ba8c0884",
         11732 => x"ba8c0c93",
         11733 => x"3d0d0481",
         11734 => x"7380dc32",
         11735 => x"70307080",
         11736 => x"25730741",
         11737 => x"555a567d",
         11738 => x"802ea138",
         11739 => x"81144280",
         11740 => x"62703355",
         11741 => x"555672af",
         11742 => x"2edd3872",
         11743 => x"80dc3270",
         11744 => x"30708025",
         11745 => x"78074054",
         11746 => x"597de138",
         11747 => x"73610c9f",
         11748 => x"7527822b",
         11749 => x"5a76812e",
         11750 => x"84f83876",
         11751 => x"822e83d1",
         11752 => x"38761759",
         11753 => x"76802ea7",
         11754 => x"38761778",
         11755 => x"11fe0570",
         11756 => x"2270a032",
         11757 => x"7030709f",
         11758 => x"2a524256",
         11759 => x"5f56597c",
         11760 => x"ae2e8438",
         11761 => x"728938ff",
         11762 => x"175776dd",
         11763 => x"38765977",
         11764 => x"19568076",
         11765 => x"2376802e",
         11766 => x"fec73880",
         11767 => x"78227083",
         11768 => x"ffff0672",
         11769 => x"585d5556",
         11770 => x"7aa02e82",
         11771 => x"e6387383",
         11772 => x"ffff0653",
         11773 => x"72ae2e82",
         11774 => x"f1387680",
         11775 => x"2eaa3877",
         11776 => x"19fe0570",
         11777 => x"225a5478",
         11778 => x"ae2e9d38",
         11779 => x"761018fe",
         11780 => x"0554ff17",
         11781 => x"5776802e",
         11782 => x"8f38fe14",
         11783 => x"70225e54",
         11784 => x"7cae2e09",
         11785 => x"8106eb38",
         11786 => x"8b0ba01d",
         11787 => x"5553a074",
         11788 => x"70810556",
         11789 => x"34ff1353",
         11790 => x"72f43872",
         11791 => x"735c5e88",
         11792 => x"78167022",
         11793 => x"81195957",
         11794 => x"545d7480",
         11795 => x"2e80ed38",
         11796 => x"74a02e83",
         11797 => x"d03874ae",
         11798 => x"32703070",
         11799 => x"8025555a",
         11800 => x"5475772e",
         11801 => x"85ce3872",
         11802 => x"83bb3872",
         11803 => x"597c7b26",
         11804 => x"83388159",
         11805 => x"75773270",
         11806 => x"30707207",
         11807 => x"8025707c",
         11808 => x"07515154",
         11809 => x"5472802e",
         11810 => x"83e0387c",
         11811 => x"8b2e8683",
         11812 => x"3875772e",
         11813 => x"8a387983",
         11814 => x"075a7577",
         11815 => x"269e3876",
         11816 => x"56885b8b",
         11817 => x"7e822b81",
         11818 => x"fc067718",
         11819 => x"575f5d77",
         11820 => x"15702281",
         11821 => x"18585653",
         11822 => x"74ff9538",
         11823 => x"a01c3357",
         11824 => x"7681e52e",
         11825 => x"8384387c",
         11826 => x"882e82e3",
         11827 => x"387d8c06",
         11828 => x"58778c2e",
         11829 => x"82ed387d",
         11830 => x"83065574",
         11831 => x"832e82e3",
         11832 => x"3879812a",
         11833 => x"81065675",
         11834 => x"9d387d81",
         11835 => x"065d7c80",
         11836 => x"2e853879",
         11837 => x"90075a7d",
         11838 => x"822a8106",
         11839 => x"5e7d802e",
         11840 => x"85387988",
         11841 => x"075a79ab",
         11842 => x"1d347b51",
         11843 => x"e4ec3f84",
         11844 => x"ba8c08ab",
         11845 => x"1d335654",
         11846 => x"84ba8c08",
         11847 => x"802e81ac",
         11848 => x"3884ba8c",
         11849 => x"08842e09",
         11850 => x"8106fbf7",
         11851 => x"3874852a",
         11852 => x"81065a79",
         11853 => x"802e84f0",
         11854 => x"3874822a",
         11855 => x"81065978",
         11856 => x"8298387b",
         11857 => x"08655556",
         11858 => x"73428c16",
         11859 => x"08588057",
         11860 => x"f9ce3981",
         11861 => x"16701179",
         11862 => x"11702240",
         11863 => x"4056567c",
         11864 => x"a02ef038",
         11865 => x"75802efd",
         11866 => x"85387983",
         11867 => x"075afd8a",
         11868 => x"39821822",
         11869 => x"5675ae2e",
         11870 => x"098106fc",
         11871 => x"ac387722",
         11872 => x"5473ae2e",
         11873 => x"098106fc",
         11874 => x"a0387610",
         11875 => x"185b807b",
         11876 => x"23800ba0",
         11877 => x"1d5653ae",
         11878 => x"54767326",
         11879 => x"8338a054",
         11880 => x"73757081",
         11881 => x"05573481",
         11882 => x"13538a73",
         11883 => x"27e93879",
         11884 => x"a0075877",
         11885 => x"ab1d347b",
         11886 => x"51e3bf3f",
         11887 => x"84ba8c08",
         11888 => x"ab1d3356",
         11889 => x"5484ba8c",
         11890 => x"08fed638",
         11891 => x"74822a81",
         11892 => x"065877fa",
         11893 => x"ce38861c",
         11894 => x"3370842a",
         11895 => x"8106565d",
         11896 => x"74802e83",
         11897 => x"cd38901c",
         11898 => x"0883ff06",
         11899 => x"600580d3",
         11900 => x"113380d2",
         11901 => x"12337188",
         11902 => x"2b076233",
         11903 => x"41575454",
         11904 => x"7d832e82",
         11905 => x"d8387488",
         11906 => x"1d0c7b08",
         11907 => x"655556fe",
         11908 => x"b7397722",
         11909 => x"5574ae2e",
         11910 => x"fef03876",
         11911 => x"175976fb",
         11912 => x"8838fbab",
         11913 => x"39798307",
         11914 => x"7617565a",
         11915 => x"fd81397d",
         11916 => x"822b81fc",
         11917 => x"06708c06",
         11918 => x"595e778c",
         11919 => x"2e098106",
         11920 => x"fd953879",
         11921 => x"82075afd",
         11922 => x"9839850b",
         11923 => x"a01d347c",
         11924 => x"882e0981",
         11925 => x"06fcf638",
         11926 => x"d639ff80",
         11927 => x"0bab1d34",
         11928 => x"800b84ba",
         11929 => x"8c0c933d",
         11930 => x"0d047480",
         11931 => x"ff269d38",
         11932 => x"81ff7527",
         11933 => x"80c938ff",
         11934 => x"1d59787b",
         11935 => x"2681f738",
         11936 => x"7983077d",
         11937 => x"7718575c",
         11938 => x"5afca439",
         11939 => x"7982075a",
         11940 => x"83b55274",
         11941 => x"518185f6",
         11942 => x"3f84ba8c",
         11943 => x"0883ffff",
         11944 => x"0670872a",
         11945 => x"81065a55",
         11946 => x"78802ec4",
         11947 => x"387480ff",
         11948 => x"0683e69c",
         11949 => x"11335654",
         11950 => x"7481ff26",
         11951 => x"ffb93874",
         11952 => x"802e8185",
         11953 => x"3883e5b4",
         11954 => x"0b83e5b4",
         11955 => x"337081ff",
         11956 => x"06565459",
         11957 => x"73802e80",
         11958 => x"e0387375",
         11959 => x"2e8f3881",
         11960 => x"19703370",
         11961 => x"81ff0656",
         11962 => x"545973ee",
         11963 => x"387281ff",
         11964 => x"06597880",
         11965 => x"d438ffbf",
         11966 => x"15547399",
         11967 => x"268a387d",
         11968 => x"82077081",
         11969 => x"ff065f53",
         11970 => x"ff9f1559",
         11971 => x"78992693",
         11972 => x"387d8107",
         11973 => x"7081ff06",
         11974 => x"e0177083",
         11975 => x"ffff0658",
         11976 => x"565f537b",
         11977 => x"1ba00559",
         11978 => x"74793481",
         11979 => x"1b5b7516",
         11980 => x"55fafc39",
         11981 => x"8053fab3",
         11982 => x"3983e5b4",
         11983 => x"337081ff",
         11984 => x"065a5378",
         11985 => x"802effae",
         11986 => x"3880df7a",
         11987 => x"83077d1d",
         11988 => x"a0055b5b",
         11989 => x"55747934",
         11990 => x"811b5bd2",
         11991 => x"3980cd14",
         11992 => x"3380cc15",
         11993 => x"3371982b",
         11994 => x"71902b07",
         11995 => x"7707881f",
         11996 => x"0c5a57fd",
         11997 => x"95397b1b",
         11998 => x"a0057588",
         11999 => x"2a545472",
         12000 => x"7434811b",
         12001 => x"7c11a005",
         12002 => x"5a5b7479",
         12003 => x"34811b5b",
         12004 => x"ff9c3979",
         12005 => x"8307a01d",
         12006 => x"33585a76",
         12007 => x"81e52e09",
         12008 => x"8106faa3",
         12009 => x"38fda339",
         12010 => x"74822a81",
         12011 => x"065c7bf6",
         12012 => x"f238850b",
         12013 => x"84ba8c0c",
         12014 => x"933d0d04",
         12015 => x"eb3d0d67",
         12016 => x"69028805",
         12017 => x"80e70533",
         12018 => x"42425e80",
         12019 => x"610cff7e",
         12020 => x"0870595b",
         12021 => x"4279802e",
         12022 => x"85d73879",
         12023 => x"7081055b",
         12024 => x"33709f26",
         12025 => x"565675ba",
         12026 => x"2e85d038",
         12027 => x"74ed3875",
         12028 => x"ba2e85c7",
         12029 => x"3884d1e8",
         12030 => x"33568076",
         12031 => x"2485b238",
         12032 => x"75101084",
         12033 => x"d1d40570",
         12034 => x"08585a8c",
         12035 => x"5876802e",
         12036 => x"85963876",
         12037 => x"610c7f81",
         12038 => x"fe067733",
         12039 => x"5d597b80",
         12040 => x"2e9b3881",
         12041 => x"173351ff",
         12042 => x"bbb03f84",
         12043 => x"ba8c0881",
         12044 => x"ff067081",
         12045 => x"065e587c",
         12046 => x"802e8696",
         12047 => x"38807734",
         12048 => x"75165d84",
         12049 => x"ba801d33",
         12050 => x"81183481",
         12051 => x"52811733",
         12052 => x"51ffbba4",
         12053 => x"3f84ba8c",
         12054 => x"0881ff06",
         12055 => x"70810641",
         12056 => x"5683587f",
         12057 => x"84c23878",
         12058 => x"802e8d38",
         12059 => x"75822a81",
         12060 => x"06418a58",
         12061 => x"6084b138",
         12062 => x"805b7a83",
         12063 => x"1834ff0b",
         12064 => x"b4180c7a",
         12065 => x"7b5a5581",
         12066 => x"547a53b8",
         12067 => x"17705381",
         12068 => x"18335258",
         12069 => x"ffbb953f",
         12070 => x"84ba8c08",
         12071 => x"7b2e8538",
         12072 => x"ff558159",
         12073 => x"74b4180c",
         12074 => x"84567899",
         12075 => x"3884b717",
         12076 => x"3384b618",
         12077 => x"3371882b",
         12078 => x"07565683",
         12079 => x"567482d4",
         12080 => x"d52e85a5",
         12081 => x"38758126",
         12082 => x"8b3884ba",
         12083 => x"811d3342",
         12084 => x"6185bf38",
         12085 => x"81587584",
         12086 => x"2e83cd38",
         12087 => x"8d587581",
         12088 => x"2683c538",
         12089 => x"80c41733",
         12090 => x"80c31833",
         12091 => x"71882b07",
         12092 => x"5e597c84",
         12093 => x"802e0981",
         12094 => x"0683ad38",
         12095 => x"80cf1733",
         12096 => x"80ce1833",
         12097 => x"71882b07",
         12098 => x"575a75a4",
         12099 => x"3880dc17",
         12100 => x"83113382",
         12101 => x"12337190",
         12102 => x"2b71882b",
         12103 => x"07811433",
         12104 => x"70720788",
         12105 => x"2b753371",
         12106 => x"07565a45",
         12107 => x"435e5f56",
         12108 => x"75a0180c",
         12109 => x"80c81733",
         12110 => x"82183480",
         12111 => x"c81733ff",
         12112 => x"117081ff",
         12113 => x"065f4059",
         12114 => x"8d587c81",
         12115 => x"2682d938",
         12116 => x"7881ff06",
         12117 => x"76712980",
         12118 => x"c519335a",
         12119 => x"5f5a778a",
         12120 => x"18237759",
         12121 => x"77802e87",
         12122 => x"c438ff18",
         12123 => x"78064261",
         12124 => x"87bb3880",
         12125 => x"ca173380",
         12126 => x"c9183371",
         12127 => x"882b0756",
         12128 => x"40748818",
         12129 => x"2374758f",
         12130 => x"065e5a8d",
         12131 => x"587c8298",
         12132 => x"3880cc17",
         12133 => x"3380cb18",
         12134 => x"3371882b",
         12135 => x"07565c74",
         12136 => x"a43880d8",
         12137 => x"17831133",
         12138 => x"82123371",
         12139 => x"902b7188",
         12140 => x"2b078114",
         12141 => x"33707207",
         12142 => x"882b7533",
         12143 => x"71075344",
         12144 => x"5a584242",
         12145 => x"4280c717",
         12146 => x"3380c618",
         12147 => x"3371882b",
         12148 => x"075d588d",
         12149 => x"587b802e",
         12150 => x"81ce387d",
         12151 => x"1c7a842a",
         12152 => x"055a7975",
         12153 => x"2681c138",
         12154 => x"7852747a",
         12155 => x"3151fded",
         12156 => x"b43f84ba",
         12157 => x"8c085684",
         12158 => x"ba8c0880",
         12159 => x"2e81a938",
         12160 => x"84ba8c08",
         12161 => x"80ffffff",
         12162 => x"f5268338",
         12163 => x"835d7583",
         12164 => x"fff52683",
         12165 => x"38825d75",
         12166 => x"9ff52685",
         12167 => x"eb38815d",
         12168 => x"8216709c",
         12169 => x"190c7ba4",
         12170 => x"190c7b1d",
         12171 => x"70a81a0c",
         12172 => x"7b1db01a",
         12173 => x"0c57597c",
         12174 => x"832e8a87",
         12175 => x"38881722",
         12176 => x"5c8d587b",
         12177 => x"802e80e0",
         12178 => x"387d16ac",
         12179 => x"180c7819",
         12180 => x"557c822e",
         12181 => x"8d387810",
         12182 => x"1970812a",
         12183 => x"7a810605",
         12184 => x"565a83ff",
         12185 => x"15892a59",
         12186 => x"8d5878a0",
         12187 => x"180826b8",
         12188 => x"38ff0b94",
         12189 => x"180cff0b",
         12190 => x"90180cff",
         12191 => x"800b8418",
         12192 => x"347c832e",
         12193 => x"8696387c",
         12194 => x"773484d1",
         12195 => x"e4228105",
         12196 => x"5d7c84d1",
         12197 => x"e4237c86",
         12198 => x"182384d1",
         12199 => x"ec0b8c18",
         12200 => x"0c800b98",
         12201 => x"180c8058",
         12202 => x"7784ba8c",
         12203 => x"0c973d0d",
         12204 => x"048b0b84",
         12205 => x"ba8c0c97",
         12206 => x"3d0d0476",
         12207 => x"33d01170",
         12208 => x"81ff0657",
         12209 => x"57587489",
         12210 => x"26913882",
         12211 => x"177881ff",
         12212 => x"06d0055d",
         12213 => x"59787a2e",
         12214 => x"87fe3880",
         12215 => x"7e0883e5",
         12216 => x"fc5f405c",
         12217 => x"7c087f5a",
         12218 => x"5b7a7081",
         12219 => x"055c3379",
         12220 => x"7081055b",
         12221 => x"33ff9f12",
         12222 => x"5a585677",
         12223 => x"99268938",
         12224 => x"e0167081",
         12225 => x"ff065755",
         12226 => x"ff9f1758",
         12227 => x"77992689",
         12228 => x"38e01770",
         12229 => x"81ff0658",
         12230 => x"55753070",
         12231 => x"9f2a5955",
         12232 => x"75772e09",
         12233 => x"81068538",
         12234 => x"77ffbe38",
         12235 => x"787a3270",
         12236 => x"30707207",
         12237 => x"9f2a7a07",
         12238 => x"5d58557a",
         12239 => x"802e8798",
         12240 => x"38811c84",
         12241 => x"1e5e5c83",
         12242 => x"7c25ff98",
         12243 => x"386156f9",
         12244 => x"a9397880",
         12245 => x"2efecf38",
         12246 => x"77822a81",
         12247 => x"065e8a58",
         12248 => x"7dfec538",
         12249 => x"8058fec0",
         12250 => x"397a7833",
         12251 => x"57597581",
         12252 => x"e92e0981",
         12253 => x"06833881",
         12254 => x"597581eb",
         12255 => x"32703070",
         12256 => x"80257b07",
         12257 => x"5a5b5c77",
         12258 => x"83ad3875",
         12259 => x"81e82e83",
         12260 => x"a638933d",
         12261 => x"77575a83",
         12262 => x"5983fa16",
         12263 => x"3370595b",
         12264 => x"7a802ea5",
         12265 => x"38848116",
         12266 => x"33848017",
         12267 => x"3371902b",
         12268 => x"71882b07",
         12269 => x"83ff1933",
         12270 => x"70720788",
         12271 => x"2b83fe1b",
         12272 => x"33710752",
         12273 => x"595b4040",
         12274 => x"40777a70",
         12275 => x"84055c0c",
         12276 => x"ff199017",
         12277 => x"57597880",
         12278 => x"25ffbe38",
         12279 => x"84ba811d",
         12280 => x"33703070",
         12281 => x"9f2a7271",
         12282 => x"319b3d71",
         12283 => x"101005f0",
         12284 => x"0584b61c",
         12285 => x"445d5243",
         12286 => x"5b427808",
         12287 => x"5b83567a",
         12288 => x"802e80fb",
         12289 => x"38800b83",
         12290 => x"1834ff0b",
         12291 => x"b4180c7a",
         12292 => x"5580567a",
         12293 => x"ff2ea538",
         12294 => x"81547a53",
         12295 => x"b8175281",
         12296 => x"173351ff",
         12297 => x"b4863f84",
         12298 => x"ba8c0876",
         12299 => x"2e8538ff",
         12300 => x"55815674",
         12301 => x"b4180c84",
         12302 => x"5875bf38",
         12303 => x"811f337f",
         12304 => x"3371882b",
         12305 => x"075d5e83",
         12306 => x"587b82d4",
         12307 => x"d52e0981",
         12308 => x"06a83880",
         12309 => x"0bb81833",
         12310 => x"57587581",
         12311 => x"e92e82b7",
         12312 => x"387581eb",
         12313 => x"32703070",
         12314 => x"80257a07",
         12315 => x"4242427f",
         12316 => x"bc387581",
         12317 => x"e82eb638",
         12318 => x"82587781",
         12319 => x"ff065680",
         12320 => x"0b84ba81",
         12321 => x"1e335d58",
         12322 => x"7b782e09",
         12323 => x"81068338",
         12324 => x"81588176",
         12325 => x"27f8bd38",
         12326 => x"77802ef8",
         12327 => x"b738811a",
         12328 => x"841a5a5a",
         12329 => x"837a27fe",
         12330 => x"d138f8a8",
         12331 => x"39830b80",
         12332 => x"ee1883e5",
         12333 => x"bc405d58",
         12334 => x"7b708105",
         12335 => x"5d337e70",
         12336 => x"81054033",
         12337 => x"717131ff",
         12338 => x"1b5b5256",
         12339 => x"5677802e",
         12340 => x"80c53875",
         12341 => x"802ee138",
         12342 => x"850b818a",
         12343 => x"1883e5c0",
         12344 => x"405d587b",
         12345 => x"7081055d",
         12346 => x"337e7081",
         12347 => x"05403371",
         12348 => x"7131ff1b",
         12349 => x"5b584240",
         12350 => x"77802e85",
         12351 => x"8e387580",
         12352 => x"2ee13882",
         12353 => x"58fef339",
         12354 => x"8d587cfa",
         12355 => x"93387784",
         12356 => x"ba8c0c97",
         12357 => x"3d0d0475",
         12358 => x"5875802e",
         12359 => x"fedc3885",
         12360 => x"0b818a18",
         12361 => x"83e5c040",
         12362 => x"5d58ffb7",
         12363 => x"398d0b84",
         12364 => x"ba8c0c97",
         12365 => x"3d0d0483",
         12366 => x"0b80ee18",
         12367 => x"83e5bc5c",
         12368 => x"5a587870",
         12369 => x"81055a33",
         12370 => x"7a708105",
         12371 => x"5c337171",
         12372 => x"31ff1b5b",
         12373 => x"575f5f77",
         12374 => x"802e83d1",
         12375 => x"3874802e",
         12376 => x"e138850b",
         12377 => x"818a1883",
         12378 => x"e5c05c5a",
         12379 => x"58787081",
         12380 => x"055a337a",
         12381 => x"7081055c",
         12382 => x"33717131",
         12383 => x"ff1b5b58",
         12384 => x"42407780",
         12385 => x"2e849138",
         12386 => x"75802ee1",
         12387 => x"38933d77",
         12388 => x"575a8359",
         12389 => x"fc833981",
         12390 => x"58fdc639",
         12391 => x"80e91733",
         12392 => x"80e81833",
         12393 => x"71882b07",
         12394 => x"57557581",
         12395 => x"2e098106",
         12396 => x"f9d53881",
         12397 => x"1b58805a",
         12398 => x"b4170878",
         12399 => x"2eb13883",
         12400 => x"17335b7a",
         12401 => x"7a2e0981",
         12402 => x"06829b38",
         12403 => x"81547753",
         12404 => x"b8175281",
         12405 => x"173351ff",
         12406 => x"b0d23f84",
         12407 => x"ba8c0880",
         12408 => x"2e8538ff",
         12409 => x"58815a77",
         12410 => x"b4180c79",
         12411 => x"f9993879",
         12412 => x"84183484",
         12413 => x"b7173384",
         12414 => x"b6183371",
         12415 => x"882b0757",
         12416 => x"5e7582d4",
         12417 => x"d52e0981",
         12418 => x"06f8fc38",
         12419 => x"b8178311",
         12420 => x"33821233",
         12421 => x"71902b71",
         12422 => x"882b0781",
         12423 => x"14337072",
         12424 => x"07882b75",
         12425 => x"3371075e",
         12426 => x"41594542",
         12427 => x"5c597784",
         12428 => x"8b85a4d2",
         12429 => x"2e098106",
         12430 => x"f8cd3884",
         12431 => x"9c178311",
         12432 => x"33821233",
         12433 => x"71902b71",
         12434 => x"882b0781",
         12435 => x"14337072",
         12436 => x"07882b75",
         12437 => x"33710747",
         12438 => x"44405b5c",
         12439 => x"5a5e6086",
         12440 => x"8a85e4f2",
         12441 => x"2e098106",
         12442 => x"f89d3884",
         12443 => x"a0178311",
         12444 => x"33821233",
         12445 => x"71902b71",
         12446 => x"882b0781",
         12447 => x"14337072",
         12448 => x"07882b75",
         12449 => x"33710794",
         12450 => x"1e0c5d84",
         12451 => x"a41c8311",
         12452 => x"33821233",
         12453 => x"71902b71",
         12454 => x"882b0781",
         12455 => x"14337072",
         12456 => x"07882b75",
         12457 => x"33710762",
         12458 => x"90050c59",
         12459 => x"4449465c",
         12460 => x"4540455b",
         12461 => x"565a7c77",
         12462 => x"3484d1e4",
         12463 => x"2281055d",
         12464 => x"7c84d1e4",
         12465 => x"237c8618",
         12466 => x"2384d1ec",
         12467 => x"0b8c180c",
         12468 => x"800b9818",
         12469 => x"0cf7cf39",
         12470 => x"7b8324f8",
         12471 => x"f0387b7a",
         12472 => x"7f0c56f2",
         12473 => x"95397554",
         12474 => x"b4170853",
         12475 => x"b8177053",
         12476 => x"81183352",
         12477 => x"59ffafb3",
         12478 => x"3f84ba8c",
         12479 => x"087a2e09",
         12480 => x"810681a4",
         12481 => x"3884ba8c",
         12482 => x"08831834",
         12483 => x"b41708a8",
         12484 => x"18083140",
         12485 => x"7fa01808",
         12486 => x"278b3882",
         12487 => x"17334160",
         12488 => x"822e818d",
         12489 => x"3884ba8c",
         12490 => x"085afda0",
         12491 => x"39745674",
         12492 => x"802ef391",
         12493 => x"38850b81",
         12494 => x"8a1883e5",
         12495 => x"c05c5a58",
         12496 => x"fcab3980",
         12497 => x"e3173380",
         12498 => x"e2183371",
         12499 => x"882b075f",
         12500 => x"5a8d587d",
         12501 => x"f6d23888",
         12502 => x"17224261",
         12503 => x"f6ca3880",
         12504 => x"e4178311",
         12505 => x"33821233",
         12506 => x"71902b71",
         12507 => x"882b0781",
         12508 => x"14337072",
         12509 => x"07882b75",
         12510 => x"337107ac",
         12511 => x"1e0c5a7d",
         12512 => x"822b5a43",
         12513 => x"44405940",
         12514 => x"f5d83975",
         12515 => x"5875802e",
         12516 => x"f9e83882",
         12517 => x"58f9e339",
         12518 => x"75802ef2",
         12519 => x"a838933d",
         12520 => x"77575a83",
         12521 => x"59f7f239",
         12522 => x"755a79f5",
         12523 => x"da38fcbf",
         12524 => x"397554b4",
         12525 => x"1708a018",
         12526 => x"08055378",
         12527 => x"52811733",
         12528 => x"51ffade7",
         12529 => x"3ffc8539",
         12530 => x"f03d0d02",
         12531 => x"80d30533",
         12532 => x"64704393",
         12533 => x"3d41575d",
         12534 => x"ff765a40",
         12535 => x"75802e80",
         12536 => x"e9387870",
         12537 => x"81055a33",
         12538 => x"709f2655",
         12539 => x"5574ba2e",
         12540 => x"80e23873",
         12541 => x"ed3874ba",
         12542 => x"2e80d938",
         12543 => x"84d1e833",
         12544 => x"54807424",
         12545 => x"80c43873",
         12546 => x"101084d1",
         12547 => x"d4057008",
         12548 => x"55557380",
         12549 => x"2e843880",
         12550 => x"74346254",
         12551 => x"73802e86",
         12552 => x"38807434",
         12553 => x"62547375",
         12554 => x"0c7c547c",
         12555 => x"802e9238",
         12556 => x"8053933d",
         12557 => x"70538405",
         12558 => x"51ef813f",
         12559 => x"84ba8c08",
         12560 => x"547384ba",
         12561 => x"8c0c923d",
         12562 => x"0d048b0b",
         12563 => x"84ba8c0c",
         12564 => x"923d0d04",
         12565 => x"7533d011",
         12566 => x"7081ff06",
         12567 => x"56565773",
         12568 => x"89269138",
         12569 => x"82167781",
         12570 => x"ff06d005",
         12571 => x"5c587779",
         12572 => x"2e80f738",
         12573 => x"807f0883",
         12574 => x"e5fc5e5f",
         12575 => x"5b7b087e",
         12576 => x"595a7970",
         12577 => x"81055b33",
         12578 => x"78708105",
         12579 => x"5a33ff9f",
         12580 => x"12595755",
         12581 => x"76992689",
         12582 => x"38e01570",
         12583 => x"81ff0656",
         12584 => x"54ff9f16",
         12585 => x"57769926",
         12586 => x"8938e016",
         12587 => x"7081ff06",
         12588 => x"57547430",
         12589 => x"709f2a58",
         12590 => x"5474762e",
         12591 => x"09810685",
         12592 => x"3876ffbe",
         12593 => x"38777932",
         12594 => x"70307072",
         12595 => x"079f2a79",
         12596 => x"075c5754",
         12597 => x"79802e92",
         12598 => x"38811b84",
         12599 => x"1d5d5b83",
         12600 => x"7b25ff99",
         12601 => x"387f54fe",
         12602 => x"98397a83",
         12603 => x"24f7387a",
         12604 => x"79600c54",
         12605 => x"fe8b39e6",
         12606 => x"3d0d6c02",
         12607 => x"840580fb",
         12608 => x"05335659",
         12609 => x"89567880",
         12610 => x"2ea63874",
         12611 => x"bf067054",
         12612 => x"9d3dcc05",
         12613 => x"539e3d84",
         12614 => x"055258ed",
         12615 => x"9f3f84ba",
         12616 => x"8c085784",
         12617 => x"ba8c0880",
         12618 => x"2e8f3880",
         12619 => x"790c7656",
         12620 => x"7584ba8c",
         12621 => x"0c9c3d0d",
         12622 => x"047e406d",
         12623 => x"52903d70",
         12624 => x"525ae19a",
         12625 => x"3f84ba8c",
         12626 => x"085784ba",
         12627 => x"8c08802e",
         12628 => x"81ba3877",
         12629 => x"9c065d7c",
         12630 => x"802e81ca",
         12631 => x"3876802e",
         12632 => x"83c13876",
         12633 => x"842e83ea",
         12634 => x"38778807",
         12635 => x"5876ffbb",
         12636 => x"3877832a",
         12637 => x"81065b7a",
         12638 => x"802e81d1",
         12639 => x"38669b11",
         12640 => x"339a1233",
         12641 => x"71882b07",
         12642 => x"61703342",
         12643 => x"585e5e56",
         12644 => x"7d832e84",
         12645 => x"e938800b",
         12646 => x"8e173480",
         12647 => x"0b8f1734",
         12648 => x"a10b9017",
         12649 => x"3480cc0b",
         12650 => x"91173466",
         12651 => x"56a00b8b",
         12652 => x"17347e67",
         12653 => x"575e800b",
         12654 => x"9a173480",
         12655 => x"0b9b1734",
         12656 => x"7d335d7c",
         12657 => x"832e84a9",
         12658 => x"38665b80",
         12659 => x"0b9c1c34",
         12660 => x"800b9d1c",
         12661 => x"34800b9e",
         12662 => x"1c34800b",
         12663 => x"9f1c347e",
         12664 => x"55810b83",
         12665 => x"16347b80",
         12666 => x"2e80e238",
         12667 => x"7eb41108",
         12668 => x"7d7c0853",
         12669 => x"575f5781",
         12670 => x"7c278938",
         12671 => x"9c17087c",
         12672 => x"26838a38",
         12673 => x"82578079",
         12674 => x"0cfea339",
         12675 => x"0280e705",
         12676 => x"3370982b",
         12677 => x"5d5b7b80",
         12678 => x"25feb838",
         12679 => x"86789c06",
         12680 => x"5e577cfe",
         12681 => x"b83876fe",
         12682 => x"82380280",
         12683 => x"c2053370",
         12684 => x"842a8106",
         12685 => x"5d567b82",
         12686 => x"91387781",
         12687 => x"2a81065e",
         12688 => x"7d802e89",
         12689 => x"38758106",
         12690 => x"5a7981f6",
         12691 => x"3877832a",
         12692 => x"81065675",
         12693 => x"802e8638",
         12694 => x"7780c007",
         12695 => x"587eb411",
         12696 => x"08a01b0c",
         12697 => x"67a41b0c",
         12698 => x"679b1133",
         12699 => x"9a123371",
         12700 => x"882b0773",
         12701 => x"33405e40",
         12702 => x"575a7b83",
         12703 => x"2e81f138",
         12704 => x"7a881a0c",
         12705 => x"9c168311",
         12706 => x"33821233",
         12707 => x"71902b71",
         12708 => x"882b0781",
         12709 => x"14337072",
         12710 => x"07882b75",
         12711 => x"33710770",
         12712 => x"608c050c",
         12713 => x"60600c51",
         12714 => x"52415957",
         12715 => x"5d5e861a",
         12716 => x"22841a23",
         12717 => x"77901a34",
         12718 => x"800b911a",
         12719 => x"34800b9c",
         12720 => x"1a0c7785",
         12721 => x"2a810655",
         12722 => x"74802e84",
         12723 => x"ac387580",
         12724 => x"2e84f138",
         12725 => x"75941a0c",
         12726 => x"8a1a2270",
         12727 => x"892b7c52",
         12728 => x"5b587630",
         12729 => x"70780780",
         12730 => x"25565b79",
         12731 => x"76278492",
         12732 => x"38817076",
         12733 => x"065f5b7d",
         12734 => x"802e8486",
         12735 => x"38775278",
         12736 => x"51ffacdb",
         12737 => x"3f84ba8c",
         12738 => x"085884ba",
         12739 => x"8c088126",
         12740 => x"83388257",
         12741 => x"84ba8c08",
         12742 => x"ff2e80cb",
         12743 => x"38757a31",
         12744 => x"56c03902",
         12745 => x"80c20533",
         12746 => x"91065e7d",
         12747 => x"95387782",
         12748 => x"2a810655",
         12749 => x"74802efc",
         12750 => x"b8388857",
         12751 => x"80790cfb",
         12752 => x"ed398757",
         12753 => x"80790cfb",
         12754 => x"e5398457",
         12755 => x"80790cfb",
         12756 => x"dd397951",
         12757 => x"cdca3f84",
         12758 => x"ba8c0878",
         12759 => x"88075957",
         12760 => x"76fbc838",
         12761 => x"fc8b397a",
         12762 => x"767b3157",
         12763 => x"57fef339",
         12764 => x"95163394",
         12765 => x"17337198",
         12766 => x"2b71902b",
         12767 => x"077d075d",
         12768 => x"5e5cfdfc",
         12769 => x"397c557c",
         12770 => x"7b2781bd",
         12771 => x"38745279",
         12772 => x"51ffabcb",
         12773 => x"3f84ba8c",
         12774 => x"085d84ba",
         12775 => x"8c08802e",
         12776 => x"81a73884",
         12777 => x"ba8c0881",
         12778 => x"2efcd938",
         12779 => x"84ba8c08",
         12780 => x"ff2e8399",
         12781 => x"38805374",
         12782 => x"527651ff",
         12783 => x"b2823f84",
         12784 => x"ba8c0883",
         12785 => x"90389c17",
         12786 => x"08fe1194",
         12787 => x"19085856",
         12788 => x"5b757527",
         12789 => x"ffaf3881",
         12790 => x"1694180c",
         12791 => x"84173381",
         12792 => x"07557484",
         12793 => x"18347c55",
         12794 => x"7a7d26ff",
         12795 => x"a03880d9",
         12796 => x"39800b94",
         12797 => x"1734800b",
         12798 => x"951734fb",
         12799 => x"cc399516",
         12800 => x"33941733",
         12801 => x"71982b71",
         12802 => x"902b077e",
         12803 => x"075e565b",
         12804 => x"800b8e17",
         12805 => x"34800b8f",
         12806 => x"1734a10b",
         12807 => x"90173480",
         12808 => x"cc0b9117",
         12809 => x"346656a0",
         12810 => x"0b8b1734",
         12811 => x"7e67575e",
         12812 => x"800b9a17",
         12813 => x"34800b9b",
         12814 => x"17347d33",
         12815 => x"5d7c832e",
         12816 => x"098106fb",
         12817 => x"8438ffa9",
         12818 => x"39807f7f",
         12819 => x"725e5957",
         12820 => x"5db41608",
         12821 => x"7e2eae38",
         12822 => x"8316335a",
         12823 => x"797d2e09",
         12824 => x"8106b538",
         12825 => x"81547d53",
         12826 => x"b8165281",
         12827 => x"163351ff",
         12828 => x"a3ba3f84",
         12829 => x"ba8c0880",
         12830 => x"2e8538ff",
         12831 => x"57815b76",
         12832 => x"b4170c7e",
         12833 => x"567aff1d",
         12834 => x"90180c57",
         12835 => x"7a802efb",
         12836 => x"bc388079",
         12837 => x"0cf99739",
         12838 => x"8154b416",
         12839 => x"0853b816",
         12840 => x"70538117",
         12841 => x"33525aff",
         12842 => x"a4813f84",
         12843 => x"ba8c087d",
         12844 => x"2e098106",
         12845 => x"81aa3884",
         12846 => x"ba8c0883",
         12847 => x"1734b416",
         12848 => x"08a81708",
         12849 => x"3184ba8c",
         12850 => x"085c5574",
         12851 => x"a0170827",
         12852 => x"ff923882",
         12853 => x"16335574",
         12854 => x"822e0981",
         12855 => x"06ff8538",
         12856 => x"8154b416",
         12857 => x"08a01708",
         12858 => x"05537952",
         12859 => x"81163351",
         12860 => x"ffa3b83f",
         12861 => x"7c5bfeec",
         12862 => x"3974941a",
         12863 => x"0c7656f8",
         12864 => x"af397798",
         12865 => x"1a0c76f8",
         12866 => x"a2387583",
         12867 => x"ff065a79",
         12868 => x"802ef89a",
         12869 => x"387efe19",
         12870 => x"9c1208fe",
         12871 => x"055f595a",
         12872 => x"777d27f9",
         12873 => x"df388a1a",
         12874 => x"22787129",
         12875 => x"b01c0805",
         12876 => x"565c7480",
         12877 => x"2ef9cd38",
         12878 => x"75892a15",
         12879 => x"9c1a0c76",
         12880 => x"56f7ed39",
         12881 => x"75941a0c",
         12882 => x"7656f7e4",
         12883 => x"39815780",
         12884 => x"790cf7da",
         12885 => x"3984ba8c",
         12886 => x"08578079",
         12887 => x"0cf7cf39",
         12888 => x"817f575b",
         12889 => x"fe9f39f0",
         12890 => x"3d0d6265",
         12891 => x"67664040",
         12892 => x"5d5a807e",
         12893 => x"0c895779",
         12894 => x"802e9f38",
         12895 => x"79085675",
         12896 => x"802e9738",
         12897 => x"75335574",
         12898 => x"802e8f38",
         12899 => x"86162284",
         12900 => x"1b225959",
         12901 => x"78782e84",
         12902 => x"b7388055",
         12903 => x"74417655",
         12904 => x"76828c38",
         12905 => x"911a3355",
         12906 => x"74828438",
         12907 => x"901a3381",
         12908 => x"06578756",
         12909 => x"76802e81",
         12910 => x"ed38941a",
         12911 => x"088c1b08",
         12912 => x"71315656",
         12913 => x"7b752681",
         12914 => x"ef387b80",
         12915 => x"2e81d538",
         12916 => x"60597583",
         12917 => x"ff065b7a",
         12918 => x"81e3388a",
         12919 => x"1922ff05",
         12920 => x"76892a06",
         12921 => x"5b7a9b38",
         12922 => x"7583d338",
         12923 => x"881a0855",
         12924 => x"81752784",
         12925 => x"853874ff",
         12926 => x"2e83f038",
         12927 => x"74981b0c",
         12928 => x"6059981a",
         12929 => x"08fe059c",
         12930 => x"1a08fe05",
         12931 => x"41577660",
         12932 => x"2783e738",
         12933 => x"8a192270",
         12934 => x"7829b01b",
         12935 => x"08055656",
         12936 => x"74802e83",
         12937 => x"d5387a15",
         12938 => x"7c892a59",
         12939 => x"5777802e",
         12940 => x"83813877",
         12941 => x"1b557575",
         12942 => x"27853875",
         12943 => x"7b315877",
         12944 => x"5476537c",
         12945 => x"52811933",
         12946 => x"51ff9fe0",
         12947 => x"3f84ba8c",
         12948 => x"08839838",
         12949 => x"60831133",
         12950 => x"57597580",
         12951 => x"2ea938b4",
         12952 => x"19087731",
         12953 => x"56757827",
         12954 => x"9e388480",
         12955 => x"7671291e",
         12956 => x"b81b5858",
         12957 => x"55757081",
         12958 => x"05573377",
         12959 => x"70810559",
         12960 => x"34ff1555",
         12961 => x"74ef3877",
         12962 => x"892b587b",
         12963 => x"78317e08",
         12964 => x"197f0c78",
         12965 => x"1e941c08",
         12966 => x"1a705994",
         12967 => x"1d0c5e5c",
         12968 => x"7bfeaf38",
         12969 => x"80567584",
         12970 => x"ba8c0c92",
         12971 => x"3d0d0474",
         12972 => x"84ba8c0c",
         12973 => x"923d0d04",
         12974 => x"745cfe8e",
         12975 => x"399c1a08",
         12976 => x"577583ff",
         12977 => x"06848071",
         12978 => x"31595b7b",
         12979 => x"78278338",
         12980 => x"7b587656",
         12981 => x"b4190877",
         12982 => x"2eb63880",
         12983 => x"0b831a33",
         12984 => x"715d415f",
         12985 => x"7f7f2e09",
         12986 => x"810680e4",
         12987 => x"38815476",
         12988 => x"53b81952",
         12989 => x"81193351",
         12990 => x"ff9eb13f",
         12991 => x"84ba8c08",
         12992 => x"802e8538",
         12993 => x"ff56815b",
         12994 => x"75b41a0c",
         12995 => x"7a81dc38",
         12996 => x"60941b08",
         12997 => x"83ff0611",
         12998 => x"797f5a58",
         12999 => x"b8055659",
         13000 => x"77802efe",
         13001 => x"e6387470",
         13002 => x"81055633",
         13003 => x"77708105",
         13004 => x"5934ff16",
         13005 => x"5675802e",
         13006 => x"fed13874",
         13007 => x"70810556",
         13008 => x"33777081",
         13009 => x"055934ff",
         13010 => x"165675da",
         13011 => x"38febc39",
         13012 => x"8154b419",
         13013 => x"0853b819",
         13014 => x"7053811a",
         13015 => x"335240ff",
         13016 => x"9ec93f81",
         13017 => x"5b84ba8c",
         13018 => x"087f2e09",
         13019 => x"8106ff9c",
         13020 => x"3884ba8c",
         13021 => x"08831a34",
         13022 => x"b41908a8",
         13023 => x"1a083184",
         13024 => x"ba8c085c",
         13025 => x"5574a01a",
         13026 => x"0827fee1",
         13027 => x"38821933",
         13028 => x"5574822e",
         13029 => x"098106fe",
         13030 => x"d4388154",
         13031 => x"b41908a0",
         13032 => x"1a080553",
         13033 => x"7f528119",
         13034 => x"3351ff9d",
         13035 => x"fe3f7e5b",
         13036 => x"febb3976",
         13037 => x"9c1b0c94",
         13038 => x"1a0856fe",
         13039 => x"8439981a",
         13040 => x"08527951",
         13041 => x"ffa3983f",
         13042 => x"84ba8c08",
         13043 => x"55fca139",
         13044 => x"81163351",
         13045 => x"ff9c833f",
         13046 => x"84ba8c08",
         13047 => x"81065574",
         13048 => x"fbb83874",
         13049 => x"7a085657",
         13050 => x"fbb23981",
         13051 => x"0b911b34",
         13052 => x"810b84ba",
         13053 => x"8c0c923d",
         13054 => x"0d04820b",
         13055 => x"911b3482",
         13056 => x"0b84ba8c",
         13057 => x"0c923d0d",
         13058 => x"04f03d0d",
         13059 => x"62656766",
         13060 => x"40405c5a",
         13061 => x"807e0c89",
         13062 => x"5779802e",
         13063 => x"9f387908",
         13064 => x"5675802e",
         13065 => x"97387533",
         13066 => x"5574802e",
         13067 => x"8f388616",
         13068 => x"22841b22",
         13069 => x"59597878",
         13070 => x"2e85fd38",
         13071 => x"80557441",
         13072 => x"76557682",
         13073 => x"c438911a",
         13074 => x"33557482",
         13075 => x"bc38901a",
         13076 => x"3370812a",
         13077 => x"81065858",
         13078 => x"87567680",
         13079 => x"2e82a138",
         13080 => x"941a087b",
         13081 => x"115d577b",
         13082 => x"77278438",
         13083 => x"76095b7a",
         13084 => x"802e8281",
         13085 => x"387683ff",
         13086 => x"065f7e82",
         13087 => x"a238608a",
         13088 => x"1122ff05",
         13089 => x"78892a06",
         13090 => x"5a5678aa",
         13091 => x"3876849e",
         13092 => x"38881a08",
         13093 => x"5574802e",
         13094 => x"84b13874",
         13095 => x"812e86a1",
         13096 => x"3874ff2e",
         13097 => x"868c3874",
         13098 => x"981b0c88",
         13099 => x"1a088538",
         13100 => x"74881b0c",
         13101 => x"6056b416",
         13102 => x"089c1b08",
         13103 => x"2e81d338",
         13104 => x"981a08fe",
         13105 => x"059c1708",
         13106 => x"fe055858",
         13107 => x"77772785",
         13108 => x"f0388a16",
         13109 => x"22707929",
         13110 => x"b0180805",
         13111 => x"56577480",
         13112 => x"2e85de38",
         13113 => x"78157b89",
         13114 => x"2a595c77",
         13115 => x"802e8398",
         13116 => x"3877195f",
         13117 => x"767f2785",
         13118 => x"38767931",
         13119 => x"5877547b",
         13120 => x"537c5281",
         13121 => x"163351ff",
         13122 => x"9ba13f84",
         13123 => x"ba8c0885",
         13124 => x"a13860b4",
         13125 => x"11087d31",
         13126 => x"56577478",
         13127 => x"27a53884",
         13128 => x"800bb818",
         13129 => x"7672291f",
         13130 => x"57585674",
         13131 => x"70810556",
         13132 => x"33777081",
         13133 => x"055934ff",
         13134 => x"165675ef",
         13135 => x"38605975",
         13136 => x"831a3477",
         13137 => x"892b597a",
         13138 => x"79317e08",
         13139 => x"1a7f0c79",
         13140 => x"1e941c08",
         13141 => x"1b707194",
         13142 => x"1f0c8c1e",
         13143 => x"085a5a57",
         13144 => x"5e5b7575",
         13145 => x"27833874",
         13146 => x"56758c1b",
         13147 => x"0c7afe85",
         13148 => x"38901a33",
         13149 => x"587780c0",
         13150 => x"075b7a90",
         13151 => x"1b348056",
         13152 => x"7584ba8c",
         13153 => x"0c923d0d",
         13154 => x"047484ba",
         13155 => x"8c0c923d",
         13156 => x"0d048316",
         13157 => x"33557482",
         13158 => x"c8386056",
         13159 => x"fea23960",
         13160 => x"9c1b0859",
         13161 => x"567683ff",
         13162 => x"06848071",
         13163 => x"315a5c7a",
         13164 => x"79278338",
         13165 => x"7a597757",
         13166 => x"b4160878",
         13167 => x"2eb63880",
         13168 => x"0b831733",
         13169 => x"715e415f",
         13170 => x"7f7f2e09",
         13171 => x"810680d5",
         13172 => x"38815477",
         13173 => x"53b81652",
         13174 => x"81163351",
         13175 => x"ff98cd3f",
         13176 => x"84ba8c08",
         13177 => x"802e8538",
         13178 => x"ff57815c",
         13179 => x"76b4170c",
         13180 => x"7b83bf38",
         13181 => x"60941b08",
         13182 => x"83ff0611",
         13183 => x"7a58b805",
         13184 => x"7e595658",
         13185 => x"78802e95",
         13186 => x"38767081",
         13187 => x"05583375",
         13188 => x"70810557",
         13189 => x"34ff1656",
         13190 => x"75ef3860",
         13191 => x"58810b83",
         13192 => x"1934fea3",
         13193 => x"398154b4",
         13194 => x"160853b8",
         13195 => x"16705381",
         13196 => x"17335240",
         13197 => x"ff98f43f",
         13198 => x"815c84ba",
         13199 => x"8c087f2e",
         13200 => x"098106ff",
         13201 => x"ab3884ba",
         13202 => x"8c088317",
         13203 => x"34b41608",
         13204 => x"a8170831",
         13205 => x"84ba8c08",
         13206 => x"5d5574a0",
         13207 => x"170827fe",
         13208 => x"f0388216",
         13209 => x"33557482",
         13210 => x"2e098106",
         13211 => x"fee33881",
         13212 => x"54b41608",
         13213 => x"a0170805",
         13214 => x"537f5281",
         13215 => x"163351ff",
         13216 => x"98a93f7e",
         13217 => x"5cfeca39",
         13218 => x"941a0857",
         13219 => x"8c1a0877",
         13220 => x"26933883",
         13221 => x"1633407f",
         13222 => x"81b93860",
         13223 => x"7cb4120c",
         13224 => x"941b0858",
         13225 => x"567b7c9c",
         13226 => x"1c0c58fd",
         13227 => x"f839981a",
         13228 => x"08527951",
         13229 => x"ffabe73f",
         13230 => x"84ba8c08",
         13231 => x"5584ba8c",
         13232 => x"08fbd838",
         13233 => x"901a3358",
         13234 => x"fdab3976",
         13235 => x"527951ff",
         13236 => x"abcc3f84",
         13237 => x"ba8c0855",
         13238 => x"84ba8c08",
         13239 => x"fbbd38e4",
         13240 => x"398154b4",
         13241 => x"160853b8",
         13242 => x"16705381",
         13243 => x"17335257",
         13244 => x"ff97b83f",
         13245 => x"84ba8c08",
         13246 => x"81b83884",
         13247 => x"ba8c0883",
         13248 => x"1734b416",
         13249 => x"08a81708",
         13250 => x"315877a0",
         13251 => x"170827fd",
         13252 => x"89388216",
         13253 => x"335c7b82",
         13254 => x"2e098106",
         13255 => x"fcfc3881",
         13256 => x"54b41608",
         13257 => x"a0170805",
         13258 => x"53765281",
         13259 => x"163351ff",
         13260 => x"96f93f60",
         13261 => x"56fb8939",
         13262 => x"81163351",
         13263 => x"ff959b3f",
         13264 => x"84ba8c08",
         13265 => x"81065574",
         13266 => x"f9f23874",
         13267 => x"7a085657",
         13268 => x"f9ec3981",
         13269 => x"54b41608",
         13270 => x"53b81670",
         13271 => x"53811733",
         13272 => x"5257ff96",
         13273 => x"c63f84ba",
         13274 => x"8c0880c6",
         13275 => x"3884ba8c",
         13276 => x"08831734",
         13277 => x"b41608a8",
         13278 => x"17083155",
         13279 => x"74a01708",
         13280 => x"27fe9838",
         13281 => x"82163358",
         13282 => x"77822e09",
         13283 => x"8106fe8b",
         13284 => x"388154b4",
         13285 => x"1608a017",
         13286 => x"08055376",
         13287 => x"52811633",
         13288 => x"51ff9687",
         13289 => x"3f607cb4",
         13290 => x"120c941b",
         13291 => x"085856fd",
         13292 => x"f439810b",
         13293 => x"911b3481",
         13294 => x"0b84ba8c",
         13295 => x"0c923d0d",
         13296 => x"04820b91",
         13297 => x"1b34820b",
         13298 => x"84ba8c0c",
         13299 => x"923d0d04",
         13300 => x"f53d0d7d",
         13301 => x"58895a77",
         13302 => x"802e9f38",
         13303 => x"77085675",
         13304 => x"802e9738",
         13305 => x"75335574",
         13306 => x"802e8f38",
         13307 => x"86162284",
         13308 => x"19225859",
         13309 => x"78772e83",
         13310 => x"b5388055",
         13311 => x"745c7956",
         13312 => x"7981d838",
         13313 => x"90183370",
         13314 => x"862a8106",
         13315 => x"5c577a80",
         13316 => x"2e81c838",
         13317 => x"7ba01908",
         13318 => x"5a57b417",
         13319 => x"08792eac",
         13320 => x"38831733",
         13321 => x"5b7a81bc",
         13322 => x"38815478",
         13323 => x"53b81752",
         13324 => x"81173351",
         13325 => x"ff93f53f",
         13326 => x"84ba8c08",
         13327 => x"802e8538",
         13328 => x"ff598156",
         13329 => x"78b4180c",
         13330 => x"75819038",
         13331 => x"a418088b",
         13332 => x"1133a007",
         13333 => x"5a57788b",
         13334 => x"18347708",
         13335 => x"88190870",
         13336 => x"83ffff06",
         13337 => x"5d5a567a",
         13338 => x"9a18347a",
         13339 => x"882a5a79",
         13340 => x"9b18349c",
         13341 => x"17763396",
         13342 => x"195c565b",
         13343 => x"74832e81",
         13344 => x"c1388c18",
         13345 => x"0855747b",
         13346 => x"3474882a",
         13347 => x"5b7a9d18",
         13348 => x"3474902a",
         13349 => x"56759e18",
         13350 => x"3474982a",
         13351 => x"59789f18",
         13352 => x"34807a34",
         13353 => x"800b9718",
         13354 => x"34a10b98",
         13355 => x"183480cc",
         13356 => x"0b991834",
         13357 => x"800b9218",
         13358 => x"34800b93",
         13359 => x"18347b5b",
         13360 => x"810b831c",
         13361 => x"347b51ff",
         13362 => x"96943f84",
         13363 => x"ba8c0890",
         13364 => x"193381bf",
         13365 => x"065b5679",
         13366 => x"90193475",
         13367 => x"84ba8c0c",
         13368 => x"8d3d0d04",
         13369 => x"8154b417",
         13370 => x"0853b817",
         13371 => x"70538118",
         13372 => x"33525bff",
         13373 => x"93b53f81",
         13374 => x"5684ba8c",
         13375 => x"08fec938",
         13376 => x"84ba8c08",
         13377 => x"831834b4",
         13378 => x"1708a818",
         13379 => x"083184ba",
         13380 => x"8c085755",
         13381 => x"74a01808",
         13382 => x"27fe8e38",
         13383 => x"82173355",
         13384 => x"74822e09",
         13385 => x"8106fe81",
         13386 => x"388154b4",
         13387 => x"1708a018",
         13388 => x"0805537a",
         13389 => x"52811733",
         13390 => x"51ff92ef",
         13391 => x"3f7956fd",
         13392 => x"e8397890",
         13393 => x"2a557494",
         13394 => x"18347488",
         13395 => x"2a567595",
         13396 => x"18348c18",
         13397 => x"0855747b",
         13398 => x"3474882a",
         13399 => x"5b7a9d18",
         13400 => x"3474902a",
         13401 => x"56759e18",
         13402 => x"3474982a",
         13403 => x"59789f18",
         13404 => x"34807a34",
         13405 => x"800b9718",
         13406 => x"34a10b98",
         13407 => x"183480cc",
         13408 => x"0b991834",
         13409 => x"800b9218",
         13410 => x"34800b93",
         13411 => x"18347b5b",
         13412 => x"810b831c",
         13413 => x"347b51ff",
         13414 => x"94c43f84",
         13415 => x"ba8c0890",
         13416 => x"193381bf",
         13417 => x"065b5679",
         13418 => x"901934fe",
         13419 => x"ae398116",
         13420 => x"3351ff90",
         13421 => x"a53f84ba",
         13422 => x"8c088106",
         13423 => x"5574fcba",
         13424 => x"38747808",
         13425 => x"565afcb4",
         13426 => x"39f93d0d",
         13427 => x"79705255",
         13428 => x"fbfe3f84",
         13429 => x"ba8c0854",
         13430 => x"84ba8c08",
         13431 => x"b1388956",
         13432 => x"74802e9e",
         13433 => x"38740853",
         13434 => x"72802e96",
         13435 => x"38723352",
         13436 => x"71802e8e",
         13437 => x"38861322",
         13438 => x"84162258",
         13439 => x"5271772e",
         13440 => x"96388052",
         13441 => x"71587554",
         13442 => x"75843875",
         13443 => x"750c7384",
         13444 => x"ba8c0c89",
         13445 => x"3d0d0481",
         13446 => x"133351ff",
         13447 => x"8fbc3f84",
         13448 => x"ba8c0881",
         13449 => x"065372da",
         13450 => x"38737508",
         13451 => x"5356d539",
         13452 => x"f63d0dff",
         13453 => x"7d705b57",
         13454 => x"5b75802e",
         13455 => x"b2387570",
         13456 => x"81055733",
         13457 => x"709f2652",
         13458 => x"5271ba2e",
         13459 => x"ac3870ee",
         13460 => x"3871ba2e",
         13461 => x"a43884d1",
         13462 => x"e8335180",
         13463 => x"71249038",
         13464 => x"7084d1e8",
         13465 => x"34800b84",
         13466 => x"ba8c0c8c",
         13467 => x"3d0d048b",
         13468 => x"0b84ba8c",
         13469 => x"0c8c3d0d",
         13470 => x"047833d0",
         13471 => x"117081ff",
         13472 => x"06535353",
         13473 => x"70892691",
         13474 => x"38821973",
         13475 => x"81ff06d0",
         13476 => x"05595473",
         13477 => x"762e80f5",
         13478 => x"38800b83",
         13479 => x"e5fc5b58",
         13480 => x"79087956",
         13481 => x"57767081",
         13482 => x"05583375",
         13483 => x"70810557",
         13484 => x"33ff9f12",
         13485 => x"53545270",
         13486 => x"99268938",
         13487 => x"e0127081",
         13488 => x"ff065354",
         13489 => x"ff9f1351",
         13490 => x"70992689",
         13491 => x"38e01370",
         13492 => x"81ff0654",
         13493 => x"54713070",
         13494 => x"9f2a5551",
         13495 => x"71732e09",
         13496 => x"81068538",
         13497 => x"73ffbe38",
         13498 => x"74763270",
         13499 => x"30707207",
         13500 => x"9f2a7607",
         13501 => x"59525276",
         13502 => x"802e9238",
         13503 => x"8118841b",
         13504 => x"5b588378",
         13505 => x"25ff9938",
         13506 => x"7a51fecf",
         13507 => x"39778324",
         13508 => x"f7387776",
         13509 => x"5e51fec3",
         13510 => x"39ea3d0d",
         13511 => x"8053983d",
         13512 => x"cc055299",
         13513 => x"3d51d194",
         13514 => x"3f84ba8c",
         13515 => x"085584ba",
         13516 => x"8c08802e",
         13517 => x"8a387484",
         13518 => x"ba8c0c98",
         13519 => x"3d0d047a",
         13520 => x"5c685298",
         13521 => x"3dd00551",
         13522 => x"c5943f84",
         13523 => x"ba8c0855",
         13524 => x"84ba8c08",
         13525 => x"80c63802",
         13526 => x"80d70533",
         13527 => x"70982b58",
         13528 => x"5a807724",
         13529 => x"80e23802",
         13530 => x"b2053370",
         13531 => x"842a8106",
         13532 => x"57597580",
         13533 => x"2eb2387a",
         13534 => x"639b1133",
         13535 => x"9a123371",
         13536 => x"882b0773",
         13537 => x"335e5a5b",
         13538 => x"57587983",
         13539 => x"2ea43876",
         13540 => x"98190c74",
         13541 => x"84ba8c0c",
         13542 => x"983d0d04",
         13543 => x"84ba8c08",
         13544 => x"842e0981",
         13545 => x"06ff8f38",
         13546 => x"850b84ba",
         13547 => x"8c0c983d",
         13548 => x"0d049516",
         13549 => x"33941733",
         13550 => x"71982b71",
         13551 => x"902b0779",
         13552 => x"07981b0c",
         13553 => x"5b54cc39",
         13554 => x"7a7e9812",
         13555 => x"0c587484",
         13556 => x"ba8c0c98",
         13557 => x"3d0d04ff",
         13558 => x"9e3d0d80",
         13559 => x"e63d0880",
         13560 => x"e63d085d",
         13561 => x"40807c34",
         13562 => x"805380e4",
         13563 => x"3dfdb405",
         13564 => x"5280e53d",
         13565 => x"51cfc53f",
         13566 => x"84ba8c08",
         13567 => x"5984ba8c",
         13568 => x"0883c838",
         13569 => x"6080d93d",
         13570 => x"0c7f6198",
         13571 => x"110880dd",
         13572 => x"3d0c5880",
         13573 => x"db3d085b",
         13574 => x"5879802e",
         13575 => x"82cc3880",
         13576 => x"d83d983d",
         13577 => x"405ba052",
         13578 => x"7a51ffa4",
         13579 => x"aa3f84ba",
         13580 => x"8c085984",
         13581 => x"ba8c0883",
         13582 => x"92386080",
         13583 => x"df3d0858",
         13584 => x"56b41608",
         13585 => x"772eb138",
         13586 => x"84ba8c08",
         13587 => x"8317335f",
         13588 => x"5d7d83c7",
         13589 => x"38815476",
         13590 => x"53b81652",
         13591 => x"81163351",
         13592 => x"ff8bc93f",
         13593 => x"84ba8c08",
         13594 => x"802e8538",
         13595 => x"ff578159",
         13596 => x"76b4170c",
         13597 => x"7882d438",
         13598 => x"80df3d08",
         13599 => x"9b11339a",
         13600 => x"12337188",
         13601 => x"2b076370",
         13602 => x"335d4059",
         13603 => x"56567883",
         13604 => x"2e82da38",
         13605 => x"7680db3d",
         13606 => x"0c80527a",
         13607 => x"51ffa3b7",
         13608 => x"3f84ba8c",
         13609 => x"085984ba",
         13610 => x"8c08829f",
         13611 => x"3880527a",
         13612 => x"51ffa8f5",
         13613 => x"3f84ba8c",
         13614 => x"085984ba",
         13615 => x"8c08bb38",
         13616 => x"80df3d08",
         13617 => x"9b11339a",
         13618 => x"12337188",
         13619 => x"2b076370",
         13620 => x"33425859",
         13621 => x"5e567d83",
         13622 => x"2e81fd38",
         13623 => x"767a2ea4",
         13624 => x"3884ba8c",
         13625 => x"08527a51",
         13626 => x"ffa4e23f",
         13627 => x"84ba8c08",
         13628 => x"5984ba8c",
         13629 => x"08802eff",
         13630 => x"b4387884",
         13631 => x"2e83d838",
         13632 => x"7881c838",
         13633 => x"80e43dfd",
         13634 => x"b805527a",
         13635 => x"51ffbd89",
         13636 => x"3f787f82",
         13637 => x"05335b57",
         13638 => x"79802e90",
         13639 => x"38821f56",
         13640 => x"81178117",
         13641 => x"70335f57",
         13642 => x"577cf538",
         13643 => x"81175675",
         13644 => x"78268195",
         13645 => x"3876802e",
         13646 => x"9c387e17",
         13647 => x"820556ff",
         13648 => x"1880e63d",
         13649 => x"0811ff19",
         13650 => x"ff195959",
         13651 => x"56587533",
         13652 => x"753476eb",
         13653 => x"38ff1880",
         13654 => x"e63d0811",
         13655 => x"5f58af7e",
         13656 => x"3480da3d",
         13657 => x"085a79fd",
         13658 => x"bd387760",
         13659 => x"2e828a38",
         13660 => x"800b84d1",
         13661 => x"e8337010",
         13662 => x"1083e5fc",
         13663 => x"05700870",
         13664 => x"33435959",
         13665 => x"5e5a7e7a",
         13666 => x"2e8d3881",
         13667 => x"1a701770",
         13668 => x"33575f5a",
         13669 => x"74f53882",
         13670 => x"1a5b7a78",
         13671 => x"26ab3880",
         13672 => x"57767a27",
         13673 => x"94387616",
         13674 => x"5f7e337c",
         13675 => x"7081055e",
         13676 => x"34811757",
         13677 => x"797726ee",
         13678 => x"38ba7c70",
         13679 => x"81055e34",
         13680 => x"76ff2e09",
         13681 => x"810681df",
         13682 => x"38915980",
         13683 => x"7c347884",
         13684 => x"ba8c0c80",
         13685 => x"e43d0d04",
         13686 => x"95163394",
         13687 => x"17337198",
         13688 => x"2b71902b",
         13689 => x"07790759",
         13690 => x"565efdf0",
         13691 => x"39951633",
         13692 => x"94173371",
         13693 => x"982b7190",
         13694 => x"2b077907",
         13695 => x"80dd3d0c",
         13696 => x"5a5d8052",
         13697 => x"7a51ffa0",
         13698 => x"ce3f84ba",
         13699 => x"8c085984",
         13700 => x"ba8c0880",
         13701 => x"2efd9638",
         13702 => x"ffb13981",
         13703 => x"54b41608",
         13704 => x"53b81670",
         13705 => x"53811733",
         13706 => x"525eff88",
         13707 => x"fe3f8159",
         13708 => x"84ba8c08",
         13709 => x"fcbe3884",
         13710 => x"ba8c0883",
         13711 => x"1734b416",
         13712 => x"08a81708",
         13713 => x"3184ba8c",
         13714 => x"085a5574",
         13715 => x"a0170827",
         13716 => x"fc833882",
         13717 => x"16335574",
         13718 => x"822e0981",
         13719 => x"06fbf638",
         13720 => x"8154b416",
         13721 => x"08a01708",
         13722 => x"05537d52",
         13723 => x"81163351",
         13724 => x"ff88b83f",
         13725 => x"7c59fbdd",
         13726 => x"39ff1880",
         13727 => x"e63d0811",
         13728 => x"5c58af7b",
         13729 => x"34800b84",
         13730 => x"d1e83370",
         13731 => x"101083e5",
         13732 => x"fc057008",
         13733 => x"70334359",
         13734 => x"595e5a7e",
         13735 => x"7a2e0981",
         13736 => x"06fde838",
         13737 => x"fdf13980",
         13738 => x"e53d0818",
         13739 => x"8119595a",
         13740 => x"79337c70",
         13741 => x"81055e34",
         13742 => x"776027fe",
         13743 => x"8e3880e5",
         13744 => x"3d081881",
         13745 => x"19595a79",
         13746 => x"337c7081",
         13747 => x"055e347f",
         13748 => x"7826d438",
         13749 => x"fdf53982",
         13750 => x"59807c34",
         13751 => x"7884ba8c",
         13752 => x"0c80e43d",
         13753 => x"0d04f73d",
         13754 => x"0d7b7d58",
         13755 => x"55895674",
         13756 => x"802e9f38",
         13757 => x"74085473",
         13758 => x"802e9738",
         13759 => x"73335372",
         13760 => x"802e8f38",
         13761 => x"86142284",
         13762 => x"16225959",
         13763 => x"78782e83",
         13764 => x"a0388053",
         13765 => x"725a7553",
         13766 => x"7581c238",
         13767 => x"91153353",
         13768 => x"7281ba38",
         13769 => x"8c150856",
         13770 => x"76762681",
         13771 => x"b9389415",
         13772 => x"08548058",
         13773 => x"76782e81",
         13774 => x"cc38798a",
         13775 => x"11227089",
         13776 => x"2b525a56",
         13777 => x"73782e81",
         13778 => x"f7387552",
         13779 => x"ff1751fd",
         13780 => x"bad33f84",
         13781 => x"ba8c08ff",
         13782 => x"15775470",
         13783 => x"535553fd",
         13784 => x"bac33f84",
         13785 => x"ba8c0873",
         13786 => x"2681d538",
         13787 => x"75307406",
         13788 => x"7094170c",
         13789 => x"77713198",
         13790 => x"17085658",
         13791 => x"5973802e",
         13792 => x"82983875",
         13793 => x"772781d9",
         13794 => x"38767631",
         13795 => x"94160817",
         13796 => x"94170c90",
         13797 => x"16337081",
         13798 => x"2a810651",
         13799 => x"5a577880",
         13800 => x"2e81fe38",
         13801 => x"73527451",
         13802 => x"ff99f33f",
         13803 => x"84ba8c08",
         13804 => x"5484ba8c",
         13805 => x"08802e81",
         13806 => x"a33873ff",
         13807 => x"2e983881",
         13808 => x"742782b4",
         13809 => x"38795373",
         13810 => x"9c140827",
         13811 => x"82aa3873",
         13812 => x"98160cff",
         13813 => x"ae39810b",
         13814 => x"91163481",
         13815 => x"537284ba",
         13816 => x"8c0c8b3d",
         13817 => x"0d049015",
         13818 => x"3370812a",
         13819 => x"81065558",
         13820 => x"73febb38",
         13821 => x"75941608",
         13822 => x"55578058",
         13823 => x"76782e09",
         13824 => x"8106feb6",
         13825 => x"38779416",
         13826 => x"0c941508",
         13827 => x"54757427",
         13828 => x"9038738c",
         13829 => x"160c9015",
         13830 => x"3380c007",
         13831 => x"57769016",
         13832 => x"347383ff",
         13833 => x"06597880",
         13834 => x"2e8c389c",
         13835 => x"1508782e",
         13836 => x"8538779c",
         13837 => x"160c800b",
         13838 => x"84ba8c0c",
         13839 => x"8b3d0d04",
         13840 => x"800b9416",
         13841 => x"0c881508",
         13842 => x"5473802e",
         13843 => x"80fe3873",
         13844 => x"98160c73",
         13845 => x"802e80c2",
         13846 => x"38fea839",
         13847 => x"84ba8c08",
         13848 => x"57941508",
         13849 => x"1794160c",
         13850 => x"7683ff06",
         13851 => x"5675802e",
         13852 => x"a93879fe",
         13853 => x"159c1208",
         13854 => x"fe055a55",
         13855 => x"56737827",
         13856 => x"80f6388a",
         13857 => x"16227471",
         13858 => x"29b01808",
         13859 => x"0578892a",
         13860 => x"115a5a53",
         13861 => x"78802e80",
         13862 => x"df388c15",
         13863 => x"0856fee9",
         13864 => x"39735274",
         13865 => x"51ff89b7",
         13866 => x"3f84ba8c",
         13867 => x"0854fe8a",
         13868 => x"39811433",
         13869 => x"51ff82a2",
         13870 => x"3f84ba8c",
         13871 => x"08810653",
         13872 => x"72fccf38",
         13873 => x"72750854",
         13874 => x"56fcc939",
         13875 => x"73527451",
         13876 => x"ff97cb3f",
         13877 => x"84ba8c08",
         13878 => x"5484ba8c",
         13879 => x"08812e98",
         13880 => x"3884ba8c",
         13881 => x"08ff2efd",
         13882 => x"ed3884ba",
         13883 => x"8c088816",
         13884 => x"0c739816",
         13885 => x"0cfedc39",
         13886 => x"820b9116",
         13887 => x"34820b84",
         13888 => x"ba8c0c8b",
         13889 => x"3d0d04f6",
         13890 => x"3d0d7c56",
         13891 => x"89547580",
         13892 => x"2ea23880",
         13893 => x"538c3dfc",
         13894 => x"05528d3d",
         13895 => x"840551c5",
         13896 => x"9b3f84ba",
         13897 => x"8c085584",
         13898 => x"ba8c0880",
         13899 => x"2e8f3880",
         13900 => x"760c7454",
         13901 => x"7384ba8c",
         13902 => x"0c8c3d0d",
         13903 => x"047a760c",
         13904 => x"7d527551",
         13905 => x"ffb9973f",
         13906 => x"84ba8c08",
         13907 => x"5584ba8c",
         13908 => x"0880d138",
         13909 => x"ab163370",
         13910 => x"982b5959",
         13911 => x"807824af",
         13912 => x"38861633",
         13913 => x"70842a81",
         13914 => x"065b5479",
         13915 => x"802e80c5",
         13916 => x"389c1608",
         13917 => x"9b11339a",
         13918 => x"12337188",
         13919 => x"2b077d70",
         13920 => x"335d5d5a",
         13921 => x"55577883",
         13922 => x"2eb33877",
         13923 => x"88170c7a",
         13924 => x"58861822",
         13925 => x"84172374",
         13926 => x"527551ff",
         13927 => x"99b93f84",
         13928 => x"ba8c0855",
         13929 => x"74842e8d",
         13930 => x"3874802e",
         13931 => x"ff843880",
         13932 => x"760cfefe",
         13933 => x"39855580",
         13934 => x"760cfef6",
         13935 => x"39951733",
         13936 => x"94183371",
         13937 => x"982b7190",
         13938 => x"2b077a07",
         13939 => x"88190c5a",
         13940 => x"5affbc39",
         13941 => x"fa3d0d78",
         13942 => x"55895474",
         13943 => x"802e9e38",
         13944 => x"74085372",
         13945 => x"802e9638",
         13946 => x"72335271",
         13947 => x"802e8e38",
         13948 => x"86132284",
         13949 => x"16225752",
         13950 => x"71762e94",
         13951 => x"38805271",
         13952 => x"57738438",
         13953 => x"73750c73",
         13954 => x"84ba8c0c",
         13955 => x"883d0d04",
         13956 => x"81133351",
         13957 => x"feffc33f",
         13958 => x"84ba8c08",
         13959 => x"81065271",
         13960 => x"dc387175",
         13961 => x"085354d7",
         13962 => x"39f83d0d",
         13963 => x"7a7c5855",
         13964 => x"89567480",
         13965 => x"2e9f3874",
         13966 => x"08547380",
         13967 => x"2e973873",
         13968 => x"33537280",
         13969 => x"2e8f3886",
         13970 => x"14228416",
         13971 => x"22595372",
         13972 => x"782e8197",
         13973 => x"38805372",
         13974 => x"59755375",
         13975 => x"80c73876",
         13976 => x"802e80f3",
         13977 => x"38755274",
         13978 => x"51ff9dbd",
         13979 => x"3f84ba8c",
         13980 => x"085384ba",
         13981 => x"8c08842e",
         13982 => x"b53884ba",
         13983 => x"8c08a638",
         13984 => x"76527451",
         13985 => x"ffb2923f",
         13986 => x"72527451",
         13987 => x"ff99be3f",
         13988 => x"84ba8c08",
         13989 => x"84327030",
         13990 => x"7072079f",
         13991 => x"2c84ba8c",
         13992 => x"08065557",
         13993 => x"547284ba",
         13994 => x"8c0c8a3d",
         13995 => x"0d047577",
         13996 => x"53755253",
         13997 => x"ffb1e23f",
         13998 => x"72527451",
         13999 => x"ff998e3f",
         14000 => x"84ba8c08",
         14001 => x"84327030",
         14002 => x"7072079f",
         14003 => x"2c84ba8c",
         14004 => x"08065557",
         14005 => x"54cf3975",
         14006 => x"527451ff",
         14007 => x"96f93f84",
         14008 => x"ba8c0884",
         14009 => x"ba8c0c8a",
         14010 => x"3d0d0481",
         14011 => x"143351fe",
         14012 => x"fde83f84",
         14013 => x"ba8c0881",
         14014 => x"065372fe",
         14015 => x"d8387275",
         14016 => x"085456fe",
         14017 => x"d239ed3d",
         14018 => x"0d665780",
         14019 => x"53893d70",
         14020 => x"53973d52",
         14021 => x"56c1a53f",
         14022 => x"84ba8c08",
         14023 => x"5584ba8c",
         14024 => x"08802e8a",
         14025 => x"387484ba",
         14026 => x"8c0c953d",
         14027 => x"0d046552",
         14028 => x"7551ffb5",
         14029 => x"a93f84ba",
         14030 => x"8c085584",
         14031 => x"ba8c08e5",
         14032 => x"380280cb",
         14033 => x"05337098",
         14034 => x"2b555880",
         14035 => x"74249738",
         14036 => x"76802ed1",
         14037 => x"38765275",
         14038 => x"51ffb0bd",
         14039 => x"3f7484ba",
         14040 => x"8c0c953d",
         14041 => x"0d04860b",
         14042 => x"84ba8c0c",
         14043 => x"953d0d04",
         14044 => x"ed3d0d66",
         14045 => x"68565f80",
         14046 => x"53953dec",
         14047 => x"0552963d",
         14048 => x"51c0b93f",
         14049 => x"84ba8c08",
         14050 => x"5a84ba8c",
         14051 => x"089a387f",
         14052 => x"750c7408",
         14053 => x"9c1108fe",
         14054 => x"11941308",
         14055 => x"59575957",
         14056 => x"7575268d",
         14057 => x"38757f0c",
         14058 => x"7984ba8c",
         14059 => x"0c953d0d",
         14060 => x"0484ba8c",
         14061 => x"0877335a",
         14062 => x"5b78812e",
         14063 => x"82933877",
         14064 => x"a8180884",
         14065 => x"ba8c085a",
         14066 => x"5d597780",
         14067 => x"c1387b81",
         14068 => x"1d715c5d",
         14069 => x"56b41708",
         14070 => x"762e82ef",
         14071 => x"38831733",
         14072 => x"785f5d7c",
         14073 => x"818d3881",
         14074 => x"547553b8",
         14075 => x"17528117",
         14076 => x"3351fefc",
         14077 => x"b73f84ba",
         14078 => x"8c08802e",
         14079 => x"8538ff5a",
         14080 => x"815e79b4",
         14081 => x"180c7f7e",
         14082 => x"5b577d80",
         14083 => x"cc387633",
         14084 => x"5e7d822e",
         14085 => x"828d3877",
         14086 => x"17b80583",
         14087 => x"11338212",
         14088 => x"3371902b",
         14089 => x"71882b07",
         14090 => x"81143370",
         14091 => x"7207882b",
         14092 => x"75337180",
         14093 => x"fffffe80",
         14094 => x"06077030",
         14095 => x"70802563",
         14096 => x"05608405",
         14097 => x"83ff0662",
         14098 => x"ff054341",
         14099 => x"43535452",
         14100 => x"5358405e",
         14101 => x"5678fef2",
         14102 => x"387a7f0c",
         14103 => x"7a94180c",
         14104 => x"84173381",
         14105 => x"07587784",
         14106 => x"18347984",
         14107 => x"ba8c0c95",
         14108 => x"3d0d0481",
         14109 => x"54b41708",
         14110 => x"53b81770",
         14111 => x"53811833",
         14112 => x"525dfefc",
         14113 => x"a63f815e",
         14114 => x"84ba8c08",
         14115 => x"fef83884",
         14116 => x"ba8c0883",
         14117 => x"1834b417",
         14118 => x"08a81808",
         14119 => x"3184ba8c",
         14120 => x"085f5574",
         14121 => x"a0180827",
         14122 => x"febd3882",
         14123 => x"17335574",
         14124 => x"822e0981",
         14125 => x"06feb038",
         14126 => x"8154b417",
         14127 => x"08a01808",
         14128 => x"05537c52",
         14129 => x"81173351",
         14130 => x"fefbe03f",
         14131 => x"775efe97",
         14132 => x"39827742",
         14133 => x"923d5956",
         14134 => x"75527751",
         14135 => x"ff81803f",
         14136 => x"84ba8c08",
         14137 => x"ff2e80e8",
         14138 => x"3884ba8c",
         14139 => x"08812e80",
         14140 => x"f73884ba",
         14141 => x"8c083070",
         14142 => x"84ba8c08",
         14143 => x"0780257c",
         14144 => x"05811862",
         14145 => x"5a585c5c",
         14146 => x"9c170876",
         14147 => x"26ca387a",
         14148 => x"7f0c7a94",
         14149 => x"180c8417",
         14150 => x"33810758",
         14151 => x"77841834",
         14152 => x"fec83977",
         14153 => x"17b80581",
         14154 => x"11337133",
         14155 => x"71882b07",
         14156 => x"70307080",
         14157 => x"251f821d",
         14158 => x"83ff06ff",
         14159 => x"1f5f5d5f",
         14160 => x"595f5f55",
         14161 => x"78fd8338",
         14162 => x"fe8f3977",
         14163 => x"5afdbf39",
         14164 => x"8160585a",
         14165 => x"7a7f0c7a",
         14166 => x"94180c84",
         14167 => x"17338107",
         14168 => x"58778418",
         14169 => x"34fe8339",
         14170 => x"8260585a",
         14171 => x"e739f73d",
         14172 => x"0d7b5789",
         14173 => x"5676802e",
         14174 => x"9f387608",
         14175 => x"5574802e",
         14176 => x"97387433",
         14177 => x"5473802e",
         14178 => x"8f388615",
         14179 => x"22841822",
         14180 => x"59597878",
         14181 => x"2e81da38",
         14182 => x"8054735a",
         14183 => x"7580dc38",
         14184 => x"91173356",
         14185 => x"7580d438",
         14186 => x"90173370",
         14187 => x"812a8106",
         14188 => x"55588755",
         14189 => x"73802e80",
         14190 => x"c4389417",
         14191 => x"0854738c",
         14192 => x"180827b7",
         14193 => x"387381d5",
         14194 => x"38881708",
         14195 => x"77085754",
         14196 => x"81742788",
         14197 => x"389c1608",
         14198 => x"7426b338",
         14199 => x"8256800b",
         14200 => x"88180c94",
         14201 => x"17088c18",
         14202 => x"0c7780c0",
         14203 => x"07597890",
         14204 => x"18347580",
         14205 => x"2e853875",
         14206 => x"91183475",
         14207 => x"557484ba",
         14208 => x"8c0c8b3d",
         14209 => x"0d047854",
         14210 => x"78782780",
         14211 => x"ff387352",
         14212 => x"7651fefe",
         14213 => x"ca3f84ba",
         14214 => x"8c085984",
         14215 => x"ba8c0880",
         14216 => x"2e80e938",
         14217 => x"84ba8c08",
         14218 => x"812e82d8",
         14219 => x"3884ba8c",
         14220 => x"08ff2e82",
         14221 => x"e5388053",
         14222 => x"73527551",
         14223 => x"ff85813f",
         14224 => x"84ba8c08",
         14225 => x"82c8389c",
         14226 => x"1608fe11",
         14227 => x"94180857",
         14228 => x"55587474",
         14229 => x"27ffaf38",
         14230 => x"81159417",
         14231 => x"0c841633",
         14232 => x"81075473",
         14233 => x"84173478",
         14234 => x"54777926",
         14235 => x"ffa0389c",
         14236 => x"39811533",
         14237 => x"51fef6e2",
         14238 => x"3f84ba8c",
         14239 => x"08810654",
         14240 => x"73fe9538",
         14241 => x"73770855",
         14242 => x"56fe8f39",
         14243 => x"800b9018",
         14244 => x"33595473",
         14245 => x"56800b88",
         14246 => x"180cfec7",
         14247 => x"39981708",
         14248 => x"527651fe",
         14249 => x"fdb93f84",
         14250 => x"ba8c08ff",
         14251 => x"2e81c238",
         14252 => x"84ba8c08",
         14253 => x"812e81be",
         14254 => x"387581ae",
         14255 => x"38795884",
         14256 => x"ba8c089c",
         14257 => x"19082781",
         14258 => x"a13884ba",
         14259 => x"8c089818",
         14260 => x"08780858",
         14261 => x"5654810b",
         14262 => x"84ba8c08",
         14263 => x"2781a138",
         14264 => x"84ba8c08",
         14265 => x"9c170827",
         14266 => x"81963874",
         14267 => x"802e9738",
         14268 => x"ff537452",
         14269 => x"7551ff83",
         14270 => x"c73f84ba",
         14271 => x"8c085584",
         14272 => x"ba8c0880",
         14273 => x"e3387352",
         14274 => x"7651fefc",
         14275 => x"d23f84ba",
         14276 => x"8c085984",
         14277 => x"ba8c0880",
         14278 => x"2e80cb38",
         14279 => x"84ba8c08",
         14280 => x"812e80dc",
         14281 => x"3884ba8c",
         14282 => x"08ff2e80",
         14283 => x"fe388053",
         14284 => x"73527551",
         14285 => x"ff83893f",
         14286 => x"84ba8c08",
         14287 => x"80e6389c",
         14288 => x"1608fe11",
         14289 => x"94180857",
         14290 => x"55587474",
         14291 => x"27903881",
         14292 => x"1594170c",
         14293 => x"84163381",
         14294 => x"07547384",
         14295 => x"17347854",
         14296 => x"777926ff",
         14297 => x"a1388055",
         14298 => x"74569017",
         14299 => x"3358fcf3",
         14300 => x"398156fe",
         14301 => x"bb39820b",
         14302 => x"90183359",
         14303 => x"56fce439",
         14304 => x"8256e739",
         14305 => x"820b9018",
         14306 => x"335954fe",
         14307 => x"863984ba",
         14308 => x"8c089018",
         14309 => x"335954fd",
         14310 => x"fa39810b",
         14311 => x"90183359",
         14312 => x"54fdf039",
         14313 => x"84ba8c08",
         14314 => x"56c03981",
         14315 => x"56ffbb39",
         14316 => x"db3d0d82",
         14317 => x"53a73dff",
         14318 => x"9c0552a8",
         14319 => x"3d51ffb7",
         14320 => x"fb3f84ba",
         14321 => x"8c085684",
         14322 => x"ba8c0880",
         14323 => x"2e8a3875",
         14324 => x"84ba8c0c",
         14325 => x"a73d0d04",
         14326 => x"7d4ba83d",
         14327 => x"08529b3d",
         14328 => x"705259ff",
         14329 => x"abf83f84",
         14330 => x"ba8c0856",
         14331 => x"84ba8c08",
         14332 => x"de380281",
         14333 => x"93053370",
         14334 => x"852a8106",
         14335 => x"59578656",
         14336 => x"77cd3876",
         14337 => x"982b5b80",
         14338 => x"7b24c438",
         14339 => x"0280ee05",
         14340 => x"33708106",
         14341 => x"5d578756",
         14342 => x"7bffb438",
         14343 => x"7da33d08",
         14344 => x"9b11339a",
         14345 => x"12337188",
         14346 => x"2b077333",
         14347 => x"415e5c57",
         14348 => x"587c832e",
         14349 => x"80d53876",
         14350 => x"842a8106",
         14351 => x"5776802e",
         14352 => x"80ed3887",
         14353 => x"56981808",
         14354 => x"7b2eff83",
         14355 => x"38775f7a",
         14356 => x"4184ba8c",
         14357 => x"08528f3d",
         14358 => x"705255ff",
         14359 => x"8bf93f84",
         14360 => x"ba8c0856",
         14361 => x"84ba8c08",
         14362 => x"fee53884",
         14363 => x"ba8c0852",
         14364 => x"7451ff91",
         14365 => x"b43f84ba",
         14366 => x"8c085684",
         14367 => x"ba8c08a0",
         14368 => x"38870b84",
         14369 => x"ba8c0ca7",
         14370 => x"3d0d0495",
         14371 => x"16339417",
         14372 => x"3371982b",
         14373 => x"71902b07",
         14374 => x"7d075d5d",
         14375 => x"5dff9839",
         14376 => x"84ba8c08",
         14377 => x"842e8838",
         14378 => x"84ba8c08",
         14379 => x"fea13878",
         14380 => x"086fa83d",
         14381 => x"08575d57",
         14382 => x"74ff2e80",
         14383 => x"d3387452",
         14384 => x"7851ff8b",
         14385 => x"923f84ba",
         14386 => x"8c085684",
         14387 => x"ba8c0880",
         14388 => x"2ebe3875",
         14389 => x"30707707",
         14390 => x"8025565a",
         14391 => x"7a802e9a",
         14392 => x"3874802e",
         14393 => x"95387a79",
         14394 => x"08585581",
         14395 => x"7b278938",
         14396 => x"9c17087b",
         14397 => x"2681fd38",
         14398 => x"825675fd",
         14399 => x"d2387d51",
         14400 => x"fef5db3f",
         14401 => x"84ba8c08",
         14402 => x"84ba8c0c",
         14403 => x"a73d0d04",
         14404 => x"b8175d98",
         14405 => x"19085680",
         14406 => x"5ab41708",
         14407 => x"762e82b9",
         14408 => x"38831733",
         14409 => x"7a595574",
         14410 => x"7a2e0981",
         14411 => x"0680dd38",
         14412 => x"81547553",
         14413 => x"b8175281",
         14414 => x"173351fe",
         14415 => x"f1ee3f84",
         14416 => x"ba8c0880",
         14417 => x"2e8538ff",
         14418 => x"56815875",
         14419 => x"b4180c77",
         14420 => x"5677ab38",
         14421 => x"9c190858",
         14422 => x"e5783481",
         14423 => x"0b831834",
         14424 => x"9019087c",
         14425 => x"27feec38",
         14426 => x"80527851",
         14427 => x"ff8bde3f",
         14428 => x"84ba8c08",
         14429 => x"5684ba8c",
         14430 => x"08802eff",
         14431 => x"96387584",
         14432 => x"2e098106",
         14433 => x"fecd3882",
         14434 => x"56fec839",
         14435 => x"8154b417",
         14436 => x"08537c52",
         14437 => x"81173351",
         14438 => x"fef2903f",
         14439 => x"815884ba",
         14440 => x"8c087a2e",
         14441 => x"098106ff",
         14442 => x"a63884ba",
         14443 => x"8c088318",
         14444 => x"34b41708",
         14445 => x"a8180831",
         14446 => x"84ba8c08",
         14447 => x"595574a0",
         14448 => x"180827fe",
         14449 => x"eb388217",
         14450 => x"33557482",
         14451 => x"2e098106",
         14452 => x"fede3881",
         14453 => x"54b41708",
         14454 => x"a0180805",
         14455 => x"537c5281",
         14456 => x"173351fe",
         14457 => x"f1c53f79",
         14458 => x"58fec539",
         14459 => x"79557978",
         14460 => x"2780e138",
         14461 => x"74527851",
         14462 => x"fef6e43f",
         14463 => x"84ba8c08",
         14464 => x"5a84ba8c",
         14465 => x"08802e80",
         14466 => x"cb3884ba",
         14467 => x"8c08812e",
         14468 => x"fde63884",
         14469 => x"ba8c08ff",
         14470 => x"2e80cb38",
         14471 => x"80537452",
         14472 => x"7651fefd",
         14473 => x"9b3f84ba",
         14474 => x"8c08b338",
         14475 => x"9c1708fe",
         14476 => x"11941908",
         14477 => x"585c5875",
         14478 => x"7b27ffb0",
         14479 => x"38811694",
         14480 => x"180c8417",
         14481 => x"3381075c",
         14482 => x"7b841834",
         14483 => x"7955777a",
         14484 => x"26ffa138",
         14485 => x"8056fda2",
         14486 => x"397956fd",
         14487 => x"f73984ba",
         14488 => x"8c0856fd",
         14489 => x"95398156",
         14490 => x"fd9039e3",
         14491 => x"3d0d8253",
         14492 => x"9f3dffbc",
         14493 => x"0552a03d",
         14494 => x"51ffb2c0",
         14495 => x"3f84ba8c",
         14496 => x"085684ba",
         14497 => x"8c08802e",
         14498 => x"8a387584",
         14499 => x"ba8c0c9f",
         14500 => x"3d0d047d",
         14501 => x"436f5293",
         14502 => x"3d70525a",
         14503 => x"ffa6bf3f",
         14504 => x"84ba8c08",
         14505 => x"5684ba8c",
         14506 => x"088b3888",
         14507 => x"0b84ba8c",
         14508 => x"0c9f3d0d",
         14509 => x"0484ba8c",
         14510 => x"08842e09",
         14511 => x"8106cb38",
         14512 => x"0280f305",
         14513 => x"3370852a",
         14514 => x"81065658",
         14515 => x"865674ff",
         14516 => x"b9387d5f",
         14517 => x"74528f3d",
         14518 => x"70525dff",
         14519 => x"83c03f84",
         14520 => x"ba8c0875",
         14521 => x"575c84ba",
         14522 => x"8c088338",
         14523 => x"875684ba",
         14524 => x"8c08812e",
         14525 => x"80f93884",
         14526 => x"ba8c08ff",
         14527 => x"2e81cb38",
         14528 => x"7581c938",
         14529 => x"7d84ba8c",
         14530 => x"08831233",
         14531 => x"5d5a577a",
         14532 => x"80e238fe",
         14533 => x"199c1808",
         14534 => x"fe055a56",
         14535 => x"805b7579",
         14536 => x"278d388a",
         14537 => x"17227671",
         14538 => x"29b01908",
         14539 => x"055c587a",
         14540 => x"b4180cb8",
         14541 => x"17598480",
         14542 => x"79575580",
         14543 => x"76708105",
         14544 => x"5834ff15",
         14545 => x"5574f438",
         14546 => x"74588a17",
         14547 => x"22557775",
         14548 => x"2781f938",
         14549 => x"8154771b",
         14550 => x"53785281",
         14551 => x"173351fe",
         14552 => x"eec93f84",
         14553 => x"ba8c0881",
         14554 => x"df388118",
         14555 => x"58dc3982",
         14556 => x"56ff8439",
         14557 => x"8154b417",
         14558 => x"0853b817",
         14559 => x"70538118",
         14560 => x"335258fe",
         14561 => x"eea53f81",
         14562 => x"5684ba8c",
         14563 => x"08be3884",
         14564 => x"ba8c0883",
         14565 => x"1834b417",
         14566 => x"08a81808",
         14567 => x"315574a0",
         14568 => x"180827fe",
         14569 => x"ee388217",
         14570 => x"335b7a82",
         14571 => x"2e098106",
         14572 => x"fee13875",
         14573 => x"54b41708",
         14574 => x"a0180805",
         14575 => x"53775281",
         14576 => x"173351fe",
         14577 => x"ede53ffe",
         14578 => x"ca398156",
         14579 => x"7b7d0858",
         14580 => x"55817c27",
         14581 => x"fdb4387b",
         14582 => x"9c180827",
         14583 => x"fdac3874",
         14584 => x"527c51fe",
         14585 => x"f2f93f84",
         14586 => x"ba8c085a",
         14587 => x"84ba8c08",
         14588 => x"802efd96",
         14589 => x"3884ba8c",
         14590 => x"08812efd",
         14591 => x"8d3884ba",
         14592 => x"8c08ff2e",
         14593 => x"fd843880",
         14594 => x"53745276",
         14595 => x"51fef9b0",
         14596 => x"3f84ba8c",
         14597 => x"08fcf338",
         14598 => x"9c1708fe",
         14599 => x"11941908",
         14600 => x"5a5c5977",
         14601 => x"7b279038",
         14602 => x"81189418",
         14603 => x"0c841733",
         14604 => x"81075c7b",
         14605 => x"84183479",
         14606 => x"55787a26",
         14607 => x"ffa13875",
         14608 => x"84ba8c0c",
         14609 => x"9f3d0d04",
         14610 => x"8a172255",
         14611 => x"7483ffff",
         14612 => x"06578156",
         14613 => x"76782e09",
         14614 => x"8106fef0",
         14615 => x"388b0bb8",
         14616 => x"1f5656a0",
         14617 => x"75708105",
         14618 => x"5734ff16",
         14619 => x"5675f438",
         14620 => x"7d57ae0b",
         14621 => x"b818347d",
         14622 => x"58900b80",
         14623 => x"c319347d",
         14624 => x"597580ce",
         14625 => x"1a347580",
         14626 => x"cf1a34a1",
         14627 => x"0b80d01a",
         14628 => x"3480cc0b",
         14629 => x"80d11a34",
         14630 => x"7d7c83ff",
         14631 => x"ff065956",
         14632 => x"7780d217",
         14633 => x"3477882a",
         14634 => x"5b7a80d3",
         14635 => x"17347533",
         14636 => x"5574832e",
         14637 => x"81cc387d",
         14638 => x"59a00b80",
         14639 => x"d81ab81b",
         14640 => x"57585674",
         14641 => x"70810556",
         14642 => x"33777081",
         14643 => x"055934ff",
         14644 => x"165675ef",
         14645 => x"387d56ae",
         14646 => x"0b80d917",
         14647 => x"34647e71",
         14648 => x"83ffff06",
         14649 => x"5b575778",
         14650 => x"80f21734",
         14651 => x"78882a5b",
         14652 => x"7a80f317",
         14653 => x"34753355",
         14654 => x"74832e80",
         14655 => x"f0387d5b",
         14656 => x"810b831c",
         14657 => x"347951ff",
         14658 => x"92963f84",
         14659 => x"ba8c0856",
         14660 => x"84ba8c08",
         14661 => x"fdb63869",
         14662 => x"5684ba8c",
         14663 => x"08961734",
         14664 => x"84ba8c08",
         14665 => x"971734a1",
         14666 => x"0b981734",
         14667 => x"80cc0b99",
         14668 => x"17347d6a",
         14669 => x"585d779a",
         14670 => x"18347788",
         14671 => x"2a59789b",
         14672 => x"18347c33",
         14673 => x"5a79832e",
         14674 => x"80d93869",
         14675 => x"55900b8b",
         14676 => x"16347d57",
         14677 => x"810b8318",
         14678 => x"347d51fe",
         14679 => x"ed803f84",
         14680 => x"ba8c0856",
         14681 => x"7584ba8c",
         14682 => x"0c9f3d0d",
         14683 => x"0476902a",
         14684 => x"557480ec",
         14685 => x"17347488",
         14686 => x"2a577680",
         14687 => x"ed1734fe",
         14688 => x"fd397b90",
         14689 => x"2a5b7a80",
         14690 => x"cc17347a",
         14691 => x"882a5574",
         14692 => x"80cd1734",
         14693 => x"7d59a00b",
         14694 => x"80d81ab8",
         14695 => x"1b575856",
         14696 => x"fea1397b",
         14697 => x"902a5877",
         14698 => x"94183477",
         14699 => x"882a5c7b",
         14700 => x"95183469",
         14701 => x"55900b8b",
         14702 => x"16347d57",
         14703 => x"810b8318",
         14704 => x"347d51fe",
         14705 => x"ec983f84",
         14706 => x"ba8c0856",
         14707 => x"ff9639d1",
         14708 => x"3d0db33d",
         14709 => x"b43d0870",
         14710 => x"595b5f79",
         14711 => x"802e9b38",
         14712 => x"79708105",
         14713 => x"5b33709f",
         14714 => x"26565675",
         14715 => x"ba2e81b8",
         14716 => x"3874ed38",
         14717 => x"75ba2e81",
         14718 => x"af388253",
         14719 => x"b13dfefc",
         14720 => x"0552b23d",
         14721 => x"51ffabb4",
         14722 => x"3f84ba8c",
         14723 => x"085684ba",
         14724 => x"8c08802e",
         14725 => x"8a387584",
         14726 => x"ba8c0cb1",
         14727 => x"3d0d047f",
         14728 => x"a63d0cb2",
         14729 => x"3d0852a5",
         14730 => x"3d705259",
         14731 => x"ff9faf3f",
         14732 => x"84ba8c08",
         14733 => x"5684ba8c",
         14734 => x"08dc3802",
         14735 => x"81bb0533",
         14736 => x"81a0065d",
         14737 => x"86567cce",
         14738 => x"38a00b92",
         14739 => x"3dae3d08",
         14740 => x"58585575",
         14741 => x"70810557",
         14742 => x"33777081",
         14743 => x"055934ff",
         14744 => x"155574ef",
         14745 => x"38993d58",
         14746 => x"b0787a58",
         14747 => x"58557570",
         14748 => x"81055733",
         14749 => x"77708105",
         14750 => x"5934ff15",
         14751 => x"5574ef38",
         14752 => x"b33d0852",
         14753 => x"7751ff9e",
         14754 => x"d53f84ba",
         14755 => x"8c085684",
         14756 => x"ba8c0885",
         14757 => x"d8386aa8",
         14758 => x"3d082e81",
         14759 => x"cb38880b",
         14760 => x"84ba8c0c",
         14761 => x"b13d0d04",
         14762 => x"7633d011",
         14763 => x"7081ff06",
         14764 => x"57575874",
         14765 => x"89269138",
         14766 => x"82177881",
         14767 => x"ff06d005",
         14768 => x"5d59787a",
         14769 => x"2e80fa38",
         14770 => x"807f0883",
         14771 => x"e5fc7008",
         14772 => x"725d5e5f",
         14773 => x"5f5c7a70",
         14774 => x"81055c33",
         14775 => x"79708105",
         14776 => x"5b33ff9f",
         14777 => x"125a5856",
         14778 => x"77992689",
         14779 => x"38e01670",
         14780 => x"81ff0657",
         14781 => x"55ff9f17",
         14782 => x"58779926",
         14783 => x"8938e017",
         14784 => x"7081ff06",
         14785 => x"58557530",
         14786 => x"709f2a59",
         14787 => x"5575772e",
         14788 => x"09810685",
         14789 => x"3877ffbe",
         14790 => x"38787a32",
         14791 => x"70307072",
         14792 => x"079f2a7a",
         14793 => x"075d5855",
         14794 => x"7a802e95",
         14795 => x"38811c84",
         14796 => x"1e5e5c7b",
         14797 => x"8324fdc2",
         14798 => x"387c087e",
         14799 => x"5a5bff96",
         14800 => x"397b8324",
         14801 => x"fdb43879",
         14802 => x"7f0c8253",
         14803 => x"b13dfefc",
         14804 => x"0552b23d",
         14805 => x"51ffa8e4",
         14806 => x"3f84ba8c",
         14807 => x"085684ba",
         14808 => x"8c08fdb2",
         14809 => x"38fdb839",
         14810 => x"6caa3d08",
         14811 => x"2e098106",
         14812 => x"feac3877",
         14813 => x"51ff8da8",
         14814 => x"3f84ba8c",
         14815 => x"085684ba",
         14816 => x"8c08fd92",
         14817 => x"386f5893",
         14818 => x"0b8d1902",
         14819 => x"880580cd",
         14820 => x"0558565a",
         14821 => x"75708105",
         14822 => x"57337570",
         14823 => x"81055734",
         14824 => x"ff1a5a79",
         14825 => x"ef380280",
         14826 => x"cb05338b",
         14827 => x"19348b18",
         14828 => x"3370842a",
         14829 => x"81064056",
         14830 => x"7e893875",
         14831 => x"a0075776",
         14832 => x"8b19347f",
         14833 => x"5d810b83",
         14834 => x"1e348b18",
         14835 => x"3370842a",
         14836 => x"8106575c",
         14837 => x"75802e81",
         14838 => x"c538a73d",
         14839 => x"086b2e81",
         14840 => x"bd387f9b",
         14841 => x"19339a1a",
         14842 => x"3371882b",
         14843 => x"07723341",
         14844 => x"585c577d",
         14845 => x"832e82e0",
         14846 => x"38fe169c",
         14847 => x"1808fe05",
         14848 => x"5e56757d",
         14849 => x"2782c738",
         14850 => x"8a172276",
         14851 => x"7129b019",
         14852 => x"0805575e",
         14853 => x"75802e82",
         14854 => x"b538757a",
         14855 => x"5d58b417",
         14856 => x"08762eaa",
         14857 => x"38831733",
         14858 => x"5f7e83bc",
         14859 => x"38815475",
         14860 => x"53b81752",
         14861 => x"81173351",
         14862 => x"fee3f13f",
         14863 => x"84ba8c08",
         14864 => x"802e8538",
         14865 => x"ff58815c",
         14866 => x"77b4180c",
         14867 => x"7f577b80",
         14868 => x"d8185656",
         14869 => x"7bfbbf38",
         14870 => x"8115335a",
         14871 => x"79ae2e09",
         14872 => x"8106bb38",
         14873 => x"6a7083ff",
         14874 => x"ff065d56",
         14875 => x"7b80f218",
         14876 => x"347b882a",
         14877 => x"587780f3",
         14878 => x"18347633",
         14879 => x"5b7a832e",
         14880 => x"09810693",
         14881 => x"3875902a",
         14882 => x"5e7d80ec",
         14883 => x"18347d88",
         14884 => x"2a567580",
         14885 => x"ed18347f",
         14886 => x"57810b83",
         14887 => x"18347808",
         14888 => x"aa3d08b2",
         14889 => x"3d08575c",
         14890 => x"5674ff2e",
         14891 => x"95387452",
         14892 => x"7851fefb",
         14893 => x"a23f84ba",
         14894 => x"8c085584",
         14895 => x"ba8c0880",
         14896 => x"f538b816",
         14897 => x"5c981908",
         14898 => x"57805ab4",
         14899 => x"1608772e",
         14900 => x"b4388316",
         14901 => x"337a595f",
         14902 => x"7e7a2e09",
         14903 => x"810681a8",
         14904 => x"38815476",
         14905 => x"53b81652",
         14906 => x"81163351",
         14907 => x"fee2bd3f",
         14908 => x"84ba8c08",
         14909 => x"802e8538",
         14910 => x"ff578158",
         14911 => x"76b4170c",
         14912 => x"775577aa",
         14913 => x"389c1908",
         14914 => x"5ae57a34",
         14915 => x"810b8317",
         14916 => x"34901908",
         14917 => x"7b27a538",
         14918 => x"80527851",
         14919 => x"fefcae3f",
         14920 => x"84ba8c08",
         14921 => x"5584ba8c",
         14922 => x"08802eff",
         14923 => x"98388256",
         14924 => x"74842ef9",
         14925 => x"e1387456",
         14926 => x"74f9db38",
         14927 => x"7f51fee5",
         14928 => x"9d3f84ba",
         14929 => x"8c0884ba",
         14930 => x"8c0cb13d",
         14931 => x"0d04820b",
         14932 => x"84ba8c0c",
         14933 => x"b13d0d04",
         14934 => x"95183394",
         14935 => x"19337198",
         14936 => x"2b71902b",
         14937 => x"07780758",
         14938 => x"565cfd8d",
         14939 => x"3984ba8c",
         14940 => x"08842efb",
         14941 => x"fe3884ba",
         14942 => x"8c08802e",
         14943 => x"fea03875",
         14944 => x"84ba8c0c",
         14945 => x"b13d0d04",
         14946 => x"8154b416",
         14947 => x"08537b52",
         14948 => x"81163351",
         14949 => x"fee2943f",
         14950 => x"815884ba",
         14951 => x"8c087a2e",
         14952 => x"098106fe",
         14953 => x"db3884ba",
         14954 => x"8c088317",
         14955 => x"34b41608",
         14956 => x"a8170831",
         14957 => x"84ba8c08",
         14958 => x"595574a0",
         14959 => x"170827fe",
         14960 => x"a0388216",
         14961 => x"335d7c82",
         14962 => x"2e098106",
         14963 => x"fe933881",
         14964 => x"54b41608",
         14965 => x"a0170805",
         14966 => x"537b5281",
         14967 => x"163351fe",
         14968 => x"e1c93f79",
         14969 => x"58fdfa39",
         14970 => x"8154b417",
         14971 => x"0853b817",
         14972 => x"70538118",
         14973 => x"33525bfe",
         14974 => x"e1b13f81",
         14975 => x"5c84ba8c",
         14976 => x"08fcc938",
         14977 => x"84ba8c08",
         14978 => x"831834b4",
         14979 => x"1708a818",
         14980 => x"083184ba",
         14981 => x"8c085d55",
         14982 => x"74a01808",
         14983 => x"27fc8e38",
         14984 => x"8217335d",
         14985 => x"7c822e09",
         14986 => x"8106fc81",
         14987 => x"388154b4",
         14988 => x"1708a018",
         14989 => x"0805537a",
         14990 => x"52811733",
         14991 => x"51fee0eb",
         14992 => x"3f795cfb",
         14993 => x"e839ec3d",
         14994 => x"0d0280df",
         14995 => x"05330284",
         14996 => x"0580e305",
         14997 => x"33565782",
         14998 => x"53963dcc",
         14999 => x"0552973d",
         15000 => x"51ffa2d8",
         15001 => x"3f84ba8c",
         15002 => x"085684ba",
         15003 => x"8c08802e",
         15004 => x"8a387584",
         15005 => x"ba8c0c96",
         15006 => x"3d0d0478",
         15007 => x"5a665296",
         15008 => x"3dd00551",
         15009 => x"ff96d73f",
         15010 => x"84ba8c08",
         15011 => x"5684ba8c",
         15012 => x"08e03802",
         15013 => x"80cf0533",
         15014 => x"81a00654",
         15015 => x"865673d2",
         15016 => x"3874a706",
         15017 => x"6171098b",
         15018 => x"12337106",
         15019 => x"7a740607",
         15020 => x"51565755",
         15021 => x"738b1734",
         15022 => x"7855810b",
         15023 => x"83163478",
         15024 => x"51fee29a",
         15025 => x"3f84ba8c",
         15026 => x"0884ba8c",
         15027 => x"0c963d0d",
         15028 => x"04ec3d0d",
         15029 => x"67578253",
         15030 => x"963dcc05",
         15031 => x"52973d51",
         15032 => x"ffa1d93f",
         15033 => x"84ba8c08",
         15034 => x"5584ba8c",
         15035 => x"08802e8a",
         15036 => x"387484ba",
         15037 => x"8c0c963d",
         15038 => x"0d04785a",
         15039 => x"6652963d",
         15040 => x"d00551ff",
         15041 => x"95d83f84",
         15042 => x"ba8c0855",
         15043 => x"84ba8c08",
         15044 => x"e0380280",
         15045 => x"cf053381",
         15046 => x"a0065686",
         15047 => x"5575d238",
         15048 => x"60841822",
         15049 => x"86192271",
         15050 => x"902b0759",
         15051 => x"59567696",
         15052 => x"17347688",
         15053 => x"2a557497",
         15054 => x"17347690",
         15055 => x"2a587798",
         15056 => x"17347698",
         15057 => x"2a547399",
         15058 => x"17347857",
         15059 => x"810b8318",
         15060 => x"347851fe",
         15061 => x"e1883f84",
         15062 => x"ba8c0884",
         15063 => x"ba8c0c96",
         15064 => x"3d0d04e8",
         15065 => x"3d0d6b6d",
         15066 => x"5d5b8053",
         15067 => x"9a3dcc05",
         15068 => x"529b3d51",
         15069 => x"ffa0c53f",
         15070 => x"84ba8c08",
         15071 => x"84ba8c08",
         15072 => x"307084ba",
         15073 => x"8c080780",
         15074 => x"25515657",
         15075 => x"7a802e8b",
         15076 => x"38817076",
         15077 => x"065a5678",
         15078 => x"81a43876",
         15079 => x"30707807",
         15080 => x"8025565b",
         15081 => x"7b802e81",
         15082 => x"8c388170",
         15083 => x"76065a58",
         15084 => x"78802e81",
         15085 => x"80387ca4",
         15086 => x"11085856",
         15087 => x"805ab416",
         15088 => x"08772e82",
         15089 => x"f6388316",
         15090 => x"337a5a55",
         15091 => x"747a2e09",
         15092 => x"81068198",
         15093 => x"38815476",
         15094 => x"53b81652",
         15095 => x"81163351",
         15096 => x"fedcc93f",
         15097 => x"84ba8c08",
         15098 => x"802e8538",
         15099 => x"ff578159",
         15100 => x"76b4170c",
         15101 => x"785778bd",
         15102 => x"387c7033",
         15103 => x"565880c3",
         15104 => x"5674832e",
         15105 => x"8b3880e4",
         15106 => x"5674842e",
         15107 => x"8338a756",
         15108 => x"7518b805",
         15109 => x"83113382",
         15110 => x"12337190",
         15111 => x"2b71882b",
         15112 => x"07811433",
         15113 => x"70720788",
         15114 => x"2b753371",
         15115 => x"07620c5f",
         15116 => x"5d5e5759",
         15117 => x"567684ba",
         15118 => x"8c0c9a3d",
         15119 => x"0d047c5e",
         15120 => x"80408052",
         15121 => x"8e3d7052",
         15122 => x"55fef48b",
         15123 => x"3f84ba8c",
         15124 => x"085784ba",
         15125 => x"8c08802e",
         15126 => x"818d3876",
         15127 => x"842e0981",
         15128 => x"06feb838",
         15129 => x"807b3480",
         15130 => x"57feb039",
         15131 => x"7754b416",
         15132 => x"0853b816",
         15133 => x"70538117",
         15134 => x"33525bfe",
         15135 => x"dcad3f77",
         15136 => x"5984ba8c",
         15137 => x"087a2e09",
         15138 => x"8106fee8",
         15139 => x"3884ba8c",
         15140 => x"08831734",
         15141 => x"b41608a8",
         15142 => x"17083184",
         15143 => x"ba8c085a",
         15144 => x"5574a017",
         15145 => x"0827fead",
         15146 => x"38821633",
         15147 => x"5574822e",
         15148 => x"098106fe",
         15149 => x"a0387754",
         15150 => x"b41608a0",
         15151 => x"17080553",
         15152 => x"7a528116",
         15153 => x"3351fedb",
         15154 => x"e23f7959",
         15155 => x"81547653",
         15156 => x"b8165281",
         15157 => x"163351fe",
         15158 => x"dad23f84",
         15159 => x"ba8c0880",
         15160 => x"2efe8d38",
         15161 => x"fe863975",
         15162 => x"527451fe",
         15163 => x"f8bb3f84",
         15164 => x"ba8c0857",
         15165 => x"84ba8c08",
         15166 => x"fee13884",
         15167 => x"ba8c0884",
         15168 => x"ba8c0866",
         15169 => x"5c595979",
         15170 => x"1881197c",
         15171 => x"1b575956",
         15172 => x"75337534",
         15173 => x"8119598a",
         15174 => x"7827ec38",
         15175 => x"8b701c57",
         15176 => x"58807634",
         15177 => x"77802efc",
         15178 => x"f238ff18",
         15179 => x"7b117033",
         15180 => x"5c575879",
         15181 => x"a02eea38",
         15182 => x"fce13979",
         15183 => x"57fdba39",
         15184 => x"e13d0d82",
         15185 => x"53a13dff",
         15186 => x"b40552a2",
         15187 => x"3d51ff9c",
         15188 => x"eb3f84ba",
         15189 => x"8c085684",
         15190 => x"ba8c0882",
         15191 => x"a6388f3d",
         15192 => x"5d8b7d57",
         15193 => x"55a07670",
         15194 => x"81055834",
         15195 => x"ff155574",
         15196 => x"f43874a3",
         15197 => x"3d087033",
         15198 => x"7081ff06",
         15199 => x"5b58585a",
         15200 => x"9f782781",
         15201 => x"b738a23d",
         15202 => x"903d5c5c",
         15203 => x"7581ff06",
         15204 => x"81185755",
         15205 => x"7481f538",
         15206 => x"757c0c74",
         15207 => x"83ffff26",
         15208 => x"81ff3874",
         15209 => x"51a1953f",
         15210 => x"83b55284",
         15211 => x"ba8c0851",
         15212 => x"9fdc3f84",
         15213 => x"ba8c0883",
         15214 => x"ffff0657",
         15215 => x"76802e81",
         15216 => x"e03883e7",
         15217 => x"9c0b83e7",
         15218 => x"9c337081",
         15219 => x"ff065b56",
         15220 => x"5878802e",
         15221 => x"81d63874",
         15222 => x"5678772e",
         15223 => x"99388118",
         15224 => x"70337081",
         15225 => x"ff065757",
         15226 => x"5874802e",
         15227 => x"89387477",
         15228 => x"2e098106",
         15229 => x"e9387581",
         15230 => x"ff065978",
         15231 => x"81a33881",
         15232 => x"ff772781",
         15233 => x"f8387989",
         15234 => x"26819638",
         15235 => x"81ff7727",
         15236 => x"8f387688",
         15237 => x"2a55747b",
         15238 => x"7081055d",
         15239 => x"34811a5a",
         15240 => x"767b7081",
         15241 => x"055d3481",
         15242 => x"1aa33d08",
         15243 => x"70337081",
         15244 => x"ff065b58",
         15245 => x"585a779f",
         15246 => x"26fed138",
         15247 => x"8f3d3357",
         15248 => x"86567681",
         15249 => x"e52ebc38",
         15250 => x"79802e99",
         15251 => x"3802b705",
         15252 => x"56791670",
         15253 => x"335c5c7a",
         15254 => x"a02e0981",
         15255 => x"068738ff",
         15256 => x"1a5a79ed",
         15257 => x"387d4580",
         15258 => x"47805295",
         15259 => x"3d705256",
         15260 => x"feefe43f",
         15261 => x"84ba8c08",
         15262 => x"5584ba8c",
         15263 => x"08802eb4",
         15264 => x"38745675",
         15265 => x"84ba8c0c",
         15266 => x"a13d0d04",
         15267 => x"83b55274",
         15268 => x"519ee73f",
         15269 => x"84ba8c08",
         15270 => x"83ffff06",
         15271 => x"5574fdf8",
         15272 => x"38865675",
         15273 => x"84ba8c0c",
         15274 => x"a13d0d04",
         15275 => x"83e79c33",
         15276 => x"56fec339",
         15277 => x"81527551",
         15278 => x"fef4ee3f",
         15279 => x"84ba8c08",
         15280 => x"5584ba8c",
         15281 => x"0880c138",
         15282 => x"79802e82",
         15283 => x"c4388b6c",
         15284 => x"7e595755",
         15285 => x"76708105",
         15286 => x"58337670",
         15287 => x"81055834",
         15288 => x"ff155574",
         15289 => x"ef387d5d",
         15290 => x"810b831e",
         15291 => x"347d51fe",
         15292 => x"d9ec3f84",
         15293 => x"ba8c0855",
         15294 => x"7456ff87",
         15295 => x"398a7a27",
         15296 => x"fe8a3886",
         15297 => x"56ff9c39",
         15298 => x"84ba8c08",
         15299 => x"842e0981",
         15300 => x"06feee38",
         15301 => x"80557975",
         15302 => x"2efee638",
         15303 => x"75087553",
         15304 => x"765258fe",
         15305 => x"eeb13f84",
         15306 => x"ba8c0857",
         15307 => x"84ba8c08",
         15308 => x"752e0981",
         15309 => x"06818438",
         15310 => x"84ba8c08",
         15311 => x"b8195c5a",
         15312 => x"98160857",
         15313 => x"8059b418",
         15314 => x"08772eb2",
         15315 => x"38831833",
         15316 => x"5574792e",
         15317 => x"09810681",
         15318 => x"d7388154",
         15319 => x"7653b818",
         15320 => x"52811833",
         15321 => x"51fed5c4",
         15322 => x"3f84ba8c",
         15323 => x"08802e85",
         15324 => x"38ff5781",
         15325 => x"5976b419",
         15326 => x"0c785778",
         15327 => x"be38789c",
         15328 => x"17087033",
         15329 => x"575a5774",
         15330 => x"81e52e81",
         15331 => x"9e387430",
         15332 => x"70802578",
         15333 => x"07565c74",
         15334 => x"802e81d7",
         15335 => x"38811a5a",
         15336 => x"79812ea5",
         15337 => x"38815275",
         15338 => x"51feefa1",
         15339 => x"3f84ba8c",
         15340 => x"085784ba",
         15341 => x"8c08802e",
         15342 => x"ff863887",
         15343 => x"5576842e",
         15344 => x"fdbf3876",
         15345 => x"5576fdb9",
         15346 => x"38a06c57",
         15347 => x"55807670",
         15348 => x"81055834",
         15349 => x"ff155574",
         15350 => x"f4386b56",
         15351 => x"880b8b17",
         15352 => x"348b6c7e",
         15353 => x"59575576",
         15354 => x"70810558",
         15355 => x"33767081",
         15356 => x"055834ff",
         15357 => x"15557480",
         15358 => x"2efdeb38",
         15359 => x"76708105",
         15360 => x"58337670",
         15361 => x"81055834",
         15362 => x"ff155574",
         15363 => x"da38fdd6",
         15364 => x"396b5ae5",
         15365 => x"7a347d5d",
         15366 => x"810b831e",
         15367 => x"347d51fe",
         15368 => x"d7bc3f84",
         15369 => x"ba8c0855",
         15370 => x"fdce3981",
         15371 => x"57fedf39",
         15372 => x"8154b418",
         15373 => x"08537a52",
         15374 => x"81183351",
         15375 => x"fed4ec3f",
         15376 => x"84ba8c08",
         15377 => x"792e0981",
         15378 => x"0680c338",
         15379 => x"84ba8c08",
         15380 => x"831934b4",
         15381 => x"1808a819",
         15382 => x"08315c7b",
         15383 => x"a0190827",
         15384 => x"8a388218",
         15385 => x"33557482",
         15386 => x"2eb13884",
         15387 => x"ba8c0859",
         15388 => x"fde83974",
         15389 => x"5a815275",
         15390 => x"51feedd1",
         15391 => x"3f84ba8c",
         15392 => x"085784ba",
         15393 => x"8c08802e",
         15394 => x"fdb638fe",
         15395 => x"ae398170",
         15396 => x"58597880",
         15397 => x"2efde738",
         15398 => x"fea13981",
         15399 => x"54b41808",
         15400 => x"a0190805",
         15401 => x"537a5281",
         15402 => x"183351fe",
         15403 => x"d3fd3ffd",
         15404 => x"a939f23d",
         15405 => x"0d606202",
         15406 => x"880580cb",
         15407 => x"05335e5b",
         15408 => x"57895676",
         15409 => x"802e9f38",
         15410 => x"76085574",
         15411 => x"802e9738",
         15412 => x"74335473",
         15413 => x"802e8f38",
         15414 => x"86152284",
         15415 => x"18225959",
         15416 => x"78782e81",
         15417 => x"c2388054",
         15418 => x"735f7581",
         15419 => x"a5389117",
         15420 => x"33567581",
         15421 => x"9d387980",
         15422 => x"2e81a238",
         15423 => x"8c170881",
         15424 => x"9c389017",
         15425 => x"3370812a",
         15426 => x"8106565d",
         15427 => x"74802e81",
         15428 => x"8c387e8a",
         15429 => x"11227089",
         15430 => x"2b70557c",
         15431 => x"54575c59",
         15432 => x"fd87823f",
         15433 => x"ff157a06",
         15434 => x"70307072",
         15435 => x"079f2a84",
         15436 => x"ba8c0805",
         15437 => x"901c0879",
         15438 => x"42535f55",
         15439 => x"58817827",
         15440 => x"88389c19",
         15441 => x"08782683",
         15442 => x"38825877",
         15443 => x"78565b80",
         15444 => x"59745276",
         15445 => x"51fed887",
         15446 => x"3f81157f",
         15447 => x"55559c14",
         15448 => x"08752683",
         15449 => x"38825584",
         15450 => x"ba8c0881",
         15451 => x"2e81dc38",
         15452 => x"84ba8c08",
         15453 => x"ff2e81d8",
         15454 => x"3884ba8c",
         15455 => x"0881c538",
         15456 => x"81195978",
         15457 => x"7d2ebb38",
         15458 => x"74782e09",
         15459 => x"8106c238",
         15460 => x"87567554",
         15461 => x"7384ba8c",
         15462 => x"0c903d0d",
         15463 => x"04870b84",
         15464 => x"ba8c0c90",
         15465 => x"3d0d0481",
         15466 => x"153351fe",
         15467 => x"d0ac3f84",
         15468 => x"ba8c0881",
         15469 => x"065473fe",
         15470 => x"ad387377",
         15471 => x"085556fe",
         15472 => x"a7397b80",
         15473 => x"2e818e38",
         15474 => x"7a7d5658",
         15475 => x"7c802eab",
         15476 => x"38811854",
         15477 => x"74812e80",
         15478 => x"e6387353",
         15479 => x"77527e51",
         15480 => x"fedddd3f",
         15481 => x"84ba8c08",
         15482 => x"5684ba8c",
         15483 => x"08ffa338",
         15484 => x"778119ff",
         15485 => x"1757595e",
         15486 => x"74d7387e",
         15487 => x"7e90120c",
         15488 => x"557b802e",
         15489 => x"ff8c387a",
         15490 => x"88180c79",
         15491 => x"8c180c90",
         15492 => x"173380c0",
         15493 => x"075c7b90",
         15494 => x"18349c15",
         15495 => x"08fe0594",
         15496 => x"1608585a",
         15497 => x"767a26fe",
         15498 => x"e938767d",
         15499 => x"3194160c",
         15500 => x"84153381",
         15501 => x"075d7c84",
         15502 => x"16347554",
         15503 => x"fed639ff",
         15504 => x"54ff9739",
         15505 => x"745b8059",
         15506 => x"febe3982",
         15507 => x"54fec539",
         15508 => x"8154fec0",
         15509 => x"39ff1b5e",
         15510 => x"ffa13984",
         15511 => x"ba9808e3",
         15512 => x"3d0da33d",
         15513 => x"08a53d08",
         15514 => x"02880581",
         15515 => x"87053344",
         15516 => x"425fff0b",
         15517 => x"a23d0870",
         15518 => x"5f5b4079",
         15519 => x"802e858a",
         15520 => x"38797081",
         15521 => x"055b3370",
         15522 => x"9f265656",
         15523 => x"75ba2e85",
         15524 => x"9b3874ed",
         15525 => x"3875ba2e",
         15526 => x"85923884",
         15527 => x"d1e83356",
         15528 => x"80762484",
         15529 => x"e5387510",
         15530 => x"1084d1d4",
         15531 => x"05700856",
         15532 => x"5a74802e",
         15533 => x"84388075",
         15534 => x"34751684",
         15535 => x"ba801133",
         15536 => x"84ba8112",
         15537 => x"33405b5d",
         15538 => x"81527951",
         15539 => x"fecea93f",
         15540 => x"84ba8c08",
         15541 => x"81ff0670",
         15542 => x"81065d56",
         15543 => x"83577b84",
         15544 => x"ab387582",
         15545 => x"2a810640",
         15546 => x"8a577f84",
         15547 => x"9f389f3d",
         15548 => x"fc055383",
         15549 => x"527951fe",
         15550 => x"d0b03f84",
         15551 => x"ba8c0884",
         15552 => x"98386d55",
         15553 => x"74802e84",
         15554 => x"90387482",
         15555 => x"80802684",
         15556 => x"8838ff15",
         15557 => x"75065574",
         15558 => x"83ff387e",
         15559 => x"802e8838",
         15560 => x"84807f26",
         15561 => x"83f8387e",
         15562 => x"81800a26",
         15563 => x"83f038ff",
         15564 => x"1f7f0655",
         15565 => x"7483e738",
         15566 => x"7e892aa6",
         15567 => x"3d08892a",
         15568 => x"70892b77",
         15569 => x"594c475b",
         15570 => x"60802e85",
         15571 => x"ab386530",
         15572 => x"70802577",
         15573 => x"07565f91",
         15574 => x"577483b0",
         15575 => x"387d802e",
         15576 => x"84df3881",
         15577 => x"54745360",
         15578 => x"527951fe",
         15579 => x"cdbe3f81",
         15580 => x"5784ba8c",
         15581 => x"08839538",
         15582 => x"6083ff05",
         15583 => x"336183fe",
         15584 => x"05337188",
         15585 => x"2b075956",
         15586 => x"8e577782",
         15587 => x"d4d52e09",
         15588 => x"810682f8",
         15589 => x"387d9029",
         15590 => x"610583b2",
         15591 => x"11334458",
         15592 => x"62802e82",
         15593 => x"e73883b6",
         15594 => x"18831133",
         15595 => x"82123371",
         15596 => x"902b7188",
         15597 => x"2b078114",
         15598 => x"33707207",
         15599 => x"882b7533",
         15600 => x"710783ba",
         15601 => x"1f831133",
         15602 => x"82123371",
         15603 => x"902b7188",
         15604 => x"2b078114",
         15605 => x"33707207",
         15606 => x"882b7533",
         15607 => x"71075ca2",
         15608 => x"3d0c42a3",
         15609 => x"3d0ca33d",
         15610 => x"0c444e54",
         15611 => x"45594f41",
         15612 => x"5a4b784d",
         15613 => x"8e5780ff",
         15614 => x"79278290",
         15615 => x"3893577a",
         15616 => x"81802682",
         15617 => x"87386181",
         15618 => x"2a708106",
         15619 => x"45496380",
         15620 => x"2e83f938",
         15621 => x"61870645",
         15622 => x"64822e89",
         15623 => x"38618106",
         15624 => x"476683f4",
         15625 => x"38836e70",
         15626 => x"304a4643",
         15627 => x"7a586283",
         15628 => x"2e8ac238",
         15629 => x"7aae3878",
         15630 => x"8c2a5781",
         15631 => x"0b83e7b0",
         15632 => x"22565874",
         15633 => x"802e9d38",
         15634 => x"74772698",
         15635 => x"3883e7b0",
         15636 => x"56771082",
         15637 => x"17702257",
         15638 => x"57587480",
         15639 => x"2e863876",
         15640 => x"7527ee38",
         15641 => x"77527851",
         15642 => x"fd80ba3f",
         15643 => x"84ba8c08",
         15644 => x"10840555",
         15645 => x"84ba8c08",
         15646 => x"9ff52696",
         15647 => x"38810b84",
         15648 => x"ba8c0810",
         15649 => x"84ba8c08",
         15650 => x"05711172",
         15651 => x"2a830557",
         15652 => x"4c4383ff",
         15653 => x"15892a5d",
         15654 => x"815ca047",
         15655 => x"7b1f7d11",
         15656 => x"68056611",
         15657 => x"ff05706b",
         15658 => x"06723158",
         15659 => x"4e574462",
         15660 => x"832e89b8",
         15661 => x"38741d5d",
         15662 => x"77902916",
         15663 => x"70603156",
         15664 => x"57747926",
         15665 => x"82f23878",
         15666 => x"7c317d31",
         15667 => x"78537068",
         15668 => x"315256fc",
         15669 => x"ffcf3f84",
         15670 => x"ba8c0840",
         15671 => x"62832e89",
         15672 => x"f6386282",
         15673 => x"2e098106",
         15674 => x"82dd3883",
         15675 => x"fff50b84",
         15676 => x"ba8c0827",
         15677 => x"82ac387a",
         15678 => x"89f93877",
         15679 => x"18557480",
         15680 => x"c02689ef",
         15681 => x"38745bfe",
         15682 => x"a3398b57",
         15683 => x"7684ba8c",
         15684 => x"0c9f3d0d",
         15685 => x"84ba980c",
         15686 => x"04814efb",
         15687 => x"fe39930b",
         15688 => x"84ba8c0c",
         15689 => x"9f3d0d84",
         15690 => x"ba980c04",
         15691 => x"7c33d011",
         15692 => x"7081ff06",
         15693 => x"57575774",
         15694 => x"89269138",
         15695 => x"821d7781",
         15696 => x"ff06d005",
         15697 => x"5d58777a",
         15698 => x"2e81b238",
         15699 => x"800b83e5",
         15700 => x"fc5f5c7d",
         15701 => x"087d575b",
         15702 => x"7a708105",
         15703 => x"5c337670",
         15704 => x"81055833",
         15705 => x"ff9f1245",
         15706 => x"59576299",
         15707 => x"268938e0",
         15708 => x"177081ff",
         15709 => x"065844ff",
         15710 => x"9f184564",
         15711 => x"99268938",
         15712 => x"e0187081",
         15713 => x"ff065946",
         15714 => x"7630709f",
         15715 => x"2a5a4776",
         15716 => x"782e0981",
         15717 => x"06853878",
         15718 => x"ffbe3875",
         15719 => x"7a327030",
         15720 => x"7072079f",
         15721 => x"2a7b075d",
         15722 => x"4a4a7a80",
         15723 => x"2e80ce38",
         15724 => x"811c841f",
         15725 => x"5f5c837c",
         15726 => x"25ff9838",
         15727 => x"7f56f9e0",
         15728 => x"399f3df8",
         15729 => x"05538152",
         15730 => x"7951feca",
         15731 => x"dd3f8157",
         15732 => x"84ba8c08",
         15733 => x"feb63861",
         15734 => x"832a7706",
         15735 => x"84ba8c08",
         15736 => x"40567583",
         15737 => x"38bf5f6c",
         15738 => x"558e577e",
         15739 => x"7526fe9c",
         15740 => x"38747f31",
         15741 => x"59fbfb39",
         15742 => x"8156fad2",
         15743 => x"397b8324",
         15744 => x"ffba387b",
         15745 => x"7aa33d0c",
         15746 => x"56f99539",
         15747 => x"61810648",
         15748 => x"93576780",
         15749 => x"2efdf538",
         15750 => x"826e7030",
         15751 => x"4a4643fc",
         15752 => x"8b3984ba",
         15753 => x"8c089ff5",
         15754 => x"269d387a",
         15755 => x"8b387718",
         15756 => x"5b81807b",
         15757 => x"27fbf538",
         15758 => x"8e577684",
         15759 => x"ba8c0c9f",
         15760 => x"3d0d84ba",
         15761 => x"980c0480",
         15762 => x"5562812e",
         15763 => x"8699389f",
         15764 => x"f560278b",
         15765 => x"38748106",
         15766 => x"5b8e577a",
         15767 => x"fdae3884",
         15768 => x"80615755",
         15769 => x"80767081",
         15770 => x"055834ff",
         15771 => x"155574f4",
         15772 => x"388b6183",
         15773 => x"e5c85957",
         15774 => x"55767081",
         15775 => x"05583376",
         15776 => x"70810558",
         15777 => x"34ff1555",
         15778 => x"74ef3860",
         15779 => x"8b054574",
         15780 => x"65348261",
         15781 => x"8c053477",
         15782 => x"618d0534",
         15783 => x"7b83ffff",
         15784 => x"064b6a61",
         15785 => x"8e05346a",
         15786 => x"882a5c7b",
         15787 => x"618f0534",
         15788 => x"81619005",
         15789 => x"34628332",
         15790 => x"70305a48",
         15791 => x"80619105",
         15792 => x"34789e2a",
         15793 => x"82064968",
         15794 => x"61920534",
         15795 => x"6c567583",
         15796 => x"ffff2686",
         15797 => x"ad387583",
         15798 => x"ffff0655",
         15799 => x"74619305",
         15800 => x"3474882a",
         15801 => x"4c6b6194",
         15802 => x"0534f861",
         15803 => x"950534bf",
         15804 => x"61980534",
         15805 => x"80619905",
         15806 => x"34ff619a",
         15807 => x"05348061",
         15808 => x"9b05347e",
         15809 => x"619c0534",
         15810 => x"7e882a48",
         15811 => x"67619d05",
         15812 => x"347e902a",
         15813 => x"4c6b619e",
         15814 => x"05347e98",
         15815 => x"2a84ba98",
         15816 => x"0c84ba98",
         15817 => x"08619f05",
         15818 => x"3462832e",
         15819 => x"85f73880",
         15820 => x"61a70534",
         15821 => x"8061a805",
         15822 => x"34a161a9",
         15823 => x"053480cc",
         15824 => x"61aa0534",
         15825 => x"7c83ffff",
         15826 => x"06557461",
         15827 => x"96053474",
         15828 => x"882a4b6a",
         15829 => x"61970534",
         15830 => x"ff8061a4",
         15831 => x"0534a961",
         15832 => x"a6053493",
         15833 => x"61ab0583",
         15834 => x"e5d45957",
         15835 => x"55767081",
         15836 => x"05583376",
         15837 => x"70810558",
         15838 => x"34ff1555",
         15839 => x"74ef3860",
         15840 => x"83fe0549",
         15841 => x"80d56934",
         15842 => x"6083ff05",
         15843 => x"4bffaa6b",
         15844 => x"3481547e",
         15845 => x"53605279",
         15846 => x"51fec68f",
         15847 => x"3f815784",
         15848 => x"ba8c08fa",
         15849 => x"e7386017",
         15850 => x"5c62832e",
         15851 => x"879c3869",
         15852 => x"61575580",
         15853 => x"76708105",
         15854 => x"5834ff15",
         15855 => x"5574f438",
         15856 => x"6375415b",
         15857 => x"62832e86",
         15858 => x"c03887ff",
         15859 => x"fff85762",
         15860 => x"812e8338",
         15861 => x"f8577661",
         15862 => x"3476882a",
         15863 => x"7c455574",
         15864 => x"64708105",
         15865 => x"46347690",
         15866 => x"2a597864",
         15867 => x"70810546",
         15868 => x"3476982a",
         15869 => x"56756434",
         15870 => x"7c576559",
         15871 => x"76662683",
         15872 => x"38765978",
         15873 => x"547a5360",
         15874 => x"527951fe",
         15875 => x"c59d3f84",
         15876 => x"ba8c0885",
         15877 => x"e6388480",
         15878 => x"61575580",
         15879 => x"76708105",
         15880 => x"5834ff15",
         15881 => x"5574f438",
         15882 => x"781b777a",
         15883 => x"31585b76",
         15884 => x"c9387f81",
         15885 => x"05407f80",
         15886 => x"2eff8938",
         15887 => x"77566283",
         15888 => x"2e833866",
         15889 => x"56655575",
         15890 => x"66268338",
         15891 => x"75557454",
         15892 => x"7a536052",
         15893 => x"7951fec4",
         15894 => x"d23f84ba",
         15895 => x"8c08859b",
         15896 => x"38741b76",
         15897 => x"7631575b",
         15898 => x"75db388c",
         15899 => x"5862832e",
         15900 => x"93388658",
         15901 => x"6c83ffff",
         15902 => x"268a3884",
         15903 => x"5862822e",
         15904 => x"83388158",
         15905 => x"7d84c138",
         15906 => x"61832a81",
         15907 => x"065e7d81",
         15908 => x"b3388480",
         15909 => x"61565980",
         15910 => x"75708105",
         15911 => x"5734ff19",
         15912 => x"5978f438",
         15913 => x"80d56934",
         15914 => x"ffaa6b34",
         15915 => x"6083be05",
         15916 => x"47786734",
         15917 => x"81678105",
         15918 => x"34816782",
         15919 => x"05347867",
         15920 => x"83053477",
         15921 => x"67840534",
         15922 => x"6c4380fd",
         15923 => x"c152621f",
         15924 => x"51fcf7d1",
         15925 => x"3ffe6785",
         15926 => x"053484ba",
         15927 => x"8c08822a",
         15928 => x"bf075776",
         15929 => x"67860534",
         15930 => x"84ba8c08",
         15931 => x"67870534",
         15932 => x"7e6183c6",
         15933 => x"05346761",
         15934 => x"83c70534",
         15935 => x"6b6183c8",
         15936 => x"053484ba",
         15937 => x"98086183",
         15938 => x"c9053462",
         15939 => x"6183ca05",
         15940 => x"3462882a",
         15941 => x"45646183",
         15942 => x"cb053462",
         15943 => x"902a5877",
         15944 => x"6183cc05",
         15945 => x"3462982a",
         15946 => x"5f7e6183",
         15947 => x"cd053481",
         15948 => x"54785360",
         15949 => x"527951fe",
         15950 => x"c2f13f81",
         15951 => x"5784ba8c",
         15952 => x"08f7c938",
         15953 => x"80538052",
         15954 => x"7951fec3",
         15955 => x"dd3f8157",
         15956 => x"84ba8c08",
         15957 => x"f7b63884",
         15958 => x"ba8c0884",
         15959 => x"ba8c0c9f",
         15960 => x"3d0d84ba",
         15961 => x"980c0462",
         15962 => x"55f9e439",
         15963 => x"741c6416",
         15964 => x"455cf6c4",
         15965 => x"397aae38",
         15966 => x"78912a57",
         15967 => x"810b83e7",
         15968 => x"c0225658",
         15969 => x"74802e9d",
         15970 => x"38747726",
         15971 => x"983883e7",
         15972 => x"c0567710",
         15973 => x"82177022",
         15974 => x"57575874",
         15975 => x"802e8638",
         15976 => x"767527ee",
         15977 => x"38775278",
         15978 => x"51fcf5f9",
         15979 => x"3f84ba8c",
         15980 => x"08101084",
         15981 => x"87057089",
         15982 => x"2a5e5ca0",
         15983 => x"5c800b84",
         15984 => x"ba8c08fc",
         15985 => x"808a0558",
         15986 => x"47fdfff0",
         15987 => x"0a7727f5",
         15988 => x"cb388e57",
         15989 => x"f8e43984",
         15990 => x"ba8c0883",
         15991 => x"fff526f8",
         15992 => x"e6387af8",
         15993 => x"d3387781",
         15994 => x"2a5b7af4",
         15995 => x"bf388e57",
         15996 => x"f8c83968",
         15997 => x"81064463",
         15998 => x"802ef8af",
         15999 => x"388343f4",
         16000 => x"ab397561",
         16001 => x"a0053475",
         16002 => x"882a4968",
         16003 => x"61a10534",
         16004 => x"75902a5b",
         16005 => x"7a61a205",
         16006 => x"3475982a",
         16007 => x"577661a3",
         16008 => x"0534f9c6",
         16009 => x"39806180",
         16010 => x"c3053480",
         16011 => x"6180c405",
         16012 => x"34a16180",
         16013 => x"c5053480",
         16014 => x"cc6180c6",
         16015 => x"05347c61",
         16016 => x"a405347c",
         16017 => x"882a5c7b",
         16018 => x"61a50534",
         16019 => x"7c902a59",
         16020 => x"7861a605",
         16021 => x"347c982a",
         16022 => x"567561a7",
         16023 => x"05348261",
         16024 => x"ac053480",
         16025 => x"61ad0534",
         16026 => x"8061ae05",
         16027 => x"348061af",
         16028 => x"05348161",
         16029 => x"b0053480",
         16030 => x"61b10534",
         16031 => x"8661b205",
         16032 => x"348061b3",
         16033 => x"0534ff80",
         16034 => x"6180c005",
         16035 => x"34a96180",
         16036 => x"c2053493",
         16037 => x"6180c705",
         16038 => x"83e5e859",
         16039 => x"57557670",
         16040 => x"81055833",
         16041 => x"76708105",
         16042 => x"5834ff15",
         16043 => x"5574802e",
         16044 => x"f9cd3876",
         16045 => x"70810558",
         16046 => x"33767081",
         16047 => x"055834ff",
         16048 => x"155574da",
         16049 => x"38f9b839",
         16050 => x"81548053",
         16051 => x"60527951",
         16052 => x"febed93f",
         16053 => x"815784ba",
         16054 => x"8c08f4b0",
         16055 => x"387d9029",
         16056 => x"61054277",
         16057 => x"6283b205",
         16058 => x"34765484",
         16059 => x"ba8c0853",
         16060 => x"60527951",
         16061 => x"febfb43f",
         16062 => x"fcc33981",
         16063 => x"0b84ba8c",
         16064 => x"0c9f3d0d",
         16065 => x"84ba980c",
         16066 => x"04f86134",
         16067 => x"7b4aff6a",
         16068 => x"7081054c",
         16069 => x"34ff6a70",
         16070 => x"81054c34",
         16071 => x"ff6a34ff",
         16072 => x"61840534",
         16073 => x"ff618505",
         16074 => x"34ff6186",
         16075 => x"0534ff61",
         16076 => x"870534ff",
         16077 => x"61880534",
         16078 => x"ff618905",
         16079 => x"34ff618a",
         16080 => x"05348f65",
         16081 => x"347c57f9",
         16082 => x"b1397654",
         16083 => x"861f5360",
         16084 => x"527951fe",
         16085 => x"bed53f84",
         16086 => x"80615657",
         16087 => x"80757081",
         16088 => x"055734ff",
         16089 => x"175776f4",
         16090 => x"38605c80",
         16091 => x"d27c7081",
         16092 => x"055e347b",
         16093 => x"5580d275",
         16094 => x"70810557",
         16095 => x"3480e175",
         16096 => x"70810557",
         16097 => x"3480c175",
         16098 => x"3480f261",
         16099 => x"83e40534",
         16100 => x"80f26183",
         16101 => x"e5053480",
         16102 => x"c16183e6",
         16103 => x"053480e1",
         16104 => x"6183e705",
         16105 => x"347fff05",
         16106 => x"5b7a6183",
         16107 => x"e805347a",
         16108 => x"882a5978",
         16109 => x"6183e905",
         16110 => x"347a902a",
         16111 => x"56756183",
         16112 => x"ea05347a",
         16113 => x"982a407f",
         16114 => x"6183eb05",
         16115 => x"34826183",
         16116 => x"ec053476",
         16117 => x"6183ed05",
         16118 => x"34766183",
         16119 => x"ee053476",
         16120 => x"6183ef05",
         16121 => x"3480d569",
         16122 => x"34ffaa6b",
         16123 => x"34815487",
         16124 => x"1f536052",
         16125 => x"7951febd",
         16126 => x"b23f8154",
         16127 => x"811f5360",
         16128 => x"527951fe",
         16129 => x"bda53f69",
         16130 => x"615755f7",
         16131 => x"a639f43d",
         16132 => x"0d7e615b",
         16133 => x"5b807b61",
         16134 => x"ff055a57",
         16135 => x"57767825",
         16136 => x"b8388d3d",
         16137 => x"598e3df8",
         16138 => x"05548153",
         16139 => x"78527951",
         16140 => x"ff9ab43f",
         16141 => x"7b812e09",
         16142 => x"81069e38",
         16143 => x"8d3d3355",
         16144 => x"748d2e90",
         16145 => x"38747670",
         16146 => x"81055834",
         16147 => x"81175774",
         16148 => x"8a2e8638",
         16149 => x"777724cd",
         16150 => x"38807634",
         16151 => x"7a557683",
         16152 => x"38765574",
         16153 => x"84ba8c0c",
         16154 => x"8e3d0d04",
         16155 => x"f73d0d7b",
         16156 => x"028405b3",
         16157 => x"05335957",
         16158 => x"778a2e80",
         16159 => x"d5388417",
         16160 => x"08568076",
         16161 => x"249e3888",
         16162 => x"17087717",
         16163 => x"8c055659",
         16164 => x"77753481",
         16165 => x"165574bb",
         16166 => x"248e3874",
         16167 => x"84180c81",
         16168 => x"1988180c",
         16169 => x"8b3d0d04",
         16170 => x"8b3dfc05",
         16171 => x"5474538c",
         16172 => x"17527608",
         16173 => x"51ff9ed1",
         16174 => x"3f747a32",
         16175 => x"70307072",
         16176 => x"079f2a70",
         16177 => x"30841b0c",
         16178 => x"811c881b",
         16179 => x"0c5a5656",
         16180 => x"d3398d52",
         16181 => x"7651ff94",
         16182 => x"3fffa339",
         16183 => x"e33d0d02",
         16184 => x"80ff0533",
         16185 => x"8d3d5858",
         16186 => x"80cc7757",
         16187 => x"55807670",
         16188 => x"81055834",
         16189 => x"ff155574",
         16190 => x"f438a13d",
         16191 => x"08770c77",
         16192 => x"8a2e80f7",
         16193 => x"387c5680",
         16194 => x"762480c0",
         16195 => x"387d7717",
         16196 => x"8c055659",
         16197 => x"77753481",
         16198 => x"165574bb",
         16199 => x"24b83874",
         16200 => x"84180c81",
         16201 => x"1988180c",
         16202 => x"7c558075",
         16203 => x"249e389f",
         16204 => x"3dffac11",
         16205 => x"557554c0",
         16206 => x"05527608",
         16207 => x"51ff9dc9",
         16208 => x"3f84ba8c",
         16209 => x"0886387c",
         16210 => x"7a2eba38",
         16211 => x"ff0b84ba",
         16212 => x"8c0c9f3d",
         16213 => x"0d049f3d",
         16214 => x"ffb01155",
         16215 => x"7554c005",
         16216 => x"52760851",
         16217 => x"ff9da23f",
         16218 => x"747b3270",
         16219 => x"30707207",
         16220 => x"9f2a7030",
         16221 => x"525a5656",
         16222 => x"ffa5398d",
         16223 => x"527651fd",
         16224 => x"eb3fff81",
         16225 => x"397d84ba",
         16226 => x"8c0c9f3d",
         16227 => x"0d04fd3d",
         16228 => x"0d750284",
         16229 => x"059a0522",
         16230 => x"52538052",
         16231 => x"7280ff26",
         16232 => x"90387283",
         16233 => x"ffff0652",
         16234 => x"7184ba8c",
         16235 => x"0c853d0d",
         16236 => x"0483ffff",
         16237 => x"73275470",
         16238 => x"83b52e09",
         16239 => x"8106e938",
         16240 => x"73802ee4",
         16241 => x"3883e7d0",
         16242 => x"22517271",
         16243 => x"2e9c3881",
         16244 => x"127083ff",
         16245 => x"ff065354",
         16246 => x"7180ff26",
         16247 => x"8d387110",
         16248 => x"83e7d005",
         16249 => x"70225151",
         16250 => x"e1398180",
         16251 => x"127081ff",
         16252 => x"0684ba8c",
         16253 => x"0c53853d",
         16254 => x"0d04fe3d",
         16255 => x"0d029205",
         16256 => x"22028405",
         16257 => x"96052253",
         16258 => x"51805370",
         16259 => x"80ff268c",
         16260 => x"38705372",
         16261 => x"84ba8c0c",
         16262 => x"843d0d04",
         16263 => x"7183b52e",
         16264 => x"098106ef",
         16265 => x"387081ff",
         16266 => x"26e93870",
         16267 => x"1083e5d0",
         16268 => x"05702284",
         16269 => x"ba8c0c51",
         16270 => x"843d0d04",
         16271 => x"fb3d0d77",
         16272 => x"517083ff",
         16273 => x"ff2680e1",
         16274 => x"387083ff",
         16275 => x"ff0683e9",
         16276 => x"d0565675",
         16277 => x"9fff2680",
         16278 => x"d9387470",
         16279 => x"82055622",
         16280 => x"75713070",
         16281 => x"8025737a",
         16282 => x"26075456",
         16283 => x"535370b7",
         16284 => x"38717082",
         16285 => x"05532272",
         16286 => x"71882a54",
         16287 => x"5681ff06",
         16288 => x"70145254",
         16289 => x"707624b1",
         16290 => x"3871cf38",
         16291 => x"73101570",
         16292 => x"70820552",
         16293 => x"22547330",
         16294 => x"70802575",
         16295 => x"79260753",
         16296 => x"55527080",
         16297 => x"2ecb3875",
         16298 => x"517084ba",
         16299 => x"8c0c873d",
         16300 => x"0d0483ed",
         16301 => x"c455ffa2",
         16302 => x"39718826",
         16303 => x"ea387110",
         16304 => x"1083caa8",
         16305 => x"05547308",
         16306 => x"04c7a016",
         16307 => x"7083ffff",
         16308 => x"06575175",
         16309 => x"51d339ff",
         16310 => x"b0167083",
         16311 => x"ffff0657",
         16312 => x"51f13988",
         16313 => x"167083ff",
         16314 => x"ff065751",
         16315 => x"e639e616",
         16316 => x"7083ffff",
         16317 => x"065751db",
         16318 => x"39d01670",
         16319 => x"83ffff06",
         16320 => x"5751d039",
         16321 => x"e0167083",
         16322 => x"ffff0657",
         16323 => x"51c539f0",
         16324 => x"167083ff",
         16325 => x"ff065751",
         16326 => x"ffb93975",
         16327 => x"73318106",
         16328 => x"76713170",
         16329 => x"83ffff06",
         16330 => x"585255ff",
         16331 => x"a6397573",
         16332 => x"31107505",
         16333 => x"70225252",
         16334 => x"feef3900",
         16335 => x"00ffffff",
         16336 => x"ff00ffff",
         16337 => x"ffff00ff",
         16338 => x"ffffff00",
         16339 => x"0000198b",
         16340 => x"00001980",
         16341 => x"00001975",
         16342 => x"0000196a",
         16343 => x"0000195f",
         16344 => x"00001954",
         16345 => x"00001949",
         16346 => x"0000193e",
         16347 => x"00001933",
         16348 => x"00001928",
         16349 => x"0000191d",
         16350 => x"00001912",
         16351 => x"00001907",
         16352 => x"000018fc",
         16353 => x"000018f1",
         16354 => x"000018e6",
         16355 => x"000018db",
         16356 => x"000018d0",
         16357 => x"000018c5",
         16358 => x"000018ba",
         16359 => x"00001ebf",
         16360 => x"00001f59",
         16361 => x"00001f59",
         16362 => x"00001f59",
         16363 => x"00001f59",
         16364 => x"00001f59",
         16365 => x"00001f59",
         16366 => x"00001f59",
         16367 => x"00001f59",
         16368 => x"00001f59",
         16369 => x"00001f59",
         16370 => x"00001f59",
         16371 => x"00001f59",
         16372 => x"00001f59",
         16373 => x"00001f59",
         16374 => x"00001f59",
         16375 => x"00001f59",
         16376 => x"00001f59",
         16377 => x"00001f59",
         16378 => x"00001f59",
         16379 => x"00001f59",
         16380 => x"00001f59",
         16381 => x"00001f59",
         16382 => x"00001f59",
         16383 => x"00001f59",
         16384 => x"00001f59",
         16385 => x"00001f59",
         16386 => x"00001f59",
         16387 => x"00001f59",
         16388 => x"00001f59",
         16389 => x"00001f59",
         16390 => x"00001f59",
         16391 => x"00001f59",
         16392 => x"00001f59",
         16393 => x"00001f59",
         16394 => x"00001f59",
         16395 => x"00001f59",
         16396 => x"00001f59",
         16397 => x"00001f59",
         16398 => x"00001f59",
         16399 => x"00001f59",
         16400 => x"00001f59",
         16401 => x"00001f59",
         16402 => x"0000247b",
         16403 => x"00001f59",
         16404 => x"00001f59",
         16405 => x"00001f59",
         16406 => x"00001f59",
         16407 => x"00001f59",
         16408 => x"00001f59",
         16409 => x"00001f59",
         16410 => x"00001f59",
         16411 => x"00001f59",
         16412 => x"00001f59",
         16413 => x"00001f59",
         16414 => x"00001f59",
         16415 => x"00001f59",
         16416 => x"00001f59",
         16417 => x"00001f59",
         16418 => x"00001f59",
         16419 => x"00002411",
         16420 => x"00002310",
         16421 => x"00001f59",
         16422 => x"00002294",
         16423 => x"000024b2",
         16424 => x"00002371",
         16425 => x"00002236",
         16426 => x"000021d8",
         16427 => x"00001f59",
         16428 => x"00001f59",
         16429 => x"00001f59",
         16430 => x"00001f59",
         16431 => x"00001f59",
         16432 => x"00001f59",
         16433 => x"00001f59",
         16434 => x"00001f59",
         16435 => x"00001f59",
         16436 => x"00001f59",
         16437 => x"00001f59",
         16438 => x"00001f59",
         16439 => x"00001f59",
         16440 => x"00001f59",
         16441 => x"00001f59",
         16442 => x"00001f59",
         16443 => x"00001f59",
         16444 => x"00001f59",
         16445 => x"00001f59",
         16446 => x"00001f59",
         16447 => x"00001f59",
         16448 => x"00001f59",
         16449 => x"00001f59",
         16450 => x"00001f59",
         16451 => x"00001f59",
         16452 => x"00001f59",
         16453 => x"00001f59",
         16454 => x"00001f59",
         16455 => x"00001f59",
         16456 => x"00001f59",
         16457 => x"00001f59",
         16458 => x"00001f59",
         16459 => x"00001f59",
         16460 => x"00001f59",
         16461 => x"00001f59",
         16462 => x"00001f59",
         16463 => x"00001f59",
         16464 => x"00001f59",
         16465 => x"00001f59",
         16466 => x"00001f59",
         16467 => x"00001f59",
         16468 => x"00001f59",
         16469 => x"00001f59",
         16470 => x"00001f59",
         16471 => x"00001f59",
         16472 => x"00001f59",
         16473 => x"00001f59",
         16474 => x"00001f59",
         16475 => x"00001f59",
         16476 => x"00001f59",
         16477 => x"00001f59",
         16478 => x"00001f59",
         16479 => x"000021b5",
         16480 => x"0000217a",
         16481 => x"00001f59",
         16482 => x"00001f59",
         16483 => x"00001f59",
         16484 => x"00001f59",
         16485 => x"00001f59",
         16486 => x"00001f59",
         16487 => x"00001f59",
         16488 => x"00001f59",
         16489 => x"0000216d",
         16490 => x"00002162",
         16491 => x"00001f59",
         16492 => x"0000214b",
         16493 => x"00001f59",
         16494 => x"0000215b",
         16495 => x"00002151",
         16496 => x"00002144",
         16497 => x"0000321c",
         16498 => x"00003234",
         16499 => x"00003240",
         16500 => x"0000324c",
         16501 => x"00003258",
         16502 => x"00003228",
         16503 => x"00003b91",
         16504 => x"00003a7f",
         16505 => x"000038fb",
         16506 => x"00003649",
         16507 => x"00003a1b",
         16508 => x"000034d8",
         16509 => x"00003795",
         16510 => x"0000366e",
         16511 => x"000039c5",
         16512 => x"0000369d",
         16513 => x"0000370c",
         16514 => x"00003924",
         16515 => x"000034d8",
         16516 => x"000038fb",
         16517 => x"00003805",
         16518 => x"00003795",
         16519 => x"000034d8",
         16520 => x"000034d8",
         16521 => x"0000370c",
         16522 => x"0000369d",
         16523 => x"0000366e",
         16524 => x"00003649",
         16525 => x"00004676",
         16526 => x"0000468f",
         16527 => x"000046b4",
         16528 => x"000046d5",
         16529 => x"00004636",
         16530 => x"000046fa",
         16531 => x"0000464f",
         16532 => x"0000479f",
         16533 => x"0000475c",
         16534 => x"0000475c",
         16535 => x"0000475c",
         16536 => x"0000475c",
         16537 => x"0000475c",
         16538 => x"0000475c",
         16539 => x"00004735",
         16540 => x"0000475c",
         16541 => x"0000475c",
         16542 => x"0000475c",
         16543 => x"0000475c",
         16544 => x"0000475c",
         16545 => x"0000475c",
         16546 => x"0000475c",
         16547 => x"0000475c",
         16548 => x"0000475c",
         16549 => x"0000475c",
         16550 => x"0000475c",
         16551 => x"0000475c",
         16552 => x"0000475c",
         16553 => x"0000475c",
         16554 => x"0000475c",
         16555 => x"0000475c",
         16556 => x"0000475c",
         16557 => x"0000475c",
         16558 => x"0000475c",
         16559 => x"0000475c",
         16560 => x"0000475c",
         16561 => x"0000475c",
         16562 => x"00004874",
         16563 => x"00004862",
         16564 => x"0000484f",
         16565 => x"0000483c",
         16566 => x"00004766",
         16567 => x"0000482a",
         16568 => x"00004817",
         16569 => x"0000477f",
         16570 => x"0000475c",
         16571 => x"0000477f",
         16572 => x"00004807",
         16573 => x"00004884",
         16574 => x"000047b0",
         16575 => x"0000478e",
         16576 => x"000047f5",
         16577 => x"000047e3",
         16578 => x"000047d1",
         16579 => x"000047c2",
         16580 => x"0000475c",
         16581 => x"00004766",
         16582 => x"00005402",
         16583 => x"00005571",
         16584 => x"00005543",
         16585 => x"0000549a",
         16586 => x"00005477",
         16587 => x"00005456",
         16588 => x"0000542c",
         16589 => x"000055fc",
         16590 => x"00005283",
         16591 => x"000055d6",
         16592 => x"000057c5",
         16593 => x"00005283",
         16594 => x"00005283",
         16595 => x"00005283",
         16596 => x"00005283",
         16597 => x"00005283",
         16598 => x"00005283",
         16599 => x"0000559f",
         16600 => x"000057ad",
         16601 => x"00005664",
         16602 => x"00005283",
         16603 => x"00005283",
         16604 => x"00005283",
         16605 => x"00005283",
         16606 => x"00005283",
         16607 => x"00005283",
         16608 => x"00005283",
         16609 => x"00005283",
         16610 => x"00005283",
         16611 => x"00005283",
         16612 => x"00005283",
         16613 => x"00005283",
         16614 => x"00005283",
         16615 => x"00005283",
         16616 => x"00005283",
         16617 => x"00005283",
         16618 => x"00005283",
         16619 => x"00005283",
         16620 => x"00005283",
         16621 => x"00005521",
         16622 => x"00005283",
         16623 => x"00005283",
         16624 => x"00005283",
         16625 => x"000054c4",
         16626 => x"000053d3",
         16627 => x"00005375",
         16628 => x"00005283",
         16629 => x"00005283",
         16630 => x"00005283",
         16631 => x"00005283",
         16632 => x"0000535a",
         16633 => x"00005283",
         16634 => x"0000533d",
         16635 => x"000059a6",
         16636 => x"0000591b",
         16637 => x"0000591b",
         16638 => x"0000591b",
         16639 => x"0000591b",
         16640 => x"0000591b",
         16641 => x"0000591b",
         16642 => x"000058f6",
         16643 => x"0000591b",
         16644 => x"0000591b",
         16645 => x"0000591b",
         16646 => x"0000591b",
         16647 => x"0000591b",
         16648 => x"0000591b",
         16649 => x"0000591b",
         16650 => x"0000591b",
         16651 => x"0000591b",
         16652 => x"0000591b",
         16653 => x"0000591b",
         16654 => x"0000591b",
         16655 => x"0000591b",
         16656 => x"0000591b",
         16657 => x"0000591b",
         16658 => x"0000591b",
         16659 => x"0000591b",
         16660 => x"0000591b",
         16661 => x"0000591b",
         16662 => x"0000591b",
         16663 => x"0000591b",
         16664 => x"0000591b",
         16665 => x"000059b8",
         16666 => x"00005a00",
         16667 => x"000059ed",
         16668 => x"000059da",
         16669 => x"000059c8",
         16670 => x"00005a8b",
         16671 => x"00005a78",
         16672 => x"00005a68",
         16673 => x"0000591b",
         16674 => x"00005a58",
         16675 => x"00005a48",
         16676 => x"00005a36",
         16677 => x"00005a24",
         16678 => x"00005a12",
         16679 => x"00005983",
         16680 => x"00005972",
         16681 => x"00005961",
         16682 => x"0000594a",
         16683 => x"0000591b",
         16684 => x"00005994",
         16685 => x"00006375",
         16686 => x"000061d1",
         16687 => x"000061d1",
         16688 => x"000061d1",
         16689 => x"000061d1",
         16690 => x"000061d1",
         16691 => x"000061d1",
         16692 => x"000061d1",
         16693 => x"000061d1",
         16694 => x"000061d1",
         16695 => x"000061d1",
         16696 => x"000061d1",
         16697 => x"000061d1",
         16698 => x"000061d1",
         16699 => x"00005ef3",
         16700 => x"000061d1",
         16701 => x"000061d1",
         16702 => x"000061d1",
         16703 => x"000061d1",
         16704 => x"000061d1",
         16705 => x"000061d1",
         16706 => x"000063bf",
         16707 => x"000061d1",
         16708 => x"000061d1",
         16709 => x"0000634a",
         16710 => x"000061d1",
         16711 => x"00006361",
         16712 => x"00005ed2",
         16713 => x"00006333",
         16714 => x"0000df2e",
         16715 => x"0000df1b",
         16716 => x"0000df0f",
         16717 => x"0000df04",
         16718 => x"0000def9",
         16719 => x"0000deee",
         16720 => x"0000dee3",
         16721 => x"0000ded7",
         16722 => x"0000dec9",
         16723 => x"00000e01",
         16724 => x"00000bfd",
         16725 => x"00000bfd",
         16726 => x"00000f49",
         16727 => x"00000bfd",
         16728 => x"00000bfd",
         16729 => x"00000bfd",
         16730 => x"00000bfd",
         16731 => x"00000bfd",
         16732 => x"00000bfd",
         16733 => x"00000bfd",
         16734 => x"00000dfd",
         16735 => x"00000bfd",
         16736 => x"00000f7f",
         16737 => x"00000f0d",
         16738 => x"00000bfd",
         16739 => x"00000bfd",
         16740 => x"00000bfd",
         16741 => x"00000bfd",
         16742 => x"00000bfd",
         16743 => x"00000bfd",
         16744 => x"00000bfd",
         16745 => x"00000bfd",
         16746 => x"00000bfd",
         16747 => x"00000bfd",
         16748 => x"00000bfd",
         16749 => x"00000bfd",
         16750 => x"00000bfd",
         16751 => x"00000bfd",
         16752 => x"00000bfd",
         16753 => x"00000bfd",
         16754 => x"00000bfd",
         16755 => x"00000bfd",
         16756 => x"00000bfd",
         16757 => x"00000bfd",
         16758 => x"00000bfd",
         16759 => x"00000bfd",
         16760 => x"00000bfd",
         16761 => x"00000bfd",
         16762 => x"00000bfd",
         16763 => x"00000bfd",
         16764 => x"00000bfd",
         16765 => x"00000bfd",
         16766 => x"00000bfd",
         16767 => x"00000bfd",
         16768 => x"00000bfd",
         16769 => x"00000bfd",
         16770 => x"00000bfd",
         16771 => x"00000bfd",
         16772 => x"00000bfd",
         16773 => x"00000bfd",
         16774 => x"00000f1d",
         16775 => x"00000bfd",
         16776 => x"00000bfd",
         16777 => x"00000bfd",
         16778 => x"00000bfd",
         16779 => x"00000e17",
         16780 => x"00000bfd",
         16781 => x"00000bfd",
         16782 => x"00000bfd",
         16783 => x"00000bfd",
         16784 => x"00000bfd",
         16785 => x"00000bfd",
         16786 => x"00000bfd",
         16787 => x"00000bfd",
         16788 => x"00000bfd",
         16789 => x"00000bfd",
         16790 => x"00000e2b",
         16791 => x"00000ee1",
         16792 => x"00000eb8",
         16793 => x"00000eb8",
         16794 => x"00000eb8",
         16795 => x"00000bfd",
         16796 => x"00000ee1",
         16797 => x"00000bfd",
         16798 => x"00000bfd",
         16799 => x"00000eff",
         16800 => x"00000bfd",
         16801 => x"00000bfd",
         16802 => x"00000c16",
         16803 => x"00000e0f",
         16804 => x"00000bfd",
         16805 => x"00000bfd",
         16806 => x"00000f58",
         16807 => x"00000bfd",
         16808 => x"00000c18",
         16809 => x"00000bfd",
         16810 => x"00000bfd",
         16811 => x"00000e17",
         16812 => x"64696e69",
         16813 => x"74000000",
         16814 => x"64696f63",
         16815 => x"746c0000",
         16816 => x"66696e69",
         16817 => x"74000000",
         16818 => x"666c6f61",
         16819 => x"64000000",
         16820 => x"66657865",
         16821 => x"63000000",
         16822 => x"6d636c65",
         16823 => x"61720000",
         16824 => x"6d636f70",
         16825 => x"79000000",
         16826 => x"6d646966",
         16827 => x"66000000",
         16828 => x"6d64756d",
         16829 => x"70000000",
         16830 => x"6d656200",
         16831 => x"6d656800",
         16832 => x"6d657700",
         16833 => x"68696400",
         16834 => x"68696500",
         16835 => x"68666400",
         16836 => x"68666500",
         16837 => x"63616c6c",
         16838 => x"00000000",
         16839 => x"6a6d7000",
         16840 => x"72657374",
         16841 => x"61727400",
         16842 => x"72657365",
         16843 => x"74000000",
         16844 => x"696e666f",
         16845 => x"00000000",
         16846 => x"74657374",
         16847 => x"00000000",
         16848 => x"636c7300",
         16849 => x"7a383000",
         16850 => x"74626173",
         16851 => x"69630000",
         16852 => x"6d626173",
         16853 => x"69630000",
         16854 => x"6b696c6f",
         16855 => x"00000000",
         16856 => x"65640000",
         16857 => x"556e6b6e",
         16858 => x"6f776e20",
         16859 => x"6572726f",
         16860 => x"722e0000",
         16861 => x"50617261",
         16862 => x"6d657465",
         16863 => x"72732069",
         16864 => x"6e636f72",
         16865 => x"72656374",
         16866 => x"2e000000",
         16867 => x"546f6f20",
         16868 => x"6d616e79",
         16869 => x"206f7065",
         16870 => x"6e206669",
         16871 => x"6c65732e",
         16872 => x"00000000",
         16873 => x"496e7375",
         16874 => x"66666963",
         16875 => x"69656e74",
         16876 => x"206d656d",
         16877 => x"6f72792e",
         16878 => x"00000000",
         16879 => x"46696c65",
         16880 => x"20697320",
         16881 => x"6c6f636b",
         16882 => x"65642e00",
         16883 => x"54696d65",
         16884 => x"6f75742c",
         16885 => x"206f7065",
         16886 => x"72617469",
         16887 => x"6f6e2063",
         16888 => x"616e6365",
         16889 => x"6c6c6564",
         16890 => x"2e000000",
         16891 => x"466f726d",
         16892 => x"61742061",
         16893 => x"626f7274",
         16894 => x"65642e00",
         16895 => x"4e6f2063",
         16896 => x"6f6d7061",
         16897 => x"7469626c",
         16898 => x"65206669",
         16899 => x"6c657379",
         16900 => x"7374656d",
         16901 => x"20666f75",
         16902 => x"6e64206f",
         16903 => x"6e206469",
         16904 => x"736b2e00",
         16905 => x"4469736b",
         16906 => x"206e6f74",
         16907 => x"20656e61",
         16908 => x"626c6564",
         16909 => x"2e000000",
         16910 => x"44726976",
         16911 => x"65206e75",
         16912 => x"6d626572",
         16913 => x"20697320",
         16914 => x"696e7661",
         16915 => x"6c69642e",
         16916 => x"00000000",
         16917 => x"53442069",
         16918 => x"73207772",
         16919 => x"69746520",
         16920 => x"70726f74",
         16921 => x"65637465",
         16922 => x"642e0000",
         16923 => x"46696c65",
         16924 => x"2068616e",
         16925 => x"646c6520",
         16926 => x"696e7661",
         16927 => x"6c69642e",
         16928 => x"00000000",
         16929 => x"46696c65",
         16930 => x"20616c72",
         16931 => x"65616479",
         16932 => x"20657869",
         16933 => x"7374732e",
         16934 => x"00000000",
         16935 => x"41636365",
         16936 => x"73732064",
         16937 => x"656e6965",
         16938 => x"642e0000",
         16939 => x"496e7661",
         16940 => x"6c696420",
         16941 => x"66696c65",
         16942 => x"6e616d65",
         16943 => x"2e000000",
         16944 => x"4e6f2070",
         16945 => x"61746820",
         16946 => x"666f756e",
         16947 => x"642e0000",
         16948 => x"4e6f2066",
         16949 => x"696c6520",
         16950 => x"666f756e",
         16951 => x"642e0000",
         16952 => x"4469736b",
         16953 => x"206e6f74",
         16954 => x"20726561",
         16955 => x"64792e00",
         16956 => x"496e7465",
         16957 => x"726e616c",
         16958 => x"20657272",
         16959 => x"6f722e00",
         16960 => x"4469736b",
         16961 => x"20457272",
         16962 => x"6f720000",
         16963 => x"53756363",
         16964 => x"6573732e",
         16965 => x"00000000",
         16966 => x"0a256c75",
         16967 => x"20627974",
         16968 => x"65732025",
         16969 => x"73206174",
         16970 => x"20256c75",
         16971 => x"20627974",
         16972 => x"65732f73",
         16973 => x"65632e0a",
         16974 => x"00000000",
         16975 => x"72656164",
         16976 => x"00000000",
         16977 => x"2530386c",
         16978 => x"58000000",
         16979 => x"3a202000",
         16980 => x"25303258",
         16981 => x"00000000",
         16982 => x"207c0000",
         16983 => x"7c000000",
         16984 => x"20200000",
         16985 => x"25303458",
         16986 => x"00000000",
         16987 => x"20202020",
         16988 => x"20202020",
         16989 => x"00000000",
         16990 => x"7a4f5300",
         16991 => x"2a2a2025",
         16992 => x"73202800",
         16993 => x"31312f31",
         16994 => x"322f3230",
         16995 => x"32300000",
         16996 => x"76312e31",
         16997 => x"64000000",
         16998 => x"205a5055",
         16999 => x"2c207265",
         17000 => x"76202530",
         17001 => x"32782920",
         17002 => x"25732025",
         17003 => x"73202a2a",
         17004 => x"0a0a0000",
         17005 => x"5a505520",
         17006 => x"496e7465",
         17007 => x"72727570",
         17008 => x"74204861",
         17009 => x"6e646c65",
         17010 => x"72000000",
         17011 => x"55415254",
         17012 => x"31205458",
         17013 => x"20696e74",
         17014 => x"65727275",
         17015 => x"70740000",
         17016 => x"55415254",
         17017 => x"31205258",
         17018 => x"20696e74",
         17019 => x"65727275",
         17020 => x"70740000",
         17021 => x"55415254",
         17022 => x"30205458",
         17023 => x"20696e74",
         17024 => x"65727275",
         17025 => x"70740000",
         17026 => x"55415254",
         17027 => x"30205258",
         17028 => x"20696e74",
         17029 => x"65727275",
         17030 => x"70740000",
         17031 => x"494f4354",
         17032 => x"4c205752",
         17033 => x"20696e74",
         17034 => x"65727275",
         17035 => x"70740000",
         17036 => x"494f4354",
         17037 => x"4c205244",
         17038 => x"20696e74",
         17039 => x"65727275",
         17040 => x"70740000",
         17041 => x"50533220",
         17042 => x"696e7465",
         17043 => x"72727570",
         17044 => x"74000000",
         17045 => x"54696d65",
         17046 => x"7220696e",
         17047 => x"74657272",
         17048 => x"75707400",
         17049 => x"53657474",
         17050 => x"696e6720",
         17051 => x"75702074",
         17052 => x"696d6572",
         17053 => x"2e2e2e00",
         17054 => x"456e6162",
         17055 => x"6c696e67",
         17056 => x"2074696d",
         17057 => x"65722e2e",
         17058 => x"2e000000",
         17059 => x"6175746f",
         17060 => x"65786563",
         17061 => x"2e626174",
         17062 => x"00000000",
         17063 => x"7a4f535f",
         17064 => x"7a70752e",
         17065 => x"68737400",
         17066 => x"4661696c",
         17067 => x"65642074",
         17068 => x"6f20696e",
         17069 => x"69746961",
         17070 => x"6c697365",
         17071 => x"20736420",
         17072 => x"63617264",
         17073 => x"20302c20",
         17074 => x"706c6561",
         17075 => x"73652069",
         17076 => x"6e697420",
         17077 => x"6d616e75",
         17078 => x"616c6c79",
         17079 => x"2e000000",
         17080 => x"2a200000",
         17081 => x"25643a5c",
         17082 => x"25730000",
         17083 => x"4469736b",
         17084 => x"20696e69",
         17085 => x"7469616c",
         17086 => x"69736564",
         17087 => x"00000000",
         17088 => x"303a0000",
         17089 => x"42616420",
         17090 => x"636f6d6d",
         17091 => x"616e642e",
         17092 => x"00000000",
         17093 => x"5a505500",
         17094 => x"62696e00",
         17095 => x"25643a5c",
         17096 => x"25735c25",
         17097 => x"732e2573",
         17098 => x"00000000",
         17099 => x"436f6c64",
         17100 => x"20726562",
         17101 => x"6f6f7469",
         17102 => x"6e672e2e",
         17103 => x"2e000000",
         17104 => x"52657374",
         17105 => x"61727469",
         17106 => x"6e672061",
         17107 => x"70706c69",
         17108 => x"63617469",
         17109 => x"6f6e2e2e",
         17110 => x"2e000000",
         17111 => x"43616c6c",
         17112 => x"696e6720",
         17113 => x"636f6465",
         17114 => x"20402025",
         17115 => x"30386c78",
         17116 => x"202e2e2e",
         17117 => x"0a000000",
         17118 => x"43616c6c",
         17119 => x"20726574",
         17120 => x"75726e65",
         17121 => x"6420636f",
         17122 => x"64652028",
         17123 => x"2564292e",
         17124 => x"0a000000",
         17125 => x"45786563",
         17126 => x"7574696e",
         17127 => x"6720636f",
         17128 => x"64652040",
         17129 => x"20253038",
         17130 => x"6c78202e",
         17131 => x"2e2e0a00",
         17132 => x"2530386c",
         17133 => x"58202530",
         17134 => x"386c582d",
         17135 => x"00000000",
         17136 => x"2530386c",
         17137 => x"58202530",
         17138 => x"34582d00",
         17139 => x"436f6d70",
         17140 => x"6172696e",
         17141 => x"672e2e2e",
         17142 => x"00000000",
         17143 => x"2530386c",
         17144 => x"78282530",
         17145 => x"3878292d",
         17146 => x"3e253038",
         17147 => x"6c782825",
         17148 => x"30387829",
         17149 => x"0a000000",
         17150 => x"436f7079",
         17151 => x"696e672e",
         17152 => x"2e2e0000",
         17153 => x"2530386c",
         17154 => x"58202530",
         17155 => x"32582d00",
         17156 => x"436c6561",
         17157 => x"72696e67",
         17158 => x"2e2e2e2e",
         17159 => x"00000000",
         17160 => x"44756d70",
         17161 => x"204d656d",
         17162 => x"6f727900",
         17163 => x"0a436f6d",
         17164 => x"706c6574",
         17165 => x"652e0000",
         17166 => x"25643a5c",
         17167 => x"25735c25",
         17168 => x"73000000",
         17169 => x"4d656d6f",
         17170 => x"72792065",
         17171 => x"78686175",
         17172 => x"73746564",
         17173 => x"2c206361",
         17174 => x"6e6e6f74",
         17175 => x"2070726f",
         17176 => x"63657373",
         17177 => x"20636f6d",
         17178 => x"6d616e64",
         17179 => x"2e000000",
         17180 => x"3f3f3f00",
         17181 => x"25642f25",
         17182 => x"642f2564",
         17183 => x"2025643a",
         17184 => x"25643a25",
         17185 => x"642e2564",
         17186 => x"25640a00",
         17187 => x"536f4320",
         17188 => x"436f6e66",
         17189 => x"69677572",
         17190 => x"6174696f",
         17191 => x"6e000000",
         17192 => x"3a0a4465",
         17193 => x"76696365",
         17194 => x"7320696d",
         17195 => x"706c656d",
         17196 => x"656e7465",
         17197 => x"643a0000",
         17198 => x"41646472",
         17199 => x"65737365",
         17200 => x"733a0000",
         17201 => x"20202020",
         17202 => x"43505520",
         17203 => x"52657365",
         17204 => x"74205665",
         17205 => x"63746f72",
         17206 => x"20416464",
         17207 => x"72657373",
         17208 => x"203d2025",
         17209 => x"3038580a",
         17210 => x"00000000",
         17211 => x"20202020",
         17212 => x"43505520",
         17213 => x"4d656d6f",
         17214 => x"72792053",
         17215 => x"74617274",
         17216 => x"20416464",
         17217 => x"72657373",
         17218 => x"203d2025",
         17219 => x"3038580a",
         17220 => x"00000000",
         17221 => x"20202020",
         17222 => x"53746163",
         17223 => x"6b205374",
         17224 => x"61727420",
         17225 => x"41646472",
         17226 => x"65737320",
         17227 => x"20202020",
         17228 => x"203d2025",
         17229 => x"3038580a",
         17230 => x"00000000",
         17231 => x"4d697363",
         17232 => x"3a000000",
         17233 => x"20202020",
         17234 => x"5a505520",
         17235 => x"49642020",
         17236 => x"20202020",
         17237 => x"20202020",
         17238 => x"20202020",
         17239 => x"20202020",
         17240 => x"203d2025",
         17241 => x"3034580a",
         17242 => x"00000000",
         17243 => x"20202020",
         17244 => x"53797374",
         17245 => x"656d2043",
         17246 => x"6c6f636b",
         17247 => x"20467265",
         17248 => x"71202020",
         17249 => x"20202020",
         17250 => x"203d2025",
         17251 => x"642e2530",
         17252 => x"34644d48",
         17253 => x"7a0a0000",
         17254 => x"20202020",
         17255 => x"57697368",
         17256 => x"626f6e65",
         17257 => x"20534452",
         17258 => x"414d2043",
         17259 => x"6c6f636b",
         17260 => x"20467265",
         17261 => x"713d2025",
         17262 => x"642e2530",
         17263 => x"34644d48",
         17264 => x"7a0a0000",
         17265 => x"20202020",
         17266 => x"53445241",
         17267 => x"4d20436c",
         17268 => x"6f636b20",
         17269 => x"46726571",
         17270 => x"20202020",
         17271 => x"20202020",
         17272 => x"203d2025",
         17273 => x"642e2530",
         17274 => x"34644d48",
         17275 => x"7a0a0000",
         17276 => x"20202020",
         17277 => x"53504900",
         17278 => x"20202020",
         17279 => x"50533200",
         17280 => x"20202020",
         17281 => x"494f4354",
         17282 => x"4c000000",
         17283 => x"20202020",
         17284 => x"57422049",
         17285 => x"32430000",
         17286 => x"20202020",
         17287 => x"57495348",
         17288 => x"424f4e45",
         17289 => x"20425553",
         17290 => x"00000000",
         17291 => x"20202020",
         17292 => x"494e5452",
         17293 => x"20435452",
         17294 => x"4c202843",
         17295 => x"68616e6e",
         17296 => x"656c733d",
         17297 => x"25303264",
         17298 => x"292e0a00",
         17299 => x"20202020",
         17300 => x"54494d45",
         17301 => x"52312020",
         17302 => x"20202854",
         17303 => x"696d6572",
         17304 => x"7320203d",
         17305 => x"25303264",
         17306 => x"292e0a00",
         17307 => x"20202020",
         17308 => x"53442043",
         17309 => x"41524420",
         17310 => x"20202844",
         17311 => x"65766963",
         17312 => x"6573203d",
         17313 => x"25303264",
         17314 => x"292e0a00",
         17315 => x"20202020",
         17316 => x"52414d20",
         17317 => x"20202020",
         17318 => x"20202825",
         17319 => x"3038583a",
         17320 => x"25303858",
         17321 => x"292e0a00",
         17322 => x"20202020",
         17323 => x"4252414d",
         17324 => x"20202020",
         17325 => x"20202825",
         17326 => x"3038583a",
         17327 => x"25303858",
         17328 => x"292e0a00",
         17329 => x"20202020",
         17330 => x"494e534e",
         17331 => x"20425241",
         17332 => x"4d202825",
         17333 => x"3038583a",
         17334 => x"25303858",
         17335 => x"292e0a00",
         17336 => x"20202020",
         17337 => x"53445241",
         17338 => x"4d202020",
         17339 => x"20202825",
         17340 => x"3038583a",
         17341 => x"25303858",
         17342 => x"292e0a00",
         17343 => x"20202020",
         17344 => x"57422053",
         17345 => x"4452414d",
         17346 => x"20202825",
         17347 => x"3038583a",
         17348 => x"25303858",
         17349 => x"292e0a00",
         17350 => x"20286672",
         17351 => x"6f6d2053",
         17352 => x"6f432063",
         17353 => x"6f6e6669",
         17354 => x"67290000",
         17355 => x"556e6b6e",
         17356 => x"6f776e00",
         17357 => x"45564f6d",
         17358 => x"00000000",
         17359 => x"536d616c",
         17360 => x"6c000000",
         17361 => x"4d656469",
         17362 => x"756d0000",
         17363 => x"466c6578",
         17364 => x"00000000",
         17365 => x"45564f00",
         17366 => x"0000f0b4",
         17367 => x"01000000",
         17368 => x"00000002",
         17369 => x"0000f0b0",
         17370 => x"01000000",
         17371 => x"00000003",
         17372 => x"0000f0ac",
         17373 => x"01000000",
         17374 => x"00000004",
         17375 => x"0000f0a8",
         17376 => x"01000000",
         17377 => x"00000005",
         17378 => x"0000f0a4",
         17379 => x"01000000",
         17380 => x"00000006",
         17381 => x"0000f0a0",
         17382 => x"01000000",
         17383 => x"00000007",
         17384 => x"0000f09c",
         17385 => x"01000000",
         17386 => x"00000001",
         17387 => x"0000f098",
         17388 => x"01000000",
         17389 => x"00000008",
         17390 => x"0000f094",
         17391 => x"01000000",
         17392 => x"0000000b",
         17393 => x"0000f090",
         17394 => x"01000000",
         17395 => x"00000009",
         17396 => x"0000f08c",
         17397 => x"01000000",
         17398 => x"0000000a",
         17399 => x"0000f088",
         17400 => x"04000000",
         17401 => x"0000000d",
         17402 => x"0000f084",
         17403 => x"04000000",
         17404 => x"0000000c",
         17405 => x"0000f080",
         17406 => x"04000000",
         17407 => x"0000000e",
         17408 => x"0000f07c",
         17409 => x"03000000",
         17410 => x"0000000f",
         17411 => x"0000f078",
         17412 => x"04000000",
         17413 => x"0000000f",
         17414 => x"0000f074",
         17415 => x"04000000",
         17416 => x"00000010",
         17417 => x"0000f070",
         17418 => x"04000000",
         17419 => x"00000011",
         17420 => x"0000f06c",
         17421 => x"03000000",
         17422 => x"00000012",
         17423 => x"0000f068",
         17424 => x"03000000",
         17425 => x"00000013",
         17426 => x"0000f064",
         17427 => x"03000000",
         17428 => x"00000014",
         17429 => x"0000f060",
         17430 => x"03000000",
         17431 => x"00000015",
         17432 => x"1b5b4400",
         17433 => x"1b5b4300",
         17434 => x"1b5b4200",
         17435 => x"1b5b4100",
         17436 => x"1b5b367e",
         17437 => x"1b5b357e",
         17438 => x"1b5b347e",
         17439 => x"1b304600",
         17440 => x"1b5b337e",
         17441 => x"1b5b327e",
         17442 => x"1b5b317e",
         17443 => x"10000000",
         17444 => x"0e000000",
         17445 => x"0d000000",
         17446 => x"0b000000",
         17447 => x"08000000",
         17448 => x"06000000",
         17449 => x"05000000",
         17450 => x"04000000",
         17451 => x"03000000",
         17452 => x"02000000",
         17453 => x"01000000",
         17454 => x"43616e6e",
         17455 => x"6f74206f",
         17456 => x"70656e2f",
         17457 => x"63726561",
         17458 => x"74652068",
         17459 => x"6973746f",
         17460 => x"72792066",
         17461 => x"696c652c",
         17462 => x"20646973",
         17463 => x"61626c69",
         17464 => x"6e672e00",
         17465 => x"68697374",
         17466 => x"6f727900",
         17467 => x"68697374",
         17468 => x"00000000",
         17469 => x"21000000",
         17470 => x"2530366c",
         17471 => x"75202025",
         17472 => x"730a0000",
         17473 => x"4661696c",
         17474 => x"65642074",
         17475 => x"6f207265",
         17476 => x"73657420",
         17477 => x"74686520",
         17478 => x"68697374",
         17479 => x"6f727920",
         17480 => x"66696c65",
         17481 => x"20746f20",
         17482 => x"454f462e",
         17483 => x"00000000",
         17484 => x"3e25730a",
         17485 => x"00000000",
         17486 => x"1b5b317e",
         17487 => x"00000000",
         17488 => x"1b5b4100",
         17489 => x"1b5b4200",
         17490 => x"1b5b4300",
         17491 => x"1b5b4400",
         17492 => x"1b5b3130",
         17493 => x"7e000000",
         17494 => x"1b5b3131",
         17495 => x"7e000000",
         17496 => x"1b5b3132",
         17497 => x"7e000000",
         17498 => x"1b5b3133",
         17499 => x"7e000000",
         17500 => x"1b5b3134",
         17501 => x"7e000000",
         17502 => x"1b5b3135",
         17503 => x"7e000000",
         17504 => x"1b5b3137",
         17505 => x"7e000000",
         17506 => x"1b5b3138",
         17507 => x"7e000000",
         17508 => x"1b5b3139",
         17509 => x"7e000000",
         17510 => x"1b5b3230",
         17511 => x"7e000000",
         17512 => x"1b5b327e",
         17513 => x"00000000",
         17514 => x"1b5b337e",
         17515 => x"00000000",
         17516 => x"1b5b4600",
         17517 => x"1b5b357e",
         17518 => x"00000000",
         17519 => x"1b5b367e",
         17520 => x"00000000",
         17521 => x"583a2564",
         17522 => x"2c25642c",
         17523 => x"25642c25",
         17524 => x"642c2564",
         17525 => x"2c25643a",
         17526 => x"25303278",
         17527 => x"00000000",
         17528 => x"443a2564",
         17529 => x"2d25642d",
         17530 => x"25643a25",
         17531 => x"633a2564",
         17532 => x"2c25642c",
         17533 => x"25643a00",
         17534 => x"25642c00",
         17535 => x"4b3a2564",
         17536 => x"3a000000",
         17537 => x"25303278",
         17538 => x"2c000000",
         17539 => x"25635b25",
         17540 => x"643b2564",
         17541 => x"52000000",
         17542 => x"5265706f",
         17543 => x"72742043",
         17544 => x"7572736f",
         17545 => x"723a0000",
         17546 => x"55703a25",
         17547 => x"30327820",
         17548 => x"25303278",
         17549 => x"00000000",
         17550 => x"44773a25",
         17551 => x"30327820",
         17552 => x"25303278",
         17553 => x"00000000",
         17554 => x"48643a25",
         17555 => x"30327820",
         17556 => x"00000000",
         17557 => x"42616420",
         17558 => x"65786974",
         17559 => x"2c205344",
         17560 => x"20496e69",
         17561 => x"74000000",
         17562 => x"42616420",
         17563 => x"65786974",
         17564 => x"2c205344",
         17565 => x"20526561",
         17566 => x"64000000",
         17567 => x"42616420",
         17568 => x"65786974",
         17569 => x"2c205344",
         17570 => x"20577269",
         17571 => x"74650000",
         17572 => x"4e6f2074",
         17573 => x"65737420",
         17574 => x"64656669",
         17575 => x"6e65642e",
         17576 => x"00000000",
         17577 => x"53440000",
         17578 => x"222a3a3c",
         17579 => x"3e3f7c7f",
         17580 => x"00000000",
         17581 => x"2b2c3b3d",
         17582 => x"5b5d0000",
         17583 => x"46415400",
         17584 => x"46415433",
         17585 => x"32000000",
         17586 => x"ebfe904d",
         17587 => x"53444f53",
         17588 => x"352e3000",
         17589 => x"4e4f204e",
         17590 => x"414d4520",
         17591 => x"20202046",
         17592 => x"41542020",
         17593 => x"20202000",
         17594 => x"4e4f204e",
         17595 => x"414d4520",
         17596 => x"20202046",
         17597 => x"41543332",
         17598 => x"20202000",
         17599 => x"0000f2a4",
         17600 => x"00000000",
         17601 => x"00000000",
         17602 => x"00000000",
         17603 => x"01030507",
         17604 => x"090e1012",
         17605 => x"1416181c",
         17606 => x"1e000000",
         17607 => x"809a4541",
         17608 => x"8e418f80",
         17609 => x"45454549",
         17610 => x"49498e8f",
         17611 => x"9092924f",
         17612 => x"994f5555",
         17613 => x"59999a9b",
         17614 => x"9c9d9e9f",
         17615 => x"41494f55",
         17616 => x"a5a5a6a7",
         17617 => x"a8a9aaab",
         17618 => x"acadaeaf",
         17619 => x"b0b1b2b3",
         17620 => x"b4b5b6b7",
         17621 => x"b8b9babb",
         17622 => x"bcbdbebf",
         17623 => x"c0c1c2c3",
         17624 => x"c4c5c6c7",
         17625 => x"c8c9cacb",
         17626 => x"cccdcecf",
         17627 => x"d0d1d2d3",
         17628 => x"d4d5d6d7",
         17629 => x"d8d9dadb",
         17630 => x"dcdddedf",
         17631 => x"e0e1e2e3",
         17632 => x"e4e5e6e7",
         17633 => x"e8e9eaeb",
         17634 => x"ecedeeef",
         17635 => x"f0f1f2f3",
         17636 => x"f4f5f6f7",
         17637 => x"f8f9fafb",
         17638 => x"fcfdfeff",
         17639 => x"2b2e2c3b",
         17640 => x"3d5b5d2f",
         17641 => x"5c222a3a",
         17642 => x"3c3e3f7c",
         17643 => x"7f000000",
         17644 => x"00010004",
         17645 => x"00100040",
         17646 => x"01000200",
         17647 => x"00000000",
         17648 => x"00010002",
         17649 => x"00040008",
         17650 => x"00100020",
         17651 => x"00000000",
         17652 => x"00c700fc",
         17653 => x"00e900e2",
         17654 => x"00e400e0",
         17655 => x"00e500e7",
         17656 => x"00ea00eb",
         17657 => x"00e800ef",
         17658 => x"00ee00ec",
         17659 => x"00c400c5",
         17660 => x"00c900e6",
         17661 => x"00c600f4",
         17662 => x"00f600f2",
         17663 => x"00fb00f9",
         17664 => x"00ff00d6",
         17665 => x"00dc00a2",
         17666 => x"00a300a5",
         17667 => x"20a70192",
         17668 => x"00e100ed",
         17669 => x"00f300fa",
         17670 => x"00f100d1",
         17671 => x"00aa00ba",
         17672 => x"00bf2310",
         17673 => x"00ac00bd",
         17674 => x"00bc00a1",
         17675 => x"00ab00bb",
         17676 => x"25912592",
         17677 => x"25932502",
         17678 => x"25242561",
         17679 => x"25622556",
         17680 => x"25552563",
         17681 => x"25512557",
         17682 => x"255d255c",
         17683 => x"255b2510",
         17684 => x"25142534",
         17685 => x"252c251c",
         17686 => x"2500253c",
         17687 => x"255e255f",
         17688 => x"255a2554",
         17689 => x"25692566",
         17690 => x"25602550",
         17691 => x"256c2567",
         17692 => x"25682564",
         17693 => x"25652559",
         17694 => x"25582552",
         17695 => x"2553256b",
         17696 => x"256a2518",
         17697 => x"250c2588",
         17698 => x"2584258c",
         17699 => x"25902580",
         17700 => x"03b100df",
         17701 => x"039303c0",
         17702 => x"03a303c3",
         17703 => x"00b503c4",
         17704 => x"03a60398",
         17705 => x"03a903b4",
         17706 => x"221e03c6",
         17707 => x"03b52229",
         17708 => x"226100b1",
         17709 => x"22652264",
         17710 => x"23202321",
         17711 => x"00f72248",
         17712 => x"00b02219",
         17713 => x"00b7221a",
         17714 => x"207f00b2",
         17715 => x"25a000a0",
         17716 => x"0061031a",
         17717 => x"00e00317",
         17718 => x"00f80307",
         17719 => x"00ff0001",
         17720 => x"01780100",
         17721 => x"01300132",
         17722 => x"01060139",
         17723 => x"0110014a",
         17724 => x"012e0179",
         17725 => x"01060180",
         17726 => x"004d0243",
         17727 => x"01810182",
         17728 => x"01820184",
         17729 => x"01840186",
         17730 => x"01870187",
         17731 => x"0189018a",
         17732 => x"018b018b",
         17733 => x"018d018e",
         17734 => x"018f0190",
         17735 => x"01910191",
         17736 => x"01930194",
         17737 => x"01f60196",
         17738 => x"01970198",
         17739 => x"0198023d",
         17740 => x"019b019c",
         17741 => x"019d0220",
         17742 => x"019f01a0",
         17743 => x"01a001a2",
         17744 => x"01a201a4",
         17745 => x"01a401a6",
         17746 => x"01a701a7",
         17747 => x"01a901aa",
         17748 => x"01ab01ac",
         17749 => x"01ac01ae",
         17750 => x"01af01af",
         17751 => x"01b101b2",
         17752 => x"01b301b3",
         17753 => x"01b501b5",
         17754 => x"01b701b8",
         17755 => x"01b801ba",
         17756 => x"01bb01bc",
         17757 => x"01bc01be",
         17758 => x"01f701c0",
         17759 => x"01c101c2",
         17760 => x"01c301c4",
         17761 => x"01c501c4",
         17762 => x"01c701c8",
         17763 => x"01c701ca",
         17764 => x"01cb01ca",
         17765 => x"01cd0110",
         17766 => x"01dd0001",
         17767 => x"018e01de",
         17768 => x"011201f3",
         17769 => x"000301f1",
         17770 => x"01f401f4",
         17771 => x"01f80128",
         17772 => x"02220112",
         17773 => x"023a0009",
         17774 => x"2c65023b",
         17775 => x"023b023d",
         17776 => x"2c66023f",
         17777 => x"02400241",
         17778 => x"02410246",
         17779 => x"010a0253",
         17780 => x"00400181",
         17781 => x"01860255",
         17782 => x"0189018a",
         17783 => x"0258018f",
         17784 => x"025a0190",
         17785 => x"025c025d",
         17786 => x"025e025f",
         17787 => x"01930261",
         17788 => x"02620194",
         17789 => x"02640265",
         17790 => x"02660267",
         17791 => x"01970196",
         17792 => x"026a2c62",
         17793 => x"026c026d",
         17794 => x"026e019c",
         17795 => x"02700271",
         17796 => x"019d0273",
         17797 => x"0274019f",
         17798 => x"02760277",
         17799 => x"02780279",
         17800 => x"027a027b",
         17801 => x"027c2c64",
         17802 => x"027e027f",
         17803 => x"01a60281",
         17804 => x"028201a9",
         17805 => x"02840285",
         17806 => x"02860287",
         17807 => x"01ae0244",
         17808 => x"01b101b2",
         17809 => x"0245028d",
         17810 => x"028e028f",
         17811 => x"02900291",
         17812 => x"01b7037b",
         17813 => x"000303fd",
         17814 => x"03fe03ff",
         17815 => x"03ac0004",
         17816 => x"03860388",
         17817 => x"0389038a",
         17818 => x"03b10311",
         17819 => x"03c20002",
         17820 => x"03a303a3",
         17821 => x"03c40308",
         17822 => x"03cc0003",
         17823 => x"038c038e",
         17824 => x"038f03d8",
         17825 => x"011803f2",
         17826 => x"000a03f9",
         17827 => x"03f303f4",
         17828 => x"03f503f6",
         17829 => x"03f703f7",
         17830 => x"03f903fa",
         17831 => x"03fa0430",
         17832 => x"03200450",
         17833 => x"07100460",
         17834 => x"0122048a",
         17835 => x"013604c1",
         17836 => x"010e04cf",
         17837 => x"000104c0",
         17838 => x"04d00144",
         17839 => x"05610426",
         17840 => x"00000000",
         17841 => x"1d7d0001",
         17842 => x"2c631e00",
         17843 => x"01961ea0",
         17844 => x"015a1f00",
         17845 => x"06081f10",
         17846 => x"06061f20",
         17847 => x"06081f30",
         17848 => x"06081f40",
         17849 => x"06061f51",
         17850 => x"00071f59",
         17851 => x"1f521f5b",
         17852 => x"1f541f5d",
         17853 => x"1f561f5f",
         17854 => x"1f600608",
         17855 => x"1f70000e",
         17856 => x"1fba1fbb",
         17857 => x"1fc81fc9",
         17858 => x"1fca1fcb",
         17859 => x"1fda1fdb",
         17860 => x"1ff81ff9",
         17861 => x"1fea1feb",
         17862 => x"1ffa1ffb",
         17863 => x"1f800608",
         17864 => x"1f900608",
         17865 => x"1fa00608",
         17866 => x"1fb00004",
         17867 => x"1fb81fb9",
         17868 => x"1fb21fbc",
         17869 => x"1fcc0001",
         17870 => x"1fc31fd0",
         17871 => x"06021fe0",
         17872 => x"06021fe5",
         17873 => x"00011fec",
         17874 => x"1ff30001",
         17875 => x"1ffc214e",
         17876 => x"00012132",
         17877 => x"21700210",
         17878 => x"21840001",
         17879 => x"218324d0",
         17880 => x"051a2c30",
         17881 => x"042f2c60",
         17882 => x"01022c67",
         17883 => x"01062c75",
         17884 => x"01022c80",
         17885 => x"01642d00",
         17886 => x"0826ff41",
         17887 => x"031a0000",
         17888 => x"00000000",
         17889 => x"0000e6b0",
         17890 => x"01020100",
         17891 => x"00000000",
         17892 => x"00000000",
         17893 => x"0000e6b8",
         17894 => x"01040100",
         17895 => x"00000000",
         17896 => x"00000000",
         17897 => x"0000e6c0",
         17898 => x"01140300",
         17899 => x"00000000",
         17900 => x"00000000",
         17901 => x"0000e6c8",
         17902 => x"012b0300",
         17903 => x"00000000",
         17904 => x"00000000",
         17905 => x"0000e6d0",
         17906 => x"01300300",
         17907 => x"00000000",
         17908 => x"00000000",
         17909 => x"0000e6d8",
         17910 => x"013c0400",
         17911 => x"00000000",
         17912 => x"00000000",
         17913 => x"0000e6e0",
         17914 => x"013d0400",
         17915 => x"00000000",
         17916 => x"00000000",
         17917 => x"0000e6e8",
         17918 => x"013f0400",
         17919 => x"00000000",
         17920 => x"00000000",
         17921 => x"0000e6f0",
         17922 => x"01400400",
         17923 => x"00000000",
         17924 => x"00000000",
         17925 => x"0000e6f8",
         17926 => x"01410400",
         17927 => x"00000000",
         17928 => x"00000000",
         17929 => x"0000e6fc",
         17930 => x"01420400",
         17931 => x"00000000",
         17932 => x"00000000",
         17933 => x"0000e700",
         17934 => x"01430400",
         17935 => x"00000000",
         17936 => x"00000000",
         17937 => x"0000e704",
         17938 => x"01500500",
         17939 => x"00000000",
         17940 => x"00000000",
         17941 => x"0000e708",
         17942 => x"01510500",
         17943 => x"00000000",
         17944 => x"00000000",
         17945 => x"0000e70c",
         17946 => x"01540500",
         17947 => x"00000000",
         17948 => x"00000000",
         17949 => x"0000e710",
         17950 => x"01550500",
         17951 => x"00000000",
         17952 => x"00000000",
         17953 => x"0000e714",
         17954 => x"01790700",
         17955 => x"00000000",
         17956 => x"00000000",
         17957 => x"0000e71c",
         17958 => x"01780700",
         17959 => x"00000000",
         17960 => x"00000000",
         17961 => x"0000e720",
         17962 => x"01820800",
         17963 => x"00000000",
         17964 => x"00000000",
         17965 => x"0000e728",
         17966 => x"01830800",
         17967 => x"00000000",
         17968 => x"00000000",
         17969 => x"0000e730",
         17970 => x"01850800",
         17971 => x"00000000",
         17972 => x"00000000",
         17973 => x"0000e738",
         17974 => x"01870800",
         17975 => x"00000000",
         17976 => x"00000000",
         17977 => x"0000e740",
         17978 => x"01880800",
         17979 => x"00000000",
         17980 => x"00000000",
         17981 => x"0000e744",
         17982 => x"01890800",
         17983 => x"00000000",
         17984 => x"00000000",
         17985 => x"0000e748",
         17986 => x"018c0900",
         17987 => x"00000000",
         17988 => x"00000000",
         17989 => x"0000e750",
         17990 => x"018d0900",
         17991 => x"00000000",
         17992 => x"00000000",
         17993 => x"0000e758",
         17994 => x"018e0900",
         17995 => x"00000000",
         17996 => x"00000000",
         17997 => x"0000e760",
         17998 => x"018f0900",
         17999 => x"00000000",
         18000 => x"00000000",
         18001 => x"00000000",
         18002 => x"00000000",
         18003 => x"00007fff",
         18004 => x"00000000",
         18005 => x"00007fff",
         18006 => x"00010000",
         18007 => x"00007fff",
         18008 => x"00010000",
         18009 => x"00810000",
         18010 => x"01000000",
         18011 => x"017fffff",
         18012 => x"00000000",
         18013 => x"00000000",
         18014 => x"00007800",
         18015 => x"00000000",
         18016 => x"05f5e100",
         18017 => x"05f5e100",
         18018 => x"05f5e100",
         18019 => x"00000000",
         18020 => x"01010101",
         18021 => x"01010101",
         18022 => x"01011001",
         18023 => x"01000000",
         18024 => x"00000000",
         18025 => x"00000000",
         18026 => x"00000000",
         18027 => x"00000000",
         18028 => x"00000000",
         18029 => x"00000000",
         18030 => x"00000000",
         18031 => x"00000000",
         18032 => x"00000000",
         18033 => x"00000000",
         18034 => x"00000000",
         18035 => x"00000000",
         18036 => x"00000000",
         18037 => x"00000000",
         18038 => x"00000000",
         18039 => x"00000000",
         18040 => x"00000000",
         18041 => x"00000000",
         18042 => x"00000000",
         18043 => x"00000000",
         18044 => x"00000000",
         18045 => x"00000000",
         18046 => x"00000000",
         18047 => x"00000000",
         18048 => x"0000f0e4",
         18049 => x"01000000",
         18050 => x"0000f0ec",
         18051 => x"01000000",
         18052 => x"0000f0f4",
         18053 => x"02000000",
         18054 => x"0001fd80",
         18055 => x"1bfc5ffd",
         18056 => x"f03b3a0d",
         18057 => x"797a405b",
         18058 => x"5df0f0f0",
         18059 => x"71727374",
         18060 => x"75767778",
         18061 => x"696a6b6c",
         18062 => x"6d6e6f70",
         18063 => x"61626364",
         18064 => x"65666768",
         18065 => x"31323334",
         18066 => x"35363738",
         18067 => x"5cf32d20",
         18068 => x"30392c2e",
         18069 => x"f67ff3f4",
         18070 => x"f1f23f2f",
         18071 => x"08f0f0f0",
         18072 => x"f0f0f0f0",
         18073 => x"80818283",
         18074 => x"84f0f0f0",
         18075 => x"1bfc58fd",
         18076 => x"f03a3b0d",
         18077 => x"595a405b",
         18078 => x"5df0f0f0",
         18079 => x"51525354",
         18080 => x"55565758",
         18081 => x"494a4b4c",
         18082 => x"4d4e4f50",
         18083 => x"41424344",
         18084 => x"45464748",
         18085 => x"31323334",
         18086 => x"35363738",
         18087 => x"5cf32d20",
         18088 => x"30392c2e",
         18089 => x"f67ff3f4",
         18090 => x"f1f23f2f",
         18091 => x"08f0f0f0",
         18092 => x"f0f0f0f0",
         18093 => x"80818283",
         18094 => x"84f0f0f0",
         18095 => x"1bfc58fd",
         18096 => x"f02b2a0d",
         18097 => x"595a607b",
         18098 => x"7df0f0f0",
         18099 => x"51525354",
         18100 => x"55565758",
         18101 => x"494a4b4c",
         18102 => x"4d4e4f50",
         18103 => x"41424344",
         18104 => x"45464748",
         18105 => x"21222324",
         18106 => x"25262728",
         18107 => x"7c7e3d20",
         18108 => x"20293c3e",
         18109 => x"f7e2e0e1",
         18110 => x"f9f83f2f",
         18111 => x"fbf0f0f0",
         18112 => x"f0f0f0f0",
         18113 => x"85868788",
         18114 => x"89f0f0f0",
         18115 => x"1bfe1efa",
         18116 => x"f0f0f0f0",
         18117 => x"191a001b",
         18118 => x"1df0f0f0",
         18119 => x"11121314",
         18120 => x"15161718",
         18121 => x"090a0b0c",
         18122 => x"0d0e0f10",
         18123 => x"01020304",
         18124 => x"05060708",
         18125 => x"f0f0f0f0",
         18126 => x"f0f0f0f0",
         18127 => x"f01ef0f0",
         18128 => x"f01ff0f0",
         18129 => x"f0f0f0f0",
         18130 => x"f0f0f01c",
         18131 => x"f0f0f0f0",
         18132 => x"f0f0f0f0",
         18133 => x"80818283",
         18134 => x"84f0f0f0",
         18135 => x"bff0cfc9",
         18136 => x"f0b54dcd",
         18137 => x"3577d7b3",
         18138 => x"b7f0f0f0",
         18139 => x"7c704131",
         18140 => x"39a678dd",
         18141 => x"3d5d6c56",
         18142 => x"1d33d5b1",
         18143 => x"466ed948",
         18144 => x"74434c73",
         18145 => x"3f367e3b",
         18146 => x"7a1e5fa2",
         18147 => x"d39fd100",
         18148 => x"9da3d0b9",
         18149 => x"c6c5c2c1",
         18150 => x"c3c4bbbe",
         18151 => x"f0f0f0f0",
         18152 => x"f0f0f0f0",
         18153 => x"80818283",
         18154 => x"84f0f0f0",
         18155 => x"00000000",
         18156 => x"00000000",
         18157 => x"00000000",
         18158 => x"00000000",
         18159 => x"00000000",
         18160 => x"00000000",
         18161 => x"00000000",
         18162 => x"00000000",
         18163 => x"00000000",
         18164 => x"00000000",
         18165 => x"00000000",
         18166 => x"00000000",
         18167 => x"00000000",
         18168 => x"00000000",
         18169 => x"00000000",
         18170 => x"00000000",
         18171 => x"00000000",
         18172 => x"00000000",
         18173 => x"00000000",
         18174 => x"00000000",
         18175 => x"00000000",
         18176 => x"00000000",
         18177 => x"00000000",
         18178 => x"00000000",
         18179 => x"00000000",
         18180 => x"00010000",
         18181 => x"00000000",
         18182 => x"f8000000",
         18183 => x"0000f138",
         18184 => x"f3000000",
         18185 => x"0000f140",
         18186 => x"f4000000",
         18187 => x"0000f144",
         18188 => x"f1000000",
         18189 => x"0000f148",
         18190 => x"f2000000",
         18191 => x"0000f14c",
         18192 => x"80000000",
         18193 => x"0000f150",
         18194 => x"81000000",
         18195 => x"0000f158",
         18196 => x"82000000",
         18197 => x"0000f160",
         18198 => x"83000000",
         18199 => x"0000f168",
         18200 => x"84000000",
         18201 => x"0000f170",
         18202 => x"85000000",
         18203 => x"0000f178",
         18204 => x"86000000",
         18205 => x"0000f180",
         18206 => x"87000000",
         18207 => x"0000f188",
         18208 => x"88000000",
         18209 => x"0000f190",
         18210 => x"89000000",
         18211 => x"0000f198",
         18212 => x"f6000000",
         18213 => x"0000f1a0",
         18214 => x"7f000000",
         18215 => x"0000f1a8",
         18216 => x"f9000000",
         18217 => x"0000f1b0",
         18218 => x"e0000000",
         18219 => x"0000f1b4",
         18220 => x"e1000000",
         18221 => x"0000f1bc",
         18222 => x"71000000",
         18223 => x"00000000",
         18224 => x"00000000",
         18225 => x"00000000",
         18226 => x"00000000",
         18227 => x"00000000",
         18228 => x"00000000",
         18229 => x"00000000",
         18230 => x"00000000",
         18231 => x"00000000",
         18232 => x"00000000",
         18233 => x"00000000",
         18234 => x"00000000",
         18235 => x"00000000",
         18236 => x"00000000",
         18237 => x"00000000",
         18238 => x"00000000",
         18239 => x"00000000",
         18240 => x"00000000",
         18241 => x"00000000",
         18242 => x"00000000",
         18243 => x"00000000",
         18244 => x"00000000",
         18245 => x"00000000",
         18246 => x"00000000",
         18247 => x"00000000",
         18248 => x"00000000",
         18249 => x"00000000",
         18250 => x"00000000",
         18251 => x"00000000",
         18252 => x"00000000",
         18253 => x"00000000",
         18254 => x"00000000",
         18255 => x"00000000",
         18256 => x"00000000",
         18257 => x"00000000",
         18258 => x"00000000",
         18259 => x"00000000",
         18260 => x"00000000",
         18261 => x"00000000",
         18262 => x"00000000",
         18263 => x"00000000",
         18264 => x"00000000",
         18265 => x"00000000",
         18266 => x"00000000",
         18267 => x"00000000",
         18268 => x"00000000",
         18269 => x"00000000",
         18270 => x"00000000",
         18271 => x"00000000",
         18272 => x"00000000",
         18273 => x"00000000",
         18274 => x"00000000",
         18275 => x"00000000",
         18276 => x"00000000",
         18277 => x"00000000",
         18278 => x"00000000",
         18279 => x"00000000",
         18280 => x"00000000",
         18281 => x"00000000",
         18282 => x"00000000",
         18283 => x"00000000",
         18284 => x"00000000",
         18285 => x"00000000",
         18286 => x"00000000",
         18287 => x"00000000",
         18288 => x"00000000",
         18289 => x"00000000",
         18290 => x"00000000",
         18291 => x"00000000",
         18292 => x"00000000",
         18293 => x"00000000",
         18294 => x"00000000",
         18295 => x"00000000",
         18296 => x"00000000",
         18297 => x"00000000",
         18298 => x"00000000",
         18299 => x"00000000",
         18300 => x"00000000",
         18301 => x"00000000",
         18302 => x"00000000",
         18303 => x"00000000",
         18304 => x"00000000",
         18305 => x"00000000",
         18306 => x"00000000",
         18307 => x"00000000",
         18308 => x"00000000",
         18309 => x"00000000",
         18310 => x"00000000",
         18311 => x"00000000",
         18312 => x"00000000",
         18313 => x"00000000",
         18314 => x"00000000",
         18315 => x"00000000",
         18316 => x"00000000",
         18317 => x"00000000",
         18318 => x"00000000",
         18319 => x"00000000",
         18320 => x"00000000",
         18321 => x"00000000",
         18322 => x"00000000",
         18323 => x"00000000",
         18324 => x"00000000",
         18325 => x"00000000",
         18326 => x"00000000",
         18327 => x"00000000",
         18328 => x"00000000",
         18329 => x"00000000",
         18330 => x"00000000",
         18331 => x"00000000",
         18332 => x"00000000",
         18333 => x"00000000",
         18334 => x"00000000",
         18335 => x"00000000",
         18336 => x"00000000",
         18337 => x"00000000",
         18338 => x"00000000",
         18339 => x"00000000",
         18340 => x"00000000",
         18341 => x"00000000",
         18342 => x"00000000",
         18343 => x"00000000",
         18344 => x"00000000",
         18345 => x"00000000",
         18346 => x"00000000",
         18347 => x"00000000",
         18348 => x"00000000",
         18349 => x"00000000",
         18350 => x"00000000",
         18351 => x"00000000",
         18352 => x"00000000",
         18353 => x"00000000",
         18354 => x"00000000",
         18355 => x"00000000",
         18356 => x"00000000",
         18357 => x"00000000",
         18358 => x"00000000",
         18359 => x"00000000",
         18360 => x"00000000",
         18361 => x"00000000",
         18362 => x"00000000",
         18363 => x"00000000",
         18364 => x"00000000",
         18365 => x"00000000",
         18366 => x"00000000",
         18367 => x"00000000",
         18368 => x"00000000",
         18369 => x"00000000",
         18370 => x"00000000",
         18371 => x"00000000",
         18372 => x"00000000",
         18373 => x"00000000",
         18374 => x"00000000",
         18375 => x"00000000",
         18376 => x"00000000",
         18377 => x"00000000",
         18378 => x"00000000",
         18379 => x"00000000",
         18380 => x"00000000",
         18381 => x"00000000",
         18382 => x"00000000",
         18383 => x"00000000",
         18384 => x"00000000",
         18385 => x"00000000",
         18386 => x"00000000",
         18387 => x"00000000",
         18388 => x"00000000",
         18389 => x"00000000",
         18390 => x"00000000",
         18391 => x"00000000",
         18392 => x"00000000",
         18393 => x"00000000",
         18394 => x"00000000",
         18395 => x"00000000",
         18396 => x"00000000",
         18397 => x"00000000",
         18398 => x"00000000",
         18399 => x"00000000",
         18400 => x"00000000",
         18401 => x"00000000",
         18402 => x"00000000",
         18403 => x"00000000",
         18404 => x"00000000",
         18405 => x"00000000",
         18406 => x"00000000",
         18407 => x"00000000",
         18408 => x"00000000",
         18409 => x"00000000",
         18410 => x"00000000",
         18411 => x"00000000",
         18412 => x"00000000",
         18413 => x"00000000",
         18414 => x"00000000",
         18415 => x"00000000",
         18416 => x"00000000",
         18417 => x"00000000",
         18418 => x"00000000",
         18419 => x"00000000",
         18420 => x"00000000",
         18421 => x"00000000",
         18422 => x"00000000",
         18423 => x"00000000",
         18424 => x"00000000",
         18425 => x"00000000",
         18426 => x"00000000",
         18427 => x"00000000",
         18428 => x"00000000",
         18429 => x"00000000",
         18430 => x"00000000",
         18431 => x"00000000",
         18432 => x"00000000",
         18433 => x"00000000",
         18434 => x"00000000",
         18435 => x"00000000",
         18436 => x"00000000",
         18437 => x"00000000",
         18438 => x"00000000",
         18439 => x"00000000",
         18440 => x"00000000",
         18441 => x"00000000",
         18442 => x"00000000",
         18443 => x"00000000",
         18444 => x"00000000",
         18445 => x"00000000",
         18446 => x"00000000",
         18447 => x"00000000",
         18448 => x"00000000",
         18449 => x"00000000",
         18450 => x"00000000",
         18451 => x"00000000",
         18452 => x"00000000",
         18453 => x"00000000",
         18454 => x"00000000",
         18455 => x"00000000",
         18456 => x"00000000",
         18457 => x"00000000",
         18458 => x"00000000",
         18459 => x"00000000",
         18460 => x"00000000",
         18461 => x"00000000",
         18462 => x"00000000",
         18463 => x"00000000",
         18464 => x"00000000",
         18465 => x"00000000",
         18466 => x"00000000",
         18467 => x"00000000",
         18468 => x"00000000",
         18469 => x"00000000",
         18470 => x"00000000",
         18471 => x"00000000",
         18472 => x"00000000",
         18473 => x"00000000",
         18474 => x"00000000",
         18475 => x"00000000",
         18476 => x"00000000",
         18477 => x"00000000",
         18478 => x"00000000",
         18479 => x"00000000",
         18480 => x"00000000",
         18481 => x"00000000",
         18482 => x"00000000",
         18483 => x"00000000",
         18484 => x"00000000",
         18485 => x"00000000",
         18486 => x"00000000",
         18487 => x"00000000",
         18488 => x"00000000",
         18489 => x"00000000",
         18490 => x"00000000",
         18491 => x"00000000",
         18492 => x"00000000",
         18493 => x"00000000",
         18494 => x"00000000",
         18495 => x"00000000",
         18496 => x"00000000",
         18497 => x"00000000",
         18498 => x"00000000",
         18499 => x"00000000",
         18500 => x"00000000",
         18501 => x"00000000",
         18502 => x"00000000",
         18503 => x"00000000",
         18504 => x"00000000",
         18505 => x"00000000",
         18506 => x"00000000",
         18507 => x"00000000",
         18508 => x"00000000",
         18509 => x"00000000",
         18510 => x"00000000",
         18511 => x"00000000",
         18512 => x"00000000",
         18513 => x"00000000",
         18514 => x"00000000",
         18515 => x"00000000",
         18516 => x"00000000",
         18517 => x"00000000",
         18518 => x"00000000",
         18519 => x"00000000",
         18520 => x"00000000",
         18521 => x"00000000",
         18522 => x"00000000",
         18523 => x"00000000",
         18524 => x"00000000",
         18525 => x"00000000",
         18526 => x"00000000",
         18527 => x"00000000",
         18528 => x"00000000",
         18529 => x"00000000",
         18530 => x"00000000",
         18531 => x"00000000",
         18532 => x"00000000",
         18533 => x"00000000",
         18534 => x"00000000",
         18535 => x"00000000",
         18536 => x"00000000",
         18537 => x"00000000",
         18538 => x"00000000",
         18539 => x"00000000",
         18540 => x"00000000",
         18541 => x"00000000",
         18542 => x"00000000",
         18543 => x"00000000",
         18544 => x"00000000",
         18545 => x"00000000",
         18546 => x"00000000",
         18547 => x"00000000",
         18548 => x"00000000",
         18549 => x"00000000",
         18550 => x"00000000",
         18551 => x"00000000",
         18552 => x"00000000",
         18553 => x"00000000",
         18554 => x"00000000",
         18555 => x"00000000",
         18556 => x"00000000",
         18557 => x"00000000",
         18558 => x"00000000",
         18559 => x"00000000",
         18560 => x"00000000",
         18561 => x"00000000",
         18562 => x"00000000",
         18563 => x"00000000",
         18564 => x"00000000",
         18565 => x"00000000",
         18566 => x"00000000",
         18567 => x"00000000",
         18568 => x"00000000",
         18569 => x"00000000",
         18570 => x"00000000",
         18571 => x"00000000",
         18572 => x"00000000",
         18573 => x"00000000",
         18574 => x"00000000",
         18575 => x"00000000",
         18576 => x"00000000",
         18577 => x"00000000",
         18578 => x"00000000",
         18579 => x"00000000",
         18580 => x"00000000",
         18581 => x"00000000",
         18582 => x"00000000",
         18583 => x"00000000",
         18584 => x"00000000",
         18585 => x"00000000",
         18586 => x"00000000",
         18587 => x"00000000",
         18588 => x"00000000",
         18589 => x"00000000",
         18590 => x"00000000",
         18591 => x"00000000",
         18592 => x"00000000",
         18593 => x"00000000",
         18594 => x"00000000",
         18595 => x"00000000",
         18596 => x"00000000",
         18597 => x"00000000",
         18598 => x"00000000",
         18599 => x"00000000",
         18600 => x"00000000",
         18601 => x"00000000",
         18602 => x"00000000",
         18603 => x"00000000",
         18604 => x"00000000",
         18605 => x"00000000",
         18606 => x"00000000",
         18607 => x"00000000",
         18608 => x"00000000",
         18609 => x"00000000",
         18610 => x"00000000",
         18611 => x"00000000",
         18612 => x"00000000",
         18613 => x"00000000",
         18614 => x"00000000",
         18615 => x"00000000",
         18616 => x"00000000",
         18617 => x"00000000",
         18618 => x"00000000",
         18619 => x"00000000",
         18620 => x"00000000",
         18621 => x"00000000",
         18622 => x"00000000",
         18623 => x"00000000",
         18624 => x"00000000",
         18625 => x"00000000",
         18626 => x"00000000",
         18627 => x"00000000",
         18628 => x"00000000",
         18629 => x"00000000",
         18630 => x"00000000",
         18631 => x"00000000",
         18632 => x"00000000",
         18633 => x"00000000",
         18634 => x"00000000",
         18635 => x"00000000",
         18636 => x"00000000",
         18637 => x"00000000",
         18638 => x"00000000",
         18639 => x"00000000",
         18640 => x"00000000",
         18641 => x"00000000",
         18642 => x"00000000",
         18643 => x"00000000",
         18644 => x"00000000",
         18645 => x"00000000",
         18646 => x"00000000",
         18647 => x"00000000",
         18648 => x"00000000",
         18649 => x"00000000",
         18650 => x"00000000",
         18651 => x"00000000",
         18652 => x"00000000",
         18653 => x"00000000",
         18654 => x"00000000",
         18655 => x"00000000",
         18656 => x"00000000",
         18657 => x"00000000",
         18658 => x"00000000",
         18659 => x"00000000",
         18660 => x"00000000",
         18661 => x"00000000",
         18662 => x"00000000",
         18663 => x"00000000",
         18664 => x"00000000",
         18665 => x"00000000",
         18666 => x"00000000",
         18667 => x"00000000",
         18668 => x"00000000",
         18669 => x"00000000",
         18670 => x"00000000",
         18671 => x"00000000",
         18672 => x"00000000",
         18673 => x"00000000",
         18674 => x"00000000",
         18675 => x"00000000",
         18676 => x"00000000",
         18677 => x"00000000",
         18678 => x"00000000",
         18679 => x"00000000",
         18680 => x"00000000",
         18681 => x"00000000",
         18682 => x"00000000",
         18683 => x"00000000",
         18684 => x"00000000",
         18685 => x"00000000",
         18686 => x"00000000",
         18687 => x"00000000",
         18688 => x"00000000",
         18689 => x"00000000",
         18690 => x"00000000",
         18691 => x"00000000",
         18692 => x"00000000",
         18693 => x"00000000",
         18694 => x"00000000",
         18695 => x"00000000",
         18696 => x"00000000",
         18697 => x"00000000",
         18698 => x"00000000",
         18699 => x"00000000",
         18700 => x"00000000",
         18701 => x"00000000",
         18702 => x"00000000",
         18703 => x"00000000",
         18704 => x"00000000",
         18705 => x"00000000",
         18706 => x"00000000",
         18707 => x"00000000",
         18708 => x"00000000",
         18709 => x"00000000",
         18710 => x"00000000",
         18711 => x"00000000",
         18712 => x"00000000",
         18713 => x"00000000",
         18714 => x"00000000",
         18715 => x"00000000",
         18716 => x"00000000",
         18717 => x"00000000",
         18718 => x"00000000",
         18719 => x"00000000",
         18720 => x"00000000",
         18721 => x"00000000",
         18722 => x"00000000",
         18723 => x"00000000",
         18724 => x"00000000",
         18725 => x"00000000",
         18726 => x"00000000",
         18727 => x"00000000",
         18728 => x"00000000",
         18729 => x"00000000",
         18730 => x"00000000",
         18731 => x"00000000",
         18732 => x"00000000",
         18733 => x"00000000",
         18734 => x"00000000",
         18735 => x"00000000",
         18736 => x"00000000",
         18737 => x"00000000",
         18738 => x"00000000",
         18739 => x"00000000",
         18740 => x"00000000",
         18741 => x"00000000",
         18742 => x"00000000",
         18743 => x"00000000",
         18744 => x"00000000",
         18745 => x"00000000",
         18746 => x"00000000",
         18747 => x"00000000",
         18748 => x"00000000",
         18749 => x"00000000",
         18750 => x"00000000",
         18751 => x"00000000",
         18752 => x"00000000",
         18753 => x"00000000",
         18754 => x"00000000",
         18755 => x"00000000",
         18756 => x"00000000",
         18757 => x"00000000",
         18758 => x"00000000",
         18759 => x"00000000",
         18760 => x"00000000",
         18761 => x"00000000",
         18762 => x"00000000",
         18763 => x"00000000",
         18764 => x"00000000",
         18765 => x"00000000",
         18766 => x"00000000",
         18767 => x"00000000",
         18768 => x"00000000",
         18769 => x"00000000",
         18770 => x"00000000",
         18771 => x"00000000",
         18772 => x"00000000",
         18773 => x"00000000",
         18774 => x"00000000",
         18775 => x"00000000",
         18776 => x"00000000",
         18777 => x"00000000",
         18778 => x"00000000",
         18779 => x"00000000",
         18780 => x"00000000",
         18781 => x"00000000",
         18782 => x"00000000",
         18783 => x"00000000",
         18784 => x"00000000",
         18785 => x"00000000",
         18786 => x"00000000",
         18787 => x"00000000",
         18788 => x"00000000",
         18789 => x"00000000",
         18790 => x"00000000",
         18791 => x"00000000",
         18792 => x"00000000",
         18793 => x"00000000",
         18794 => x"00000000",
         18795 => x"00000000",
         18796 => x"00000000",
         18797 => x"00000000",
         18798 => x"00000000",
         18799 => x"00000000",
         18800 => x"00000000",
         18801 => x"00000000",
         18802 => x"00000000",
         18803 => x"00000000",
         18804 => x"00000000",
         18805 => x"00000000",
         18806 => x"00000000",
         18807 => x"00000000",
         18808 => x"00000000",
         18809 => x"00000000",
         18810 => x"00000000",
         18811 => x"00000000",
         18812 => x"00000000",
         18813 => x"00000000",
         18814 => x"00000000",
         18815 => x"00000000",
         18816 => x"00000000",
         18817 => x"00000000",
         18818 => x"00000000",
         18819 => x"00000000",
         18820 => x"00000000",
         18821 => x"00000000",
         18822 => x"00000000",
         18823 => x"00000000",
         18824 => x"00000000",
         18825 => x"00000000",
         18826 => x"00000000",
         18827 => x"00000000",
         18828 => x"00000000",
         18829 => x"00000000",
         18830 => x"00000000",
         18831 => x"00000000",
         18832 => x"00000000",
         18833 => x"00000000",
         18834 => x"00000000",
         18835 => x"00000000",
         18836 => x"00000000",
         18837 => x"00000000",
         18838 => x"00000000",
         18839 => x"00000000",
         18840 => x"00000000",
         18841 => x"00000000",
         18842 => x"00000000",
         18843 => x"00000000",
         18844 => x"00000000",
         18845 => x"00000000",
         18846 => x"00000000",
         18847 => x"00000000",
         18848 => x"00000000",
         18849 => x"00000000",
         18850 => x"00000000",
         18851 => x"00000000",
         18852 => x"00000000",
         18853 => x"00000000",
         18854 => x"00000000",
         18855 => x"00000000",
         18856 => x"00000000",
         18857 => x"00000000",
         18858 => x"00000000",
         18859 => x"00000000",
         18860 => x"00000000",
         18861 => x"00000000",
         18862 => x"00000000",
         18863 => x"00000000",
         18864 => x"00000000",
         18865 => x"00000000",
         18866 => x"00000000",
         18867 => x"00000000",
         18868 => x"00000000",
         18869 => x"00000000",
         18870 => x"00000000",
         18871 => x"00000000",
         18872 => x"00000000",
         18873 => x"00000000",
         18874 => x"00000000",
         18875 => x"00000000",
         18876 => x"00000000",
         18877 => x"00000000",
         18878 => x"00000000",
         18879 => x"00000000",
         18880 => x"00000000",
         18881 => x"00000000",
         18882 => x"00000000",
         18883 => x"00000000",
         18884 => x"00000000",
         18885 => x"00000000",
         18886 => x"00000000",
         18887 => x"00000000",
         18888 => x"00000000",
         18889 => x"00000000",
         18890 => x"00000000",
         18891 => x"00000000",
         18892 => x"00000000",
         18893 => x"00000000",
         18894 => x"00000000",
         18895 => x"00000000",
         18896 => x"00000000",
         18897 => x"00000000",
         18898 => x"00000000",
         18899 => x"00000000",
         18900 => x"00000000",
         18901 => x"00000000",
         18902 => x"00000000",
         18903 => x"00000000",
         18904 => x"00000000",
         18905 => x"00000000",
         18906 => x"00000000",
         18907 => x"00000000",
         18908 => x"00000000",
         18909 => x"00000000",
         18910 => x"00000000",
         18911 => x"00000000",
         18912 => x"00000000",
         18913 => x"00000000",
         18914 => x"00000000",
         18915 => x"00000000",
         18916 => x"00000000",
         18917 => x"00000000",
         18918 => x"00000000",
         18919 => x"00000000",
         18920 => x"00000000",
         18921 => x"00000000",
         18922 => x"00000000",
         18923 => x"00000000",
         18924 => x"00000000",
         18925 => x"00000000",
         18926 => x"00000000",
         18927 => x"00000000",
         18928 => x"00000000",
         18929 => x"00000000",
         18930 => x"00000000",
         18931 => x"00000000",
         18932 => x"00000000",
         18933 => x"00000000",
         18934 => x"00000000",
         18935 => x"00000000",
         18936 => x"00000000",
         18937 => x"00000000",
         18938 => x"00000000",
         18939 => x"00000000",
         18940 => x"00000000",
         18941 => x"00000000",
         18942 => x"00000000",
         18943 => x"00000000",
         18944 => x"00000000",
         18945 => x"00000000",
         18946 => x"00000000",
         18947 => x"00000000",
         18948 => x"00000000",
         18949 => x"00000000",
         18950 => x"00000000",
         18951 => x"00000000",
         18952 => x"00000000",
         18953 => x"00000000",
         18954 => x"00000000",
         18955 => x"00000000",
         18956 => x"00000000",
         18957 => x"00000000",
         18958 => x"00000000",
         18959 => x"00000000",
         18960 => x"00000000",
         18961 => x"00000000",
         18962 => x"00000000",
         18963 => x"00000000",
         18964 => x"00000000",
         18965 => x"00000000",
         18966 => x"00000000",
         18967 => x"00000000",
         18968 => x"00000000",
         18969 => x"00000000",
         18970 => x"00000000",
         18971 => x"00000000",
         18972 => x"00000000",
         18973 => x"00000000",
         18974 => x"00000000",
         18975 => x"00000000",
         18976 => x"00000000",
         18977 => x"00000000",
         18978 => x"00000000",
         18979 => x"00000000",
         18980 => x"00000000",
         18981 => x"00000000",
         18982 => x"00000000",
         18983 => x"00000000",
         18984 => x"00000000",
         18985 => x"00000000",
         18986 => x"00000000",
         18987 => x"00000000",
         18988 => x"00000000",
         18989 => x"00000000",
         18990 => x"00000000",
         18991 => x"00000000",
         18992 => x"00000000",
         18993 => x"00000000",
         18994 => x"00000000",
         18995 => x"00000000",
         18996 => x"00000000",
         18997 => x"00000000",
         18998 => x"00000000",
         18999 => x"00000000",
         19000 => x"00000000",
         19001 => x"00000000",
         19002 => x"00000000",
         19003 => x"00000000",
         19004 => x"00000000",
         19005 => x"00000000",
         19006 => x"00000000",
         19007 => x"00000000",
         19008 => x"00000000",
         19009 => x"00000000",
         19010 => x"00000000",
         19011 => x"00000000",
         19012 => x"00000000",
         19013 => x"00000000",
         19014 => x"00000000",
         19015 => x"00000000",
         19016 => x"00000000",
         19017 => x"00000000",
         19018 => x"00000000",
         19019 => x"00000000",
         19020 => x"00000000",
         19021 => x"00000000",
         19022 => x"00000000",
         19023 => x"00000000",
         19024 => x"00000000",
         19025 => x"00000000",
         19026 => x"00000000",
         19027 => x"00000000",
         19028 => x"00000000",
         19029 => x"00000000",
         19030 => x"00000000",
         19031 => x"00000000",
         19032 => x"00000000",
         19033 => x"00000000",
         19034 => x"00000000",
         19035 => x"00000000",
         19036 => x"00000000",
         19037 => x"00000000",
         19038 => x"00000000",
         19039 => x"00000000",
         19040 => x"00000000",
         19041 => x"00000000",
         19042 => x"00000000",
         19043 => x"00000000",
         19044 => x"00000000",
         19045 => x"00000000",
         19046 => x"00000000",
         19047 => x"00000000",
         19048 => x"00000000",
         19049 => x"00000000",
         19050 => x"00000000",
         19051 => x"00000000",
         19052 => x"00000000",
         19053 => x"00000000",
         19054 => x"00000000",
         19055 => x"00000000",
         19056 => x"00000000",
         19057 => x"00000000",
         19058 => x"00000000",
         19059 => x"00000000",
         19060 => x"00000000",
         19061 => x"00000000",
         19062 => x"00000000",
         19063 => x"00000000",
         19064 => x"00000000",
         19065 => x"00000000",
         19066 => x"00000000",
         19067 => x"00000000",
         19068 => x"00000000",
         19069 => x"00000000",
         19070 => x"00000000",
         19071 => x"00000000",
         19072 => x"00000000",
         19073 => x"00000000",
         19074 => x"00000000",
         19075 => x"00000000",
         19076 => x"00000000",
         19077 => x"00000000",
         19078 => x"00000000",
         19079 => x"00000000",
         19080 => x"00000000",
         19081 => x"00000000",
         19082 => x"00000000",
         19083 => x"00000000",
         19084 => x"00000000",
         19085 => x"00000000",
         19086 => x"00000000",
         19087 => x"00000000",
         19088 => x"00000000",
         19089 => x"00000000",
         19090 => x"00000000",
         19091 => x"00000000",
         19092 => x"00000000",
         19093 => x"00000000",
         19094 => x"00000000",
         19095 => x"00000000",
         19096 => x"00000000",
         19097 => x"00000000",
         19098 => x"00000000",
         19099 => x"00000000",
         19100 => x"00000000",
         19101 => x"00000000",
         19102 => x"00000000",
         19103 => x"00000000",
         19104 => x"00000000",
         19105 => x"00000000",
         19106 => x"00000000",
         19107 => x"00000000",
         19108 => x"00000000",
         19109 => x"00000000",
         19110 => x"00000000",
         19111 => x"00000000",
         19112 => x"00000000",
         19113 => x"00000000",
         19114 => x"00000000",
         19115 => x"00000000",
         19116 => x"00000000",
         19117 => x"00000000",
         19118 => x"00000000",
         19119 => x"00000000",
         19120 => x"00000000",
         19121 => x"00000000",
         19122 => x"00000000",
         19123 => x"00000000",
         19124 => x"00000000",
         19125 => x"00000000",
         19126 => x"00000000",
         19127 => x"00000000",
         19128 => x"00000000",
         19129 => x"00000000",
         19130 => x"00000000",
         19131 => x"00000000",
         19132 => x"00000000",
         19133 => x"00000000",
         19134 => x"00000000",
         19135 => x"00000000",
         19136 => x"00000000",
         19137 => x"00000000",
         19138 => x"00000000",
         19139 => x"00000000",
         19140 => x"00000000",
         19141 => x"00000000",
         19142 => x"00000000",
         19143 => x"00000000",
         19144 => x"00000000",
         19145 => x"00000000",
         19146 => x"00000000",
         19147 => x"00000000",
         19148 => x"00000000",
         19149 => x"00000000",
         19150 => x"00000000",
         19151 => x"00000000",
         19152 => x"00000000",
         19153 => x"00000000",
         19154 => x"00000000",
         19155 => x"00000000",
         19156 => x"00000000",
         19157 => x"00000000",
         19158 => x"00000000",
         19159 => x"00000000",
         19160 => x"00000000",
         19161 => x"00000000",
         19162 => x"00000000",
         19163 => x"00000000",
         19164 => x"00000000",
         19165 => x"00000000",
         19166 => x"00000000",
         19167 => x"00000000",
         19168 => x"00000000",
         19169 => x"00000000",
         19170 => x"00000000",
         19171 => x"00000000",
         19172 => x"00000000",
         19173 => x"00000000",
         19174 => x"00000000",
         19175 => x"00000000",
         19176 => x"00000000",
         19177 => x"00000000",
         19178 => x"00000000",
         19179 => x"00000000",
         19180 => x"00000000",
         19181 => x"00000000",
         19182 => x"00000000",
         19183 => x"00000000",
         19184 => x"00000000",
         19185 => x"00000000",
         19186 => x"00000000",
         19187 => x"00000000",
         19188 => x"00000000",
         19189 => x"00000000",
         19190 => x"00000000",
         19191 => x"00000000",
         19192 => x"00000000",
         19193 => x"00000000",
         19194 => x"00000000",
         19195 => x"00000000",
         19196 => x"00000000",
         19197 => x"00000000",
         19198 => x"00000000",
         19199 => x"00000000",
         19200 => x"00000000",
         19201 => x"00000000",
         19202 => x"00000000",
         19203 => x"00000000",
         19204 => x"00000000",
         19205 => x"00000000",
         19206 => x"00000000",
         19207 => x"00000000",
         19208 => x"00000000",
         19209 => x"00000000",
         19210 => x"00000000",
         19211 => x"00000000",
         19212 => x"00000000",
         19213 => x"00000000",
         19214 => x"00000000",
         19215 => x"00000000",
         19216 => x"00000000",
         19217 => x"00000000",
         19218 => x"00000000",
         19219 => x"00000000",
         19220 => x"00000000",
         19221 => x"00000000",
         19222 => x"00000000",
         19223 => x"00000000",
         19224 => x"00000000",
         19225 => x"00000000",
         19226 => x"00000000",
         19227 => x"00000000",
         19228 => x"00000000",
         19229 => x"00000000",
         19230 => x"00000000",
         19231 => x"00000000",
         19232 => x"00000000",
         19233 => x"00000000",
         19234 => x"00000000",
         19235 => x"00000000",
         19236 => x"00000000",
         19237 => x"00000000",
         19238 => x"00000000",
         19239 => x"00000000",
         19240 => x"00000000",
         19241 => x"00000000",
         19242 => x"00000000",
         19243 => x"00000000",
         19244 => x"00000000",
         19245 => x"00000000",
         19246 => x"00000000",
         19247 => x"00000000",
         19248 => x"00000000",
         19249 => x"00000000",
         19250 => x"00000000",
         19251 => x"00000000",
         19252 => x"00000000",
         19253 => x"00000000",
         19254 => x"00000000",
         19255 => x"00000000",
         19256 => x"00000000",
         19257 => x"00000000",
         19258 => x"00000000",
         19259 => x"00000000",
         19260 => x"00000000",
         19261 => x"00000000",
         19262 => x"00000000",
         19263 => x"00000000",
         19264 => x"00000000",
         19265 => x"00000000",
         19266 => x"00000000",
         19267 => x"00000000",
         19268 => x"00000000",
         19269 => x"00000000",
         19270 => x"00000000",
         19271 => x"00000000",
         19272 => x"00000000",
         19273 => x"00000000",
         19274 => x"00000000",
         19275 => x"00000000",
         19276 => x"00000000",
         19277 => x"00000000",
         19278 => x"00000000",
         19279 => x"00000000",
         19280 => x"00000000",
         19281 => x"00000000",
         19282 => x"00000000",
         19283 => x"00000000",
         19284 => x"00000000",
         19285 => x"00000000",
         19286 => x"00000000",
         19287 => x"00000000",
         19288 => x"00000000",
         19289 => x"00000000",
         19290 => x"00000000",
         19291 => x"00000000",
         19292 => x"00000000",
         19293 => x"00000000",
         19294 => x"00000000",
         19295 => x"00000000",
         19296 => x"00000000",
         19297 => x"00000000",
         19298 => x"00000000",
         19299 => x"00000000",
         19300 => x"00000000",
         19301 => x"00000000",
         19302 => x"00000000",
         19303 => x"00000000",
         19304 => x"00000000",
         19305 => x"00000000",
         19306 => x"00000000",
         19307 => x"00000000",
         19308 => x"00000000",
         19309 => x"00000000",
         19310 => x"00000000",
         19311 => x"00000000",
         19312 => x"00000000",
         19313 => x"00000000",
         19314 => x"00000000",
         19315 => x"00000000",
         19316 => x"00000000",
         19317 => x"00000000",
         19318 => x"00000000",
         19319 => x"00000000",
         19320 => x"00000000",
         19321 => x"00000000",
         19322 => x"00000000",
         19323 => x"00000000",
         19324 => x"00000000",
         19325 => x"00000000",
         19326 => x"00000000",
         19327 => x"00000000",
         19328 => x"00000000",
         19329 => x"00000000",
         19330 => x"00000000",
         19331 => x"00000000",
         19332 => x"00000000",
         19333 => x"00000000",
         19334 => x"00000000",
         19335 => x"00000000",
         19336 => x"00000000",
         19337 => x"00000000",
         19338 => x"00000000",
         19339 => x"00000000",
         19340 => x"00000000",
         19341 => x"00000000",
         19342 => x"00000000",
         19343 => x"00000000",
         19344 => x"00000000",
         19345 => x"00000000",
         19346 => x"00000000",
         19347 => x"00000000",
         19348 => x"00000000",
         19349 => x"00000000",
         19350 => x"00000000",
         19351 => x"00000000",
         19352 => x"00000000",
         19353 => x"00000000",
         19354 => x"00000000",
         19355 => x"00000000",
         19356 => x"00000000",
         19357 => x"00000000",
         19358 => x"00000000",
         19359 => x"00000000",
         19360 => x"00000000",
         19361 => x"00000000",
         19362 => x"00000000",
         19363 => x"00000000",
         19364 => x"00000000",
         19365 => x"00000000",
         19366 => x"00000000",
         19367 => x"00000000",
         19368 => x"00000000",
         19369 => x"00000000",
         19370 => x"00000000",
         19371 => x"00000000",
         19372 => x"00000000",
         19373 => x"00000000",
         19374 => x"00000000",
         19375 => x"00000000",
         19376 => x"00000000",
         19377 => x"00000000",
         19378 => x"00000000",
         19379 => x"00000000",
         19380 => x"00000000",
         19381 => x"00000000",
         19382 => x"00000000",
         19383 => x"00000000",
         19384 => x"00000000",
         19385 => x"00000000",
         19386 => x"00000000",
         19387 => x"00000000",
         19388 => x"00000000",
         19389 => x"00000000",
         19390 => x"00000000",
         19391 => x"00000000",
         19392 => x"00000000",
         19393 => x"00000000",
         19394 => x"00000000",
         19395 => x"00000000",
         19396 => x"00000000",
         19397 => x"00000000",
         19398 => x"00000000",
         19399 => x"00000000",
         19400 => x"00000000",
         19401 => x"00000000",
         19402 => x"00000000",
         19403 => x"00000000",
         19404 => x"00000000",
         19405 => x"00000000",
         19406 => x"00000000",
         19407 => x"00000000",
         19408 => x"00000000",
         19409 => x"00000000",
         19410 => x"00000000",
         19411 => x"00000000",
         19412 => x"00000000",
         19413 => x"00000000",
         19414 => x"00000000",
         19415 => x"00000000",
         19416 => x"00000000",
         19417 => x"00000000",
         19418 => x"00000000",
         19419 => x"00000000",
         19420 => x"00000000",
         19421 => x"00000000",
         19422 => x"00000000",
         19423 => x"00000000",
         19424 => x"00000000",
         19425 => x"00000000",
         19426 => x"00000000",
         19427 => x"00000000",
         19428 => x"00000000",
         19429 => x"00000000",
         19430 => x"00000000",
         19431 => x"00000000",
         19432 => x"00000000",
         19433 => x"00000000",
         19434 => x"00000000",
         19435 => x"00000000",
         19436 => x"00000000",
         19437 => x"00000000",
         19438 => x"00000000",
         19439 => x"00000000",
         19440 => x"00000000",
         19441 => x"00000000",
         19442 => x"00000000",
         19443 => x"00000000",
         19444 => x"00000000",
         19445 => x"00000000",
         19446 => x"00000000",
         19447 => x"00000000",
         19448 => x"00000000",
         19449 => x"00000000",
         19450 => x"00000000",
         19451 => x"00000000",
         19452 => x"00000000",
         19453 => x"00000000",
         19454 => x"00000000",
         19455 => x"00000000",
         19456 => x"00000000",
         19457 => x"00000000",
         19458 => x"00000000",
         19459 => x"00000000",
         19460 => x"00000000",
         19461 => x"00000000",
         19462 => x"00000000",
         19463 => x"00000000",
         19464 => x"00000000",
         19465 => x"00000000",
         19466 => x"00000000",
         19467 => x"00000000",
         19468 => x"00000000",
         19469 => x"00000000",
         19470 => x"00000000",
         19471 => x"00000000",
         19472 => x"00000000",
         19473 => x"00000000",
         19474 => x"00000000",
         19475 => x"00000000",
         19476 => x"00000000",
         19477 => x"00000000",
         19478 => x"00000000",
         19479 => x"00000000",
         19480 => x"00000000",
         19481 => x"00000000",
         19482 => x"00000000",
         19483 => x"00000000",
         19484 => x"00000000",
         19485 => x"00000000",
         19486 => x"00000000",
         19487 => x"00000000",
         19488 => x"00000000",
         19489 => x"00000000",
         19490 => x"00000000",
         19491 => x"00000000",
         19492 => x"00000000",
         19493 => x"00000000",
         19494 => x"00000000",
         19495 => x"00000000",
         19496 => x"00000000",
         19497 => x"00000000",
         19498 => x"00000000",
         19499 => x"00000000",
         19500 => x"00000000",
         19501 => x"00000000",
         19502 => x"00000000",
         19503 => x"00000000",
         19504 => x"00000000",
         19505 => x"00000000",
         19506 => x"00000000",
         19507 => x"00000000",
         19508 => x"00000000",
         19509 => x"00000000",
         19510 => x"00000000",
         19511 => x"00000000",
         19512 => x"00000000",
         19513 => x"00000000",
         19514 => x"00000000",
         19515 => x"00000000",
         19516 => x"00000000",
         19517 => x"00000000",
         19518 => x"00000000",
         19519 => x"00000000",
         19520 => x"00000000",
         19521 => x"00000000",
         19522 => x"00000000",
         19523 => x"00000000",
         19524 => x"00000000",
         19525 => x"00000000",
         19526 => x"00000000",
         19527 => x"00000000",
         19528 => x"00000000",
         19529 => x"00000000",
         19530 => x"00000000",
         19531 => x"00000000",
         19532 => x"00000000",
         19533 => x"00000000",
         19534 => x"00000000",
         19535 => x"00000000",
         19536 => x"00000000",
         19537 => x"00000000",
         19538 => x"00000000",
         19539 => x"00000000",
         19540 => x"00000000",
         19541 => x"00000000",
         19542 => x"00000000",
         19543 => x"00000000",
         19544 => x"00000000",
         19545 => x"00000000",
         19546 => x"00000000",
         19547 => x"00000000",
         19548 => x"00000000",
         19549 => x"00000000",
         19550 => x"00000000",
         19551 => x"00000000",
         19552 => x"00000000",
         19553 => x"00000000",
         19554 => x"00000000",
         19555 => x"00000000",
         19556 => x"00000000",
         19557 => x"00000000",
         19558 => x"00000000",
         19559 => x"00000000",
         19560 => x"00000000",
         19561 => x"00000000",
         19562 => x"00000000",
         19563 => x"00000000",
         19564 => x"00000000",
         19565 => x"00000000",
         19566 => x"00000000",
         19567 => x"00000000",
         19568 => x"00000000",
         19569 => x"00000000",
         19570 => x"00000000",
         19571 => x"00000000",
         19572 => x"00000000",
         19573 => x"00000000",
         19574 => x"00000000",
         19575 => x"00000000",
         19576 => x"00000000",
         19577 => x"00000000",
         19578 => x"00000000",
         19579 => x"00000000",
         19580 => x"00000000",
         19581 => x"00000000",
         19582 => x"00000000",
         19583 => x"00000000",
         19584 => x"00000000",
         19585 => x"00000000",
         19586 => x"00000000",
         19587 => x"00000000",
         19588 => x"00000000",
         19589 => x"00000000",
         19590 => x"00000000",
         19591 => x"00000000",
         19592 => x"00000000",
         19593 => x"00000000",
         19594 => x"00000000",
         19595 => x"00000000",
         19596 => x"00000000",
         19597 => x"00000000",
         19598 => x"00000000",
         19599 => x"00000000",
         19600 => x"00000000",
         19601 => x"00000000",
         19602 => x"00000000",
         19603 => x"00000000",
         19604 => x"00000000",
         19605 => x"00000000",
         19606 => x"00000000",
         19607 => x"00000000",
         19608 => x"00000000",
         19609 => x"00000000",
         19610 => x"00000000",
         19611 => x"00000000",
         19612 => x"00000000",
         19613 => x"00000000",
         19614 => x"00000000",
         19615 => x"00000000",
         19616 => x"00000000",
         19617 => x"00000000",
         19618 => x"00000000",
         19619 => x"00000000",
         19620 => x"00000000",
         19621 => x"00000000",
         19622 => x"00000000",
         19623 => x"00000000",
         19624 => x"00000000",
         19625 => x"00000000",
         19626 => x"00000000",
         19627 => x"00000000",
         19628 => x"00000000",
         19629 => x"00000000",
         19630 => x"00000000",
         19631 => x"00000000",
         19632 => x"00000000",
         19633 => x"00000000",
         19634 => x"00000000",
         19635 => x"00000000",
         19636 => x"00000000",
         19637 => x"00000000",
         19638 => x"00000000",
         19639 => x"00000000",
         19640 => x"00000000",
         19641 => x"00000000",
         19642 => x"00000000",
         19643 => x"00000000",
         19644 => x"00000000",
         19645 => x"00000000",
         19646 => x"00000000",
         19647 => x"00000000",
         19648 => x"00000000",
         19649 => x"00000000",
         19650 => x"00000000",
         19651 => x"00000000",
         19652 => x"00000000",
         19653 => x"00000000",
         19654 => x"00000000",
         19655 => x"00000000",
         19656 => x"00000000",
         19657 => x"00000000",
         19658 => x"00000000",
         19659 => x"00000000",
         19660 => x"00000000",
         19661 => x"00000000",
         19662 => x"00000000",
         19663 => x"00000000",
         19664 => x"00000000",
         19665 => x"00000000",
         19666 => x"00000000",
         19667 => x"00000000",
         19668 => x"00000000",
         19669 => x"00000000",
         19670 => x"00000000",
         19671 => x"00000000",
         19672 => x"00000000",
         19673 => x"00000000",
         19674 => x"00000000",
         19675 => x"00000000",
         19676 => x"00000000",
         19677 => x"00000000",
         19678 => x"00000000",
         19679 => x"00000000",
         19680 => x"00000000",
         19681 => x"00000000",
         19682 => x"00000000",
         19683 => x"00000000",
         19684 => x"00000000",
         19685 => x"00000000",
         19686 => x"00000000",
         19687 => x"00000000",
         19688 => x"00000000",
         19689 => x"00000000",
         19690 => x"00000000",
         19691 => x"00000000",
         19692 => x"00000000",
         19693 => x"00000000",
         19694 => x"00000000",
         19695 => x"00000000",
         19696 => x"00000000",
         19697 => x"00000000",
         19698 => x"00000000",
         19699 => x"00000000",
         19700 => x"00000000",
         19701 => x"00000000",
         19702 => x"00000000",
         19703 => x"00000000",
         19704 => x"00000000",
         19705 => x"00000000",
         19706 => x"00000000",
         19707 => x"00000000",
         19708 => x"00000000",
         19709 => x"00000000",
         19710 => x"00000000",
         19711 => x"00000000",
         19712 => x"00000000",
         19713 => x"00000000",
         19714 => x"00000000",
         19715 => x"00000000",
         19716 => x"00000000",
         19717 => x"00000000",
         19718 => x"00000000",
         19719 => x"00000000",
         19720 => x"00000000",
         19721 => x"00000000",
         19722 => x"00000000",
         19723 => x"00000000",
         19724 => x"00000000",
         19725 => x"00000000",
         19726 => x"00000000",
         19727 => x"00000000",
         19728 => x"00000000",
         19729 => x"00000000",
         19730 => x"00000000",
         19731 => x"00000000",
         19732 => x"00000000",
         19733 => x"00000000",
         19734 => x"00000000",
         19735 => x"00000000",
         19736 => x"00000000",
         19737 => x"00000000",
         19738 => x"00000000",
         19739 => x"00000000",
         19740 => x"00000000",
         19741 => x"00000000",
         19742 => x"00000000",
         19743 => x"00000000",
         19744 => x"00000000",
         19745 => x"00000000",
         19746 => x"00000000",
         19747 => x"00000000",
         19748 => x"00000000",
         19749 => x"00000000",
         19750 => x"00000000",
         19751 => x"00000000",
         19752 => x"00000000",
         19753 => x"00000000",
         19754 => x"00000000",
         19755 => x"00000000",
         19756 => x"00000000",
         19757 => x"00000000",
         19758 => x"00000000",
         19759 => x"00000000",
         19760 => x"00000000",
         19761 => x"00000000",
         19762 => x"00000000",
         19763 => x"00000000",
         19764 => x"00000000",
         19765 => x"00000000",
         19766 => x"00000000",
         19767 => x"00000000",
         19768 => x"00000000",
         19769 => x"00000000",
         19770 => x"00000000",
         19771 => x"00000000",
         19772 => x"00000000",
         19773 => x"00000000",
         19774 => x"00000000",
         19775 => x"00000000",
         19776 => x"00000000",
         19777 => x"00000000",
         19778 => x"00000000",
         19779 => x"00000000",
         19780 => x"00000000",
         19781 => x"00000000",
         19782 => x"00000000",
         19783 => x"00000000",
         19784 => x"00000000",
         19785 => x"00000000",
         19786 => x"00000000",
         19787 => x"00000000",
         19788 => x"00000000",
         19789 => x"00000000",
         19790 => x"00000000",
         19791 => x"00000000",
         19792 => x"00000000",
         19793 => x"00000000",
         19794 => x"00000000",
         19795 => x"00000000",
         19796 => x"00000000",
         19797 => x"00000000",
         19798 => x"00000000",
         19799 => x"00000000",
         19800 => x"00000000",
         19801 => x"00000000",
         19802 => x"00000000",
         19803 => x"00000000",
         19804 => x"00000000",
         19805 => x"00000000",
         19806 => x"00000000",
         19807 => x"00000000",
         19808 => x"00000000",
         19809 => x"00000000",
         19810 => x"00000000",
         19811 => x"00000000",
         19812 => x"00000000",
         19813 => x"00000000",
         19814 => x"00000000",
         19815 => x"00000000",
         19816 => x"00000000",
         19817 => x"00000000",
         19818 => x"00000000",
         19819 => x"00000000",
         19820 => x"00000000",
         19821 => x"00000000",
         19822 => x"00000000",
         19823 => x"00000000",
         19824 => x"00000000",
         19825 => x"00000000",
         19826 => x"00000000",
         19827 => x"00000000",
         19828 => x"00000000",
         19829 => x"00000000",
         19830 => x"00000000",
         19831 => x"00000000",
         19832 => x"00000000",
         19833 => x"00000000",
         19834 => x"00000000",
         19835 => x"00000000",
         19836 => x"00000000",
         19837 => x"00000000",
         19838 => x"00000000",
         19839 => x"00000000",
         19840 => x"00000000",
         19841 => x"00000000",
         19842 => x"00000000",
         19843 => x"00000000",
         19844 => x"00000000",
         19845 => x"00000000",
         19846 => x"00000000",
         19847 => x"00000000",
         19848 => x"00000000",
         19849 => x"00000000",
         19850 => x"00000000",
         19851 => x"00000000",
         19852 => x"00000000",
         19853 => x"00000000",
         19854 => x"00000000",
         19855 => x"00000000",
         19856 => x"00000000",
         19857 => x"00000000",
         19858 => x"00000000",
         19859 => x"00000000",
         19860 => x"00000000",
         19861 => x"00000000",
         19862 => x"00000000",
         19863 => x"00000000",
         19864 => x"00000000",
         19865 => x"00000000",
         19866 => x"00000000",
         19867 => x"00000000",
         19868 => x"00000000",
         19869 => x"00000000",
         19870 => x"00000000",
         19871 => x"00000000",
         19872 => x"00000000",
         19873 => x"00000000",
         19874 => x"00000000",
         19875 => x"00000000",
         19876 => x"00000000",
         19877 => x"00000000",
         19878 => x"00000000",
         19879 => x"00000000",
         19880 => x"00000000",
         19881 => x"00000000",
         19882 => x"00000000",
         19883 => x"00000000",
         19884 => x"00000000",
         19885 => x"00000000",
         19886 => x"00000000",
         19887 => x"00000000",
         19888 => x"00000000",
         19889 => x"00000000",
         19890 => x"00000000",
         19891 => x"00000000",
         19892 => x"00000000",
         19893 => x"00000000",
         19894 => x"00000000",
         19895 => x"00000000",
         19896 => x"00000000",
         19897 => x"00000000",
         19898 => x"00000000",
         19899 => x"00000000",
         19900 => x"00000000",
         19901 => x"00000000",
         19902 => x"00000000",
         19903 => x"00000000",
         19904 => x"00000000",
         19905 => x"00000000",
         19906 => x"00000000",
         19907 => x"00000000",
         19908 => x"00000000",
         19909 => x"00000000",
         19910 => x"00000000",
         19911 => x"00000000",
         19912 => x"00000000",
         19913 => x"00000000",
         19914 => x"00000000",
         19915 => x"00000000",
         19916 => x"00000000",
         19917 => x"00000000",
         19918 => x"00000000",
         19919 => x"00000000",
         19920 => x"00000000",
         19921 => x"00000000",
         19922 => x"00000000",
         19923 => x"00000000",
         19924 => x"00000000",
         19925 => x"00000000",
         19926 => x"00000000",
         19927 => x"00000000",
         19928 => x"00000000",
         19929 => x"00000000",
         19930 => x"00000000",
         19931 => x"00000000",
         19932 => x"00000000",
         19933 => x"00000000",
         19934 => x"00000000",
         19935 => x"00000000",
         19936 => x"00000000",
         19937 => x"00000000",
         19938 => x"00000000",
         19939 => x"00000000",
         19940 => x"00000000",
         19941 => x"00000000",
         19942 => x"00000000",
         19943 => x"00000000",
         19944 => x"00000000",
         19945 => x"00000000",
         19946 => x"00000000",
         19947 => x"00000000",
         19948 => x"00000000",
         19949 => x"00000000",
         19950 => x"00000000",
         19951 => x"00000000",
         19952 => x"00000000",
         19953 => x"00000000",
         19954 => x"00000000",
         19955 => x"00000000",
         19956 => x"00000000",
         19957 => x"00000000",
         19958 => x"00000000",
         19959 => x"00000000",
         19960 => x"00000000",
         19961 => x"00000000",
         19962 => x"00000000",
         19963 => x"00000000",
         19964 => x"00000000",
         19965 => x"00000000",
         19966 => x"00000000",
         19967 => x"00000000",
         19968 => x"00000000",
         19969 => x"00000000",
         19970 => x"00000000",
         19971 => x"00000000",
         19972 => x"00000000",
         19973 => x"00000000",
         19974 => x"00000000",
         19975 => x"00000000",
         19976 => x"00000000",
         19977 => x"00000000",
         19978 => x"00000000",
         19979 => x"00000000",
         19980 => x"00000000",
         19981 => x"00000000",
         19982 => x"00000000",
         19983 => x"00000000",
         19984 => x"00000000",
         19985 => x"00000000",
         19986 => x"00000000",
         19987 => x"00000000",
         19988 => x"00000000",
         19989 => x"00000000",
         19990 => x"00000000",
         19991 => x"00000000",
         19992 => x"00000000",
         19993 => x"00000000",
         19994 => x"00000000",
         19995 => x"00000000",
         19996 => x"00000000",
         19997 => x"00000000",
         19998 => x"00000000",
         19999 => x"00000000",
         20000 => x"00000000",
         20001 => x"00000000",
         20002 => x"00000000",
         20003 => x"00000000",
         20004 => x"00000000",
         20005 => x"00000000",
         20006 => x"00000000",
         20007 => x"00000000",
         20008 => x"00000000",
         20009 => x"00000000",
         20010 => x"00000000",
         20011 => x"00000000",
         20012 => x"00000000",
         20013 => x"00000000",
         20014 => x"00000000",
         20015 => x"00000000",
         20016 => x"00000000",
         20017 => x"00000000",
         20018 => x"00000000",
         20019 => x"00000000",
         20020 => x"00000000",
         20021 => x"00000000",
         20022 => x"00000000",
         20023 => x"00000000",
         20024 => x"00000000",
         20025 => x"00000000",
         20026 => x"00000000",
         20027 => x"00000000",
         20028 => x"00000000",
         20029 => x"00000000",
         20030 => x"00000000",
         20031 => x"00000000",
         20032 => x"00000000",
         20033 => x"00000000",
         20034 => x"00000000",
         20035 => x"00000000",
         20036 => x"00000000",
         20037 => x"00000000",
         20038 => x"00000000",
         20039 => x"00000000",
         20040 => x"00000000",
         20041 => x"00000000",
         20042 => x"00000000",
         20043 => x"00000000",
         20044 => x"00000000",
         20045 => x"00000000",
         20046 => x"00000000",
         20047 => x"00000000",
         20048 => x"00000000",
         20049 => x"00000000",
         20050 => x"00000000",
         20051 => x"00000000",
         20052 => x"00000000",
         20053 => x"00000000",
         20054 => x"00000000",
         20055 => x"00000000",
         20056 => x"00000000",
         20057 => x"00000000",
         20058 => x"00000000",
         20059 => x"00000000",
         20060 => x"00000000",
         20061 => x"00000000",
         20062 => x"00000000",
         20063 => x"00000000",
         20064 => x"00000000",
         20065 => x"00000000",
         20066 => x"00000000",
         20067 => x"00000000",
         20068 => x"00000000",
         20069 => x"00000000",
         20070 => x"00000000",
         20071 => x"00000000",
         20072 => x"00000000",
         20073 => x"00000000",
         20074 => x"00000000",
         20075 => x"00000000",
         20076 => x"00000000",
         20077 => x"00000000",
         20078 => x"00000000",
         20079 => x"00000000",
         20080 => x"00000000",
         20081 => x"00000000",
         20082 => x"00000000",
         20083 => x"00000000",
         20084 => x"00000000",
         20085 => x"00000000",
         20086 => x"00000000",
         20087 => x"00000000",
         20088 => x"00000000",
         20089 => x"00000000",
         20090 => x"00000000",
         20091 => x"00000000",
         20092 => x"00000000",
         20093 => x"00000000",
         20094 => x"00000000",
         20095 => x"00000000",
         20096 => x"00000000",
         20097 => x"00000000",
         20098 => x"00000000",
         20099 => x"00000000",
         20100 => x"00000000",
         20101 => x"00000000",
         20102 => x"00000000",
         20103 => x"00000000",
         20104 => x"00000000",
         20105 => x"00000000",
         20106 => x"00000000",
         20107 => x"00000000",
         20108 => x"00000000",
         20109 => x"00000000",
         20110 => x"00000000",
         20111 => x"00000000",
         20112 => x"00000000",
         20113 => x"00000000",
         20114 => x"00000000",
         20115 => x"00000000",
         20116 => x"00000000",
         20117 => x"00000000",
         20118 => x"00000000",
         20119 => x"00000000",
         20120 => x"00000000",
         20121 => x"00000000",
         20122 => x"00000000",
         20123 => x"00000000",
         20124 => x"00000000",
         20125 => x"00000000",
         20126 => x"00000000",
         20127 => x"00000000",
         20128 => x"00000000",
         20129 => x"00000000",
         20130 => x"00000000",
         20131 => x"00000000",
         20132 => x"00000000",
         20133 => x"00000000",
         20134 => x"00000000",
         20135 => x"00000000",
         20136 => x"00000000",
         20137 => x"00000000",
         20138 => x"00000000",
         20139 => x"00000000",
         20140 => x"00000000",
         20141 => x"00000000",
         20142 => x"00000000",
         20143 => x"00000000",
         20144 => x"00000000",
         20145 => x"00000000",
         20146 => x"00000000",
         20147 => x"00000000",
         20148 => x"00000000",
         20149 => x"00000000",
         20150 => x"00000000",
         20151 => x"00000000",
         20152 => x"00000000",
         20153 => x"00000000",
         20154 => x"00000000",
         20155 => x"00000000",
         20156 => x"00000000",
         20157 => x"00000000",
         20158 => x"00000000",
         20159 => x"00000000",
         20160 => x"00000000",
         20161 => x"00000000",
         20162 => x"00000000",
         20163 => x"00000000",
         20164 => x"00000000",
         20165 => x"00000000",
         20166 => x"00000000",
         20167 => x"00000000",
         20168 => x"00000000",
         20169 => x"00000000",
         20170 => x"00000000",
         20171 => x"00000000",
         20172 => x"00000000",
         20173 => x"00000000",
         20174 => x"00000000",
         20175 => x"00000000",
         20176 => x"00000000",
         20177 => x"00000000",
         20178 => x"00000000",
         20179 => x"00000000",
         20180 => x"00000000",
         20181 => x"00000000",
         20182 => x"00000000",
         20183 => x"00000000",
         20184 => x"00000000",
         20185 => x"00000000",
         20186 => x"00000000",
         20187 => x"00000000",
         20188 => x"00000000",
         20189 => x"00000000",
         20190 => x"00000000",
         20191 => x"00000000",
         20192 => x"00000000",
         20193 => x"00000000",
         20194 => x"00000000",
         20195 => x"00000000",
         20196 => x"00000000",
         20197 => x"00000000",
         20198 => x"00000000",
         20199 => x"00000000",
         20200 => x"00000000",
         20201 => x"00000000",
         20202 => x"00000000",
         20203 => x"00000000",
         20204 => x"00000000",
         20205 => x"00000000",
         20206 => x"00000000",
         20207 => x"00000000",
         20208 => x"00000000",
         20209 => x"00000000",
         20210 => x"00000000",
         20211 => x"00000000",
         20212 => x"00000000",
         20213 => x"00000000",
         20214 => x"00000000",
         20215 => x"00000000",
         20216 => x"00000000",
         20217 => x"00000000",
         20218 => x"00000000",
         20219 => x"00000000",
         20220 => x"00000000",
         20221 => x"00000000",
         20222 => x"00000000",
         20223 => x"00003219",
         20224 => x"50000101",
         20225 => x"00000000",
         20226 => x"cce0f2f3",
         20227 => x"cecff6f7",
         20228 => x"f8f9fafb",
         20229 => x"fcfdfeff",
         20230 => x"e1c1c2c3",
         20231 => x"c4c5c6e2",
         20232 => x"e3e4e5e6",
         20233 => x"ebeeeff4",
         20234 => x"00616263",
         20235 => x"64656667",
         20236 => x"68696b6a",
         20237 => x"2f2a2e2d",
         20238 => x"20212223",
         20239 => x"24252627",
         20240 => x"28294f2c",
         20241 => x"512b5749",
         20242 => x"55010203",
         20243 => x"04050607",
         20244 => x"08090a0b",
         20245 => x"0c0d0e0f",
         20246 => x"10111213",
         20247 => x"14151617",
         20248 => x"18191a52",
         20249 => x"5954be3c",
         20250 => x"c7818283",
         20251 => x"84858687",
         20252 => x"88898a8b",
         20253 => x"8c8d8e8f",
         20254 => x"90919293",
         20255 => x"94959697",
         20256 => x"98999abc",
         20257 => x"8040a5c0",
         20258 => x"00000000",
         20259 => x"00000000",
         20260 => x"00000000",
         20261 => x"00000000",
         20262 => x"00000000",
         20263 => x"00000000",
         20264 => x"00000000",
         20265 => x"00000000",
         20266 => x"00000000",
         20267 => x"00000000",
         20268 => x"00000000",
         20269 => x"00000000",
         20270 => x"00000000",
         20271 => x"00000000",
         20272 => x"00000000",
         20273 => x"00000000",
         20274 => x"00000000",
         20275 => x"00000000",
         20276 => x"00000000",
         20277 => x"00000000",
         20278 => x"00000000",
         20279 => x"00000000",
         20280 => x"00000000",
         20281 => x"00000000",
         20282 => x"00000000",
         20283 => x"00000000",
         20284 => x"00000000",
         20285 => x"00000000",
         20286 => x"00000000",
         20287 => x"00000000",
         20288 => x"00020003",
         20289 => x"00040101",
         20290 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

