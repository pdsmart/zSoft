-- Byte Addressed 32bit/64bit BRAM module for the ZPU Evo implementation.
--
-- This template provides a 32bit wide bus on port A and a 64bit bus
-- on port B. This is typically used for the ZPU Boot BRAM where port B
-- is used exclusively for instruction storage.
--
-- Copyright 2018-2021 - Philip Smart for the ZPU Evo implementation.
-- History:
--   20190618  - Initial 32 bit dual port BRAM described by inference rather than
--               using an IP Megacore. This was to make it more portable but also
--               to allow 8/16/32 bit writes to the memory.
--   20210108  - Updated to 64bit on Port B to allow for the 64bit decoder on the ZPU.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPort3264BootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 3);
        memBWrite            : in  std_logic_vector(WORD_64BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_64BIT_RANGE)
    );
end DualPort3264BootBRAM;

architecture arch of DualPort3264BootBRAM is

    -- Declare 8 byte wide arrays for byte level addressing.
    type ramArray is array(natural range 0 to (2**(addrbits-3))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"fa",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"05",
            10 => x"52",
            11 => x"00",
            12 => x"08",
            13 => x"81",
            14 => x"06",
            15 => x"0b",
            16 => x"05",
            17 => x"06",
            18 => x"06",
            19 => x"00",
            20 => x"73",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"09",
            25 => x"72",
            26 => x"31",
            27 => x"51",
            28 => x"73",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"93",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"2b",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"06",
            45 => x"b0",
            46 => x"00",
            47 => x"00",
            48 => x"ff",
            49 => x"0a",
            50 => x"51",
            51 => x"00",
            52 => x"51",
            53 => x"05",
            54 => x"72",
            55 => x"00",
            56 => x"05",
            57 => x"06",
            58 => x"00",
            59 => x"00",
            60 => x"05",
            61 => x"06",
            62 => x"00",
            63 => x"00",
            64 => x"05",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"81",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"06",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"08",
            77 => x"05",
            78 => x"52",
            79 => x"00",
            80 => x"08",
            81 => x"06",
            82 => x"0b",
            83 => x"00",
            84 => x"08",
            85 => x"ac",
            86 => x"90",
            87 => x"00",
            88 => x"08",
            89 => x"ab",
            90 => x"90",
            91 => x"00",
            92 => x"81",
            93 => x"05",
            94 => x"74",
            95 => x"51",
            96 => x"81",
            97 => x"ff",
            98 => x"72",
            99 => x"51",
           100 => x"04",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"52",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"72",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"ff",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"8c",
           133 => x"04",
           134 => x"0b",
           135 => x"8c",
           136 => x"04",
           137 => x"0b",
           138 => x"8c",
           139 => x"04",
           140 => x"0b",
           141 => x"8d",
           142 => x"04",
           143 => x"0b",
           144 => x"8d",
           145 => x"04",
           146 => x"0b",
           147 => x"8e",
           148 => x"04",
           149 => x"0b",
           150 => x"8f",
           151 => x"04",
           152 => x"0b",
           153 => x"8f",
           154 => x"04",
           155 => x"0b",
           156 => x"90",
           157 => x"04",
           158 => x"0b",
           159 => x"90",
           160 => x"04",
           161 => x"0b",
           162 => x"91",
           163 => x"04",
           164 => x"0b",
           165 => x"91",
           166 => x"04",
           167 => x"0b",
           168 => x"92",
           169 => x"04",
           170 => x"0b",
           171 => x"92",
           172 => x"04",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"81",
           193 => x"ec",
           194 => x"80",
           195 => x"ee",
           196 => x"80",
           197 => x"f3",
           198 => x"80",
           199 => x"e0",
           200 => x"80",
           201 => x"a3",
           202 => x"80",
           203 => x"f6",
           204 => x"80",
           205 => x"86",
           206 => x"80",
           207 => x"82",
           208 => x"80",
           209 => x"88",
           210 => x"80",
           211 => x"a8",
           212 => x"80",
           213 => x"d1",
           214 => x"80",
           215 => x"8a",
           216 => x"80",
           217 => x"d4",
           218 => x"c0",
           219 => x"80",
           220 => x"80",
           221 => x"0c",
           222 => x"08",
           223 => x"f0",
           224 => x"f0",
           225 => x"b8",
           226 => x"b8",
           227 => x"84",
           228 => x"84",
           229 => x"04",
           230 => x"2d",
           231 => x"90",
           232 => x"af",
           233 => x"80",
           234 => x"ed",
           235 => x"c0",
           236 => x"82",
           237 => x"80",
           238 => x"0c",
           239 => x"08",
           240 => x"f0",
           241 => x"f0",
           242 => x"b8",
           243 => x"b8",
           244 => x"84",
           245 => x"84",
           246 => x"04",
           247 => x"2d",
           248 => x"90",
           249 => x"d6",
           250 => x"80",
           251 => x"8a",
           252 => x"c0",
           253 => x"82",
           254 => x"80",
           255 => x"0c",
           256 => x"08",
           257 => x"f0",
           258 => x"f0",
           259 => x"b8",
           260 => x"b8",
           261 => x"84",
           262 => x"84",
           263 => x"04",
           264 => x"2d",
           265 => x"90",
           266 => x"96",
           267 => x"80",
           268 => x"96",
           269 => x"c0",
           270 => x"83",
           271 => x"80",
           272 => x"0c",
           273 => x"08",
           274 => x"f0",
           275 => x"f0",
           276 => x"b8",
           277 => x"b8",
           278 => x"84",
           279 => x"84",
           280 => x"04",
           281 => x"2d",
           282 => x"90",
           283 => x"d2",
           284 => x"80",
           285 => x"f4",
           286 => x"c0",
           287 => x"81",
           288 => x"80",
           289 => x"0c",
           290 => x"08",
           291 => x"f0",
           292 => x"f0",
           293 => x"b8",
           294 => x"b8",
           295 => x"84",
           296 => x"b8",
           297 => x"84",
           298 => x"84",
           299 => x"04",
           300 => x"2d",
           301 => x"90",
           302 => x"ac",
           303 => x"80",
           304 => x"d5",
           305 => x"c0",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"00",
           311 => x"06",
           312 => x"10",
           313 => x"51",
           314 => x"ff",
           315 => x"52",
           316 => x"38",
           317 => x"e4",
           318 => x"80",
           319 => x"0b",
           320 => x"80",
           321 => x"87",
           322 => x"56",
           323 => x"51",
           324 => x"fa",
           325 => x"33",
           326 => x"07",
           327 => x"72",
           328 => x"ff",
           329 => x"70",
           330 => x"56",
           331 => x"80",
           332 => x"3f",
           333 => x"e4",
           334 => x"e4",
           335 => x"ff",
           336 => x"72",
           337 => x"73",
           338 => x"76",
           339 => x"3d",
           340 => x"0c",
           341 => x"7d",
           342 => x"34",
           343 => x"88",
           344 => x"05",
           345 => x"74",
           346 => x"0d",
           347 => x"75",
           348 => x"f1",
           349 => x"5d",
           350 => x"33",
           351 => x"55",
           352 => x"09",
           353 => x"57",
           354 => x"1c",
           355 => x"2e",
           356 => x"89",
           357 => x"70",
           358 => x"78",
           359 => x"7a",
           360 => x"40",
           361 => x"82",
           362 => x"ff",
           363 => x"84",
           364 => x"7a",
           365 => x"79",
           366 => x"2c",
           367 => x"0a",
           368 => x"56",
           369 => x"73",
           370 => x"78",
           371 => x"38",
           372 => x"81",
           373 => x"5a",
           374 => x"fe",
           375 => x"76",
           376 => x"76",
           377 => x"83",
           378 => x"8a",
           379 => x"7e",
           380 => x"d8",
           381 => x"c9",
           382 => x"e0",
           383 => x"eb",
           384 => x"3f",
           385 => x"86",
           386 => x"fe",
           387 => x"05",
           388 => x"5e",
           389 => x"79",
           390 => x"b8",
           391 => x"e4",
           392 => x"89",
           393 => x"b0",
           394 => x"40",
           395 => x"3f",
           396 => x"e4",
           397 => x"31",
           398 => x"7e",
           399 => x"80",
           400 => x"2c",
           401 => x"06",
           402 => x"77",
           403 => x"05",
           404 => x"84",
           405 => x"53",
           406 => x"70",
           407 => x"9e",
           408 => x"06",
           409 => x"38",
           410 => x"2a",
           411 => x"81",
           412 => x"38",
           413 => x"2c",
           414 => x"73",
           415 => x"2a",
           416 => x"7a",
           417 => x"98",
           418 => x"73",
           419 => x"73",
           420 => x"06",
           421 => x"78",
           422 => x"05",
           423 => x"74",
           424 => x"88",
           425 => x"29",
           426 => x"5a",
           427 => x"74",
           428 => x"38",
           429 => x"ff",
           430 => x"55",
           431 => x"b0",
           432 => x"80",
           433 => x"98",
           434 => x"e5",
           435 => x"5c",
           436 => x"76",
           437 => x"80",
           438 => x"d3",
           439 => x"f4",
           440 => x"70",
           441 => x"84",
           442 => x"38",
           443 => x"fc",
           444 => x"29",
           445 => x"5a",
           446 => x"38",
           447 => x"e2",
           448 => x"07",
           449 => x"38",
           450 => x"5b",
           451 => x"05",
           452 => x"5f",
           453 => x"7f",
           454 => x"06",
           455 => x"07",
           456 => x"80",
           457 => x"56",
           458 => x"81",
           459 => x"77",
           460 => x"80",
           461 => x"80",
           462 => x"a0",
           463 => x"1a",
           464 => x"79",
           465 => x"7c",
           466 => x"51",
           467 => x"70",
           468 => x"83",
           469 => x"52",
           470 => x"85",
           471 => x"06",
           472 => x"80",
           473 => x"2c",
           474 => x"2a",
           475 => x"fd",
           476 => x"84",
           477 => x"56",
           478 => x"83",
           479 => x"5e",
           480 => x"33",
           481 => x"ca",
           482 => x"33",
           483 => x"ba",
           484 => x"77",
           485 => x"82",
           486 => x"84",
           487 => x"78",
           488 => x"90",
           489 => x"c0",
           490 => x"be",
           491 => x"05",
           492 => x"41",
           493 => x"87",
           494 => x"ff",
           495 => x"54",
           496 => x"7c",
           497 => x"f7",
           498 => x"29",
           499 => x"5a",
           500 => x"38",
           501 => x"e2",
           502 => x"3f",
           503 => x"e3",
           504 => x"3f",
           505 => x"80",
           506 => x"75",
           507 => x"70",
           508 => x"5a",
           509 => x"a2",
           510 => x"3f",
           511 => x"fa",
           512 => x"75",
           513 => x"81",
           514 => x"38",
           515 => x"2b",
           516 => x"39",
           517 => x"c8",
           518 => x"3f",
           519 => x"88",
           520 => x"ff",
           521 => x"54",
           522 => x"7e",
           523 => x"57",
           524 => x"84",
           525 => x"51",
           526 => x"fa",
           527 => x"d4",
           528 => x"2a",
           529 => x"58",
           530 => x"09",
           531 => x"81",
           532 => x"b0",
           533 => x"51",
           534 => x"b8",
           535 => x"57",
           536 => x"72",
           537 => x"08",
           538 => x"54",
           539 => x"90",
           540 => x"e4",
           541 => x"76",
           542 => x"3d",
           543 => x"56",
           544 => x"81",
           545 => x"55",
           546 => x"09",
           547 => x"05",
           548 => x"81",
           549 => x"b8",
           550 => x"70",
           551 => x"2e",
           552 => x"15",
           553 => x"08",
           554 => x"81",
           555 => x"38",
           556 => x"c8",
           557 => x"3d",
           558 => x"85",
           559 => x"81",
           560 => x"72",
           561 => x"54",
           562 => x"08",
           563 => x"38",
           564 => x"08",
           565 => x"53",
           566 => x"75",
           567 => x"04",
           568 => x"90",
           569 => x"84",
           570 => x"08",
           571 => x"d7",
           572 => x"33",
           573 => x"81",
           574 => x"71",
           575 => x"52",
           576 => x"06",
           577 => x"75",
           578 => x"2e",
           579 => x"8c",
           580 => x"71",
           581 => x"e4",
           582 => x"bf",
           583 => x"16",
           584 => x"16",
           585 => x"0d",
           586 => x"74",
           587 => x"b8",
           588 => x"85",
           589 => x"84",
           590 => x"71",
           591 => x"ff",
           592 => x"3d",
           593 => x"85",
           594 => x"3d",
           595 => x"71",
           596 => x"f7",
           597 => x"05",
           598 => x"05",
           599 => x"b8",
           600 => x"3d",
           601 => x"52",
           602 => x"72",
           603 => x"38",
           604 => x"70",
           605 => x"70",
           606 => x"86",
           607 => x"75",
           608 => x"53",
           609 => x"33",
           610 => x"2e",
           611 => x"53",
           612 => x"70",
           613 => x"74",
           614 => x"53",
           615 => x"70",
           616 => x"84",
           617 => x"77",
           618 => x"05",
           619 => x"05",
           620 => x"b8",
           621 => x"3d",
           622 => x"52",
           623 => x"70",
           624 => x"05",
           625 => x"38",
           626 => x"0d",
           627 => x"55",
           628 => x"73",
           629 => x"52",
           630 => x"9a",
           631 => x"b7",
           632 => x"80",
           633 => x"3d",
           634 => x"73",
           635 => x"e9",
           636 => x"71",
           637 => x"84",
           638 => x"71",
           639 => x"04",
           640 => x"52",
           641 => x"08",
           642 => x"55",
           643 => x"08",
           644 => x"9b",
           645 => x"80",
           646 => x"b8",
           647 => x"b8",
           648 => x"0c",
           649 => x"75",
           650 => x"71",
           651 => x"05",
           652 => x"38",
           653 => x"81",
           654 => x"31",
           655 => x"85",
           656 => x"77",
           657 => x"80",
           658 => x"05",
           659 => x"38",
           660 => x"0d",
           661 => x"54",
           662 => x"76",
           663 => x"08",
           664 => x"8d",
           665 => x"84",
           666 => x"72",
           667 => x"72",
           668 => x"74",
           669 => x"2b",
           670 => x"76",
           671 => x"2a",
           672 => x"31",
           673 => x"7b",
           674 => x"5c",
           675 => x"74",
           676 => x"71",
           677 => x"04",
           678 => x"80",
           679 => x"25",
           680 => x"71",
           681 => x"30",
           682 => x"31",
           683 => x"70",
           684 => x"71",
           685 => x"1b",
           686 => x"80",
           687 => x"2a",
           688 => x"06",
           689 => x"19",
           690 => x"54",
           691 => x"55",
           692 => x"58",
           693 => x"fd",
           694 => x"53",
           695 => x"e4",
           696 => x"b8",
           697 => x"fa",
           698 => x"53",
           699 => x"fe",
           700 => x"e0",
           701 => x"73",
           702 => x"e4",
           703 => x"26",
           704 => x"2e",
           705 => x"a0",
           706 => x"54",
           707 => x"38",
           708 => x"10",
           709 => x"9f",
           710 => x"75",
           711 => x"52",
           712 => x"72",
           713 => x"04",
           714 => x"9f",
           715 => x"9f",
           716 => x"74",
           717 => x"56",
           718 => x"b8",
           719 => x"b8",
           720 => x"3d",
           721 => x"7b",
           722 => x"59",
           723 => x"38",
           724 => x"55",
           725 => x"ad",
           726 => x"81",
           727 => x"77",
           728 => x"80",
           729 => x"80",
           730 => x"70",
           731 => x"70",
           732 => x"27",
           733 => x"06",
           734 => x"38",
           735 => x"76",
           736 => x"70",
           737 => x"ff",
           738 => x"75",
           739 => x"75",
           740 => x"04",
           741 => x"33",
           742 => x"81",
           743 => x"78",
           744 => x"e2",
           745 => x"f8",
           746 => x"27",
           747 => x"88",
           748 => x"75",
           749 => x"04",
           750 => x"70",
           751 => x"39",
           752 => x"3d",
           753 => x"5b",
           754 => x"70",
           755 => x"09",
           756 => x"78",
           757 => x"2e",
           758 => x"38",
           759 => x"14",
           760 => x"db",
           761 => x"27",
           762 => x"89",
           763 => x"55",
           764 => x"51",
           765 => x"13",
           766 => x"73",
           767 => x"81",
           768 => x"16",
           769 => x"56",
           770 => x"80",
           771 => x"7a",
           772 => x"0c",
           773 => x"70",
           774 => x"73",
           775 => x"38",
           776 => x"55",
           777 => x"90",
           778 => x"81",
           779 => x"14",
           780 => x"27",
           781 => x"0c",
           782 => x"15",
           783 => x"80",
           784 => x"b8",
           785 => x"d6",
           786 => x"ff",
           787 => x"3d",
           788 => x"38",
           789 => x"52",
           790 => x"ef",
           791 => x"ce",
           792 => x"0d",
           793 => x"3f",
           794 => x"51",
           795 => x"83",
           796 => x"3d",
           797 => x"87",
           798 => x"94",
           799 => x"04",
           800 => x"83",
           801 => x"ee",
           802 => x"cf",
           803 => x"0d",
           804 => x"3f",
           805 => x"51",
           806 => x"83",
           807 => x"3d",
           808 => x"af",
           809 => x"d4",
           810 => x"04",
           811 => x"83",
           812 => x"ee",
           813 => x"d1",
           814 => x"0d",
           815 => x"3f",
           816 => x"51",
           817 => x"83",
           818 => x"3d",
           819 => x"84",
           820 => x"80",
           821 => x"25",
           822 => x"87",
           823 => x"77",
           824 => x"93",
           825 => x"77",
           826 => x"95",
           827 => x"84",
           828 => x"38",
           829 => x"30",
           830 => x"70",
           831 => x"58",
           832 => x"98",
           833 => x"80",
           834 => x"29",
           835 => x"08",
           836 => x"83",
           837 => x"84",
           838 => x"84",
           839 => x"0c",
           840 => x"d4",
           841 => x"77",
           842 => x"e4",
           843 => x"88",
           844 => x"80",
           845 => x"d5",
           846 => x"b1",
           847 => x"51",
           848 => x"54",
           849 => x"d1",
           850 => x"39",
           851 => x"b7",
           852 => x"53",
           853 => x"84",
           854 => x"2e",
           855 => x"77",
           856 => x"04",
           857 => x"55",
           858 => x"52",
           859 => x"08",
           860 => x"04",
           861 => x"8c",
           862 => x"15",
           863 => x"5e",
           864 => x"52",
           865 => x"83",
           866 => x"54",
           867 => x"2e",
           868 => x"a8",
           869 => x"81",
           870 => x"f8",
           871 => x"d4",
           872 => x"aa",
           873 => x"d2",
           874 => x"75",
           875 => x"70",
           876 => x"27",
           877 => x"74",
           878 => x"06",
           879 => x"80",
           880 => x"81",
           881 => x"a0",
           882 => x"78",
           883 => x"51",
           884 => x"5c",
           885 => x"b8",
           886 => x"58",
           887 => x"76",
           888 => x"57",
           889 => x"0b",
           890 => x"04",
           891 => x"81",
           892 => x"a0",
           893 => x"fe",
           894 => x"98",
           895 => x"d4",
           896 => x"ea",
           897 => x"73",
           898 => x"72",
           899 => x"ec",
           900 => x"53",
           901 => x"74",
           902 => x"d2",
           903 => x"84",
           904 => x"ea",
           905 => x"38",
           906 => x"38",
           907 => x"db",
           908 => x"08",
           909 => x"78",
           910 => x"84",
           911 => x"f2",
           912 => x"80",
           913 => x"81",
           914 => x"2e",
           915 => x"d0",
           916 => x"90",
           917 => x"a5",
           918 => x"70",
           919 => x"72",
           920 => x"73",
           921 => x"57",
           922 => x"38",
           923 => x"e4",
           924 => x"a0",
           925 => x"30",
           926 => x"51",
           927 => x"73",
           928 => x"80",
           929 => x"0d",
           930 => x"80",
           931 => x"9c",
           932 => x"fe",
           933 => x"81",
           934 => x"82",
           935 => x"06",
           936 => x"83",
           937 => x"81",
           938 => x"06",
           939 => x"85",
           940 => x"80",
           941 => x"06",
           942 => x"87",
           943 => x"a9",
           944 => x"72",
           945 => x"0d",
           946 => x"d2",
           947 => x"9b",
           948 => x"0d",
           949 => x"d3",
           950 => x"9b",
           951 => x"53",
           952 => x"81",
           953 => x"51",
           954 => x"3f",
           955 => x"52",
           956 => x"39",
           957 => x"b0",
           958 => x"96",
           959 => x"51",
           960 => x"ff",
           961 => x"83",
           962 => x"51",
           963 => x"81",
           964 => x"c2",
           965 => x"de",
           966 => x"3f",
           967 => x"2a",
           968 => x"2e",
           969 => x"51",
           970 => x"9a",
           971 => x"72",
           972 => x"71",
           973 => x"39",
           974 => x"fc",
           975 => x"8e",
           976 => x"51",
           977 => x"ff",
           978 => x"41",
           979 => x"42",
           980 => x"3f",
           981 => x"9b",
           982 => x"b1",
           983 => x"3f",
           984 => x"d6",
           985 => x"80",
           986 => x"0b",
           987 => x"06",
           988 => x"38",
           989 => x"81",
           990 => x"c1",
           991 => x"2e",
           992 => x"a0",
           993 => x"1a",
           994 => x"f6",
           995 => x"38",
           996 => x"70",
           997 => x"b8",
           998 => x"7a",
           999 => x"3f",
          1000 => x"1b",
          1001 => x"38",
          1002 => x"5b",
          1003 => x"33",
          1004 => x"80",
          1005 => x"84",
          1006 => x"08",
          1007 => x"e4",
          1008 => x"51",
          1009 => x"60",
          1010 => x"81",
          1011 => x"e7",
          1012 => x"26",
          1013 => x"5e",
          1014 => x"7a",
          1015 => x"2e",
          1016 => x"83",
          1017 => x"3f",
          1018 => x"57",
          1019 => x"80",
          1020 => x"51",
          1021 => x"84",
          1022 => x"72",
          1023 => x"80",
          1024 => x"5a",
          1025 => x"8d",
          1026 => x"5c",
          1027 => x"32",
          1028 => x"ee",
          1029 => x"7d",
          1030 => x"88",
          1031 => x"f8",
          1032 => x"3f",
          1033 => x"81",
          1034 => x"38",
          1035 => x"cf",
          1036 => x"b8",
          1037 => x"0b",
          1038 => x"f4",
          1039 => x"f6",
          1040 => x"2e",
          1041 => x"df",
          1042 => x"33",
          1043 => x"82",
          1044 => x"91",
          1045 => x"c3",
          1046 => x"d8",
          1047 => x"52",
          1048 => x"5a",
          1049 => x"7c",
          1050 => x"78",
          1051 => x"10",
          1052 => x"08",
          1053 => x"7e",
          1054 => x"52",
          1055 => x"3f",
          1056 => x"81",
          1057 => x"3d",
          1058 => x"d5",
          1059 => x"81",
          1060 => x"d5",
          1061 => x"54",
          1062 => x"51",
          1063 => x"8c",
          1064 => x"3f",
          1065 => x"bf",
          1066 => x"c5",
          1067 => x"51",
          1068 => x"83",
          1069 => x"fd",
          1070 => x"84",
          1071 => x"8a",
          1072 => x"fa",
          1073 => x"51",
          1074 => x"84",
          1075 => x"38",
          1076 => x"8c",
          1077 => x"b8",
          1078 => x"05",
          1079 => x"08",
          1080 => x"83",
          1081 => x"59",
          1082 => x"53",
          1083 => x"84",
          1084 => x"38",
          1085 => x"80",
          1086 => x"e4",
          1087 => x"08",
          1088 => x"d0",
          1089 => x"80",
          1090 => x"7e",
          1091 => x"f9",
          1092 => x"38",
          1093 => x"39",
          1094 => x"80",
          1095 => x"e4",
          1096 => x"3d",
          1097 => x"51",
          1098 => x"86",
          1099 => x"78",
          1100 => x"3f",
          1101 => x"52",
          1102 => x"7e",
          1103 => x"38",
          1104 => x"82",
          1105 => x"3d",
          1106 => x"51",
          1107 => x"80",
          1108 => x"fc",
          1109 => x"da",
          1110 => x"f8",
          1111 => x"53",
          1112 => x"84",
          1113 => x"38",
          1114 => x"68",
          1115 => x"8d",
          1116 => x"5c",
          1117 => x"55",
          1118 => x"83",
          1119 => x"66",
          1120 => x"59",
          1121 => x"53",
          1122 => x"84",
          1123 => x"38",
          1124 => x"80",
          1125 => x"e4",
          1126 => x"3d",
          1127 => x"51",
          1128 => x"80",
          1129 => x"51",
          1130 => x"27",
          1131 => x"81",
          1132 => x"05",
          1133 => x"11",
          1134 => x"3f",
          1135 => x"c3",
          1136 => x"ff",
          1137 => x"b8",
          1138 => x"54",
          1139 => x"3f",
          1140 => x"52",
          1141 => x"7e",
          1142 => x"38",
          1143 => x"81",
          1144 => x"80",
          1145 => x"05",
          1146 => x"ff",
          1147 => x"b8",
          1148 => x"68",
          1149 => x"34",
          1150 => x"fc",
          1151 => x"8a",
          1152 => x"38",
          1153 => x"11",
          1154 => x"3f",
          1155 => x"a3",
          1156 => x"ff",
          1157 => x"b8",
          1158 => x"b8",
          1159 => x"05",
          1160 => x"08",
          1161 => x"83",
          1162 => x"67",
          1163 => x"65",
          1164 => x"0c",
          1165 => x"d9",
          1166 => x"ff",
          1167 => x"b8",
          1168 => x"52",
          1169 => x"b8",
          1170 => x"3f",
          1171 => x"a3",
          1172 => x"f6",
          1173 => x"84",
          1174 => x"d2",
          1175 => x"83",
          1176 => x"83",
          1177 => x"b8",
          1178 => x"05",
          1179 => x"08",
          1180 => x"79",
          1181 => x"a4",
          1182 => x"53",
          1183 => x"84",
          1184 => x"80",
          1185 => x"38",
          1186 => x"70",
          1187 => x"5f",
          1188 => x"a0",
          1189 => x"b4",
          1190 => x"54",
          1191 => x"a8",
          1192 => x"3f",
          1193 => x"59",
          1194 => x"f0",
          1195 => x"a6",
          1196 => x"f2",
          1197 => x"64",
          1198 => x"11",
          1199 => x"3f",
          1200 => x"bb",
          1201 => x"22",
          1202 => x"45",
          1203 => x"80",
          1204 => x"e4",
          1205 => x"5e",
          1206 => x"82",
          1207 => x"fe",
          1208 => x"e1",
          1209 => x"b9",
          1210 => x"fc",
          1211 => x"aa",
          1212 => x"81",
          1213 => x"05",
          1214 => x"fb",
          1215 => x"53",
          1216 => x"84",
          1217 => x"38",
          1218 => x"05",
          1219 => x"83",
          1220 => x"7b",
          1221 => x"83",
          1222 => x"3f",
          1223 => x"da",
          1224 => x"d8",
          1225 => x"b8",
          1226 => x"05",
          1227 => x"08",
          1228 => x"80",
          1229 => x"5b",
          1230 => x"f1",
          1231 => x"cf",
          1232 => x"ea",
          1233 => x"80",
          1234 => x"49",
          1235 => x"d3",
          1236 => x"83",
          1237 => x"59",
          1238 => x"59",
          1239 => x"b0",
          1240 => x"84",
          1241 => x"83",
          1242 => x"9b",
          1243 => x"92",
          1244 => x"80",
          1245 => x"49",
          1246 => x"5e",
          1247 => x"bc",
          1248 => x"e6",
          1249 => x"83",
          1250 => x"83",
          1251 => x"94",
          1252 => x"ca",
          1253 => x"05",
          1254 => x"08",
          1255 => x"3d",
          1256 => x"87",
          1257 => x"87",
          1258 => x"3f",
          1259 => x"08",
          1260 => x"51",
          1261 => x"08",
          1262 => x"70",
          1263 => x"74",
          1264 => x"08",
          1265 => x"84",
          1266 => x"74",
          1267 => x"8c",
          1268 => x"0c",
          1269 => x"94",
          1270 => x"e0",
          1271 => x"34",
          1272 => x"3d",
          1273 => x"84",
          1274 => x"89",
          1275 => x"51",
          1276 => x"83",
          1277 => x"f1",
          1278 => x"3f",
          1279 => x"53",
          1280 => x"51",
          1281 => x"82",
          1282 => x"70",
          1283 => x"74",
          1284 => x"70",
          1285 => x"2e",
          1286 => x"70",
          1287 => x"55",
          1288 => x"ff",
          1289 => x"38",
          1290 => x"38",
          1291 => x"53",
          1292 => x"81",
          1293 => x"80",
          1294 => x"39",
          1295 => x"70",
          1296 => x"81",
          1297 => x"80",
          1298 => x"80",
          1299 => x"05",
          1300 => x"70",
          1301 => x"04",
          1302 => x"2e",
          1303 => x"72",
          1304 => x"54",
          1305 => x"e0",
          1306 => x"53",
          1307 => x"f8",
          1308 => x"53",
          1309 => x"b8",
          1310 => x"3d",
          1311 => x"3f",
          1312 => x"38",
          1313 => x"0d",
          1314 => x"33",
          1315 => x"8b",
          1316 => x"ff",
          1317 => x"81",
          1318 => x"52",
          1319 => x"13",
          1320 => x"80",
          1321 => x"52",
          1322 => x"13",
          1323 => x"26",
          1324 => x"87",
          1325 => x"38",
          1326 => x"72",
          1327 => x"13",
          1328 => x"13",
          1329 => x"13",
          1330 => x"13",
          1331 => x"13",
          1332 => x"87",
          1333 => x"98",
          1334 => x"9c",
          1335 => x"0c",
          1336 => x"7f",
          1337 => x"7d",
          1338 => x"7d",
          1339 => x"5c",
          1340 => x"b4",
          1341 => x"c0",
          1342 => x"34",
          1343 => x"85",
          1344 => x"5c",
          1345 => x"a4",
          1346 => x"c0",
          1347 => x"23",
          1348 => x"06",
          1349 => x"86",
          1350 => x"84",
          1351 => x"82",
          1352 => x"06",
          1353 => x"bc",
          1354 => x"0d",
          1355 => x"2e",
          1356 => x"3f",
          1357 => x"98",
          1358 => x"81",
          1359 => x"38",
          1360 => x"0d",
          1361 => x"84",
          1362 => x"2c",
          1363 => x"06",
          1364 => x"3f",
          1365 => x"98",
          1366 => x"38",
          1367 => x"54",
          1368 => x"80",
          1369 => x"98",
          1370 => x"ff",
          1371 => x"14",
          1372 => x"71",
          1373 => x"04",
          1374 => x"83",
          1375 => x"53",
          1376 => x"38",
          1377 => x"2a",
          1378 => x"80",
          1379 => x"81",
          1380 => x"81",
          1381 => x"8a",
          1382 => x"71",
          1383 => x"87",
          1384 => x"86",
          1385 => x"72",
          1386 => x"3d",
          1387 => x"06",
          1388 => x"32",
          1389 => x"38",
          1390 => x"80",
          1391 => x"08",
          1392 => x"54",
          1393 => x"3d",
          1394 => x"70",
          1395 => x"f1",
          1396 => x"3d",
          1397 => x"56",
          1398 => x"38",
          1399 => x"81",
          1400 => x"2e",
          1401 => x"08",
          1402 => x"54",
          1403 => x"91",
          1404 => x"e3",
          1405 => x"72",
          1406 => x"81",
          1407 => x"ff",
          1408 => x"70",
          1409 => x"90",
          1410 => x"33",
          1411 => x"84",
          1412 => x"71",
          1413 => x"70",
          1414 => x"53",
          1415 => x"2a",
          1416 => x"b5",
          1417 => x"96",
          1418 => x"70",
          1419 => x"87",
          1420 => x"8a",
          1421 => x"ab",
          1422 => x"f1",
          1423 => x"83",
          1424 => x"08",
          1425 => x"98",
          1426 => x"9e",
          1427 => x"c0",
          1428 => x"87",
          1429 => x"0c",
          1430 => x"bc",
          1431 => x"f1",
          1432 => x"83",
          1433 => x"08",
          1434 => x"c0",
          1435 => x"9e",
          1436 => x"c0",
          1437 => x"d4",
          1438 => x"f1",
          1439 => x"83",
          1440 => x"08",
          1441 => x"f1",
          1442 => x"90",
          1443 => x"52",
          1444 => x"f1",
          1445 => x"90",
          1446 => x"52",
          1447 => x"52",
          1448 => x"87",
          1449 => x"0a",
          1450 => x"83",
          1451 => x"34",
          1452 => x"70",
          1453 => x"70",
          1454 => x"83",
          1455 => x"9e",
          1456 => x"51",
          1457 => x"81",
          1458 => x"0b",
          1459 => x"80",
          1460 => x"2e",
          1461 => x"ea",
          1462 => x"08",
          1463 => x"52",
          1464 => x"71",
          1465 => x"c0",
          1466 => x"06",
          1467 => x"38",
          1468 => x"80",
          1469 => x"81",
          1470 => x"80",
          1471 => x"f1",
          1472 => x"90",
          1473 => x"52",
          1474 => x"52",
          1475 => x"87",
          1476 => x"06",
          1477 => x"38",
          1478 => x"87",
          1479 => x"70",
          1480 => x"f0",
          1481 => x"08",
          1482 => x"70",
          1483 => x"83",
          1484 => x"08",
          1485 => x"51",
          1486 => x"87",
          1487 => x"51",
          1488 => x"81",
          1489 => x"c0",
          1490 => x"83",
          1491 => x"81",
          1492 => x"83",
          1493 => x"83",
          1494 => x"38",
          1495 => x"83",
          1496 => x"38",
          1497 => x"d1",
          1498 => x"85",
          1499 => x"74",
          1500 => x"54",
          1501 => x"33",
          1502 => x"f3",
          1503 => x"f1",
          1504 => x"83",
          1505 => x"38",
          1506 => x"b1",
          1507 => x"83",
          1508 => x"75",
          1509 => x"54",
          1510 => x"51",
          1511 => x"52",
          1512 => x"3f",
          1513 => x"80",
          1514 => x"d0",
          1515 => x"b5",
          1516 => x"8f",
          1517 => x"d9",
          1518 => x"f1",
          1519 => x"75",
          1520 => x"08",
          1521 => x"54",
          1522 => x"da",
          1523 => x"f1",
          1524 => x"83",
          1525 => x"8a",
          1526 => x"04",
          1527 => x"c0",
          1528 => x"b8",
          1529 => x"71",
          1530 => x"52",
          1531 => x"3f",
          1532 => x"0d",
          1533 => x"84",
          1534 => x"84",
          1535 => x"76",
          1536 => x"08",
          1537 => x"fc",
          1538 => x"80",
          1539 => x"83",
          1540 => x"d8",
          1541 => x"c8",
          1542 => x"b3",
          1543 => x"83",
          1544 => x"83",
          1545 => x"51",
          1546 => x"51",
          1547 => x"52",
          1548 => x"3f",
          1549 => x"c0",
          1550 => x"b8",
          1551 => x"71",
          1552 => x"52",
          1553 => x"3f",
          1554 => x"2e",
          1555 => x"db",
          1556 => x"f1",
          1557 => x"84",
          1558 => x"51",
          1559 => x"33",
          1560 => x"d6",
          1561 => x"a7",
          1562 => x"80",
          1563 => x"db",
          1564 => x"f1",
          1565 => x"a9",
          1566 => x"52",
          1567 => x"3f",
          1568 => x"2e",
          1569 => x"f4",
          1570 => x"b1",
          1571 => x"74",
          1572 => x"83",
          1573 => x"51",
          1574 => x"33",
          1575 => x"cd",
          1576 => x"b4",
          1577 => x"51",
          1578 => x"33",
          1579 => x"c7",
          1580 => x"ac",
          1581 => x"51",
          1582 => x"33",
          1583 => x"c1",
          1584 => x"a4",
          1585 => x"51",
          1586 => x"33",
          1587 => x"c1",
          1588 => x"bc",
          1589 => x"51",
          1590 => x"33",
          1591 => x"c1",
          1592 => x"c4",
          1593 => x"51",
          1594 => x"33",
          1595 => x"c1",
          1596 => x"a4",
          1597 => x"87",
          1598 => x"80",
          1599 => x"3d",
          1600 => x"85",
          1601 => x"c2",
          1602 => x"dd",
          1603 => x"3d",
          1604 => x"af",
          1605 => x"dd",
          1606 => x"3d",
          1607 => x"af",
          1608 => x"dd",
          1609 => x"3d",
          1610 => x"af",
          1611 => x"88",
          1612 => x"96",
          1613 => x"87",
          1614 => x"0d",
          1615 => x"5a",
          1616 => x"f2",
          1617 => x"84",
          1618 => x"3d",
          1619 => x"54",
          1620 => x"d2",
          1621 => x"2e",
          1622 => x"84",
          1623 => x"80",
          1624 => x"38",
          1625 => x"18",
          1626 => x"70",
          1627 => x"55",
          1628 => x"ff",
          1629 => x"11",
          1630 => x"84",
          1631 => x"2e",
          1632 => x"a9",
          1633 => x"ff",
          1634 => x"81",
          1635 => x"c0",
          1636 => x"ab",
          1637 => x"76",
          1638 => x"ff",
          1639 => x"e4",
          1640 => x"0d",
          1641 => x"72",
          1642 => x"73",
          1643 => x"8d",
          1644 => x"83",
          1645 => x"ff",
          1646 => x"53",
          1647 => x"3f",
          1648 => x"14",
          1649 => x"38",
          1650 => x"70",
          1651 => x"27",
          1652 => x"e4",
          1653 => x"5a",
          1654 => x"80",
          1655 => x"e4",
          1656 => x"53",
          1657 => x"84",
          1658 => x"73",
          1659 => x"81",
          1660 => x"fe",
          1661 => x"77",
          1662 => x"38",
          1663 => x"55",
          1664 => x"d5",
          1665 => x"0b",
          1666 => x"73",
          1667 => x"d0",
          1668 => x"84",
          1669 => x"f2",
          1670 => x"51",
          1671 => x"08",
          1672 => x"bd",
          1673 => x"80",
          1674 => x"38",
          1675 => x"19",
          1676 => x"75",
          1677 => x"56",
          1678 => x"09",
          1679 => x"84",
          1680 => x"ce",
          1681 => x"08",
          1682 => x"0b",
          1683 => x"83",
          1684 => x"38",
          1685 => x"74",
          1686 => x"2e",
          1687 => x"5a",
          1688 => x"2e",
          1689 => x"5f",
          1690 => x"b8",
          1691 => x"5b",
          1692 => x"81",
          1693 => x"98",
          1694 => x"33",
          1695 => x"98",
          1696 => x"ec",
          1697 => x"53",
          1698 => x"59",
          1699 => x"38",
          1700 => x"81",
          1701 => x"70",
          1702 => x"81",
          1703 => x"2b",
          1704 => x"16",
          1705 => x"38",
          1706 => x"33",
          1707 => x"38",
          1708 => x"d0",
          1709 => x"81",
          1710 => x"70",
          1711 => x"98",
          1712 => x"05",
          1713 => x"33",
          1714 => x"57",
          1715 => x"84",
          1716 => x"57",
          1717 => x"0a",
          1718 => x"2c",
          1719 => x"76",
          1720 => x"16",
          1721 => x"83",
          1722 => x"61",
          1723 => x"08",
          1724 => x"2e",
          1725 => x"bc",
          1726 => x"80",
          1727 => x"81",
          1728 => x"fe",
          1729 => x"76",
          1730 => x"76",
          1731 => x"fd",
          1732 => x"84",
          1733 => x"f4",
          1734 => x"d0",
          1735 => x"34",
          1736 => x"75",
          1737 => x"c8",
          1738 => x"3f",
          1739 => x"76",
          1740 => x"84",
          1741 => x"84",
          1742 => x"79",
          1743 => x"08",
          1744 => x"a8",
          1745 => x"ff",
          1746 => x"93",
          1747 => x"83",
          1748 => x"75",
          1749 => x"34",
          1750 => x"84",
          1751 => x"2e",
          1752 => x"88",
          1753 => x"c8",
          1754 => x"3f",
          1755 => x"ff",
          1756 => x"ff",
          1757 => x"7a",
          1758 => x"7b",
          1759 => x"d0",
          1760 => x"38",
          1761 => x"9e",
          1762 => x"05",
          1763 => x"f9",
          1764 => x"fb",
          1765 => x"3f",
          1766 => x"34",
          1767 => x"81",
          1768 => x"b8",
          1769 => x"d0",
          1770 => x"ff",
          1771 => x"88",
          1772 => x"c8",
          1773 => x"3f",
          1774 => x"ff",
          1775 => x"ff",
          1776 => x"74",
          1777 => x"d0",
          1778 => x"d0",
          1779 => x"27",
          1780 => x"52",
          1781 => x"34",
          1782 => x"b3",
          1783 => x"81",
          1784 => x"57",
          1785 => x"84",
          1786 => x"76",
          1787 => x"33",
          1788 => x"d0",
          1789 => x"d0",
          1790 => x"26",
          1791 => x"d0",
          1792 => x"56",
          1793 => x"15",
          1794 => x"98",
          1795 => x"06",
          1796 => x"ef",
          1797 => x"51",
          1798 => x"33",
          1799 => x"d0",
          1800 => x"77",
          1801 => x"08",
          1802 => x"74",
          1803 => x"05",
          1804 => x"5d",
          1805 => x"38",
          1806 => x"ff",
          1807 => x"29",
          1808 => x"84",
          1809 => x"75",
          1810 => x"7b",
          1811 => x"84",
          1812 => x"ff",
          1813 => x"29",
          1814 => x"84",
          1815 => x"79",
          1816 => x"81",
          1817 => x"08",
          1818 => x"3f",
          1819 => x"0a",
          1820 => x"33",
          1821 => x"a7",
          1822 => x"33",
          1823 => x"84",
          1824 => x"b0",
          1825 => x"05",
          1826 => x"81",
          1827 => x"a4",
          1828 => x"84",
          1829 => x"b0",
          1830 => x"51",
          1831 => x"81",
          1832 => x"84",
          1833 => x"80",
          1834 => x"10",
          1835 => x"57",
          1836 => x"82",
          1837 => x"05",
          1838 => x"e7",
          1839 => x"0c",
          1840 => x"83",
          1841 => x"41",
          1842 => x"08",
          1843 => x"f2",
          1844 => x"bc",
          1845 => x"80",
          1846 => x"b8",
          1847 => x"d0",
          1848 => x"38",
          1849 => x"ff",
          1850 => x"52",
          1851 => x"d4",
          1852 => x"8a",
          1853 => x"56",
          1854 => x"ff",
          1855 => x"e0",
          1856 => x"84",
          1857 => x"a4",
          1858 => x"80",
          1859 => x"33",
          1860 => x"d4",
          1861 => x"c2",
          1862 => x"51",
          1863 => x"08",
          1864 => x"84",
          1865 => x"84",
          1866 => x"55",
          1867 => x"ff",
          1868 => x"a8",
          1869 => x"7b",
          1870 => x"04",
          1871 => x"06",
          1872 => x"38",
          1873 => x"78",
          1874 => x"77",
          1875 => x"08",
          1876 => x"84",
          1877 => x"98",
          1878 => x"5b",
          1879 => x"84",
          1880 => x"ad",
          1881 => x"98",
          1882 => x"33",
          1883 => x"f3",
          1884 => x"88",
          1885 => x"80",
          1886 => x"98",
          1887 => x"55",
          1888 => x"d4",
          1889 => x"e2",
          1890 => x"80",
          1891 => x"a4",
          1892 => x"ff",
          1893 => x"57",
          1894 => x"c8",
          1895 => x"b2",
          1896 => x"80",
          1897 => x"a4",
          1898 => x"fe",
          1899 => x"33",
          1900 => x"76",
          1901 => x"81",
          1902 => x"70",
          1903 => x"57",
          1904 => x"fe",
          1905 => x"81",
          1906 => x"f2",
          1907 => x"76",
          1908 => x"70",
          1909 => x"a1",
          1910 => x"1c",
          1911 => x"ff",
          1912 => x"a8",
          1913 => x"e1",
          1914 => x"a8",
          1915 => x"5a",
          1916 => x"a4",
          1917 => x"81",
          1918 => x"75",
          1919 => x"80",
          1920 => x"98",
          1921 => x"5c",
          1922 => x"77",
          1923 => x"ff",
          1924 => x"f1",
          1925 => x"88",
          1926 => x"80",
          1927 => x"98",
          1928 => x"41",
          1929 => x"d4",
          1930 => x"9a",
          1931 => x"80",
          1932 => x"a4",
          1933 => x"ff",
          1934 => x"fc",
          1935 => x"38",
          1936 => x"b8",
          1937 => x"b8",
          1938 => x"53",
          1939 => x"3f",
          1940 => x"33",
          1941 => x"38",
          1942 => x"ff",
          1943 => x"52",
          1944 => x"d4",
          1945 => x"a2",
          1946 => x"5b",
          1947 => x"ff",
          1948 => x"e1",
          1949 => x"f2",
          1950 => x"a5",
          1951 => x"ef",
          1952 => x"c8",
          1953 => x"58",
          1954 => x"0a",
          1955 => x"2c",
          1956 => x"76",
          1957 => x"33",
          1958 => x"81",
          1959 => x"7a",
          1960 => x"83",
          1961 => x"38",
          1962 => x"08",
          1963 => x"18",
          1964 => x"80",
          1965 => x"d0",
          1966 => x"38",
          1967 => x"f2",
          1968 => x"80",
          1969 => x"b4",
          1970 => x"51",
          1971 => x"ff",
          1972 => x"25",
          1973 => x"51",
          1974 => x"08",
          1975 => x"08",
          1976 => x"52",
          1977 => x"0b",
          1978 => x"33",
          1979 => x"97",
          1980 => x"51",
          1981 => x"08",
          1982 => x"84",
          1983 => x"a6",
          1984 => x"05",
          1985 => x"81",
          1986 => x"34",
          1987 => x"0b",
          1988 => x"e4",
          1989 => x"ff",
          1990 => x"84",
          1991 => x"81",
          1992 => x"7b",
          1993 => x"70",
          1994 => x"84",
          1995 => x"74",
          1996 => x"c8",
          1997 => x"3f",
          1998 => x"ff",
          1999 => x"52",
          2000 => x"d0",
          2001 => x"d0",
          2002 => x"c7",
          2003 => x"84",
          2004 => x"84",
          2005 => x"05",
          2006 => x"b6",
          2007 => x"84",
          2008 => x"58",
          2009 => x"a7",
          2010 => x"51",
          2011 => x"08",
          2012 => x"84",
          2013 => x"a5",
          2014 => x"05",
          2015 => x"81",
          2016 => x"80",
          2017 => x"70",
          2018 => x"fc",
          2019 => x"56",
          2020 => x"08",
          2021 => x"10",
          2022 => x"57",
          2023 => x"38",
          2024 => x"a8",
          2025 => x"05",
          2026 => x"79",
          2027 => x"d4",
          2028 => x"f8",
          2029 => x"51",
          2030 => x"08",
          2031 => x"83",
          2032 => x"3f",
          2033 => x"0b",
          2034 => x"e4",
          2035 => x"77",
          2036 => x"c9",
          2037 => x"a5",
          2038 => x"5c",
          2039 => x"f8",
          2040 => x"84",
          2041 => x"08",
          2042 => x"38",
          2043 => x"cc",
          2044 => x"0b",
          2045 => x"38",
          2046 => x"1b",
          2047 => x"ff",
          2048 => x"10",
          2049 => x"40",
          2050 => x"82",
          2051 => x"05",
          2052 => x"da",
          2053 => x"0c",
          2054 => x"83",
          2055 => x"41",
          2056 => x"ff",
          2057 => x"38",
          2058 => x"06",
          2059 => x"f9",
          2060 => x"51",
          2061 => x"33",
          2062 => x"57",
          2063 => x"0b",
          2064 => x"74",
          2065 => x"d4",
          2066 => x"83",
          2067 => x"52",
          2068 => x"b8",
          2069 => x"33",
          2070 => x"70",
          2071 => x"ff",
          2072 => x"f2",
          2073 => x"f2",
          2074 => x"cc",
          2075 => x"eb",
          2076 => x"02",
          2077 => x"80",
          2078 => x"26",
          2079 => x"8b",
          2080 => x"72",
          2081 => x"a0",
          2082 => x"5e",
          2083 => x"76",
          2084 => x"34",
          2085 => x"f8",
          2086 => x"98",
          2087 => x"2b",
          2088 => x"56",
          2089 => x"74",
          2090 => x"70",
          2091 => x"ee",
          2092 => x"f8",
          2093 => x"78",
          2094 => x"e0",
          2095 => x"56",
          2096 => x"90",
          2097 => x"0b",
          2098 => x"11",
          2099 => x"11",
          2100 => x"86",
          2101 => x"33",
          2102 => x"33",
          2103 => x"22",
          2104 => x"29",
          2105 => x"5d",
          2106 => x"31",
          2107 => x"7e",
          2108 => x"7a",
          2109 => x"06",
          2110 => x"57",
          2111 => x"83",
          2112 => x"70",
          2113 => x"06",
          2114 => x"78",
          2115 => x"c1",
          2116 => x"34",
          2117 => x"05",
          2118 => x"80",
          2119 => x"b6",
          2120 => x"b6",
          2121 => x"f8",
          2122 => x"5d",
          2123 => x"27",
          2124 => x"73",
          2125 => x"5a",
          2126 => x"38",
          2127 => x"0b",
          2128 => x"33",
          2129 => x"71",
          2130 => x"56",
          2131 => x"ae",
          2132 => x"38",
          2133 => x"06",
          2134 => x"33",
          2135 => x"80",
          2136 => x"86",
          2137 => x"d8",
          2138 => x"d7",
          2139 => x"92",
          2140 => x"75",
          2141 => x"58",
          2142 => x"8b",
          2143 => x"29",
          2144 => x"74",
          2145 => x"83",
          2146 => x"70",
          2147 => x"55",
          2148 => x"29",
          2149 => x"06",
          2150 => x"83",
          2151 => x"f2",
          2152 => x"fe",
          2153 => x"80",
          2154 => x"73",
          2155 => x"86",
          2156 => x"34",
          2157 => x"98",
          2158 => x"86",
          2159 => x"80",
          2160 => x"52",
          2161 => x"87",
          2162 => x"56",
          2163 => x"84",
          2164 => x"08",
          2165 => x"51",
          2166 => x"cc",
          2167 => x"53",
          2168 => x"08",
          2169 => x"75",
          2170 => x"34",
          2171 => x"3d",
          2172 => x"b8",
          2173 => x"af",
          2174 => x"33",
          2175 => x"81",
          2176 => x"84",
          2177 => x"83",
          2178 => x"86",
          2179 => x"22",
          2180 => x"05",
          2181 => x"ea",
          2182 => x"2e",
          2183 => x"76",
          2184 => x"83",
          2185 => x"ff",
          2186 => x"55",
          2187 => x"19",
          2188 => x"f8",
          2189 => x"84",
          2190 => x"74",
          2191 => x"33",
          2192 => x"72",
          2193 => x"b6",
          2194 => x"33",
          2195 => x"05",
          2196 => x"34",
          2197 => x"27",
          2198 => x"38",
          2199 => x"15",
          2200 => x"34",
          2201 => x"81",
          2202 => x"38",
          2203 => x"75",
          2204 => x"81",
          2205 => x"54",
          2206 => x"72",
          2207 => x"33",
          2208 => x"55",
          2209 => x"b0",
          2210 => x"ff",
          2211 => x"54",
          2212 => x"97",
          2213 => x"53",
          2214 => x"81",
          2215 => x"55",
          2216 => x"81",
          2217 => x"d7",
          2218 => x"5a",
          2219 => x"53",
          2220 => x"0d",
          2221 => x"f8",
          2222 => x"84",
          2223 => x"7a",
          2224 => x"fe",
          2225 => x"05",
          2226 => x"75",
          2227 => x"73",
          2228 => x"33",
          2229 => x"56",
          2230 => x"ae",
          2231 => x"b6",
          2232 => x"a0",
          2233 => x"70",
          2234 => x"72",
          2235 => x"e0",
          2236 => x"05",
          2237 => x"38",
          2238 => x"d8",
          2239 => x"f8",
          2240 => x"19",
          2241 => x"59",
          2242 => x"02",
          2243 => x"70",
          2244 => x"83",
          2245 => x"84",
          2246 => x"86",
          2247 => x"0b",
          2248 => x"04",
          2249 => x"f8",
          2250 => x"52",
          2251 => x"51",
          2252 => x"84",
          2253 => x"83",
          2254 => x"09",
          2255 => x"53",
          2256 => x"39",
          2257 => x"b6",
          2258 => x"70",
          2259 => x"83",
          2260 => x"e4",
          2261 => x"95",
          2262 => x"9f",
          2263 => x"70",
          2264 => x"b8",
          2265 => x"f8",
          2266 => x"33",
          2267 => x"25",
          2268 => x"95",
          2269 => x"86",
          2270 => x"95",
          2271 => x"d7",
          2272 => x"25",
          2273 => x"83",
          2274 => x"3d",
          2275 => x"b1",
          2276 => x"c3",
          2277 => x"f8",
          2278 => x"84",
          2279 => x"2a",
          2280 => x"f0",
          2281 => x"f2",
          2282 => x"84",
          2283 => x"83",
          2284 => x"07",
          2285 => x"0b",
          2286 => x"04",
          2287 => x"51",
          2288 => x"83",
          2289 => x"07",
          2290 => x"39",
          2291 => x"80",
          2292 => x"0d",
          2293 => x"06",
          2294 => x"34",
          2295 => x"87",
          2296 => x"ff",
          2297 => x"fd",
          2298 => x"90",
          2299 => x"33",
          2300 => x"83",
          2301 => x"f8",
          2302 => x"51",
          2303 => x"39",
          2304 => x"51",
          2305 => x"39",
          2306 => x"80",
          2307 => x"34",
          2308 => x"81",
          2309 => x"f8",
          2310 => x"90",
          2311 => x"51",
          2312 => x"39",
          2313 => x"80",
          2314 => x"34",
          2315 => x"81",
          2316 => x"f8",
          2317 => x"90",
          2318 => x"f8",
          2319 => x"90",
          2320 => x"70",
          2321 => x"f3",
          2322 => x"84",
          2323 => x"94",
          2324 => x"95",
          2325 => x"5f",
          2326 => x"a1",
          2327 => x"81",
          2328 => x"da",
          2329 => x"7a",
          2330 => x"92",
          2331 => x"3d",
          2332 => x"06",
          2333 => x"34",
          2334 => x"0b",
          2335 => x"f8",
          2336 => x"23",
          2337 => x"84",
          2338 => x"33",
          2339 => x"83",
          2340 => x"7d",
          2341 => x"b6",
          2342 => x"7b",
          2343 => x"95",
          2344 => x"84",
          2345 => x"dc",
          2346 => x"a8",
          2347 => x"83",
          2348 => x"58",
          2349 => x"e5",
          2350 => x"53",
          2351 => x"81",
          2352 => x"33",
          2353 => x"79",
          2354 => x"53",
          2355 => x"ec",
          2356 => x"84",
          2357 => x"7a",
          2358 => x"ff",
          2359 => x"34",
          2360 => x"83",
          2361 => x"23",
          2362 => x"0d",
          2363 => x"81",
          2364 => x"83",
          2365 => x"95",
          2366 => x"83",
          2367 => x"84",
          2368 => x"51",
          2369 => x"f6",
          2370 => x"84",
          2371 => x"83",
          2372 => x"98",
          2373 => x"70",
          2374 => x"f9",
          2375 => x"05",
          2376 => x"95",
          2377 => x"29",
          2378 => x"f8",
          2379 => x"7c",
          2380 => x"83",
          2381 => x"57",
          2382 => x"75",
          2383 => x"24",
          2384 => x"85",
          2385 => x"84",
          2386 => x"83",
          2387 => x"55",
          2388 => x"86",
          2389 => x"d8",
          2390 => x"92",
          2391 => x"56",
          2392 => x"83",
          2393 => x"58",
          2394 => x"b0",
          2395 => x"70",
          2396 => x"83",
          2397 => x"57",
          2398 => x"33",
          2399 => x"70",
          2400 => x"26",
          2401 => x"58",
          2402 => x"72",
          2403 => x"33",
          2404 => x"b6",
          2405 => x"fb",
          2406 => x"89",
          2407 => x"38",
          2408 => x"8a",
          2409 => x"81",
          2410 => x"0b",
          2411 => x"83",
          2412 => x"e0",
          2413 => x"09",
          2414 => x"76",
          2415 => x"13",
          2416 => x"83",
          2417 => x"51",
          2418 => x"ff",
          2419 => x"38",
          2420 => x"34",
          2421 => x"f9",
          2422 => x"0c",
          2423 => x"2e",
          2424 => x"f8",
          2425 => x"ff",
          2426 => x"72",
          2427 => x"51",
          2428 => x"70",
          2429 => x"73",
          2430 => x"f8",
          2431 => x"83",
          2432 => x"ef",
          2433 => x"75",
          2434 => x"e6",
          2435 => x"84",
          2436 => x"2e",
          2437 => x"82",
          2438 => x"78",
          2439 => x"2e",
          2440 => x"8f",
          2441 => x"94",
          2442 => x"29",
          2443 => x"19",
          2444 => x"84",
          2445 => x"83",
          2446 => x"5a",
          2447 => x"18",
          2448 => x"29",
          2449 => x"33",
          2450 => x"84",
          2451 => x"83",
          2452 => x"72",
          2453 => x"59",
          2454 => x"1f",
          2455 => x"42",
          2456 => x"84",
          2457 => x"38",
          2458 => x"34",
          2459 => x"3d",
          2460 => x"38",
          2461 => x"b8",
          2462 => x"2e",
          2463 => x"e0",
          2464 => x"94",
          2465 => x"29",
          2466 => x"19",
          2467 => x"84",
          2468 => x"83",
          2469 => x"41",
          2470 => x"1f",
          2471 => x"29",
          2472 => x"86",
          2473 => x"d8",
          2474 => x"92",
          2475 => x"29",
          2476 => x"f8",
          2477 => x"34",
          2478 => x"41",
          2479 => x"83",
          2480 => x"e4",
          2481 => x"2e",
          2482 => x"81",
          2483 => x"fd",
          2484 => x"34",
          2485 => x"3d",
          2486 => x"38",
          2487 => x"d0",
          2488 => x"59",
          2489 => x"84",
          2490 => x"06",
          2491 => x"34",
          2492 => x"3d",
          2493 => x"38",
          2494 => x"b6",
          2495 => x"f8",
          2496 => x"40",
          2497 => x"a7",
          2498 => x"33",
          2499 => x"22",
          2500 => x"56",
          2501 => x"f8",
          2502 => x"57",
          2503 => x"80",
          2504 => x"81",
          2505 => x"f8",
          2506 => x"42",
          2507 => x"60",
          2508 => x"58",
          2509 => x"ea",
          2510 => x"34",
          2511 => x"83",
          2512 => x"83",
          2513 => x"86",
          2514 => x"22",
          2515 => x"70",
          2516 => x"33",
          2517 => x"2e",
          2518 => x"ff",
          2519 => x"76",
          2520 => x"90",
          2521 => x"80",
          2522 => x"84",
          2523 => x"e7",
          2524 => x"80",
          2525 => x"0d",
          2526 => x"cc",
          2527 => x"cd",
          2528 => x"ce",
          2529 => x"80",
          2530 => x"0d",
          2531 => x"06",
          2532 => x"84",
          2533 => x"83",
          2534 => x"72",
          2535 => x"05",
          2536 => x"7b",
          2537 => x"83",
          2538 => x"42",
          2539 => x"38",
          2540 => x"56",
          2541 => x"f8",
          2542 => x"81",
          2543 => x"72",
          2544 => x"80",
          2545 => x"84",
          2546 => x"83",
          2547 => x"5a",
          2548 => x"96",
          2549 => x"71",
          2550 => x"90",
          2551 => x"84",
          2552 => x"83",
          2553 => x"72",
          2554 => x"59",
          2555 => x"b6",
          2556 => x"06",
          2557 => x"38",
          2558 => x"d0",
          2559 => x"95",
          2560 => x"ff",
          2561 => x"39",
          2562 => x"bd",
          2563 => x"95",
          2564 => x"7e",
          2565 => x"75",
          2566 => x"10",
          2567 => x"04",
          2568 => x"52",
          2569 => x"84",
          2570 => x"83",
          2571 => x"70",
          2572 => x"70",
          2573 => x"86",
          2574 => x"22",
          2575 => x"83",
          2576 => x"46",
          2577 => x"81",
          2578 => x"81",
          2579 => x"81",
          2580 => x"58",
          2581 => x"a0",
          2582 => x"83",
          2583 => x"72",
          2584 => x"a0",
          2585 => x"f8",
          2586 => x"5e",
          2587 => x"80",
          2588 => x"81",
          2589 => x"f8",
          2590 => x"44",
          2591 => x"84",
          2592 => x"70",
          2593 => x"26",
          2594 => x"58",
          2595 => x"75",
          2596 => x"81",
          2597 => x"f7",
          2598 => x"b6",
          2599 => x"81",
          2600 => x"81",
          2601 => x"5b",
          2602 => x"33",
          2603 => x"b6",
          2604 => x"f8",
          2605 => x"41",
          2606 => x"1c",
          2607 => x"29",
          2608 => x"86",
          2609 => x"d8",
          2610 => x"92",
          2611 => x"29",
          2612 => x"f8",
          2613 => x"60",
          2614 => x"58",
          2615 => x"83",
          2616 => x"0b",
          2617 => x"b8",
          2618 => x"f8",
          2619 => x"19",
          2620 => x"70",
          2621 => x"f9",
          2622 => x"34",
          2623 => x"3d",
          2624 => x"5b",
          2625 => x"83",
          2626 => x"83",
          2627 => x"5c",
          2628 => x"9c",
          2629 => x"ff",
          2630 => x"80",
          2631 => x"33",
          2632 => x"e5",
          2633 => x"02",
          2634 => x"b8",
          2635 => x"96",
          2636 => x"33",
          2637 => x"b6",
          2638 => x"5b",
          2639 => x"33",
          2640 => x"33",
          2641 => x"84",
          2642 => x"a0",
          2643 => x"83",
          2644 => x"72",
          2645 => x"78",
          2646 => x"94",
          2647 => x"83",
          2648 => x"80",
          2649 => x"81",
          2650 => x"f8",
          2651 => x"5f",
          2652 => x"84",
          2653 => x"81",
          2654 => x"90",
          2655 => x"77",
          2656 => x"83",
          2657 => x"e0",
          2658 => x"80",
          2659 => x"33",
          2660 => x"81",
          2661 => x"b8",
          2662 => x"b8",
          2663 => x"b8",
          2664 => x"b8",
          2665 => x"23",
          2666 => x"84",
          2667 => x"84",
          2668 => x"84",
          2669 => x"b7",
          2670 => x"93",
          2671 => x"86",
          2672 => x"83",
          2673 => x"f8",
          2674 => x"83",
          2675 => x"57",
          2676 => x"ff",
          2677 => x"ff",
          2678 => x"05",
          2679 => x"76",
          2680 => x"ce",
          2681 => x"b7",
          2682 => x"06",
          2683 => x"77",
          2684 => x"33",
          2685 => x"38",
          2686 => x"5f",
          2687 => x"5e",
          2688 => x"f8",
          2689 => x"71",
          2690 => x"06",
          2691 => x"f8",
          2692 => x"e5",
          2693 => x"38",
          2694 => x"81",
          2695 => x"57",
          2696 => x"75",
          2697 => x"80",
          2698 => x"94",
          2699 => x"7b",
          2700 => x"56",
          2701 => x"39",
          2702 => x"f8",
          2703 => x"05",
          2704 => x"38",
          2705 => x"34",
          2706 => x"40",
          2707 => x"f8",
          2708 => x"71",
          2709 => x"06",
          2710 => x"f8",
          2711 => x"e5",
          2712 => x"38",
          2713 => x"2e",
          2714 => x"b6",
          2715 => x"f8",
          2716 => x"a7",
          2717 => x"43",
          2718 => x"70",
          2719 => x"08",
          2720 => x"5d",
          2721 => x"bf",
          2722 => x"fb",
          2723 => x"79",
          2724 => x"b8",
          2725 => x"06",
          2726 => x"e9",
          2727 => x"33",
          2728 => x"84",
          2729 => x"5d",
          2730 => x"11",
          2731 => x"38",
          2732 => x"fb",
          2733 => x"76",
          2734 => x"b9",
          2735 => x"05",
          2736 => x"41",
          2737 => x"57",
          2738 => x"39",
          2739 => x"3f",
          2740 => x"57",
          2741 => x"10",
          2742 => x"5a",
          2743 => x"3f",
          2744 => x"b7",
          2745 => x"82",
          2746 => x"7d",
          2747 => x"22",
          2748 => x"57",
          2749 => x"d5",
          2750 => x"e5",
          2751 => x"38",
          2752 => x"81",
          2753 => x"05",
          2754 => x"33",
          2755 => x"43",
          2756 => x"27",
          2757 => x"92",
          2758 => x"58",
          2759 => x"57",
          2760 => x"d8",
          2761 => x"27",
          2762 => x"f8",
          2763 => x"e5",
          2764 => x"38",
          2765 => x"33",
          2766 => x"38",
          2767 => x"33",
          2768 => x"33",
          2769 => x"80",
          2770 => x"71",
          2771 => x"06",
          2772 => x"59",
          2773 => x"38",
          2774 => x"31",
          2775 => x"38",
          2776 => x"27",
          2777 => x"83",
          2778 => x"70",
          2779 => x"8e",
          2780 => x"76",
          2781 => x"56",
          2782 => x"ff",
          2783 => x"80",
          2784 => x"77",
          2785 => x"71",
          2786 => x"86",
          2787 => x"80",
          2788 => x"06",
          2789 => x"5c",
          2790 => x"97",
          2791 => x"5f",
          2792 => x"81",
          2793 => x"58",
          2794 => x"81",
          2795 => x"d7",
          2796 => x"5e",
          2797 => x"e0",
          2798 => x"1f",
          2799 => x"76",
          2800 => x"81",
          2801 => x"d8",
          2802 => x"29",
          2803 => x"26",
          2804 => x"b7",
          2805 => x"e0",
          2806 => x"51",
          2807 => x"0b",
          2808 => x"b7",
          2809 => x"78",
          2810 => x"56",
          2811 => x"be",
          2812 => x"81",
          2813 => x"43",
          2814 => x"38",
          2815 => x"26",
          2816 => x"56",
          2817 => x"76",
          2818 => x"f5",
          2819 => x"90",
          2820 => x"11",
          2821 => x"80",
          2822 => x"75",
          2823 => x"76",
          2824 => x"70",
          2825 => x"88",
          2826 => x"52",
          2827 => x"80",
          2828 => x"76",
          2829 => x"26",
          2830 => x"b6",
          2831 => x"06",
          2832 => x"22",
          2833 => x"59",
          2834 => x"78",
          2835 => x"57",
          2836 => x"76",
          2837 => x"33",
          2838 => x"0b",
          2839 => x"81",
          2840 => x"76",
          2841 => x"e0",
          2842 => x"5a",
          2843 => x"d6",
          2844 => x"81",
          2845 => x"83",
          2846 => x"71",
          2847 => x"2a",
          2848 => x"2e",
          2849 => x"0b",
          2850 => x"81",
          2851 => x"83",
          2852 => x"e0",
          2853 => x"33",
          2854 => x"22",
          2855 => x"5d",
          2856 => x"87",
          2857 => x"81",
          2858 => x"f4",
          2859 => x"fd",
          2860 => x"90",
          2861 => x"81",
          2862 => x"f8",
          2863 => x"33",
          2864 => x"83",
          2865 => x"90",
          2866 => x"75",
          2867 => x"80",
          2868 => x"18",
          2869 => x"a4",
          2870 => x"06",
          2871 => x"8f",
          2872 => x"06",
          2873 => x"34",
          2874 => x"81",
          2875 => x"83",
          2876 => x"f8",
          2877 => x"07",
          2878 => x"d7",
          2879 => x"06",
          2880 => x"34",
          2881 => x"81",
          2882 => x"f8",
          2883 => x"90",
          2884 => x"75",
          2885 => x"83",
          2886 => x"07",
          2887 => x"8f",
          2888 => x"06",
          2889 => x"ff",
          2890 => x"07",
          2891 => x"ef",
          2892 => x"07",
          2893 => x"df",
          2894 => x"06",
          2895 => x"90",
          2896 => x"33",
          2897 => x"83",
          2898 => x"0b",
          2899 => x"51",
          2900 => x"b8",
          2901 => x"b8",
          2902 => x"b8",
          2903 => x"23",
          2904 => x"c7",
          2905 => x"80",
          2906 => x"0d",
          2907 => x"f8",
          2908 => x"ff",
          2909 => x"e8",
          2910 => x"05",
          2911 => x"e4",
          2912 => x"84",
          2913 => x"e4",
          2914 => x"9c",
          2915 => x"34",
          2916 => x"81",
          2917 => x"34",
          2918 => x"80",
          2919 => x"23",
          2920 => x"39",
          2921 => x"52",
          2922 => x"95",
          2923 => x"05",
          2924 => x"f8",
          2925 => x"fb",
          2926 => x"eb",
          2927 => x"95",
          2928 => x"2c",
          2929 => x"39",
          2930 => x"b6",
          2931 => x"eb",
          2932 => x"e3",
          2933 => x"70",
          2934 => x"40",
          2935 => x"33",
          2936 => x"11",
          2937 => x"c0",
          2938 => x"b6",
          2939 => x"5c",
          2940 => x"f8",
          2941 => x"81",
          2942 => x"74",
          2943 => x"83",
          2944 => x"29",
          2945 => x"f6",
          2946 => x"5d",
          2947 => x"83",
          2948 => x"80",
          2949 => x"d7",
          2950 => x"38",
          2951 => x"23",
          2952 => x"57",
          2953 => x"b6",
          2954 => x"ec",
          2955 => x"94",
          2956 => x"92",
          2957 => x"26",
          2958 => x"7e",
          2959 => x"5e",
          2960 => x"5b",
          2961 => x"06",
          2962 => x"1d",
          2963 => x"ec",
          2964 => x"e0",
          2965 => x"1e",
          2966 => x"76",
          2967 => x"81",
          2968 => x"d8",
          2969 => x"29",
          2970 => x"27",
          2971 => x"5e",
          2972 => x"81",
          2973 => x"58",
          2974 => x"81",
          2975 => x"d7",
          2976 => x"5d",
          2977 => x"eb",
          2978 => x"5c",
          2979 => x"83",
          2980 => x"83",
          2981 => x"5f",
          2982 => x"eb",
          2983 => x"81",
          2984 => x"76",
          2985 => x"83",
          2986 => x"ff",
          2987 => x"38",
          2988 => x"84",
          2989 => x"ff",
          2990 => x"eb",
          2991 => x"95",
          2992 => x"33",
          2993 => x"11",
          2994 => x"ca",
          2995 => x"81",
          2996 => x"83",
          2997 => x"83",
          2998 => x"57",
          2999 => x"b8",
          3000 => x"75",
          3001 => x"ff",
          3002 => x"fc",
          3003 => x"83",
          3004 => x"7d",
          3005 => x"38",
          3006 => x"83",
          3007 => x"59",
          3008 => x"80",
          3009 => x"f8",
          3010 => x"34",
          3011 => x"39",
          3012 => x"92",
          3013 => x"f8",
          3014 => x"f8",
          3015 => x"83",
          3016 => x"0b",
          3017 => x"83",
          3018 => x"e0",
          3019 => x"f6",
          3020 => x"0d",
          3021 => x"33",
          3022 => x"73",
          3023 => x"b8",
          3024 => x"52",
          3025 => x"84",
          3026 => x"f3",
          3027 => x"ff",
          3028 => x"ff",
          3029 => x"55",
          3030 => x"38",
          3031 => x"34",
          3032 => x"8f",
          3033 => x"54",
          3034 => x"73",
          3035 => x"09",
          3036 => x"72",
          3037 => x"54",
          3038 => x"38",
          3039 => x"70",
          3040 => x"79",
          3041 => x"d8",
          3042 => x"94",
          3043 => x"a0",
          3044 => x"59",
          3045 => x"ff",
          3046 => x"59",
          3047 => x"38",
          3048 => x"80",
          3049 => x"0c",
          3050 => x"80",
          3051 => x"08",
          3052 => x"81",
          3053 => x"81",
          3054 => x"83",
          3055 => x"06",
          3056 => x"55",
          3057 => x"81",
          3058 => x"f6",
          3059 => x"5a",
          3060 => x"75",
          3061 => x"84",
          3062 => x"81",
          3063 => x"89",
          3064 => x"8c",
          3065 => x"58",
          3066 => x"73",
          3067 => x"32",
          3068 => x"80",
          3069 => x"f6",
          3070 => x"72",
          3071 => x"83",
          3072 => x"bd",
          3073 => x"be",
          3074 => x"f6",
          3075 => x"5e",
          3076 => x"74",
          3077 => x"ac",
          3078 => x"82",
          3079 => x"72",
          3080 => x"ac",
          3081 => x"74",
          3082 => x"2e",
          3083 => x"53",
          3084 => x"81",
          3085 => x"84",
          3086 => x"54",
          3087 => x"f6",
          3088 => x"98",
          3089 => x"83",
          3090 => x"9c",
          3091 => x"16",
          3092 => x"76",
          3093 => x"bf",
          3094 => x"9e",
          3095 => x"38",
          3096 => x"5a",
          3097 => x"54",
          3098 => x"14",
          3099 => x"7d",
          3100 => x"83",
          3101 => x"2e",
          3102 => x"ea",
          3103 => x"f6",
          3104 => x"77",
          3105 => x"17",
          3106 => x"76",
          3107 => x"83",
          3108 => x"82",
          3109 => x"38",
          3110 => x"fc",
          3111 => x"80",
          3112 => x"2e",
          3113 => x"06",
          3114 => x"ed",
          3115 => x"79",
          3116 => x"75",
          3117 => x"a1",
          3118 => x"17",
          3119 => x"fe",
          3120 => x"57",
          3121 => x"e1",
          3122 => x"05",
          3123 => x"f2",
          3124 => x"78",
          3125 => x"b8",
          3126 => x"7d",
          3127 => x"ff",
          3128 => x"ff",
          3129 => x"38",
          3130 => x"54",
          3131 => x"82",
          3132 => x"07",
          3133 => x"83",
          3134 => x"78",
          3135 => x"72",
          3136 => x"70",
          3137 => x"ba",
          3138 => x"54",
          3139 => x"b6",
          3140 => x"9a",
          3141 => x"f9",
          3142 => x"82",
          3143 => x"e4",
          3144 => x"34",
          3145 => x"81",
          3146 => x"14",
          3147 => x"ac",
          3148 => x"83",
          3149 => x"f6",
          3150 => x"a2",
          3151 => x"ff",
          3152 => x"96",
          3153 => x"81",
          3154 => x"ff",
          3155 => x"06",
          3156 => x"81",
          3157 => x"54",
          3158 => x"87",
          3159 => x"0c",
          3160 => x"39",
          3161 => x"f9",
          3162 => x"73",
          3163 => x"38",
          3164 => x"83",
          3165 => x"83",
          3166 => x"33",
          3167 => x"5e",
          3168 => x"82",
          3169 => x"7a",
          3170 => x"79",
          3171 => x"38",
          3172 => x"f0",
          3173 => x"b6",
          3174 => x"81",
          3175 => x"59",
          3176 => x"da",
          3177 => x"54",
          3178 => x"f7",
          3179 => x"08",
          3180 => x"83",
          3181 => x"b6",
          3182 => x"11",
          3183 => x"38",
          3184 => x"73",
          3185 => x"80",
          3186 => x"83",
          3187 => x"70",
          3188 => x"80",
          3189 => x"83",
          3190 => x"39",
          3191 => x"3f",
          3192 => x"fc",
          3193 => x"f6",
          3194 => x"0b",
          3195 => x"33",
          3196 => x"81",
          3197 => x"04",
          3198 => x"f0",
          3199 => x"82",
          3200 => x"80",
          3201 => x"f0",
          3202 => x"34",
          3203 => x"87",
          3204 => x"08",
          3205 => x"c0",
          3206 => x"9c",
          3207 => x"81",
          3208 => x"56",
          3209 => x"81",
          3210 => x"a4",
          3211 => x"80",
          3212 => x"80",
          3213 => x"80",
          3214 => x"9c",
          3215 => x"55",
          3216 => x"33",
          3217 => x"70",
          3218 => x"2e",
          3219 => x"55",
          3220 => x"71",
          3221 => x"57",
          3222 => x"81",
          3223 => x"74",
          3224 => x"e4",
          3225 => x"84",
          3226 => x"fa",
          3227 => x"05",
          3228 => x"f0",
          3229 => x"80",
          3230 => x"55",
          3231 => x"90",
          3232 => x"90",
          3233 => x"86",
          3234 => x"74",
          3235 => x"51",
          3236 => x"f2",
          3237 => x"15",
          3238 => x"34",
          3239 => x"f0",
          3240 => x"87",
          3241 => x"98",
          3242 => x"38",
          3243 => x"08",
          3244 => x"71",
          3245 => x"98",
          3246 => x"27",
          3247 => x"2e",
          3248 => x"08",
          3249 => x"98",
          3250 => x"08",
          3251 => x"14",
          3252 => x"52",
          3253 => x"ff",
          3254 => x"08",
          3255 => x"52",
          3256 => x"06",
          3257 => x"38",
          3258 => x"d4",
          3259 => x"56",
          3260 => x"84",
          3261 => x"27",
          3262 => x"33",
          3263 => x"71",
          3264 => x"0c",
          3265 => x"b8",
          3266 => x"51",
          3267 => x"84",
          3268 => x"0b",
          3269 => x"87",
          3270 => x"2a",
          3271 => x"15",
          3272 => x"15",
          3273 => x"15",
          3274 => x"f2",
          3275 => x"13",
          3276 => x"97",
          3277 => x"72",
          3278 => x"26",
          3279 => x"74",
          3280 => x"55",
          3281 => x"f2",
          3282 => x"15",
          3283 => x"34",
          3284 => x"f0",
          3285 => x"87",
          3286 => x"98",
          3287 => x"38",
          3288 => x"08",
          3289 => x"71",
          3290 => x"98",
          3291 => x"27",
          3292 => x"2e",
          3293 => x"08",
          3294 => x"98",
          3295 => x"08",
          3296 => x"14",
          3297 => x"52",
          3298 => x"ff",
          3299 => x"08",
          3300 => x"52",
          3301 => x"06",
          3302 => x"74",
          3303 => x"38",
          3304 => x"73",
          3305 => x"84",
          3306 => x"ff",
          3307 => x"f2",
          3308 => x"85",
          3309 => x"fe",
          3310 => x"f0",
          3311 => x"08",
          3312 => x"90",
          3313 => x"52",
          3314 => x"72",
          3315 => x"c0",
          3316 => x"27",
          3317 => x"38",
          3318 => x"53",
          3319 => x"53",
          3320 => x"c0",
          3321 => x"53",
          3322 => x"c0",
          3323 => x"f6",
          3324 => x"9c",
          3325 => x"38",
          3326 => x"c0",
          3327 => x"83",
          3328 => x"70",
          3329 => x"2e",
          3330 => x"73",
          3331 => x"0d",
          3332 => x"3f",
          3333 => x"84",
          3334 => x"2a",
          3335 => x"2b",
          3336 => x"71",
          3337 => x"11",
          3338 => x"2b",
          3339 => x"53",
          3340 => x"53",
          3341 => x"16",
          3342 => x"8b",
          3343 => x"70",
          3344 => x"71",
          3345 => x"59",
          3346 => x"38",
          3347 => x"8b",
          3348 => x"76",
          3349 => x"86",
          3350 => x"73",
          3351 => x"70",
          3352 => x"71",
          3353 => x"55",
          3354 => x"71",
          3355 => x"16",
          3356 => x"0b",
          3357 => x"53",
          3358 => x"34",
          3359 => x"81",
          3360 => x"80",
          3361 => x"52",
          3362 => x"34",
          3363 => x"87",
          3364 => x"2b",
          3365 => x"17",
          3366 => x"2a",
          3367 => x"71",
          3368 => x"84",
          3369 => x"33",
          3370 => x"83",
          3371 => x"05",
          3372 => x"88",
          3373 => x"59",
          3374 => x"13",
          3375 => x"33",
          3376 => x"81",
          3377 => x"5a",
          3378 => x"13",
          3379 => x"70",
          3380 => x"71",
          3381 => x"81",
          3382 => x"83",
          3383 => x"7b",
          3384 => x"5a",
          3385 => x"73",
          3386 => x"70",
          3387 => x"8b",
          3388 => x"70",
          3389 => x"07",
          3390 => x"5f",
          3391 => x"77",
          3392 => x"b8",
          3393 => x"83",
          3394 => x"2b",
          3395 => x"33",
          3396 => x"58",
          3397 => x"70",
          3398 => x"81",
          3399 => x"80",
          3400 => x"54",
          3401 => x"84",
          3402 => x"81",
          3403 => x"2b",
          3404 => x"15",
          3405 => x"2a",
          3406 => x"53",
          3407 => x"34",
          3408 => x"79",
          3409 => x"80",
          3410 => x"38",
          3411 => x"0d",
          3412 => x"d4",
          3413 => x"23",
          3414 => x"ff",
          3415 => x"b8",
          3416 => x"0b",
          3417 => x"54",
          3418 => x"15",
          3419 => x"86",
          3420 => x"84",
          3421 => x"ff",
          3422 => x"ff",
          3423 => x"55",
          3424 => x"17",
          3425 => x"10",
          3426 => x"05",
          3427 => x"0b",
          3428 => x"3d",
          3429 => x"84",
          3430 => x"2a",
          3431 => x"51",
          3432 => x"b8",
          3433 => x"33",
          3434 => x"5a",
          3435 => x"80",
          3436 => x"10",
          3437 => x"88",
          3438 => x"79",
          3439 => x"7a",
          3440 => x"72",
          3441 => x"85",
          3442 => x"33",
          3443 => x"57",
          3444 => x"ff",
          3445 => x"80",
          3446 => x"81",
          3447 => x"81",
          3448 => x"59",
          3449 => x"59",
          3450 => x"38",
          3451 => x"38",
          3452 => x"16",
          3453 => x"80",
          3454 => x"56",
          3455 => x"15",
          3456 => x"88",
          3457 => x"75",
          3458 => x"70",
          3459 => x"88",
          3460 => x"f8",
          3461 => x"06",
          3462 => x"59",
          3463 => x"81",
          3464 => x"84",
          3465 => x"34",
          3466 => x"08",
          3467 => x"33",
          3468 => x"74",
          3469 => x"84",
          3470 => x"b8",
          3471 => x"86",
          3472 => x"2b",
          3473 => x"59",
          3474 => x"34",
          3475 => x"11",
          3476 => x"71",
          3477 => x"5c",
          3478 => x"87",
          3479 => x"16",
          3480 => x"12",
          3481 => x"2a",
          3482 => x"34",
          3483 => x"08",
          3484 => x"e4",
          3485 => x"33",
          3486 => x"83",
          3487 => x"85",
          3488 => x"88",
          3489 => x"74",
          3490 => x"84",
          3491 => x"33",
          3492 => x"83",
          3493 => x"87",
          3494 => x"88",
          3495 => x"57",
          3496 => x"1a",
          3497 => x"33",
          3498 => x"81",
          3499 => x"57",
          3500 => x"18",
          3501 => x"05",
          3502 => x"79",
          3503 => x"80",
          3504 => x"38",
          3505 => x"0d",
          3506 => x"b8",
          3507 => x"3d",
          3508 => x"b8",
          3509 => x"d0",
          3510 => x"84",
          3511 => x"84",
          3512 => x"81",
          3513 => x"08",
          3514 => x"85",
          3515 => x"76",
          3516 => x"34",
          3517 => x"22",
          3518 => x"83",
          3519 => x"51",
          3520 => x"89",
          3521 => x"10",
          3522 => x"f8",
          3523 => x"81",
          3524 => x"80",
          3525 => x"ed",
          3526 => x"70",
          3527 => x"76",
          3528 => x"2e",
          3529 => x"d7",
          3530 => x"38",
          3531 => x"70",
          3532 => x"83",
          3533 => x"2a",
          3534 => x"2b",
          3535 => x"71",
          3536 => x"83",
          3537 => x"fc",
          3538 => x"33",
          3539 => x"70",
          3540 => x"45",
          3541 => x"48",
          3542 => x"24",
          3543 => x"16",
          3544 => x"10",
          3545 => x"71",
          3546 => x"5c",
          3547 => x"85",
          3548 => x"38",
          3549 => x"a2",
          3550 => x"60",
          3551 => x"38",
          3552 => x"f7",
          3553 => x"33",
          3554 => x"7a",
          3555 => x"98",
          3556 => x"59",
          3557 => x"24",
          3558 => x"33",
          3559 => x"83",
          3560 => x"87",
          3561 => x"2b",
          3562 => x"15",
          3563 => x"2a",
          3564 => x"53",
          3565 => x"79",
          3566 => x"70",
          3567 => x"71",
          3568 => x"05",
          3569 => x"88",
          3570 => x"5e",
          3571 => x"16",
          3572 => x"d4",
          3573 => x"71",
          3574 => x"70",
          3575 => x"79",
          3576 => x"d4",
          3577 => x"12",
          3578 => x"07",
          3579 => x"71",
          3580 => x"5c",
          3581 => x"79",
          3582 => x"d4",
          3583 => x"33",
          3584 => x"74",
          3585 => x"71",
          3586 => x"5c",
          3587 => x"82",
          3588 => x"b8",
          3589 => x"83",
          3590 => x"57",
          3591 => x"5a",
          3592 => x"c4",
          3593 => x"84",
          3594 => x"ff",
          3595 => x"26",
          3596 => x"b8",
          3597 => x"ff",
          3598 => x"80",
          3599 => x"80",
          3600 => x"fe",
          3601 => x"5e",
          3602 => x"34",
          3603 => x"1e",
          3604 => x"b8",
          3605 => x"81",
          3606 => x"08",
          3607 => x"80",
          3608 => x"70",
          3609 => x"88",
          3610 => x"b8",
          3611 => x"b8",
          3612 => x"60",
          3613 => x"34",
          3614 => x"d3",
          3615 => x"7e",
          3616 => x"7f",
          3617 => x"08",
          3618 => x"04",
          3619 => x"83",
          3620 => x"70",
          3621 => x"07",
          3622 => x"48",
          3623 => x"60",
          3624 => x"08",
          3625 => x"82",
          3626 => x"b8",
          3627 => x"12",
          3628 => x"2b",
          3629 => x"83",
          3630 => x"5c",
          3631 => x"82",
          3632 => x"60",
          3633 => x"08",
          3634 => x"1c",
          3635 => x"84",
          3636 => x"fd",
          3637 => x"ff",
          3638 => x"77",
          3639 => x"83",
          3640 => x"18",
          3641 => x"10",
          3642 => x"71",
          3643 => x"5e",
          3644 => x"80",
          3645 => x"61",
          3646 => x"24",
          3647 => x"06",
          3648 => x"fe",
          3649 => x"b8",
          3650 => x"d0",
          3651 => x"84",
          3652 => x"84",
          3653 => x"81",
          3654 => x"08",
          3655 => x"85",
          3656 => x"7e",
          3657 => x"34",
          3658 => x"22",
          3659 => x"83",
          3660 => x"56",
          3661 => x"73",
          3662 => x"22",
          3663 => x"08",
          3664 => x"82",
          3665 => x"fc",
          3666 => x"38",
          3667 => x"7b",
          3668 => x"76",
          3669 => x"ea",
          3670 => x"e4",
          3671 => x"82",
          3672 => x"2b",
          3673 => x"11",
          3674 => x"71",
          3675 => x"33",
          3676 => x"70",
          3677 => x"46",
          3678 => x"84",
          3679 => x"84",
          3680 => x"33",
          3681 => x"83",
          3682 => x"87",
          3683 => x"88",
          3684 => x"5d",
          3685 => x"64",
          3686 => x"16",
          3687 => x"2b",
          3688 => x"2a",
          3689 => x"79",
          3690 => x"70",
          3691 => x"71",
          3692 => x"05",
          3693 => x"2b",
          3694 => x"40",
          3695 => x"75",
          3696 => x"70",
          3697 => x"8b",
          3698 => x"82",
          3699 => x"2b",
          3700 => x"5b",
          3701 => x"34",
          3702 => x"08",
          3703 => x"33",
          3704 => x"56",
          3705 => x"7e",
          3706 => x"3f",
          3707 => x"78",
          3708 => x"99",
          3709 => x"d4",
          3710 => x"23",
          3711 => x"ff",
          3712 => x"b8",
          3713 => x"0b",
          3714 => x"55",
          3715 => x"16",
          3716 => x"86",
          3717 => x"84",
          3718 => x"ff",
          3719 => x"ff",
          3720 => x"44",
          3721 => x"1f",
          3722 => x"10",
          3723 => x"05",
          3724 => x"0b",
          3725 => x"3f",
          3726 => x"33",
          3727 => x"83",
          3728 => x"85",
          3729 => x"88",
          3730 => x"76",
          3731 => x"05",
          3732 => x"84",
          3733 => x"2b",
          3734 => x"14",
          3735 => x"07",
          3736 => x"59",
          3737 => x"34",
          3738 => x"d4",
          3739 => x"71",
          3740 => x"70",
          3741 => x"78",
          3742 => x"d4",
          3743 => x"33",
          3744 => x"74",
          3745 => x"88",
          3746 => x"f8",
          3747 => x"5d",
          3748 => x"7f",
          3749 => x"84",
          3750 => x"81",
          3751 => x"2b",
          3752 => x"33",
          3753 => x"06",
          3754 => x"46",
          3755 => x"60",
          3756 => x"06",
          3757 => x"87",
          3758 => x"2b",
          3759 => x"19",
          3760 => x"2a",
          3761 => x"84",
          3762 => x"b8",
          3763 => x"85",
          3764 => x"2b",
          3765 => x"15",
          3766 => x"2a",
          3767 => x"56",
          3768 => x"87",
          3769 => x"70",
          3770 => x"07",
          3771 => x"5b",
          3772 => x"81",
          3773 => x"1f",
          3774 => x"2b",
          3775 => x"33",
          3776 => x"70",
          3777 => x"05",
          3778 => x"58",
          3779 => x"34",
          3780 => x"08",
          3781 => x"71",
          3782 => x"05",
          3783 => x"2b",
          3784 => x"2a",
          3785 => x"55",
          3786 => x"84",
          3787 => x"33",
          3788 => x"83",
          3789 => x"87",
          3790 => x"2b",
          3791 => x"15",
          3792 => x"2a",
          3793 => x"53",
          3794 => x"34",
          3795 => x"08",
          3796 => x"33",
          3797 => x"74",
          3798 => x"71",
          3799 => x"42",
          3800 => x"86",
          3801 => x"b8",
          3802 => x"33",
          3803 => x"06",
          3804 => x"76",
          3805 => x"b8",
          3806 => x"83",
          3807 => x"2b",
          3808 => x"33",
          3809 => x"41",
          3810 => x"79",
          3811 => x"b8",
          3812 => x"12",
          3813 => x"07",
          3814 => x"33",
          3815 => x"41",
          3816 => x"79",
          3817 => x"84",
          3818 => x"33",
          3819 => x"66",
          3820 => x"52",
          3821 => x"fe",
          3822 => x"1e",
          3823 => x"83",
          3824 => x"d5",
          3825 => x"71",
          3826 => x"05",
          3827 => x"88",
          3828 => x"5d",
          3829 => x"34",
          3830 => x"d4",
          3831 => x"12",
          3832 => x"07",
          3833 => x"33",
          3834 => x"5b",
          3835 => x"73",
          3836 => x"05",
          3837 => x"33",
          3838 => x"81",
          3839 => x"5f",
          3840 => x"16",
          3841 => x"70",
          3842 => x"71",
          3843 => x"81",
          3844 => x"83",
          3845 => x"63",
          3846 => x"5e",
          3847 => x"7b",
          3848 => x"70",
          3849 => x"8b",
          3850 => x"70",
          3851 => x"07",
          3852 => x"47",
          3853 => x"7f",
          3854 => x"83",
          3855 => x"7e",
          3856 => x"b8",
          3857 => x"80",
          3858 => x"84",
          3859 => x"3f",
          3860 => x"61",
          3861 => x"39",
          3862 => x"b8",
          3863 => x"b7",
          3864 => x"84",
          3865 => x"77",
          3866 => x"08",
          3867 => x"e6",
          3868 => x"e4",
          3869 => x"84",
          3870 => x"84",
          3871 => x"a0",
          3872 => x"80",
          3873 => x"51",
          3874 => x"08",
          3875 => x"16",
          3876 => x"84",
          3877 => x"84",
          3878 => x"34",
          3879 => x"d4",
          3880 => x"fe",
          3881 => x"06",
          3882 => x"74",
          3883 => x"84",
          3884 => x"84",
          3885 => x"55",
          3886 => x"15",
          3887 => x"c6",
          3888 => x"02",
          3889 => x"72",
          3890 => x"33",
          3891 => x"3d",
          3892 => x"05",
          3893 => x"9d",
          3894 => x"b8",
          3895 => x"87",
          3896 => x"84",
          3897 => x"b8",
          3898 => x"3d",
          3899 => x"af",
          3900 => x"54",
          3901 => x"e0",
          3902 => x"83",
          3903 => x"0b",
          3904 => x"75",
          3905 => x"b8",
          3906 => x"80",
          3907 => x"08",
          3908 => x"d6",
          3909 => x"73",
          3910 => x"55",
          3911 => x"0d",
          3912 => x"81",
          3913 => x"26",
          3914 => x"0d",
          3915 => x"05",
          3916 => x"76",
          3917 => x"17",
          3918 => x"55",
          3919 => x"87",
          3920 => x"52",
          3921 => x"e4",
          3922 => x"2e",
          3923 => x"54",
          3924 => x"38",
          3925 => x"80",
          3926 => x"74",
          3927 => x"04",
          3928 => x"ff",
          3929 => x"ff",
          3930 => x"78",
          3931 => x"88",
          3932 => x"81",
          3933 => x"b8",
          3934 => x"54",
          3935 => x"87",
          3936 => x"73",
          3937 => x"38",
          3938 => x"72",
          3939 => x"04",
          3940 => x"b8",
          3941 => x"80",
          3942 => x"0c",
          3943 => x"87",
          3944 => x"cd",
          3945 => x"06",
          3946 => x"87",
          3947 => x"38",
          3948 => x"ca",
          3949 => x"8c",
          3950 => x"73",
          3951 => x"82",
          3952 => x"39",
          3953 => x"83",
          3954 => x"77",
          3955 => x"33",
          3956 => x"80",
          3957 => x"fe",
          3958 => x"2e",
          3959 => x"e4",
          3960 => x"b4",
          3961 => x"81",
          3962 => x"81",
          3963 => x"09",
          3964 => x"08",
          3965 => x"a8",
          3966 => x"b8",
          3967 => x"76",
          3968 => x"55",
          3969 => x"8e",
          3970 => x"52",
          3971 => x"76",
          3972 => x"09",
          3973 => x"33",
          3974 => x"fe",
          3975 => x"7a",
          3976 => x"57",
          3977 => x"80",
          3978 => x"aa",
          3979 => x"7a",
          3980 => x"80",
          3981 => x"0b",
          3982 => x"9c",
          3983 => x"19",
          3984 => x"34",
          3985 => x"94",
          3986 => x"34",
          3987 => x"19",
          3988 => x"a2",
          3989 => x"84",
          3990 => x"7a",
          3991 => x"55",
          3992 => x"2a",
          3993 => x"98",
          3994 => x"a4",
          3995 => x"0c",
          3996 => x"81",
          3997 => x"84",
          3998 => x"18",
          3999 => x"e4",
          4000 => x"b2",
          4001 => x"08",
          4002 => x"38",
          4003 => x"81",
          4004 => x"3d",
          4005 => x"74",
          4006 => x"24",
          4007 => x"81",
          4008 => x"70",
          4009 => x"5a",
          4010 => x"b0",
          4011 => x"2e",
          4012 => x"54",
          4013 => x"33",
          4014 => x"08",
          4015 => x"5b",
          4016 => x"38",
          4017 => x"33",
          4018 => x"08",
          4019 => x"08",
          4020 => x"18",
          4021 => x"2e",
          4022 => x"54",
          4023 => x"33",
          4024 => x"08",
          4025 => x"5a",
          4026 => x"38",
          4027 => x"33",
          4028 => x"06",
          4029 => x"5d",
          4030 => x"06",
          4031 => x"04",
          4032 => x"59",
          4033 => x"80",
          4034 => x"5b",
          4035 => x"c2",
          4036 => x"52",
          4037 => x"84",
          4038 => x"ff",
          4039 => x"79",
          4040 => x"06",
          4041 => x"71",
          4042 => x"e4",
          4043 => x"74",
          4044 => x"38",
          4045 => x"59",
          4046 => x"80",
          4047 => x"5b",
          4048 => x"81",
          4049 => x"52",
          4050 => x"84",
          4051 => x"ff",
          4052 => x"79",
          4053 => x"fc",
          4054 => x"33",
          4055 => x"88",
          4056 => x"07",
          4057 => x"ff",
          4058 => x"0c",
          4059 => x"3d",
          4060 => x"53",
          4061 => x"52",
          4062 => x"b8",
          4063 => x"fe",
          4064 => x"18",
          4065 => x"31",
          4066 => x"a0",
          4067 => x"17",
          4068 => x"06",
          4069 => x"08",
          4070 => x"81",
          4071 => x"5a",
          4072 => x"08",
          4073 => x"33",
          4074 => x"e4",
          4075 => x"81",
          4076 => x"34",
          4077 => x"5d",
          4078 => x"82",
          4079 => x"cb",
          4080 => x"de",
          4081 => x"b8",
          4082 => x"5c",
          4083 => x"e4",
          4084 => x"ff",
          4085 => x"34",
          4086 => x"84",
          4087 => x"18",
          4088 => x"33",
          4089 => x"fd",
          4090 => x"a0",
          4091 => x"17",
          4092 => x"fd",
          4093 => x"53",
          4094 => x"52",
          4095 => x"b8",
          4096 => x"fb",
          4097 => x"18",
          4098 => x"31",
          4099 => x"a0",
          4100 => x"17",
          4101 => x"06",
          4102 => x"08",
          4103 => x"81",
          4104 => x"5a",
          4105 => x"08",
          4106 => x"81",
          4107 => x"86",
          4108 => x"fa",
          4109 => x"64",
          4110 => x"27",
          4111 => x"95",
          4112 => x"96",
          4113 => x"74",
          4114 => x"b8",
          4115 => x"88",
          4116 => x"0b",
          4117 => x"2e",
          4118 => x"5b",
          4119 => x"83",
          4120 => x"19",
          4121 => x"3f",
          4122 => x"38",
          4123 => x"0c",
          4124 => x"10",
          4125 => x"ff",
          4126 => x"34",
          4127 => x"34",
          4128 => x"b8",
          4129 => x"83",
          4130 => x"75",
          4131 => x"80",
          4132 => x"78",
          4133 => x"7c",
          4134 => x"06",
          4135 => x"b8",
          4136 => x"8e",
          4137 => x"85",
          4138 => x"1a",
          4139 => x"75",
          4140 => x"b8",
          4141 => x"8f",
          4142 => x"41",
          4143 => x"88",
          4144 => x"90",
          4145 => x"98",
          4146 => x"0b",
          4147 => x"81",
          4148 => x"08",
          4149 => x"76",
          4150 => x"1a",
          4151 => x"2e",
          4152 => x"54",
          4153 => x"33",
          4154 => x"08",
          4155 => x"5c",
          4156 => x"fd",
          4157 => x"b8",
          4158 => x"5f",
          4159 => x"38",
          4160 => x"33",
          4161 => x"77",
          4162 => x"89",
          4163 => x"0b",
          4164 => x"2e",
          4165 => x"b8",
          4166 => x"57",
          4167 => x"e4",
          4168 => x"c7",
          4169 => x"34",
          4170 => x"31",
          4171 => x"5b",
          4172 => x"38",
          4173 => x"82",
          4174 => x"52",
          4175 => x"84",
          4176 => x"ff",
          4177 => x"77",
          4178 => x"19",
          4179 => x"7c",
          4180 => x"81",
          4181 => x"5c",
          4182 => x"34",
          4183 => x"b8",
          4184 => x"5d",
          4185 => x"e4",
          4186 => x"88",
          4187 => x"34",
          4188 => x"31",
          4189 => x"5d",
          4190 => x"ca",
          4191 => x"2e",
          4192 => x"54",
          4193 => x"33",
          4194 => x"aa",
          4195 => x"70",
          4196 => x"ad",
          4197 => x"7d",
          4198 => x"84",
          4199 => x"19",
          4200 => x"1b",
          4201 => x"56",
          4202 => x"82",
          4203 => x"81",
          4204 => x"1f",
          4205 => x"ed",
          4206 => x"81",
          4207 => x"81",
          4208 => x"81",
          4209 => x"09",
          4210 => x"e4",
          4211 => x"70",
          4212 => x"84",
          4213 => x"7e",
          4214 => x"33",
          4215 => x"fa",
          4216 => x"76",
          4217 => x"3f",
          4218 => x"79",
          4219 => x"51",
          4220 => x"39",
          4221 => x"05",
          4222 => x"58",
          4223 => x"5a",
          4224 => x"7e",
          4225 => x"2b",
          4226 => x"83",
          4227 => x"06",
          4228 => x"5f",
          4229 => x"2a",
          4230 => x"2a",
          4231 => x"2a",
          4232 => x"39",
          4233 => x"5b",
          4234 => x"19",
          4235 => x"38",
          4236 => x"38",
          4237 => x"80",
          4238 => x"81",
          4239 => x"9c",
          4240 => x"56",
          4241 => x"52",
          4242 => x"e4",
          4243 => x"58",
          4244 => x"38",
          4245 => x"70",
          4246 => x"51",
          4247 => x"75",
          4248 => x"38",
          4249 => x"8c",
          4250 => x"39",
          4251 => x"7a",
          4252 => x"55",
          4253 => x"38",
          4254 => x"e4",
          4255 => x"08",
          4256 => x"7a",
          4257 => x"9c",
          4258 => x"56",
          4259 => x"80",
          4260 => x"81",
          4261 => x"70",
          4262 => x"7b",
          4263 => x"51",
          4264 => x"b8",
          4265 => x"19",
          4266 => x"38",
          4267 => x"38",
          4268 => x"75",
          4269 => x"75",
          4270 => x"b8",
          4271 => x"70",
          4272 => x"56",
          4273 => x"80",
          4274 => x"19",
          4275 => x"58",
          4276 => x"94",
          4277 => x"5a",
          4278 => x"84",
          4279 => x"80",
          4280 => x"0d",
          4281 => x"da",
          4282 => x"75",
          4283 => x"3f",
          4284 => x"39",
          4285 => x"0c",
          4286 => x"81",
          4287 => x"b6",
          4288 => x"08",
          4289 => x"26",
          4290 => x"72",
          4291 => x"88",
          4292 => x"76",
          4293 => x"38",
          4294 => x"18",
          4295 => x"38",
          4296 => x"94",
          4297 => x"56",
          4298 => x"2a",
          4299 => x"06",
          4300 => x"56",
          4301 => x"0d",
          4302 => x"8a",
          4303 => x"74",
          4304 => x"22",
          4305 => x"27",
          4306 => x"15",
          4307 => x"73",
          4308 => x"71",
          4309 => x"78",
          4310 => x"52",
          4311 => x"e4",
          4312 => x"2e",
          4313 => x"08",
          4314 => x"53",
          4315 => x"91",
          4316 => x"27",
          4317 => x"84",
          4318 => x"f3",
          4319 => x"08",
          4320 => x"0a",
          4321 => x"18",
          4322 => x"74",
          4323 => x"06",
          4324 => x"18",
          4325 => x"85",
          4326 => x"76",
          4327 => x"0c",
          4328 => x"05",
          4329 => x"b8",
          4330 => x"98",
          4331 => x"7a",
          4332 => x"75",
          4333 => x"b8",
          4334 => x"84",
          4335 => x"56",
          4336 => x"38",
          4337 => x"26",
          4338 => x"98",
          4339 => x"f9",
          4340 => x"87",
          4341 => x"ff",
          4342 => x"08",
          4343 => x"84",
          4344 => x"38",
          4345 => x"5f",
          4346 => x"9c",
          4347 => x"5c",
          4348 => x"22",
          4349 => x"5d",
          4350 => x"58",
          4351 => x"70",
          4352 => x"74",
          4353 => x"55",
          4354 => x"54",
          4355 => x"33",
          4356 => x"08",
          4357 => x"39",
          4358 => x"b8",
          4359 => x"54",
          4360 => x"53",
          4361 => x"3f",
          4362 => x"84",
          4363 => x"19",
          4364 => x"a0",
          4365 => x"19",
          4366 => x"06",
          4367 => x"08",
          4368 => x"81",
          4369 => x"c5",
          4370 => x"ff",
          4371 => x"81",
          4372 => x"fe",
          4373 => x"56",
          4374 => x"38",
          4375 => x"1b",
          4376 => x"f8",
          4377 => x"8f",
          4378 => x"66",
          4379 => x"81",
          4380 => x"5e",
          4381 => x"19",
          4382 => x"08",
          4383 => x"33",
          4384 => x"81",
          4385 => x"53",
          4386 => x"e1",
          4387 => x"2e",
          4388 => x"b4",
          4389 => x"38",
          4390 => x"76",
          4391 => x"33",
          4392 => x"41",
          4393 => x"32",
          4394 => x"72",
          4395 => x"45",
          4396 => x"7a",
          4397 => x"81",
          4398 => x"38",
          4399 => x"fa",
          4400 => x"84",
          4401 => x"1c",
          4402 => x"84",
          4403 => x"81",
          4404 => x"81",
          4405 => x"57",
          4406 => x"81",
          4407 => x"08",
          4408 => x"1a",
          4409 => x"5b",
          4410 => x"38",
          4411 => x"09",
          4412 => x"b4",
          4413 => x"7e",
          4414 => x"3f",
          4415 => x"2e",
          4416 => x"86",
          4417 => x"93",
          4418 => x"06",
          4419 => x"0c",
          4420 => x"38",
          4421 => x"39",
          4422 => x"06",
          4423 => x"80",
          4424 => x"e4",
          4425 => x"fd",
          4426 => x"77",
          4427 => x"19",
          4428 => x"71",
          4429 => x"ff",
          4430 => x"06",
          4431 => x"76",
          4432 => x"78",
          4433 => x"88",
          4434 => x"2e",
          4435 => x"ff",
          4436 => x"5c",
          4437 => x"81",
          4438 => x"77",
          4439 => x"57",
          4440 => x"fe",
          4441 => x"05",
          4442 => x"81",
          4443 => x"75",
          4444 => x"ff",
          4445 => x"7c",
          4446 => x"81",
          4447 => x"5a",
          4448 => x"06",
          4449 => x"38",
          4450 => x"0b",
          4451 => x"0c",
          4452 => x"63",
          4453 => x"51",
          4454 => x"5a",
          4455 => x"81",
          4456 => x"1d",
          4457 => x"56",
          4458 => x"82",
          4459 => x"55",
          4460 => x"df",
          4461 => x"52",
          4462 => x"84",
          4463 => x"ff",
          4464 => x"76",
          4465 => x"08",
          4466 => x"84",
          4467 => x"70",
          4468 => x"1d",
          4469 => x"38",
          4470 => x"8f",
          4471 => x"38",
          4472 => x"aa",
          4473 => x"74",
          4474 => x"78",
          4475 => x"05",
          4476 => x"56",
          4477 => x"80",
          4478 => x"57",
          4479 => x"59",
          4480 => x"78",
          4481 => x"31",
          4482 => x"80",
          4483 => x"e1",
          4484 => x"1d",
          4485 => x"3f",
          4486 => x"e4",
          4487 => x"84",
          4488 => x"81",
          4489 => x"81",
          4490 => x"57",
          4491 => x"81",
          4492 => x"08",
          4493 => x"1c",
          4494 => x"59",
          4495 => x"38",
          4496 => x"09",
          4497 => x"b4",
          4498 => x"7d",
          4499 => x"3f",
          4500 => x"fd",
          4501 => x"2a",
          4502 => x"38",
          4503 => x"80",
          4504 => x"81",
          4505 => x"ac",
          4506 => x"2e",
          4507 => x"80",
          4508 => x"b8",
          4509 => x"80",
          4510 => x"75",
          4511 => x"5d",
          4512 => x"39",
          4513 => x"09",
          4514 => x"9b",
          4515 => x"2b",
          4516 => x"38",
          4517 => x"f3",
          4518 => x"83",
          4519 => x"11",
          4520 => x"52",
          4521 => x"38",
          4522 => x"76",
          4523 => x"e4",
          4524 => x"53",
          4525 => x"f6",
          4526 => x"09",
          4527 => x"81",
          4528 => x"38",
          4529 => x"56",
          4530 => x"80",
          4531 => x"70",
          4532 => x"ff",
          4533 => x"fe",
          4534 => x"0c",
          4535 => x"ff",
          4536 => x"fe",
          4537 => x"08",
          4538 => x"58",
          4539 => x"b5",
          4540 => x"57",
          4541 => x"81",
          4542 => x"56",
          4543 => x"1f",
          4544 => x"55",
          4545 => x"70",
          4546 => x"74",
          4547 => x"70",
          4548 => x"82",
          4549 => x"34",
          4550 => x"1c",
          4551 => x"5a",
          4552 => x"33",
          4553 => x"15",
          4554 => x"80",
          4555 => x"74",
          4556 => x"5a",
          4557 => x"10",
          4558 => x"ff",
          4559 => x"58",
          4560 => x"76",
          4561 => x"58",
          4562 => x"55",
          4563 => x"80",
          4564 => x"bf",
          4565 => x"87",
          4566 => x"ff",
          4567 => x"76",
          4568 => x"79",
          4569 => x"27",
          4570 => x"2e",
          4571 => x"27",
          4572 => x"56",
          4573 => x"ea",
          4574 => x"87",
          4575 => x"ec",
          4576 => x"41",
          4577 => x"f4",
          4578 => x"b8",
          4579 => x"80",
          4580 => x"56",
          4581 => x"84",
          4582 => x"08",
          4583 => x"38",
          4584 => x"34",
          4585 => x"05",
          4586 => x"06",
          4587 => x"38",
          4588 => x"c1",
          4589 => x"80",
          4590 => x"b8",
          4591 => x"81",
          4592 => x"19",
          4593 => x"57",
          4594 => x"38",
          4595 => x"09",
          4596 => x"75",
          4597 => x"51",
          4598 => x"80",
          4599 => x"75",
          4600 => x"38",
          4601 => x"74",
          4602 => x"30",
          4603 => x"74",
          4604 => x"59",
          4605 => x"52",
          4606 => x"e4",
          4607 => x"2e",
          4608 => x"2e",
          4609 => x"83",
          4610 => x"38",
          4611 => x"77",
          4612 => x"57",
          4613 => x"76",
          4614 => x"51",
          4615 => x"80",
          4616 => x"76",
          4617 => x"c3",
          4618 => x"55",
          4619 => x"ff",
          4620 => x"9c",
          4621 => x"70",
          4622 => x"05",
          4623 => x"38",
          4624 => x"06",
          4625 => x"0b",
          4626 => x"b8",
          4627 => x"75",
          4628 => x"40",
          4629 => x"81",
          4630 => x"b8",
          4631 => x"80",
          4632 => x"81",
          4633 => x"81",
          4634 => x"b8",
          4635 => x"83",
          4636 => x"19",
          4637 => x"31",
          4638 => x"38",
          4639 => x"84",
          4640 => x"fd",
          4641 => x"08",
          4642 => x"e9",
          4643 => x"b8",
          4644 => x"b8",
          4645 => x"81",
          4646 => x"70",
          4647 => x"70",
          4648 => x"5d",
          4649 => x"b8",
          4650 => x"80",
          4651 => x"38",
          4652 => x"09",
          4653 => x"76",
          4654 => x"51",
          4655 => x"80",
          4656 => x"76",
          4657 => x"83",
          4658 => x"61",
          4659 => x"8d",
          4660 => x"75",
          4661 => x"75",
          4662 => x"05",
          4663 => x"ff",
          4664 => x"70",
          4665 => x"e4",
          4666 => x"75",
          4667 => x"2a",
          4668 => x"83",
          4669 => x"78",
          4670 => x"2e",
          4671 => x"22",
          4672 => x"38",
          4673 => x"34",
          4674 => x"84",
          4675 => x"08",
          4676 => x"7f",
          4677 => x"54",
          4678 => x"53",
          4679 => x"3f",
          4680 => x"83",
          4681 => x"34",
          4682 => x"84",
          4683 => x"1d",
          4684 => x"33",
          4685 => x"fb",
          4686 => x"a0",
          4687 => x"1c",
          4688 => x"fb",
          4689 => x"33",
          4690 => x"09",
          4691 => x"39",
          4692 => x"fa",
          4693 => x"c0",
          4694 => x"b4",
          4695 => x"33",
          4696 => x"08",
          4697 => x"84",
          4698 => x"1c",
          4699 => x"a0",
          4700 => x"33",
          4701 => x"b8",
          4702 => x"ff",
          4703 => x"98",
          4704 => x"f7",
          4705 => x"80",
          4706 => x"81",
          4707 => x"05",
          4708 => x"ce",
          4709 => x"b4",
          4710 => x"7c",
          4711 => x"3f",
          4712 => x"61",
          4713 => x"96",
          4714 => x"82",
          4715 => x"80",
          4716 => x"05",
          4717 => x"58",
          4718 => x"74",
          4719 => x"56",
          4720 => x"14",
          4721 => x"76",
          4722 => x"79",
          4723 => x"55",
          4724 => x"80",
          4725 => x"5e",
          4726 => x"82",
          4727 => x"57",
          4728 => x"81",
          4729 => x"b2",
          4730 => x"75",
          4731 => x"80",
          4732 => x"90",
          4733 => x"77",
          4734 => x"58",
          4735 => x"81",
          4736 => x"38",
          4737 => x"81",
          4738 => x"a5",
          4739 => x"96",
          4740 => x"05",
          4741 => x"1c",
          4742 => x"89",
          4743 => x"08",
          4744 => x"9c",
          4745 => x"82",
          4746 => x"2b",
          4747 => x"88",
          4748 => x"59",
          4749 => x"88",
          4750 => x"56",
          4751 => x"15",
          4752 => x"07",
          4753 => x"3d",
          4754 => x"39",
          4755 => x"31",
          4756 => x"90",
          4757 => x"3f",
          4758 => x"06",
          4759 => x"81",
          4760 => x"2a",
          4761 => x"34",
          4762 => x"1f",
          4763 => x"70",
          4764 => x"38",
          4765 => x"70",
          4766 => x"07",
          4767 => x"74",
          4768 => x"0b",
          4769 => x"72",
          4770 => x"77",
          4771 => x"1e",
          4772 => x"ff",
          4773 => x"a4",
          4774 => x"54",
          4775 => x"84",
          4776 => x"80",
          4777 => x"ff",
          4778 => x"81",
          4779 => x"81",
          4780 => x"59",
          4781 => x"b4",
          4782 => x"80",
          4783 => x"73",
          4784 => x"39",
          4785 => x"42",
          4786 => x"55",
          4787 => x"53",
          4788 => x"72",
          4789 => x"08",
          4790 => x"94",
          4791 => x"82",
          4792 => x"58",
          4793 => x"52",
          4794 => x"72",
          4795 => x"38",
          4796 => x"76",
          4797 => x"17",
          4798 => x"af",
          4799 => x"80",
          4800 => x"82",
          4801 => x"89",
          4802 => x"83",
          4803 => x"70",
          4804 => x"80",
          4805 => x"8f",
          4806 => x"ff",
          4807 => x"72",
          4808 => x"38",
          4809 => x"76",
          4810 => x"17",
          4811 => x"56",
          4812 => x"38",
          4813 => x"32",
          4814 => x"51",
          4815 => x"38",
          4816 => x"33",
          4817 => x"72",
          4818 => x"25",
          4819 => x"38",
          4820 => x"3d",
          4821 => x"26",
          4822 => x"52",
          4823 => x"b8",
          4824 => x"73",
          4825 => x"b8",
          4826 => x"e4",
          4827 => x"53",
          4828 => x"39",
          4829 => x"52",
          4830 => x"e4",
          4831 => x"0d",
          4832 => x"30",
          4833 => x"5a",
          4834 => x"14",
          4835 => x"56",
          4836 => x"dc",
          4837 => x"07",
          4838 => x"61",
          4839 => x"76",
          4840 => x"2e",
          4841 => x"80",
          4842 => x"fe",
          4843 => x"30",
          4844 => x"56",
          4845 => x"89",
          4846 => x"76",
          4847 => x"76",
          4848 => x"22",
          4849 => x"5d",
          4850 => x"38",
          4851 => x"ae",
          4852 => x"aa",
          4853 => x"5a",
          4854 => x"10",
          4855 => x"76",
          4856 => x"22",
          4857 => x"06",
          4858 => x"53",
          4859 => x"ff",
          4860 => x"5c",
          4861 => x"19",
          4862 => x"80",
          4863 => x"38",
          4864 => x"25",
          4865 => x"ce",
          4866 => x"7c",
          4867 => x"77",
          4868 => x"25",
          4869 => x"72",
          4870 => x"2e",
          4871 => x"38",
          4872 => x"9e",
          4873 => x"82",
          4874 => x"5f",
          4875 => x"58",
          4876 => x"1c",
          4877 => x"84",
          4878 => x"7d",
          4879 => x"ed",
          4880 => x"2e",
          4881 => x"06",
          4882 => x"5d",
          4883 => x"07",
          4884 => x"7d",
          4885 => x"5a",
          4886 => x"ec",
          4887 => x"33",
          4888 => x"2e",
          4889 => x"84",
          4890 => x"74",
          4891 => x"2e",
          4892 => x"06",
          4893 => x"65",
          4894 => x"58",
          4895 => x"70",
          4896 => x"56",
          4897 => x"80",
          4898 => x"5a",
          4899 => x"75",
          4900 => x"38",
          4901 => x"81",
          4902 => x"5b",
          4903 => x"56",
          4904 => x"38",
          4905 => x"57",
          4906 => x"e9",
          4907 => x"1d",
          4908 => x"b8",
          4909 => x"84",
          4910 => x"82",
          4911 => x"38",
          4912 => x"06",
          4913 => x"38",
          4914 => x"05",
          4915 => x"33",
          4916 => x"57",
          4917 => x"38",
          4918 => x"55",
          4919 => x"74",
          4920 => x"59",
          4921 => x"79",
          4922 => x"81",
          4923 => x"70",
          4924 => x"09",
          4925 => x"07",
          4926 => x"1d",
          4927 => x"fc",
          4928 => x"ab",
          4929 => x"0c",
          4930 => x"26",
          4931 => x"c9",
          4932 => x"81",
          4933 => x"18",
          4934 => x"82",
          4935 => x"81",
          4936 => x"83",
          4937 => x"06",
          4938 => x"74",
          4939 => x"33",
          4940 => x"b9",
          4941 => x"83",
          4942 => x"70",
          4943 => x"80",
          4944 => x"8f",
          4945 => x"ff",
          4946 => x"72",
          4947 => x"38",
          4948 => x"8a",
          4949 => x"06",
          4950 => x"99",
          4951 => x"81",
          4952 => x"ff",
          4953 => x"a0",
          4954 => x"5b",
          4955 => x"53",
          4956 => x"70",
          4957 => x"2e",
          4958 => x"07",
          4959 => x"74",
          4960 => x"80",
          4961 => x"71",
          4962 => x"07",
          4963 => x"39",
          4964 => x"54",
          4965 => x"11",
          4966 => x"81",
          4967 => x"07",
          4968 => x"e5",
          4969 => x"fd",
          4970 => x"5c",
          4971 => x"b8",
          4972 => x"3d",
          4973 => x"e7",
          4974 => x"0c",
          4975 => x"79",
          4976 => x"81",
          4977 => x"56",
          4978 => x"ed",
          4979 => x"84",
          4980 => x"85",
          4981 => x"ac",
          4982 => x"76",
          4983 => x"0c",
          4984 => x"59",
          4985 => x"33",
          4986 => x"e4",
          4987 => x"5e",
          4988 => x"80",
          4989 => x"d8",
          4990 => x"81",
          4991 => x"84",
          4992 => x"81",
          4993 => x"c2",
          4994 => x"82",
          4995 => x"84",
          4996 => x"34",
          4997 => x"5a",
          4998 => x"70",
          4999 => x"bb",
          5000 => x"2e",
          5001 => x"b4",
          5002 => x"84",
          5003 => x"71",
          5004 => x"74",
          5005 => x"75",
          5006 => x"1d",
          5007 => x"58",
          5008 => x"58",
          5009 => x"c4",
          5010 => x"88",
          5011 => x"2e",
          5012 => x"cf",
          5013 => x"88",
          5014 => x"80",
          5015 => x"33",
          5016 => x"81",
          5017 => x"75",
          5018 => x"5e",
          5019 => x"c8",
          5020 => x"17",
          5021 => x"5f",
          5022 => x"82",
          5023 => x"71",
          5024 => x"5a",
          5025 => x"80",
          5026 => x"06",
          5027 => x"17",
          5028 => x"2b",
          5029 => x"74",
          5030 => x"7c",
          5031 => x"80",
          5032 => x"56",
          5033 => x"83",
          5034 => x"2b",
          5035 => x"70",
          5036 => x"07",
          5037 => x"80",
          5038 => x"71",
          5039 => x"7b",
          5040 => x"7a",
          5041 => x"81",
          5042 => x"51",
          5043 => x"08",
          5044 => x"81",
          5045 => x"ff",
          5046 => x"5d",
          5047 => x"82",
          5048 => x"38",
          5049 => x"0c",
          5050 => x"a8",
          5051 => x"57",
          5052 => x"88",
          5053 => x"2e",
          5054 => x"0c",
          5055 => x"38",
          5056 => x"81",
          5057 => x"89",
          5058 => x"08",
          5059 => x"0c",
          5060 => x"0b",
          5061 => x"96",
          5062 => x"22",
          5063 => x"23",
          5064 => x"0b",
          5065 => x"0c",
          5066 => x"97",
          5067 => x"e4",
          5068 => x"d0",
          5069 => x"58",
          5070 => x"78",
          5071 => x"78",
          5072 => x"08",
          5073 => x"08",
          5074 => x"5c",
          5075 => x"ff",
          5076 => x"26",
          5077 => x"06",
          5078 => x"99",
          5079 => x"ff",
          5080 => x"2a",
          5081 => x"06",
          5082 => x"7a",
          5083 => x"2a",
          5084 => x"2e",
          5085 => x"5e",
          5086 => x"61",
          5087 => x"fe",
          5088 => x"5e",
          5089 => x"58",
          5090 => x"59",
          5091 => x"83",
          5092 => x"70",
          5093 => x"5b",
          5094 => x"e8",
          5095 => x"57",
          5096 => x"70",
          5097 => x"84",
          5098 => x"71",
          5099 => x"ff",
          5100 => x"83",
          5101 => x"5b",
          5102 => x"05",
          5103 => x"59",
          5104 => x"b8",
          5105 => x"2a",
          5106 => x"10",
          5107 => x"5d",
          5108 => x"83",
          5109 => x"80",
          5110 => x"18",
          5111 => x"2e",
          5112 => x"17",
          5113 => x"86",
          5114 => x"85",
          5115 => x"18",
          5116 => x"1f",
          5117 => x"5d",
          5118 => x"2e",
          5119 => x"b8",
          5120 => x"2e",
          5121 => x"70",
          5122 => x"42",
          5123 => x"2e",
          5124 => x"06",
          5125 => x"33",
          5126 => x"06",
          5127 => x"f8",
          5128 => x"38",
          5129 => x"7a",
          5130 => x"83",
          5131 => x"40",
          5132 => x"33",
          5133 => x"71",
          5134 => x"77",
          5135 => x"2e",
          5136 => x"83",
          5137 => x"81",
          5138 => x"40",
          5139 => x"58",
          5140 => x"38",
          5141 => x"fe",
          5142 => x"38",
          5143 => x"0d",
          5144 => x"dc",
          5145 => x"e4",
          5146 => x"8d",
          5147 => x"0d",
          5148 => x"e4",
          5149 => x"05",
          5150 => x"33",
          5151 => x"5f",
          5152 => x"74",
          5153 => x"8a",
          5154 => x"78",
          5155 => x"81",
          5156 => x"1b",
          5157 => x"84",
          5158 => x"93",
          5159 => x"83",
          5160 => x"e9",
          5161 => x"88",
          5162 => x"09",
          5163 => x"58",
          5164 => x"b1",
          5165 => x"2e",
          5166 => x"54",
          5167 => x"33",
          5168 => x"e4",
          5169 => x"81",
          5170 => x"99",
          5171 => x"17",
          5172 => x"2b",
          5173 => x"2e",
          5174 => x"17",
          5175 => x"90",
          5176 => x"33",
          5177 => x"71",
          5178 => x"59",
          5179 => x"09",
          5180 => x"17",
          5181 => x"90",
          5182 => x"33",
          5183 => x"71",
          5184 => x"5e",
          5185 => x"09",
          5186 => x"17",
          5187 => x"90",
          5188 => x"33",
          5189 => x"71",
          5190 => x"1c",
          5191 => x"90",
          5192 => x"33",
          5193 => x"71",
          5194 => x"49",
          5195 => x"5a",
          5196 => x"81",
          5197 => x"7c",
          5198 => x"8c",
          5199 => x"f7",
          5200 => x"38",
          5201 => x"39",
          5202 => x"17",
          5203 => x"ff",
          5204 => x"7a",
          5205 => x"84",
          5206 => x"17",
          5207 => x"a0",
          5208 => x"33",
          5209 => x"84",
          5210 => x"74",
          5211 => x"85",
          5212 => x"5c",
          5213 => x"17",
          5214 => x"2b",
          5215 => x"d2",
          5216 => x"ca",
          5217 => x"82",
          5218 => x"2b",
          5219 => x"88",
          5220 => x"0c",
          5221 => x"40",
          5222 => x"75",
          5223 => x"f9",
          5224 => x"38",
          5225 => x"f7",
          5226 => x"38",
          5227 => x"08",
          5228 => x"81",
          5229 => x"fc",
          5230 => x"d3",
          5231 => x"41",
          5232 => x"80",
          5233 => x"05",
          5234 => x"74",
          5235 => x"38",
          5236 => x"d0",
          5237 => x"c4",
          5238 => x"05",
          5239 => x"84",
          5240 => x"80",
          5241 => x"54",
          5242 => x"2e",
          5243 => x"53",
          5244 => x"b8",
          5245 => x"0c",
          5246 => x"b8",
          5247 => x"33",
          5248 => x"56",
          5249 => x"16",
          5250 => x"58",
          5251 => x"7f",
          5252 => x"7b",
          5253 => x"05",
          5254 => x"33",
          5255 => x"99",
          5256 => x"ff",
          5257 => x"76",
          5258 => x"81",
          5259 => x"9f",
          5260 => x"81",
          5261 => x"77",
          5262 => x"9f",
          5263 => x"80",
          5264 => x"5d",
          5265 => x"7f",
          5266 => x"f7",
          5267 => x"8b",
          5268 => x"05",
          5269 => x"56",
          5270 => x"06",
          5271 => x"9e",
          5272 => x"3f",
          5273 => x"e4",
          5274 => x"0c",
          5275 => x"9c",
          5276 => x"90",
          5277 => x"84",
          5278 => x"08",
          5279 => x"06",
          5280 => x"76",
          5281 => x"2e",
          5282 => x"76",
          5283 => x"06",
          5284 => x"66",
          5285 => x"88",
          5286 => x"5e",
          5287 => x"38",
          5288 => x"8f",
          5289 => x"80",
          5290 => x"a0",
          5291 => x"5e",
          5292 => x"9b",
          5293 => x"2e",
          5294 => x"9c",
          5295 => x"80",
          5296 => x"1c",
          5297 => x"34",
          5298 => x"b4",
          5299 => x"5f",
          5300 => x"17",
          5301 => x"57",
          5302 => x"80",
          5303 => x"5b",
          5304 => x"78",
          5305 => x"38",
          5306 => x"05",
          5307 => x"56",
          5308 => x"81",
          5309 => x"75",
          5310 => x"77",
          5311 => x"2e",
          5312 => x"7e",
          5313 => x"a4",
          5314 => x"12",
          5315 => x"40",
          5316 => x"81",
          5317 => x"16",
          5318 => x"90",
          5319 => x"33",
          5320 => x"71",
          5321 => x"60",
          5322 => x"5e",
          5323 => x"90",
          5324 => x"80",
          5325 => x"81",
          5326 => x"38",
          5327 => x"94",
          5328 => x"2b",
          5329 => x"78",
          5330 => x"27",
          5331 => x"5f",
          5332 => x"77",
          5333 => x"84",
          5334 => x"08",
          5335 => x"b8",
          5336 => x"75",
          5337 => x"c2",
          5338 => x"38",
          5339 => x"80",
          5340 => x"79",
          5341 => x"79",
          5342 => x"79",
          5343 => x"ca",
          5344 => x"07",
          5345 => x"8b",
          5346 => x"fe",
          5347 => x"33",
          5348 => x"7d",
          5349 => x"7c",
          5350 => x"74",
          5351 => x"84",
          5352 => x"08",
          5353 => x"e4",
          5354 => x"b8",
          5355 => x"80",
          5356 => x"82",
          5357 => x"38",
          5358 => x"08",
          5359 => x"af",
          5360 => x"17",
          5361 => x"34",
          5362 => x"38",
          5363 => x"34",
          5364 => x"39",
          5365 => x"98",
          5366 => x"5e",
          5367 => x"80",
          5368 => x"17",
          5369 => x"66",
          5370 => x"67",
          5371 => x"80",
          5372 => x"7c",
          5373 => x"38",
          5374 => x"5e",
          5375 => x"2e",
          5376 => x"7d",
          5377 => x"54",
          5378 => x"33",
          5379 => x"e4",
          5380 => x"81",
          5381 => x"7a",
          5382 => x"80",
          5383 => x"f9",
          5384 => x"53",
          5385 => x"52",
          5386 => x"e4",
          5387 => x"aa",
          5388 => x"34",
          5389 => x"84",
          5390 => x"17",
          5391 => x"33",
          5392 => x"ff",
          5393 => x"a0",
          5394 => x"16",
          5395 => x"5b",
          5396 => x"76",
          5397 => x"0c",
          5398 => x"06",
          5399 => x"7e",
          5400 => x"5f",
          5401 => x"38",
          5402 => x"1c",
          5403 => x"f9",
          5404 => x"1a",
          5405 => x"94",
          5406 => x"81",
          5407 => x"84",
          5408 => x"f7",
          5409 => x"9f",
          5410 => x"66",
          5411 => x"89",
          5412 => x"08",
          5413 => x"33",
          5414 => x"16",
          5415 => x"78",
          5416 => x"41",
          5417 => x"1a",
          5418 => x"1a",
          5419 => x"80",
          5420 => x"8c",
          5421 => x"75",
          5422 => x"81",
          5423 => x"06",
          5424 => x"22",
          5425 => x"7a",
          5426 => x"1a",
          5427 => x"38",
          5428 => x"98",
          5429 => x"fe",
          5430 => x"57",
          5431 => x"19",
          5432 => x"05",
          5433 => x"38",
          5434 => x"77",
          5435 => x"55",
          5436 => x"31",
          5437 => x"81",
          5438 => x"84",
          5439 => x"83",
          5440 => x"a9",
          5441 => x"75",
          5442 => x"71",
          5443 => x"75",
          5444 => x"81",
          5445 => x"ef",
          5446 => x"31",
          5447 => x"94",
          5448 => x"0c",
          5449 => x"56",
          5450 => x"0d",
          5451 => x"3d",
          5452 => x"9c",
          5453 => x"84",
          5454 => x"27",
          5455 => x"19",
          5456 => x"83",
          5457 => x"7f",
          5458 => x"81",
          5459 => x"19",
          5460 => x"b8",
          5461 => x"56",
          5462 => x"81",
          5463 => x"ff",
          5464 => x"05",
          5465 => x"38",
          5466 => x"70",
          5467 => x"75",
          5468 => x"81",
          5469 => x"59",
          5470 => x"fe",
          5471 => x"53",
          5472 => x"52",
          5473 => x"84",
          5474 => x"06",
          5475 => x"83",
          5476 => x"08",
          5477 => x"74",
          5478 => x"82",
          5479 => x"81",
          5480 => x"19",
          5481 => x"52",
          5482 => x"3f",
          5483 => x"1b",
          5484 => x"39",
          5485 => x"a3",
          5486 => x"fc",
          5487 => x"9c",
          5488 => x"06",
          5489 => x"08",
          5490 => x"91",
          5491 => x"0c",
          5492 => x"1b",
          5493 => x"92",
          5494 => x"65",
          5495 => x"7e",
          5496 => x"38",
          5497 => x"38",
          5498 => x"38",
          5499 => x"59",
          5500 => x"55",
          5501 => x"38",
          5502 => x"38",
          5503 => x"06",
          5504 => x"82",
          5505 => x"5d",
          5506 => x"09",
          5507 => x"76",
          5508 => x"38",
          5509 => x"89",
          5510 => x"76",
          5511 => x"74",
          5512 => x"2e",
          5513 => x"8c",
          5514 => x"08",
          5515 => x"56",
          5516 => x"81",
          5517 => x"9c",
          5518 => x"77",
          5519 => x"70",
          5520 => x"57",
          5521 => x"15",
          5522 => x"2e",
          5523 => x"7f",
          5524 => x"77",
          5525 => x"33",
          5526 => x"e4",
          5527 => x"08",
          5528 => x"a5",
          5529 => x"72",
          5530 => x"81",
          5531 => x"59",
          5532 => x"60",
          5533 => x"2b",
          5534 => x"7f",
          5535 => x"70",
          5536 => x"5a",
          5537 => x"83",
          5538 => x"7a",
          5539 => x"77",
          5540 => x"34",
          5541 => x"92",
          5542 => x"0c",
          5543 => x"55",
          5544 => x"a2",
          5545 => x"76",
          5546 => x"5a",
          5547 => x"59",
          5548 => x"b6",
          5549 => x"5e",
          5550 => x"06",
          5551 => x"b8",
          5552 => x"98",
          5553 => x"2e",
          5554 => x"b4",
          5555 => x"94",
          5556 => x"58",
          5557 => x"80",
          5558 => x"58",
          5559 => x"ff",
          5560 => x"81",
          5561 => x"81",
          5562 => x"70",
          5563 => x"98",
          5564 => x"08",
          5565 => x"38",
          5566 => x"b4",
          5567 => x"b8",
          5568 => x"08",
          5569 => x"55",
          5570 => x"e3",
          5571 => x"17",
          5572 => x"33",
          5573 => x"fe",
          5574 => x"1a",
          5575 => x"33",
          5576 => x"b4",
          5577 => x"7b",
          5578 => x"39",
          5579 => x"ab",
          5580 => x"84",
          5581 => x"1a",
          5582 => x"79",
          5583 => x"e4",
          5584 => x"bd",
          5585 => x"08",
          5586 => x"33",
          5587 => x"b8",
          5588 => x"e4",
          5589 => x"a8",
          5590 => x"08",
          5591 => x"5c",
          5592 => x"fc",
          5593 => x"17",
          5594 => x"33",
          5595 => x"fb",
          5596 => x"95",
          5597 => x"06",
          5598 => x"08",
          5599 => x"b4",
          5600 => x"81",
          5601 => x"3f",
          5602 => x"84",
          5603 => x"16",
          5604 => x"a0",
          5605 => x"16",
          5606 => x"06",
          5607 => x"08",
          5608 => x"81",
          5609 => x"60",
          5610 => x"58",
          5611 => x"1b",
          5612 => x"92",
          5613 => x"34",
          5614 => x"3d",
          5615 => x"89",
          5616 => x"08",
          5617 => x"33",
          5618 => x"16",
          5619 => x"77",
          5620 => x"5c",
          5621 => x"18",
          5622 => x"57",
          5623 => x"a0",
          5624 => x"79",
          5625 => x"7a",
          5626 => x"b8",
          5627 => x"93",
          5628 => x"2e",
          5629 => x"b4",
          5630 => x"18",
          5631 => x"57",
          5632 => x"19",
          5633 => x"5a",
          5634 => x"2a",
          5635 => x"76",
          5636 => x"83",
          5637 => x"55",
          5638 => x"7a",
          5639 => x"75",
          5640 => x"78",
          5641 => x"0b",
          5642 => x"34",
          5643 => x"0b",
          5644 => x"34",
          5645 => x"7b",
          5646 => x"e4",
          5647 => x"5b",
          5648 => x"b8",
          5649 => x"54",
          5650 => x"53",
          5651 => x"b5",
          5652 => x"fe",
          5653 => x"18",
          5654 => x"31",
          5655 => x"a0",
          5656 => x"17",
          5657 => x"06",
          5658 => x"08",
          5659 => x"81",
          5660 => x"79",
          5661 => x"55",
          5662 => x"56",
          5663 => x"55",
          5664 => x"7a",
          5665 => x"75",
          5666 => x"78",
          5667 => x"0b",
          5668 => x"34",
          5669 => x"0b",
          5670 => x"34",
          5671 => x"7b",
          5672 => x"e4",
          5673 => x"5b",
          5674 => x"39",
          5675 => x"3f",
          5676 => x"74",
          5677 => x"5a",
          5678 => x"70",
          5679 => x"e4",
          5680 => x"38",
          5681 => x"74",
          5682 => x"72",
          5683 => x"86",
          5684 => x"71",
          5685 => x"58",
          5686 => x"0c",
          5687 => x"0d",
          5688 => x"bc",
          5689 => x"53",
          5690 => x"56",
          5691 => x"70",
          5692 => x"38",
          5693 => x"9f",
          5694 => x"38",
          5695 => x"38",
          5696 => x"24",
          5697 => x"80",
          5698 => x"0d",
          5699 => x"8c",
          5700 => x"70",
          5701 => x"89",
          5702 => x"ff",
          5703 => x"2e",
          5704 => x"d4",
          5705 => x"76",
          5706 => x"81",
          5707 => x"54",
          5708 => x"12",
          5709 => x"9f",
          5710 => x"e0",
          5711 => x"71",
          5712 => x"73",
          5713 => x"ff",
          5714 => x"70",
          5715 => x"52",
          5716 => x"18",
          5717 => x"ff",
          5718 => x"77",
          5719 => x"51",
          5720 => x"53",
          5721 => x"51",
          5722 => x"55",
          5723 => x"38",
          5724 => x"0d",
          5725 => x"d0",
          5726 => x"e4",
          5727 => x"c6",
          5728 => x"98",
          5729 => x"e2",
          5730 => x"2a",
          5731 => x"b2",
          5732 => x"12",
          5733 => x"5e",
          5734 => x"a4",
          5735 => x"b8",
          5736 => x"b8",
          5737 => x"ff",
          5738 => x"0c",
          5739 => x"94",
          5740 => x"2b",
          5741 => x"54",
          5742 => x"58",
          5743 => x"0d",
          5744 => x"3d",
          5745 => x"80",
          5746 => x"fd",
          5747 => x"cf",
          5748 => x"84",
          5749 => x"80",
          5750 => x"08",
          5751 => x"3d",
          5752 => x"cc",
          5753 => x"5b",
          5754 => x"3f",
          5755 => x"e4",
          5756 => x"3d",
          5757 => x"2e",
          5758 => x"17",
          5759 => x"81",
          5760 => x"16",
          5761 => x"b8",
          5762 => x"57",
          5763 => x"82",
          5764 => x"11",
          5765 => x"07",
          5766 => x"56",
          5767 => x"80",
          5768 => x"ff",
          5769 => x"59",
          5770 => x"80",
          5771 => x"84",
          5772 => x"08",
          5773 => x"11",
          5774 => x"07",
          5775 => x"56",
          5776 => x"7a",
          5777 => x"52",
          5778 => x"b8",
          5779 => x"80",
          5780 => x"83",
          5781 => x"e4",
          5782 => x"ff",
          5783 => x"33",
          5784 => x"82",
          5785 => x"33",
          5786 => x"17",
          5787 => x"76",
          5788 => x"05",
          5789 => x"11",
          5790 => x"58",
          5791 => x"ff",
          5792 => x"58",
          5793 => x"5a",
          5794 => x"82",
          5795 => x"33",
          5796 => x"70",
          5797 => x"5a",
          5798 => x"70",
          5799 => x"f5",
          5800 => x"ab",
          5801 => x"38",
          5802 => x"81",
          5803 => x"77",
          5804 => x"05",
          5805 => x"06",
          5806 => x"34",
          5807 => x"3d",
          5808 => x"33",
          5809 => x"79",
          5810 => x"95",
          5811 => x"2b",
          5812 => x"dd",
          5813 => x"51",
          5814 => x"08",
          5815 => x"fd",
          5816 => x"b4",
          5817 => x"81",
          5818 => x"3f",
          5819 => x"be",
          5820 => x"34",
          5821 => x"84",
          5822 => x"17",
          5823 => x"33",
          5824 => x"fb",
          5825 => x"a0",
          5826 => x"16",
          5827 => x"59",
          5828 => x"3d",
          5829 => x"80",
          5830 => x"10",
          5831 => x"33",
          5832 => x"2e",
          5833 => x"f1",
          5834 => x"19",
          5835 => x"05",
          5836 => x"38",
          5837 => x"59",
          5838 => x"5e",
          5839 => x"f5",
          5840 => x"84",
          5841 => x"04",
          5842 => x"89",
          5843 => x"08",
          5844 => x"33",
          5845 => x"14",
          5846 => x"78",
          5847 => x"5a",
          5848 => x"15",
          5849 => x"15",
          5850 => x"38",
          5851 => x"78",
          5852 => x"22",
          5853 => x"78",
          5854 => x"17",
          5855 => x"e4",
          5856 => x"55",
          5857 => x"e4",
          5858 => x"30",
          5859 => x"71",
          5860 => x"73",
          5861 => x"27",
          5862 => x"16",
          5863 => x"33",
          5864 => x"57",
          5865 => x"52",
          5866 => x"b8",
          5867 => x"80",
          5868 => x"98",
          5869 => x"79",
          5870 => x"aa",
          5871 => x"39",
          5872 => x"72",
          5873 => x"04",
          5874 => x"06",
          5875 => x"94",
          5876 => x"78",
          5877 => x"77",
          5878 => x"75",
          5879 => x"0c",
          5880 => x"76",
          5881 => x"59",
          5882 => x"08",
          5883 => x"0c",
          5884 => x"3d",
          5885 => x"88",
          5886 => x"fe",
          5887 => x"2e",
          5888 => x"b8",
          5889 => x"94",
          5890 => x"75",
          5891 => x"9c",
          5892 => x"73",
          5893 => x"22",
          5894 => x"78",
          5895 => x"80",
          5896 => x"56",
          5897 => x"ff",
          5898 => x"54",
          5899 => x"ff",
          5900 => x"81",
          5901 => x"75",
          5902 => x"52",
          5903 => x"b8",
          5904 => x"81",
          5905 => x"ff",
          5906 => x"08",
          5907 => x"fe",
          5908 => x"82",
          5909 => x"0d",
          5910 => x"54",
          5911 => x"8c",
          5912 => x"05",
          5913 => x"08",
          5914 => x"8f",
          5915 => x"84",
          5916 => x"7a",
          5917 => x"b9",
          5918 => x"84",
          5919 => x"16",
          5920 => x"78",
          5921 => x"84",
          5922 => x"2e",
          5923 => x"11",
          5924 => x"07",
          5925 => x"57",
          5926 => x"17",
          5927 => x"17",
          5928 => x"b9",
          5929 => x"84",
          5930 => x"84",
          5931 => x"85",
          5932 => x"95",
          5933 => x"2b",
          5934 => x"19",
          5935 => x"3d",
          5936 => x"2e",
          5937 => x"2e",
          5938 => x"2e",
          5939 => x"22",
          5940 => x"80",
          5941 => x"75",
          5942 => x"3d",
          5943 => x"ff",
          5944 => x"06",
          5945 => x"53",
          5946 => x"7c",
          5947 => x"9f",
          5948 => x"97",
          5949 => x"8f",
          5950 => x"59",
          5951 => x"80",
          5952 => x"c7",
          5953 => x"75",
          5954 => x"84",
          5955 => x"08",
          5956 => x"08",
          5957 => x"b2",
          5958 => x"99",
          5959 => x"32",
          5960 => x"84",
          5961 => x"72",
          5962 => x"04",
          5963 => x"b1",
          5964 => x"99",
          5965 => x"32",
          5966 => x"84",
          5967 => x"cf",
          5968 => x"f9",
          5969 => x"e4",
          5970 => x"33",
          5971 => x"e4",
          5972 => x"38",
          5973 => x"39",
          5974 => x"89",
          5975 => x"c1",
          5976 => x"84",
          5977 => x"74",
          5978 => x"04",
          5979 => x"3f",
          5980 => x"e4",
          5981 => x"33",
          5982 => x"24",
          5983 => x"76",
          5984 => x"74",
          5985 => x"04",
          5986 => x"3d",
          5987 => x"56",
          5988 => x"52",
          5989 => x"b8",
          5990 => x"9a",
          5991 => x"11",
          5992 => x"57",
          5993 => x"75",
          5994 => x"95",
          5995 => x"77",
          5996 => x"93",
          5997 => x"e4",
          5998 => x"38",
          5999 => x"b4",
          6000 => x"83",
          6001 => x"8d",
          6002 => x"52",
          6003 => x"3f",
          6004 => x"38",
          6005 => x"0c",
          6006 => x"38",
          6007 => x"8d",
          6008 => x"33",
          6009 => x"88",
          6010 => x"07",
          6011 => x"ff",
          6012 => x"80",
          6013 => x"ff",
          6014 => x"53",
          6015 => x"78",
          6016 => x"94",
          6017 => x"58",
          6018 => x"e4",
          6019 => x"b4",
          6020 => x"81",
          6021 => x"3f",
          6022 => x"f8",
          6023 => x"34",
          6024 => x"84",
          6025 => x"18",
          6026 => x"33",
          6027 => x"fe",
          6028 => x"a0",
          6029 => x"17",
          6030 => x"5e",
          6031 => x"3d",
          6032 => x"81",
          6033 => x"2e",
          6034 => x"81",
          6035 => x"08",
          6036 => x"80",
          6037 => x"58",
          6038 => x"ca",
          6039 => x"0c",
          6040 => x"84",
          6041 => x"b8",
          6042 => x"88",
          6043 => x"1f",
          6044 => x"5f",
          6045 => x"fd",
          6046 => x"fd",
          6047 => x"7f",
          6048 => x"33",
          6049 => x"fe",
          6050 => x"39",
          6051 => x"76",
          6052 => x"74",
          6053 => x"73",
          6054 => x"84",
          6055 => x"81",
          6056 => x"80",
          6057 => x"80",
          6058 => x"2a",
          6059 => x"80",
          6060 => x"54",
          6061 => x"73",
          6062 => x"08",
          6063 => x"9c",
          6064 => x"56",
          6065 => x"08",
          6066 => x"59",
          6067 => x"85",
          6068 => x"74",
          6069 => x"04",
          6070 => x"38",
          6071 => x"3f",
          6072 => x"e4",
          6073 => x"b8",
          6074 => x"84",
          6075 => x"38",
          6076 => x"85",
          6077 => x"c8",
          6078 => x"18",
          6079 => x"ff",
          6080 => x"84",
          6081 => x"17",
          6082 => x"a0",
          6083 => x"fe",
          6084 => x"81",
          6085 => x"77",
          6086 => x"0b",
          6087 => x"80",
          6088 => x"98",
          6089 => x"b9",
          6090 => x"81",
          6091 => x"2e",
          6092 => x"79",
          6093 => x"08",
          6094 => x"08",
          6095 => x"54",
          6096 => x"81",
          6097 => x"17",
          6098 => x"2e",
          6099 => x"51",
          6100 => x"08",
          6101 => x"38",
          6102 => x"3f",
          6103 => x"e4",
          6104 => x"b8",
          6105 => x"84",
          6106 => x"38",
          6107 => x"83",
          6108 => x"e6",
          6109 => x"18",
          6110 => x"90",
          6111 => x"16",
          6112 => x"34",
          6113 => x"38",
          6114 => x"58",
          6115 => x"39",
          6116 => x"fc",
          6117 => x"0b",
          6118 => x"39",
          6119 => x"59",
          6120 => x"18",
          6121 => x"b8",
          6122 => x"ff",
          6123 => x"a7",
          6124 => x"51",
          6125 => x"08",
          6126 => x"8a",
          6127 => x"3d",
          6128 => x"52",
          6129 => x"f8",
          6130 => x"b8",
          6131 => x"05",
          6132 => x"57",
          6133 => x"2b",
          6134 => x"80",
          6135 => x"57",
          6136 => x"a3",
          6137 => x"33",
          6138 => x"5e",
          6139 => x"d5",
          6140 => x"76",
          6141 => x"98",
          6142 => x"77",
          6143 => x"52",
          6144 => x"f9",
          6145 => x"b8",
          6146 => x"e4",
          6147 => x"3f",
          6148 => x"e4",
          6149 => x"e4",
          6150 => x"33",
          6151 => x"90",
          6152 => x"ff",
          6153 => x"2e",
          6154 => x"a1",
          6155 => x"57",
          6156 => x"38",
          6157 => x"3f",
          6158 => x"e4",
          6159 => x"70",
          6160 => x"80",
          6161 => x"38",
          6162 => x"27",
          6163 => x"81",
          6164 => x"38",
          6165 => x"b8",
          6166 => x"3d",
          6167 => x"08",
          6168 => x"2e",
          6169 => x"59",
          6170 => x"80",
          6171 => x"17",
          6172 => x"ee",
          6173 => x"85",
          6174 => x"18",
          6175 => x"19",
          6176 => x"83",
          6177 => x"fe",
          6178 => x"8b",
          6179 => x"84",
          6180 => x"38",
          6181 => x"cd",
          6182 => x"54",
          6183 => x"17",
          6184 => x"58",
          6185 => x"81",
          6186 => x"08",
          6187 => x"18",
          6188 => x"55",
          6189 => x"38",
          6190 => x"09",
          6191 => x"b4",
          6192 => x"7c",
          6193 => x"c5",
          6194 => x"55",
          6195 => x"52",
          6196 => x"b8",
          6197 => x"80",
          6198 => x"08",
          6199 => x"e4",
          6200 => x"53",
          6201 => x"3f",
          6202 => x"17",
          6203 => x"5c",
          6204 => x"81",
          6205 => x"81",
          6206 => x"55",
          6207 => x"56",
          6208 => x"39",
          6209 => x"39",
          6210 => x"0d",
          6211 => x"52",
          6212 => x"84",
          6213 => x"08",
          6214 => x"e4",
          6215 => x"6f",
          6216 => x"a6",
          6217 => x"84",
          6218 => x"84",
          6219 => x"84",
          6220 => x"06",
          6221 => x"70",
          6222 => x"56",
          6223 => x"52",
          6224 => x"c0",
          6225 => x"5c",
          6226 => x"56",
          6227 => x"f9",
          6228 => x"81",
          6229 => x"84",
          6230 => x"5a",
          6231 => x"9c",
          6232 => x"5b",
          6233 => x"22",
          6234 => x"5c",
          6235 => x"59",
          6236 => x"70",
          6237 => x"74",
          6238 => x"55",
          6239 => x"54",
          6240 => x"33",
          6241 => x"e4",
          6242 => x"dc",
          6243 => x"54",
          6244 => x"53",
          6245 => x"a5",
          6246 => x"be",
          6247 => x"34",
          6248 => x"55",
          6249 => x"38",
          6250 => x"09",
          6251 => x"b4",
          6252 => x"77",
          6253 => x"e5",
          6254 => x"7d",
          6255 => x"b4",
          6256 => x"ac",
          6257 => x"f9",
          6258 => x"b8",
          6259 => x"84",
          6260 => x"38",
          6261 => x"84",
          6262 => x"fe",
          6263 => x"fc",
          6264 => x"94",
          6265 => x"27",
          6266 => x"84",
          6267 => x"18",
          6268 => x"a1",
          6269 => x"3d",
          6270 => x"83",
          6271 => x"78",
          6272 => x"8b",
          6273 => x"70",
          6274 => x"75",
          6275 => x"18",
          6276 => x"19",
          6277 => x"34",
          6278 => x"80",
          6279 => x"d1",
          6280 => x"06",
          6281 => x"77",
          6282 => x"34",
          6283 => x"cc",
          6284 => x"1a",
          6285 => x"81",
          6286 => x"59",
          6287 => x"7d",
          6288 => x"64",
          6289 => x"57",
          6290 => x"88",
          6291 => x"75",
          6292 => x"38",
          6293 => x"79",
          6294 => x"e4",
          6295 => x"b6",
          6296 => x"96",
          6297 => x"17",
          6298 => x"cc",
          6299 => x"5d",
          6300 => x"59",
          6301 => x"79",
          6302 => x"90",
          6303 => x"0b",
          6304 => x"80",
          6305 => x"84",
          6306 => x"76",
          6307 => x"34",
          6308 => x"17",
          6309 => x"5b",
          6310 => x"2a",
          6311 => x"59",
          6312 => x"57",
          6313 => x"2a",
          6314 => x"2a",
          6315 => x"90",
          6316 => x"0b",
          6317 => x"98",
          6318 => x"96",
          6319 => x"3d",
          6320 => x"2e",
          6321 => x"33",
          6322 => x"2e",
          6323 => x"ba",
          6324 => x"3d",
          6325 => x"ff",
          6326 => x"56",
          6327 => x"38",
          6328 => x"0d",
          6329 => x"08",
          6330 => x"9f",
          6331 => x"84",
          6332 => x"bb",
          6333 => x"56",
          6334 => x"ae",
          6335 => x"81",
          6336 => x"59",
          6337 => x"99",
          6338 => x"55",
          6339 => x"70",
          6340 => x"74",
          6341 => x"51",
          6342 => x"08",
          6343 => x"38",
          6344 => x"38",
          6345 => x"3d",
          6346 => x"81",
          6347 => x"26",
          6348 => x"06",
          6349 => x"80",
          6350 => x"d4",
          6351 => x"5c",
          6352 => x"70",
          6353 => x"5a",
          6354 => x"e0",
          6355 => x"ff",
          6356 => x"38",
          6357 => x"55",
          6358 => x"75",
          6359 => x"77",
          6360 => x"30",
          6361 => x"5d",
          6362 => x"81",
          6363 => x"24",
          6364 => x"5b",
          6365 => x"b4",
          6366 => x"3d",
          6367 => x"ff",
          6368 => x"56",
          6369 => x"fd",
          6370 => x"09",
          6371 => x"ff",
          6372 => x"56",
          6373 => x"6f",
          6374 => x"05",
          6375 => x"70",
          6376 => x"05",
          6377 => x"38",
          6378 => x"34",
          6379 => x"06",
          6380 => x"07",
          6381 => x"81",
          6382 => x"70",
          6383 => x"80",
          6384 => x"6b",
          6385 => x"33",
          6386 => x"72",
          6387 => x"2e",
          6388 => x"08",
          6389 => x"82",
          6390 => x"29",
          6391 => x"80",
          6392 => x"58",
          6393 => x"83",
          6394 => x"81",
          6395 => x"17",
          6396 => x"b8",
          6397 => x"58",
          6398 => x"57",
          6399 => x"fb",
          6400 => x"ae",
          6401 => x"70",
          6402 => x"80",
          6403 => x"77",
          6404 => x"7a",
          6405 => x"75",
          6406 => x"34",
          6407 => x"18",
          6408 => x"34",
          6409 => x"08",
          6410 => x"38",
          6411 => x"3f",
          6412 => x"e4",
          6413 => x"98",
          6414 => x"08",
          6415 => x"7a",
          6416 => x"06",
          6417 => x"b8",
          6418 => x"e2",
          6419 => x"2e",
          6420 => x"b4",
          6421 => x"9c",
          6422 => x"0b",
          6423 => x"27",
          6424 => x"fc",
          6425 => x"84",
          6426 => x"38",
          6427 => x"38",
          6428 => x"51",
          6429 => x"08",
          6430 => x"04",
          6431 => x"3d",
          6432 => x"33",
          6433 => x"78",
          6434 => x"84",
          6435 => x"38",
          6436 => x"a0",
          6437 => x"3d",
          6438 => x"53",
          6439 => x"e2",
          6440 => x"08",
          6441 => x"38",
          6442 => x"b4",
          6443 => x"b8",
          6444 => x"08",
          6445 => x"5d",
          6446 => x"93",
          6447 => x"17",
          6448 => x"33",
          6449 => x"fd",
          6450 => x"53",
          6451 => x"52",
          6452 => x"84",
          6453 => x"b8",
          6454 => x"08",
          6455 => x"08",
          6456 => x"fc",
          6457 => x"82",
          6458 => x"81",
          6459 => x"05",
          6460 => x"fe",
          6461 => x"39",
          6462 => x"33",
          6463 => x"56",
          6464 => x"52",
          6465 => x"84",
          6466 => x"08",
          6467 => x"e4",
          6468 => x"66",
          6469 => x"96",
          6470 => x"84",
          6471 => x"cf",
          6472 => x"56",
          6473 => x"71",
          6474 => x"74",
          6475 => x"8b",
          6476 => x"16",
          6477 => x"84",
          6478 => x"96",
          6479 => x"57",
          6480 => x"97",
          6481 => x"b8",
          6482 => x"80",
          6483 => x"0c",
          6484 => x"52",
          6485 => x"d8",
          6486 => x"b8",
          6487 => x"05",
          6488 => x"75",
          6489 => x"19",
          6490 => x"56",
          6491 => x"55",
          6492 => x"58",
          6493 => x"54",
          6494 => x"0b",
          6495 => x"88",
          6496 => x"e4",
          6497 => x"0d",
          6498 => x"3d",
          6499 => x"a0",
          6500 => x"b8",
          6501 => x"08",
          6502 => x"80",
          6503 => x"5a",
          6504 => x"70",
          6505 => x"80",
          6506 => x"06",
          6507 => x"38",
          6508 => x"5a",
          6509 => x"38",
          6510 => x"7a",
          6511 => x"81",
          6512 => x"16",
          6513 => x"b8",
          6514 => x"57",
          6515 => x"57",
          6516 => x"58",
          6517 => x"38",
          6518 => x"38",
          6519 => x"11",
          6520 => x"71",
          6521 => x"72",
          6522 => x"62",
          6523 => x"76",
          6524 => x"04",
          6525 => x"3d",
          6526 => x"84",
          6527 => x"08",
          6528 => x"2e",
          6529 => x"7b",
          6530 => x"54",
          6531 => x"53",
          6532 => x"ad",
          6533 => x"7a",
          6534 => x"84",
          6535 => x"16",
          6536 => x"e4",
          6537 => x"27",
          6538 => x"74",
          6539 => x"38",
          6540 => x"08",
          6541 => x"51",
          6542 => x"54",
          6543 => x"33",
          6544 => x"e4",
          6545 => x"86",
          6546 => x"bb",
          6547 => x"b8",
          6548 => x"e4",
          6549 => x"59",
          6550 => x"57",
          6551 => x"19",
          6552 => x"70",
          6553 => x"80",
          6554 => x"11",
          6555 => x"2e",
          6556 => x"fd",
          6557 => x"a1",
          6558 => x"51",
          6559 => x"08",
          6560 => x"38",
          6561 => x"a0",
          6562 => x"15",
          6563 => x"08",
          6564 => x"58",
          6565 => x"38",
          6566 => x"81",
          6567 => x"81",
          6568 => x"ff",
          6569 => x"a1",
          6570 => x"e4",
          6571 => x"e4",
          6572 => x"80",
          6573 => x"0b",
          6574 => x"06",
          6575 => x"d6",
          6576 => x"38",
          6577 => x"06",
          6578 => x"38",
          6579 => x"38",
          6580 => x"a3",
          6581 => x"38",
          6582 => x"ff",
          6583 => x"55",
          6584 => x"81",
          6585 => x"5d",
          6586 => x"33",
          6587 => x"5a",
          6588 => x"3d",
          6589 => x"2e",
          6590 => x"02",
          6591 => x"5c",
          6592 => x"87",
          6593 => x"7d",
          6594 => x"70",
          6595 => x"b8",
          6596 => x"80",
          6597 => x"b8",
          6598 => x"b5",
          6599 => x"b8",
          6600 => x"74",
          6601 => x"b8",
          6602 => x"e5",
          6603 => x"52",
          6604 => x"b8",
          6605 => x"80",
          6606 => x"38",
          6607 => x"70",
          6608 => x"05",
          6609 => x"38",
          6610 => x"7d",
          6611 => x"e4",
          6612 => x"8a",
          6613 => x"ff",
          6614 => x"2e",
          6615 => x"55",
          6616 => x"08",
          6617 => x"b1",
          6618 => x"b8",
          6619 => x"81",
          6620 => x"19",
          6621 => x"59",
          6622 => x"83",
          6623 => x"81",
          6624 => x"53",
          6625 => x"fe",
          6626 => x"80",
          6627 => x"76",
          6628 => x"38",
          6629 => x"5a",
          6630 => x"38",
          6631 => x"56",
          6632 => x"81",
          6633 => x"81",
          6634 => x"84",
          6635 => x"08",
          6636 => x"76",
          6637 => x"76",
          6638 => x"80",
          6639 => x"15",
          6640 => x"0b",
          6641 => x"57",
          6642 => x"76",
          6643 => x"55",
          6644 => x"70",
          6645 => x"05",
          6646 => x"38",
          6647 => x"34",
          6648 => x"7d",
          6649 => x"e4",
          6650 => x"fe",
          6651 => x"53",
          6652 => x"d4",
          6653 => x"2e",
          6654 => x"b8",
          6655 => x"08",
          6656 => x"19",
          6657 => x"55",
          6658 => x"e4",
          6659 => x"81",
          6660 => x"84",
          6661 => x"08",
          6662 => x"39",
          6663 => x"fd",
          6664 => x"b4",
          6665 => x"7a",
          6666 => x"fd",
          6667 => x"60",
          6668 => x"33",
          6669 => x"2e",
          6670 => x"2e",
          6671 => x"2e",
          6672 => x"22",
          6673 => x"38",
          6674 => x"38",
          6675 => x"38",
          6676 => x"17",
          6677 => x"70",
          6678 => x"80",
          6679 => x"22",
          6680 => x"57",
          6681 => x"15",
          6682 => x"9f",
          6683 => x"1c",
          6684 => x"81",
          6685 => x"78",
          6686 => x"56",
          6687 => x"fe",
          6688 => x"55",
          6689 => x"82",
          6690 => x"81",
          6691 => x"2e",
          6692 => x"81",
          6693 => x"2e",
          6694 => x"06",
          6695 => x"84",
          6696 => x"87",
          6697 => x"0d",
          6698 => x"ac",
          6699 => x"54",
          6700 => x"55",
          6701 => x"81",
          6702 => x"80",
          6703 => x"81",
          6704 => x"52",
          6705 => x"b8",
          6706 => x"ff",
          6707 => x"57",
          6708 => x"90",
          6709 => x"8c",
          6710 => x"18",
          6711 => x"5c",
          6712 => x"fe",
          6713 => x"7a",
          6714 => x"94",
          6715 => x"5d",
          6716 => x"d6",
          6717 => x"5b",
          6718 => x"fe",
          6719 => x"ff",
          6720 => x"f0",
          6721 => x"a5",
          6722 => x"05",
          6723 => x"3d",
          6724 => x"2e",
          6725 => x"5b",
          6726 => x"ba",
          6727 => x"75",
          6728 => x"c0",
          6729 => x"38",
          6730 => x"70",
          6731 => x"38",
          6732 => x"d8",
          6733 => x"40",
          6734 => x"ce",
          6735 => x"ff",
          6736 => x"57",
          6737 => x"81",
          6738 => x"38",
          6739 => x"79",
          6740 => x"e4",
          6741 => x"80",
          6742 => x"80",
          6743 => x"06",
          6744 => x"2e",
          6745 => x"f8",
          6746 => x"f0",
          6747 => x"83",
          6748 => x"08",
          6749 => x"4c",
          6750 => x"38",
          6751 => x"56",
          6752 => x"7d",
          6753 => x"74",
          6754 => x"be",
          6755 => x"83",
          6756 => x"61",
          6757 => x"07",
          6758 => x"d5",
          6759 => x"7d",
          6760 => x"33",
          6761 => x"38",
          6762 => x"12",
          6763 => x"07",
          6764 => x"2b",
          6765 => x"83",
          6766 => x"2b",
          6767 => x"70",
          6768 => x"07",
          6769 => x"0c",
          6770 => x"59",
          6771 => x"57",
          6772 => x"93",
          6773 => x"38",
          6774 => x"49",
          6775 => x"87",
          6776 => x"61",
          6777 => x"83",
          6778 => x"58",
          6779 => x"ae",
          6780 => x"83",
          6781 => x"2e",
          6782 => x"83",
          6783 => x"70",
          6784 => x"86",
          6785 => x"52",
          6786 => x"b8",
          6787 => x"b8",
          6788 => x"81",
          6789 => x"b8",
          6790 => x"83",
          6791 => x"89",
          6792 => x"1f",
          6793 => x"05",
          6794 => x"57",
          6795 => x"74",
          6796 => x"60",
          6797 => x"f2",
          6798 => x"53",
          6799 => x"a9",
          6800 => x"83",
          6801 => x"09",
          6802 => x"f5",
          6803 => x"ac",
          6804 => x"55",
          6805 => x"74",
          6806 => x"84",
          6807 => x"b8",
          6808 => x"39",
          6809 => x"3d",
          6810 => x"33",
          6811 => x"57",
          6812 => x"1d",
          6813 => x"58",
          6814 => x"0b",
          6815 => x"7d",
          6816 => x"33",
          6817 => x"9f",
          6818 => x"89",
          6819 => x"58",
          6820 => x"26",
          6821 => x"06",
          6822 => x"5a",
          6823 => x"85",
          6824 => x"32",
          6825 => x"7b",
          6826 => x"80",
          6827 => x"5c",
          6828 => x"56",
          6829 => x"53",
          6830 => x"3f",
          6831 => x"b6",
          6832 => x"b8",
          6833 => x"bf",
          6834 => x"26",
          6835 => x"fb",
          6836 => x"7b",
          6837 => x"a3",
          6838 => x"81",
          6839 => x"fd",
          6840 => x"46",
          6841 => x"08",
          6842 => x"38",
          6843 => x"fb",
          6844 => x"e4",
          6845 => x"0c",
          6846 => x"99",
          6847 => x"74",
          6848 => x"ae",
          6849 => x"76",
          6850 => x"55",
          6851 => x"a0",
          6852 => x"58",
          6853 => x"ff",
          6854 => x"05",
          6855 => x"05",
          6856 => x"83",
          6857 => x"05",
          6858 => x"8f",
          6859 => x"62",
          6860 => x"61",
          6861 => x"06",
          6862 => x"56",
          6863 => x"38",
          6864 => x"61",
          6865 => x"6b",
          6866 => x"05",
          6867 => x"61",
          6868 => x"34",
          6869 => x"9c",
          6870 => x"61",
          6871 => x"6b",
          6872 => x"84",
          6873 => x"61",
          6874 => x"f7",
          6875 => x"61",
          6876 => x"34",
          6877 => x"83",
          6878 => x"05",
          6879 => x"97",
          6880 => x"34",
          6881 => x"ab",
          6882 => x"76",
          6883 => x"81",
          6884 => x"ef",
          6885 => x"d5",
          6886 => x"ff",
          6887 => x"60",
          6888 => x"81",
          6889 => x"38",
          6890 => x"9c",
          6891 => x"70",
          6892 => x"74",
          6893 => x"83",
          6894 => x"f8",
          6895 => x"57",
          6896 => x"45",
          6897 => x"34",
          6898 => x"81",
          6899 => x"75",
          6900 => x"66",
          6901 => x"7a",
          6902 => x"9d",
          6903 => x"38",
          6904 => x"70",
          6905 => x"74",
          6906 => x"58",
          6907 => x"40",
          6908 => x"56",
          6909 => x"65",
          6910 => x"55",
          6911 => x"51",
          6912 => x"08",
          6913 => x"31",
          6914 => x"62",
          6915 => x"83",
          6916 => x"62",
          6917 => x"84",
          6918 => x"5e",
          6919 => x"56",
          6920 => x"34",
          6921 => x"d5",
          6922 => x"83",
          6923 => x"67",
          6924 => x"34",
          6925 => x"84",
          6926 => x"52",
          6927 => x"fe",
          6928 => x"08",
          6929 => x"86",
          6930 => x"87",
          6931 => x"34",
          6932 => x"61",
          6933 => x"08",
          6934 => x"83",
          6935 => x"64",
          6936 => x"2a",
          6937 => x"62",
          6938 => x"05",
          6939 => x"79",
          6940 => x"84",
          6941 => x"53",
          6942 => x"3f",
          6943 => x"b6",
          6944 => x"e4",
          6945 => x"0c",
          6946 => x"1c",
          6947 => x"7a",
          6948 => x"0b",
          6949 => x"80",
          6950 => x"38",
          6951 => x"17",
          6952 => x"2e",
          6953 => x"77",
          6954 => x"84",
          6955 => x"05",
          6956 => x"80",
          6957 => x"8a",
          6958 => x"77",
          6959 => x"e4",
          6960 => x"f5",
          6961 => x"38",
          6962 => x"38",
          6963 => x"06",
          6964 => x"83",
          6965 => x"05",
          6966 => x"a1",
          6967 => x"61",
          6968 => x"76",
          6969 => x"80",
          6970 => x"80",
          6971 => x"05",
          6972 => x"34",
          6973 => x"2a",
          6974 => x"90",
          6975 => x"7c",
          6976 => x"34",
          6977 => x"ad",
          6978 => x"80",
          6979 => x"05",
          6980 => x"61",
          6981 => x"34",
          6982 => x"a9",
          6983 => x"80",
          6984 => x"55",
          6985 => x"70",
          6986 => x"74",
          6987 => x"81",
          6988 => x"58",
          6989 => x"f9",
          6990 => x"52",
          6991 => x"57",
          6992 => x"7d",
          6993 => x"83",
          6994 => x"e4",
          6995 => x"bf",
          6996 => x"84",
          6997 => x"b8",
          6998 => x"4a",
          6999 => x"ff",
          7000 => x"6a",
          7001 => x"61",
          7002 => x"34",
          7003 => x"88",
          7004 => x"ff",
          7005 => x"7c",
          7006 => x"1f",
          7007 => x"d5",
          7008 => x"75",
          7009 => x"57",
          7010 => x"7c",
          7011 => x"80",
          7012 => x"80",
          7013 => x"80",
          7014 => x"e4",
          7015 => x"05",
          7016 => x"34",
          7017 => x"7f",
          7018 => x"05",
          7019 => x"83",
          7020 => x"75",
          7021 => x"2a",
          7022 => x"82",
          7023 => x"83",
          7024 => x"05",
          7025 => x"80",
          7026 => x"81",
          7027 => x"51",
          7028 => x"1f",
          7029 => x"a5",
          7030 => x"39",
          7031 => x"80",
          7032 => x"76",
          7033 => x"8e",
          7034 => x"52",
          7035 => x"81",
          7036 => x"3d",
          7037 => x"74",
          7038 => x"17",
          7039 => x"77",
          7040 => x"55",
          7041 => x"b8",
          7042 => x"3d",
          7043 => x"33",
          7044 => x"38",
          7045 => x"9e",
          7046 => x"05",
          7047 => x"55",
          7048 => x"18",
          7049 => x"3d",
          7050 => x"74",
          7051 => x"ff",
          7052 => x"30",
          7053 => x"84",
          7054 => x"5a",
          7055 => x"51",
          7056 => x"3d",
          7057 => x"3d",
          7058 => x"80",
          7059 => x"15",
          7060 => x"77",
          7061 => x"7c",
          7062 => x"7d",
          7063 => x"75",
          7064 => x"b8",
          7065 => x"88",
          7066 => x"9e",
          7067 => x"75",
          7068 => x"ff",
          7069 => x"86",
          7070 => x"0b",
          7071 => x"04",
          7072 => x"54",
          7073 => x"9d",
          7074 => x"70",
          7075 => x"5a",
          7076 => x"76",
          7077 => x"7d",
          7078 => x"04",
          7079 => x"9a",
          7080 => x"80",
          7081 => x"ff",
          7082 => x"85",
          7083 => x"27",
          7084 => x"06",
          7085 => x"83",
          7086 => x"9c",
          7087 => x"06",
          7088 => x"38",
          7089 => x"22",
          7090 => x"70",
          7091 => x"53",
          7092 => x"02",
          7093 => x"05",
          7094 => x"ff",
          7095 => x"b8",
          7096 => x"83",
          7097 => x"70",
          7098 => x"83",
          7099 => x"e4",
          7100 => x"3d",
          7101 => x"26",
          7102 => x"06",
          7103 => x"ff",
          7104 => x"05",
          7105 => x"25",
          7106 => x"53",
          7107 => x"53",
          7108 => x"81",
          7109 => x"76",
          7110 => x"10",
          7111 => x"54",
          7112 => x"26",
          7113 => x"cb",
          7114 => x"0c",
          7115 => x"55",
          7116 => x"38",
          7117 => x"54",
          7118 => x"83",
          7119 => x"d3",
          7120 => x"ff",
          7121 => x"70",
          7122 => x"39",
          7123 => x"57",
          7124 => x"ff",
          7125 => x"16",
          7126 => x"c5",
          7127 => x"06",
          7128 => x"31",
          7129 => x"ff",
          7130 => x"39",
          7131 => x"22",
          7132 => x"00",
          7133 => x"ff",
          7134 => x"00",
          7135 => x"80",
          7136 => x"6a",
          7137 => x"54",
          7138 => x"3e",
          7139 => x"28",
          7140 => x"12",
          7141 => x"fc",
          7142 => x"e6",
          7143 => x"d0",
          7144 => x"ba",
          7145 => x"59",
          7146 => x"59",
          7147 => x"59",
          7148 => x"59",
          7149 => x"59",
          7150 => x"59",
          7151 => x"59",
          7152 => x"59",
          7153 => x"59",
          7154 => x"59",
          7155 => x"59",
          7156 => x"59",
          7157 => x"59",
          7158 => x"59",
          7159 => x"59",
          7160 => x"59",
          7161 => x"59",
          7162 => x"59",
          7163 => x"59",
          7164 => x"59",
          7165 => x"59",
          7166 => x"71",
          7167 => x"59",
          7168 => x"59",
          7169 => x"59",
          7170 => x"59",
          7171 => x"59",
          7172 => x"59",
          7173 => x"59",
          7174 => x"59",
          7175 => x"06",
          7176 => x"8a",
          7177 => x"67",
          7178 => x"ce",
          7179 => x"59",
          7180 => x"59",
          7181 => x"59",
          7182 => x"59",
          7183 => x"59",
          7184 => x"59",
          7185 => x"59",
          7186 => x"59",
          7187 => x"59",
          7188 => x"59",
          7189 => x"59",
          7190 => x"59",
          7191 => x"59",
          7192 => x"59",
          7193 => x"59",
          7194 => x"59",
          7195 => x"59",
          7196 => x"59",
          7197 => x"59",
          7198 => x"59",
          7199 => x"59",
          7200 => x"59",
          7201 => x"59",
          7202 => x"59",
          7203 => x"59",
          7204 => x"59",
          7205 => x"70",
          7206 => x"59",
          7207 => x"59",
          7208 => x"59",
          7209 => x"59",
          7210 => x"58",
          7211 => x"41",
          7212 => x"51",
          7213 => x"3a",
          7214 => x"2a",
          7215 => x"42",
          7216 => x"1e",
          7217 => x"74",
          7218 => x"3e",
          7219 => x"cd",
          7220 => x"63",
          7221 => x"92",
          7222 => x"19",
          7223 => x"f0",
          7224 => x"8a",
          7225 => x"cd",
          7226 => x"92",
          7227 => x"3e",
          7228 => x"84",
          7229 => x"ca",
          7230 => x"ef",
          7231 => x"94",
          7232 => x"51",
          7233 => x"51",
          7234 => x"51",
          7235 => x"51",
          7236 => x"51",
          7237 => x"51",
          7238 => x"51",
          7239 => x"51",
          7240 => x"51",
          7241 => x"51",
          7242 => x"51",
          7243 => x"51",
          7244 => x"51",
          7245 => x"51",
          7246 => x"69",
          7247 => x"44",
          7248 => x"5b",
          7249 => x"0c",
          7250 => x"51",
          7251 => x"fc",
          7252 => x"a5",
          7253 => x"ea",
          7254 => x"c6",
          7255 => x"51",
          7256 => x"f7",
          7257 => x"38",
          7258 => x"6c",
          7259 => x"21",
          7260 => x"78",
          7261 => x"ba",
          7262 => x"78",
          7263 => x"78",
          7264 => x"78",
          7265 => x"a2",
          7266 => x"78",
          7267 => x"78",
          7268 => x"78",
          7269 => x"78",
          7270 => x"78",
          7271 => x"78",
          7272 => x"78",
          7273 => x"78",
          7274 => x"78",
          7275 => x"78",
          7276 => x"78",
          7277 => x"78",
          7278 => x"c8",
          7279 => x"78",
          7280 => x"78",
          7281 => x"4f",
          7282 => x"32",
          7283 => x"10",
          7284 => x"10",
          7285 => x"10",
          7286 => x"eb",
          7287 => x"10",
          7288 => x"10",
          7289 => x"10",
          7290 => x"10",
          7291 => x"10",
          7292 => x"10",
          7293 => x"10",
          7294 => x"10",
          7295 => x"10",
          7296 => x"10",
          7297 => x"10",
          7298 => x"f5",
          7299 => x"cf",
          7300 => x"80",
          7301 => x"5d",
          7302 => x"4d",
          7303 => x"2b",
          7304 => x"07",
          7305 => x"67",
          7306 => x"3f",
          7307 => x"89",
          7308 => x"c6",
          7309 => x"c6",
          7310 => x"c6",
          7311 => x"c6",
          7312 => x"c6",
          7313 => x"c6",
          7314 => x"c6",
          7315 => x"c6",
          7316 => x"c6",
          7317 => x"c6",
          7318 => x"b4",
          7319 => x"c6",
          7320 => x"c6",
          7321 => x"c7",
          7322 => x"d4",
          7323 => x"b5",
          7324 => x"9f",
          7325 => x"89",
          7326 => x"6f",
          7327 => x"fd",
          7328 => x"49",
          7329 => x"fd",
          7330 => x"fd",
          7331 => x"fd",
          7332 => x"fd",
          7333 => x"7f",
          7334 => x"fd",
          7335 => x"fd",
          7336 => x"fd",
          7337 => x"fd",
          7338 => x"fd",
          7339 => x"fd",
          7340 => x"fd",
          7341 => x"fd",
          7342 => x"fd",
          7343 => x"fd",
          7344 => x"fd",
          7345 => x"fd",
          7346 => x"fd",
          7347 => x"fd",
          7348 => x"fd",
          7349 => x"fd",
          7350 => x"fd",
          7351 => x"fd",
          7352 => x"1d",
          7353 => x"fd",
          7354 => x"fd",
          7355 => x"fd",
          7356 => x"fd",
          7357 => x"fd",
          7358 => x"fd",
          7359 => x"fd",
          7360 => x"2b",
          7361 => x"b8",
          7362 => x"b8",
          7363 => x"e1",
          7364 => x"fd",
          7365 => x"fd",
          7366 => x"16",
          7367 => x"fd",
          7368 => x"58",
          7369 => x"18",
          7370 => x"fd",
          7371 => x"69",
          7372 => x"63",
          7373 => x"69",
          7374 => x"61",
          7375 => x"65",
          7376 => x"65",
          7377 => x"70",
          7378 => x"66",
          7379 => x"6d",
          7380 => x"00",
          7381 => x"00",
          7382 => x"00",
          7383 => x"00",
          7384 => x"00",
          7385 => x"74",
          7386 => x"65",
          7387 => x"6f",
          7388 => x"74",
          7389 => x"00",
          7390 => x"73",
          7391 => x"73",
          7392 => x"6f",
          7393 => x"00",
          7394 => x"20",
          7395 => x"00",
          7396 => x"65",
          7397 => x"72",
          7398 => x"00",
          7399 => x"79",
          7400 => x"69",
          7401 => x"00",
          7402 => x"63",
          7403 => x"6d",
          7404 => x"00",
          7405 => x"20",
          7406 => x"00",
          7407 => x"2c",
          7408 => x"69",
          7409 => x"65",
          7410 => x"00",
          7411 => x"61",
          7412 => x"00",
          7413 => x"61",
          7414 => x"69",
          7415 => x"6d",
          7416 => x"6f",
          7417 => x"00",
          7418 => x"74",
          7419 => x"64",
          7420 => x"76",
          7421 => x"72",
          7422 => x"61",
          7423 => x"00",
          7424 => x"72",
          7425 => x"74",
          7426 => x"00",
          7427 => x"6e",
          7428 => x"61",
          7429 => x"00",
          7430 => x"72",
          7431 => x"69",
          7432 => x"00",
          7433 => x"64",
          7434 => x"00",
          7435 => x"20",
          7436 => x"65",
          7437 => x"70",
          7438 => x"6e",
          7439 => x"66",
          7440 => x"6e",
          7441 => x"6b",
          7442 => x"61",
          7443 => x"65",
          7444 => x"72",
          7445 => x"6b",
          7446 => x"00",
          7447 => x"2e",
          7448 => x"75",
          7449 => x"25",
          7450 => x"75",
          7451 => x"73",
          7452 => x"00",
          7453 => x"00",
          7454 => x"00",
          7455 => x"58",
          7456 => x"00",
          7457 => x"00",
          7458 => x"00",
          7459 => x"20",
          7460 => x"00",
          7461 => x"00",
          7462 => x"30",
          7463 => x"31",
          7464 => x"55",
          7465 => x"30",
          7466 => x"25",
          7467 => x"00",
          7468 => x"65",
          7469 => x"61",
          7470 => x"00",
          7471 => x"58",
          7472 => x"75",
          7473 => x"54",
          7474 => x"74",
          7475 => x"00",
          7476 => x"58",
          7477 => x"75",
          7478 => x"54",
          7479 => x"74",
          7480 => x"00",
          7481 => x"52",
          7482 => x"75",
          7483 => x"54",
          7484 => x"74",
          7485 => x"00",
          7486 => x"65",
          7487 => x"00",
          7488 => x"6e",
          7489 => x"00",
          7490 => x"20",
          7491 => x"72",
          7492 => x"62",
          7493 => x"6d",
          7494 => x"00",
          7495 => x"63",
          7496 => x"00",
          7497 => x"2e",
          7498 => x"6c",
          7499 => x"6e",
          7500 => x"65",
          7501 => x"64",
          7502 => x"61",
          7503 => x"20",
          7504 => x"79",
          7505 => x"00",
          7506 => x"00",
          7507 => x"20",
          7508 => x"2e",
          7509 => x"00",
          7510 => x"5c",
          7511 => x"73",
          7512 => x"64",
          7513 => x"69",
          7514 => x"00",
          7515 => x"69",
          7516 => x"69",
          7517 => x"2e",
          7518 => x"6c",
          7519 => x"65",
          7520 => x"78",
          7521 => x"00",
          7522 => x"74",
          7523 => x"6f",
          7524 => x"2e",
          7525 => x"63",
          7526 => x"6f",
          7527 => x"38",
          7528 => x"00",
          7529 => x"30",
          7530 => x"00",
          7531 => x"30",
          7532 => x"70",
          7533 => x"2e",
          7534 => x"6c",
          7535 => x"2d",
          7536 => x"25",
          7537 => x"00",
          7538 => x"2e",
          7539 => x"6c",
          7540 => x"00",
          7541 => x"67",
          7542 => x"00",
          7543 => x"6d",
          7544 => x"6d",
          7545 => x"00",
          7546 => x"25",
          7547 => x"6f",
          7548 => x"75",
          7549 => x"61",
          7550 => x"6f",
          7551 => x"6d",
          7552 => x"00",
          7553 => x"25",
          7554 => x"3a",
          7555 => x"64",
          7556 => x"20",
          7557 => x"72",
          7558 => x"00",
          7559 => x"65",
          7560 => x"6d",
          7561 => x"00",
          7562 => x"65",
          7563 => x"20",
          7564 => x"65",
          7565 => x"72",
          7566 => x"73",
          7567 => x"0a",
          7568 => x"20",
          7569 => x"6f",
          7570 => x"74",
          7571 => x"73",
          7572 => x"0a",
          7573 => x"20",
          7574 => x"74",
          7575 => x"72",
          7576 => x"20",
          7577 => x"0a",
          7578 => x"63",
          7579 => x"20",
          7580 => x"20",
          7581 => x"20",
          7582 => x"20",
          7583 => x"0a",
          7584 => x"20",
          7585 => x"43",
          7586 => x"65",
          7587 => x"20",
          7588 => x"30",
          7589 => x"00",
          7590 => x"68",
          7591 => x"52",
          7592 => x"6b",
          7593 => x"25",
          7594 => x"48",
          7595 => x"20",
          7596 => x"6c",
          7597 => x"71",
          7598 => x"20",
          7599 => x"30",
          7600 => x"00",
          7601 => x"00",
          7602 => x"00",
          7603 => x"54",
          7604 => x"20",
          7605 => x"00",
          7606 => x"48",
          7607 => x"53",
          7608 => x"20",
          7609 => x"52",
          7610 => x"6e",
          7611 => x"64",
          7612 => x"20",
          7613 => x"20",
          7614 => x"72",
          7615 => x"64",
          7616 => x"20",
          7617 => x"20",
          7618 => x"63",
          7619 => x"64",
          7620 => x"20",
          7621 => x"20",
          7622 => x"3a",
          7623 => x"00",
          7624 => x"4d",
          7625 => x"25",
          7626 => x"58",
          7627 => x"20",
          7628 => x"41",
          7629 => x"3a",
          7630 => x"00",
          7631 => x"41",
          7632 => x"25",
          7633 => x"58",
          7634 => x"20",
          7635 => x"4d",
          7636 => x"3a",
          7637 => x"00",
          7638 => x"53",
          7639 => x"69",
          7640 => x"6e",
          7641 => x"6d",
          7642 => x"6c",
          7643 => x"69",
          7644 => x"78",
          7645 => x"00",
          7646 => x"00",
          7647 => x"44",
          7648 => x"03",
          7649 => x"00",
          7650 => x"3c",
          7651 => x"05",
          7652 => x"00",
          7653 => x"34",
          7654 => x"07",
          7655 => x"00",
          7656 => x"2c",
          7657 => x"08",
          7658 => x"00",
          7659 => x"24",
          7660 => x"09",
          7661 => x"00",
          7662 => x"1c",
          7663 => x"0d",
          7664 => x"00",
          7665 => x"14",
          7666 => x"0e",
          7667 => x"00",
          7668 => x"0c",
          7669 => x"0f",
          7670 => x"00",
          7671 => x"04",
          7672 => x"11",
          7673 => x"00",
          7674 => x"fc",
          7675 => x"13",
          7676 => x"00",
          7677 => x"f4",
          7678 => x"15",
          7679 => x"00",
          7680 => x"00",
          7681 => x"7e",
          7682 => x"00",
          7683 => x"7e",
          7684 => x"00",
          7685 => x"00",
          7686 => x"00",
          7687 => x"00",
          7688 => x"00",
          7689 => x"00",
          7690 => x"6f",
          7691 => x"61",
          7692 => x"6f",
          7693 => x"2c",
          7694 => x"69",
          7695 => x"74",
          7696 => x"74",
          7697 => x"00",
          7698 => x"25",
          7699 => x"6c",
          7700 => x"65",
          7701 => x"20",
          7702 => x"20",
          7703 => x"20",
          7704 => x"00",
          7705 => x"00",
          7706 => x"00",
          7707 => x"00",
          7708 => x"00",
          7709 => x"00",
          7710 => x"00",
          7711 => x"00",
          7712 => x"00",
          7713 => x"00",
          7714 => x"00",
          7715 => x"00",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"00",
          7721 => x"7e",
          7722 => x"7e",
          7723 => x"64",
          7724 => x"25",
          7725 => x"3a",
          7726 => x"00",
          7727 => x"2d",
          7728 => x"64",
          7729 => x"00",
          7730 => x"64",
          7731 => x"78",
          7732 => x"25",
          7733 => x"00",
          7734 => x"43",
          7735 => x"00",
          7736 => x"20",
          7737 => x"00",
          7738 => x"20",
          7739 => x"00",
          7740 => x"20",
          7741 => x"74",
          7742 => x"69",
          7743 => x"00",
          7744 => x"3c",
          7745 => x"00",
          7746 => x"00",
          7747 => x"33",
          7748 => x"4d",
          7749 => x"00",
          7750 => x"20",
          7751 => x"20",
          7752 => x"4e",
          7753 => x"46",
          7754 => x"00",
          7755 => x"00",
          7756 => x"00",
          7757 => x"12",
          7758 => x"00",
          7759 => x"80",
          7760 => x"8f",
          7761 => x"55",
          7762 => x"9f",
          7763 => x"a7",
          7764 => x"af",
          7765 => x"b7",
          7766 => x"bf",
          7767 => x"c7",
          7768 => x"cf",
          7769 => x"d7",
          7770 => x"df",
          7771 => x"e7",
          7772 => x"ef",
          7773 => x"f7",
          7774 => x"ff",
          7775 => x"2f",
          7776 => x"7c",
          7777 => x"04",
          7778 => x"00",
          7779 => x"02",
          7780 => x"20",
          7781 => x"fc",
          7782 => x"e0",
          7783 => x"eb",
          7784 => x"ec",
          7785 => x"e6",
          7786 => x"f2",
          7787 => x"d6",
          7788 => x"a5",
          7789 => x"ed",
          7790 => x"d1",
          7791 => x"10",
          7792 => x"a1",
          7793 => x"92",
          7794 => x"61",
          7795 => x"63",
          7796 => x"5c",
          7797 => x"34",
          7798 => x"3c",
          7799 => x"54",
          7800 => x"50",
          7801 => x"64",
          7802 => x"52",
          7803 => x"18",
          7804 => x"8c",
          7805 => x"df",
          7806 => x"c3",
          7807 => x"98",
          7808 => x"c6",
          7809 => x"b1",
          7810 => x"21",
          7811 => x"19",
          7812 => x"b2",
          7813 => x"1a",
          7814 => x"07",
          7815 => x"00",
          7816 => x"39",
          7817 => x"79",
          7818 => x"43",
          7819 => x"84",
          7820 => x"87",
          7821 => x"8b",
          7822 => x"90",
          7823 => x"94",
          7824 => x"98",
          7825 => x"9c",
          7826 => x"a0",
          7827 => x"a4",
          7828 => x"a7",
          7829 => x"ac",
          7830 => x"af",
          7831 => x"b3",
          7832 => x"b8",
          7833 => x"bc",
          7834 => x"c0",
          7835 => x"c4",
          7836 => x"c8",
          7837 => x"ca",
          7838 => x"01",
          7839 => x"f3",
          7840 => x"f4",
          7841 => x"12",
          7842 => x"3b",
          7843 => x"3f",
          7844 => x"46",
          7845 => x"81",
          7846 => x"8a",
          7847 => x"90",
          7848 => x"5f",
          7849 => x"94",
          7850 => x"67",
          7851 => x"62",
          7852 => x"9c",
          7853 => x"73",
          7854 => x"77",
          7855 => x"7b",
          7856 => x"7f",
          7857 => x"a9",
          7858 => x"87",
          7859 => x"b2",
          7860 => x"8f",
          7861 => x"7b",
          7862 => x"ff",
          7863 => x"88",
          7864 => x"11",
          7865 => x"a3",
          7866 => x"03",
          7867 => x"d8",
          7868 => x"f9",
          7869 => x"f6",
          7870 => x"fa",
          7871 => x"50",
          7872 => x"8a",
          7873 => x"cf",
          7874 => x"44",
          7875 => x"00",
          7876 => x"00",
          7877 => x"00",
          7878 => x"20",
          7879 => x"40",
          7880 => x"59",
          7881 => x"5d",
          7882 => x"08",
          7883 => x"bb",
          7884 => x"cb",
          7885 => x"f9",
          7886 => x"fb",
          7887 => x"08",
          7888 => x"04",
          7889 => x"bc",
          7890 => x"d0",
          7891 => x"e5",
          7892 => x"01",
          7893 => x"32",
          7894 => x"01",
          7895 => x"30",
          7896 => x"67",
          7897 => x"80",
          7898 => x"41",
          7899 => x"00",
          7900 => x"00",
          7901 => x"00",
          7902 => x"00",
          7903 => x"00",
          7904 => x"00",
          7905 => x"00",
          7906 => x"00",
          7907 => x"00",
          7908 => x"00",
          7909 => x"00",
          7910 => x"00",
          7911 => x"00",
          7912 => x"00",
          7913 => x"00",
          7914 => x"00",
          7915 => x"00",
          7916 => x"00",
          7917 => x"00",
          7918 => x"00",
          7919 => x"00",
          7920 => x"00",
          7921 => x"00",
          7922 => x"00",
          7923 => x"00",
          7924 => x"00",
          7925 => x"00",
          7926 => x"00",
          7927 => x"00",
          7928 => x"00",
          7929 => x"00",
          7930 => x"00",
          7931 => x"00",
          7932 => x"00",
          7933 => x"00",
          7934 => x"00",
          7935 => x"00",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"00",
          7940 => x"00",
          7941 => x"00",
          7942 => x"00",
          7943 => x"00",
          7944 => x"00",
          7945 => x"00",
          7946 => x"00",
          7947 => x"00",
          7948 => x"00",
          7949 => x"00",
          7950 => x"00",
          7951 => x"00",
          7952 => x"00",
          7953 => x"00",
          7954 => x"00",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"00",
          7959 => x"00",
          7960 => x"00",
          7961 => x"00",
          7962 => x"00",
          7963 => x"00",
          7964 => x"00",
          7965 => x"01",
          7966 => x"01",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"78",
          7980 => x"80",
          7981 => x"88",
          7982 => x"80",
          7983 => x"0d",
          7984 => x"f0",
          7985 => x"78",
          7986 => x"70",
          7987 => x"68",
          7988 => x"38",
          7989 => x"2e",
          7990 => x"2f",
          7991 => x"f0",
          7992 => x"f0",
          7993 => x"0d",
          7994 => x"f0",
          7995 => x"58",
          7996 => x"50",
          7997 => x"48",
          7998 => x"38",
          7999 => x"2e",
          8000 => x"2f",
          8001 => x"f0",
          8002 => x"f0",
          8003 => x"0d",
          8004 => x"f0",
          8005 => x"58",
          8006 => x"50",
          8007 => x"48",
          8008 => x"28",
          8009 => x"3e",
          8010 => x"2f",
          8011 => x"f0",
          8012 => x"f0",
          8013 => x"f0",
          8014 => x"f0",
          8015 => x"18",
          8016 => x"10",
          8017 => x"08",
          8018 => x"f0",
          8019 => x"f0",
          8020 => x"1c",
          8021 => x"f0",
          8022 => x"f0",
          8023 => x"cd",
          8024 => x"f0",
          8025 => x"dd",
          8026 => x"b1",
          8027 => x"73",
          8028 => x"a2",
          8029 => x"b9",
          8030 => x"be",
          8031 => x"f0",
          8032 => x"f0",
          8033 => x"00",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"00",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"f3",
          9069 => x"fb",
          9070 => x"c3",
          9071 => x"e6",
          9072 => x"63",
          9073 => x"6a",
          9074 => x"23",
          9075 => x"2c",
          9076 => x"03",
          9077 => x"0b",
          9078 => x"13",
          9079 => x"52",
          9080 => x"83",
          9081 => x"8b",
          9082 => x"93",
          9083 => x"bc",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"03",
          9100 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"87",
             1 => x"e9",
             2 => x"00",
             3 => x"00",
             4 => x"8c",
             5 => x"90",
             6 => x"00",
             7 => x"00",
             8 => x"06",
             9 => x"82",
            10 => x"06",
            11 => x"00",
            12 => x"06",
            13 => x"09",
            14 => x"09",
            15 => x"0b",
            16 => x"81",
            17 => x"09",
            18 => x"81",
            19 => x"00",
            20 => x"24",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"05",
            26 => x"0a",
            27 => x"53",
            28 => x"26",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"9f",
            45 => x"93",
            46 => x"00",
            47 => x"00",
            48 => x"2a",
            49 => x"09",
            50 => x"53",
            51 => x"00",
            52 => x"53",
            53 => x"81",
            54 => x"07",
            55 => x"00",
            56 => x"81",
            57 => x"09",
            58 => x"00",
            59 => x"00",
            60 => x"81",
            61 => x"09",
            62 => x"04",
            63 => x"00",
            64 => x"81",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"09",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"72",
            73 => x"51",
            74 => x"00",
            75 => x"00",
            76 => x"06",
            77 => x"83",
            78 => x"06",
            79 => x"00",
            80 => x"06",
            81 => x"83",
            82 => x"0b",
            83 => x"00",
            84 => x"8c",
            85 => x"0b",
            86 => x"56",
            87 => x"04",
            88 => x"8c",
            89 => x"0b",
            90 => x"56",
            91 => x"04",
            92 => x"70",
            93 => x"ff",
            94 => x"72",
            95 => x"51",
            96 => x"70",
            97 => x"06",
            98 => x"09",
            99 => x"51",
           100 => x"05",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"05",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"05",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"05",
           125 => x"04",
           126 => x"ff",
           127 => x"ff",
           128 => x"06",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"85",
           134 => x"0b",
           135 => x"0b",
           136 => x"c6",
           137 => x"0b",
           138 => x"0b",
           139 => x"86",
           140 => x"0b",
           141 => x"0b",
           142 => x"c6",
           143 => x"0b",
           144 => x"0b",
           145 => x"8a",
           146 => x"0b",
           147 => x"0b",
           148 => x"ce",
           149 => x"0b",
           150 => x"0b",
           151 => x"92",
           152 => x"0b",
           153 => x"0b",
           154 => x"d6",
           155 => x"0b",
           156 => x"0b",
           157 => x"9a",
           158 => x"0b",
           159 => x"0b",
           160 => x"de",
           161 => x"0b",
           162 => x"0b",
           163 => x"a2",
           164 => x"0b",
           165 => x"0b",
           166 => x"e6",
           167 => x"0b",
           168 => x"0b",
           169 => x"aa",
           170 => x"0b",
           171 => x"0b",
           172 => x"ed",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"8c",
           193 => x"d5",
           194 => x"c0",
           195 => x"a2",
           196 => x"c0",
           197 => x"a0",
           198 => x"c0",
           199 => x"a0",
           200 => x"c0",
           201 => x"94",
           202 => x"c0",
           203 => x"a1",
           204 => x"c0",
           205 => x"af",
           206 => x"c0",
           207 => x"ad",
           208 => x"c0",
           209 => x"94",
           210 => x"c0",
           211 => x"95",
           212 => x"c0",
           213 => x"95",
           214 => x"c0",
           215 => x"b1",
           216 => x"c0",
           217 => x"80",
           218 => x"80",
           219 => x"0c",
           220 => x"08",
           221 => x"f0",
           222 => x"f0",
           223 => x"b8",
           224 => x"b8",
           225 => x"84",
           226 => x"84",
           227 => x"04",
           228 => x"2d",
           229 => x"90",
           230 => x"8d",
           231 => x"80",
           232 => x"d7",
           233 => x"c0",
           234 => x"82",
           235 => x"80",
           236 => x"0c",
           237 => x"08",
           238 => x"f0",
           239 => x"f0",
           240 => x"b8",
           241 => x"b8",
           242 => x"84",
           243 => x"84",
           244 => x"04",
           245 => x"2d",
           246 => x"90",
           247 => x"91",
           248 => x"80",
           249 => x"fe",
           250 => x"c0",
           251 => x"83",
           252 => x"80",
           253 => x"0c",
           254 => x"08",
           255 => x"f0",
           256 => x"f0",
           257 => x"b8",
           258 => x"b8",
           259 => x"84",
           260 => x"84",
           261 => x"04",
           262 => x"2d",
           263 => x"90",
           264 => x"fd",
           265 => x"80",
           266 => x"f6",
           267 => x"c0",
           268 => x"83",
           269 => x"80",
           270 => x"0c",
           271 => x"08",
           272 => x"f0",
           273 => x"f0",
           274 => x"b8",
           275 => x"b8",
           276 => x"84",
           277 => x"84",
           278 => x"04",
           279 => x"2d",
           280 => x"90",
           281 => x"b4",
           282 => x"80",
           283 => x"f3",
           284 => x"c0",
           285 => x"81",
           286 => x"80",
           287 => x"0c",
           288 => x"08",
           289 => x"f0",
           290 => x"f0",
           291 => x"b8",
           292 => x"b8",
           293 => x"84",
           294 => x"84",
           295 => x"04",
           296 => x"84",
           297 => x"04",
           298 => x"2d",
           299 => x"90",
           300 => x"ab",
           301 => x"80",
           302 => x"f1",
           303 => x"c0",
           304 => x"81",
           305 => x"80",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"04",
           311 => x"83",
           312 => x"10",
           313 => x"51",
           314 => x"06",
           315 => x"10",
           316 => x"ed",
           317 => x"b8",
           318 => x"38",
           319 => x"0b",
           320 => x"51",
           321 => x"0d",
           322 => x"08",
           323 => x"08",
           324 => x"04",
           325 => x"11",
           326 => x"25",
           327 => x"72",
           328 => x"38",
           329 => x"30",
           330 => x"55",
           331 => x"71",
           332 => x"fa",
           333 => x"b8",
           334 => x"b8",
           335 => x"34",
           336 => x"70",
           337 => x"54",
           338 => x"34",
           339 => x"88",
           340 => x"e4",
           341 => x"0d",
           342 => x"05",
           343 => x"3d",
           344 => x"e4",
           345 => x"80",
           346 => x"3d",
           347 => x"52",
           348 => x"04",
           349 => x"5d",
           350 => x"1e",
           351 => x"06",
           352 => x"2e",
           353 => x"33",
           354 => x"81",
           355 => x"80",
           356 => x"7e",
           357 => x"32",
           358 => x"55",
           359 => x"38",
           360 => x"06",
           361 => x"7a",
           362 => x"76",
           363 => x"73",
           364 => x"04",
           365 => x"10",
           366 => x"98",
           367 => x"8b",
           368 => x"5b",
           369 => x"38",
           370 => x"38",
           371 => x"f7",
           372 => x"09",
           373 => x"5a",
           374 => x"76",
           375 => x"52",
           376 => x"57",
           377 => x"7a",
           378 => x"78",
           379 => x"54",
           380 => x"80",
           381 => x"83",
           382 => x"73",
           383 => x"27",
           384 => x"eb",
           385 => x"fe",
           386 => x"59",
           387 => x"84",
           388 => x"06",
           389 => x"5e",
           390 => x"84",
           391 => x"b8",
           392 => x"72",
           393 => x"08",
           394 => x"05",
           395 => x"ca",
           396 => x"b8",
           397 => x"f4",
           398 => x"56",
           399 => x"80",
           400 => x"90",
           401 => x"81",
           402 => x"38",
           403 => x"80",
           404 => x"77",
           405 => x"05",
           406 => x"2a",
           407 => x"2e",
           408 => x"ff",
           409 => x"cc",
           410 => x"83",
           411 => x"74",
           412 => x"f0",
           413 => x"90",
           414 => x"53",
           415 => x"81",
           416 => x"38",
           417 => x"86",
           418 => x"54",
           419 => x"54",
           420 => x"81",
           421 => x"77",
           422 => x"80",
           423 => x"80",
           424 => x"51",
           425 => x"80",
           426 => x"2c",
           427 => x"38",
           428 => x"b2",
           429 => x"81",
           430 => x"55",
           431 => x"52",
           432 => x"81",
           433 => x"70",
           434 => x"24",
           435 => x"06",
           436 => x"38",
           437 => x"76",
           438 => x"80",
           439 => x"b8",
           440 => x"1e",
           441 => x"7d",
           442 => x"ec",
           443 => x"2e",
           444 => x"80",
           445 => x"2c",
           446 => x"91",
           447 => x"3f",
           448 => x"a0",
           449 => x"87",
           450 => x"07",
           451 => x"84",
           452 => x"06",
           453 => x"39",
           454 => x"0a",
           455 => x"72",
           456 => x"80",
           457 => x"5a",
           458 => x"70",
           459 => x"38",
           460 => x"80",
           461 => x"5f",
           462 => x"52",
           463 => x"ff",
           464 => x"57",
           465 => x"38",
           466 => x"33",
           467 => x"1a",
           468 => x"79",
           469 => x"7c",
           470 => x"51",
           471 => x"0a",
           472 => x"80",
           473 => x"90",
           474 => x"87",
           475 => x"7a",
           476 => x"60",
           477 => x"41",
           478 => x"7a",
           479 => x"f4",
           480 => x"7c",
           481 => x"f8",
           482 => x"7c",
           483 => x"f8",
           484 => x"08",
           485 => x"72",
           486 => x"3f",
           487 => x"06",
           488 => x"72",
           489 => x"80",
           490 => x"f7",
           491 => x"84",
           492 => x"58",
           493 => x"51",
           494 => x"83",
           495 => x"2b",
           496 => x"07",
           497 => x"38",
           498 => x"80",
           499 => x"2c",
           500 => x"d6",
           501 => x"3f",
           502 => x"bb",
           503 => x"fa",
           504 => x"ab",
           505 => x"7e",
           506 => x"39",
           507 => x"2b",
           508 => x"57",
           509 => x"ff",
           510 => x"fb",
           511 => x"2e",
           512 => x"52",
           513 => x"74",
           514 => x"f1",
           515 => x"98",
           516 => x"b7",
           517 => x"3f",
           518 => x"bb",
           519 => x"51",
           520 => x"83",
           521 => x"2b",
           522 => x"07",
           523 => x"52",
           524 => x"0d",
           525 => x"74",
           526 => x"04",
           527 => x"84",
           528 => x"81",
           529 => x"56",
           530 => x"2e",
           531 => x"70",
           532 => x"2e",
           533 => x"72",
           534 => x"84",
           535 => x"ff",
           536 => x"53",
           537 => x"c8",
           538 => x"08",
           539 => x"51",
           540 => x"b8",
           541 => x"57",
           542 => x"88",
           543 => x"7a",
           544 => x"70",
           545 => x"51",
           546 => x"2e",
           547 => x"81",
           548 => x"09",
           549 => x"84",
           550 => x"73",
           551 => x"80",
           552 => x"90",
           553 => x"e4",
           554 => x"70",
           555 => x"e3",
           556 => x"d4",
           557 => x"83",
           558 => x"7a",
           559 => x"32",
           560 => x"56",
           561 => x"06",
           562 => x"15",
           563 => x"91",
           564 => x"74",
           565 => x"08",
           566 => x"56",
           567 => x"0d",
           568 => x"51",
           569 => x"56",
           570 => x"15",
           571 => x"56",
           572 => x"11",
           573 => x"32",
           574 => x"54",
           575 => x"06",
           576 => x"81",
           577 => x"38",
           578 => x"80",
           579 => x"0c",
           580 => x"0c",
           581 => x"b8",
           582 => x"ff",
           583 => x"8c",
           584 => x"84",
           585 => x"3d",
           586 => x"55",
           587 => x"84",
           588 => x"38",
           589 => x"52",
           590 => x"38",
           591 => x"34",
           592 => x"87",
           593 => x"72",
           594 => x"fd",
           595 => x"54",
           596 => x"70",
           597 => x"81",
           598 => x"81",
           599 => x"84",
           600 => x"fc",
           601 => x"55",
           602 => x"73",
           603 => x"93",
           604 => x"73",
           605 => x"51",
           606 => x"0c",
           607 => x"73",
           608 => x"53",
           609 => x"71",
           610 => x"80",
           611 => x"53",
           612 => x"51",
           613 => x"0d",
           614 => x"05",
           615 => x"12",
           616 => x"51",
           617 => x"75",
           618 => x"81",
           619 => x"81",
           620 => x"84",
           621 => x"fd",
           622 => x"55",
           623 => x"71",
           624 => x"81",
           625 => x"ef",
           626 => x"3d",
           627 => x"7a",
           628 => x"38",
           629 => x"33",
           630 => x"06",
           631 => x"2e",
           632 => x"38",
           633 => x"86",
           634 => x"38",
           635 => x"2e",
           636 => x"51",
           637 => x"31",
           638 => x"04",
           639 => x"0d",
           640 => x"70",
           641 => x"e4",
           642 => x"52",
           643 => x"e4",
           644 => x"2e",
           645 => x"54",
           646 => x"84",
           647 => x"84",
           648 => x"e4",
           649 => x"0d",
           650 => x"54",
           651 => x"81",
           652 => x"8c",
           653 => x"09",
           654 => x"75",
           655 => x"0c",
           656 => x"75",
           657 => x"70",
           658 => x"81",
           659 => x"f4",
           660 => x"3d",
           661 => x"58",
           662 => x"38",
           663 => x"e4",
           664 => x"2e",
           665 => x"71",
           666 => x"52",
           667 => x"52",
           668 => x"13",
           669 => x"71",
           670 => x"74",
           671 => x"9f",
           672 => x"72",
           673 => x"06",
           674 => x"1c",
           675 => x"53",
           676 => x"52",
           677 => x"0d",
           678 => x"80",
           679 => x"80",
           680 => x"75",
           681 => x"70",
           682 => x"71",
           683 => x"06",
           684 => x"84",
           685 => x"75",
           686 => x"70",
           687 => x"71",
           688 => x"81",
           689 => x"75",
           690 => x"52",
           691 => x"55",
           692 => x"51",
           693 => x"04",
           694 => x"71",
           695 => x"b8",
           696 => x"84",
           697 => x"04",
           698 => x"a0",
           699 => x"51",
           700 => x"53",
           701 => x"38",
           702 => x"b8",
           703 => x"9f",
           704 => x"9f",
           705 => x"2a",
           706 => x"54",
           707 => x"a8",
           708 => x"74",
           709 => x"11",
           710 => x"06",
           711 => x"52",
           712 => x"38",
           713 => x"0d",
           714 => x"7a",
           715 => x"7c",
           716 => x"71",
           717 => x"59",
           718 => x"84",
           719 => x"84",
           720 => x"f7",
           721 => x"70",
           722 => x"56",
           723 => x"8f",
           724 => x"33",
           725 => x"73",
           726 => x"2e",
           727 => x"56",
           728 => x"58",
           729 => x"38",
           730 => x"14",
           731 => x"14",
           732 => x"73",
           733 => x"ff",
           734 => x"89",
           735 => x"77",
           736 => x"0c",
           737 => x"26",
           738 => x"38",
           739 => x"56",
           740 => x"0d",
           741 => x"70",
           742 => x"09",
           743 => x"70",
           744 => x"80",
           745 => x"80",
           746 => x"74",
           747 => x"56",
           748 => x"38",
           749 => x"0d",
           750 => x"0c",
           751 => x"ca",
           752 => x"8b",
           753 => x"7d",
           754 => x"08",
           755 => x"2e",
           756 => x"70",
           757 => x"a0",
           758 => x"f5",
           759 => x"d0",
           760 => x"80",
           761 => x"74",
           762 => x"27",
           763 => x"06",
           764 => x"06",
           765 => x"f9",
           766 => x"89",
           767 => x"27",
           768 => x"81",
           769 => x"56",
           770 => x"78",
           771 => x"75",
           772 => x"e4",
           773 => x"16",
           774 => x"59",
           775 => x"ff",
           776 => x"33",
           777 => x"38",
           778 => x"38",
           779 => x"d0",
           780 => x"73",
           781 => x"e4",
           782 => x"81",
           783 => x"55",
           784 => x"84",
           785 => x"80",
           786 => x"81",
           787 => x"ff",
           788 => x"8c",
           789 => x"05",
           790 => x"51",
           791 => x"83",
           792 => x"3d",
           793 => x"a8",
           794 => x"cc",
           795 => x"04",
           796 => x"83",
           797 => x"ef",
           798 => x"cf",
           799 => x"0d",
           800 => x"3f",
           801 => x"51",
           802 => x"83",
           803 => x"3d",
           804 => x"d0",
           805 => x"94",
           806 => x"04",
           807 => x"83",
           808 => x"ee",
           809 => x"d0",
           810 => x"0d",
           811 => x"3f",
           812 => x"51",
           813 => x"83",
           814 => x"3d",
           815 => x"f8",
           816 => x"a8",
           817 => x"04",
           818 => x"83",
           819 => x"02",
           820 => x"58",
           821 => x"73",
           822 => x"75",
           823 => x"74",
           824 => x"55",
           825 => x"53",
           826 => x"82",
           827 => x"57",
           828 => x"d0",
           829 => x"76",
           830 => x"30",
           831 => x"57",
           832 => x"c0",
           833 => x"26",
           834 => x"e8",
           835 => x"e4",
           836 => x"52",
           837 => x"76",
           838 => x"04",
           839 => x"88",
           840 => x"3d",
           841 => x"52",
           842 => x"b8",
           843 => x"ff",
           844 => x"ff",
           845 => x"59",
           846 => x"f4",
           847 => x"78",
           848 => x"08",
           849 => x"83",
           850 => x"97",
           851 => x"05",
           852 => x"80",
           853 => x"3f",
           854 => x"80",
           855 => x"38",
           856 => x"0d",
           857 => x"61",
           858 => x"7f",
           859 => x"e4",
           860 => x"0d",
           861 => x"02",
           862 => x"73",
           863 => x"5d",
           864 => x"7a",
           865 => x"3f",
           866 => x"80",
           867 => x"90",
           868 => x"82",
           869 => x"27",
           870 => x"d1",
           871 => x"84",
           872 => x"ec",
           873 => x"83",
           874 => x"56",
           875 => x"18",
           876 => x"7a",
           877 => x"9f",
           878 => x"73",
           879 => x"74",
           880 => x"27",
           881 => x"52",
           882 => x"56",
           883 => x"84",
           884 => x"1c",
           885 => x"84",
           886 => x"2c",
           887 => x"38",
           888 => x"1e",
           889 => x"ff",
           890 => x"0d",
           891 => x"3f",
           892 => x"54",
           893 => x"26",
           894 => x"d2",
           895 => x"84",
           896 => x"ea",
           897 => x"38",
           898 => x"38",
           899 => x"db",
           900 => x"08",
           901 => x"78",
           902 => x"83",
           903 => x"14",
           904 => x"51",
           905 => x"ff",
           906 => x"df",
           907 => x"51",
           908 => x"c8",
           909 => x"3f",
           910 => x"39",
           911 => x"e9",
           912 => x"39",
           913 => x"08",
           914 => x"a8",
           915 => x"80",
           916 => x"38",
           917 => x"9b",
           918 => x"2b",
           919 => x"30",
           920 => x"07",
           921 => x"59",
           922 => x"e8",
           923 => x"b8",
           924 => x"70",
           925 => x"70",
           926 => x"06",
           927 => x"80",
           928 => x"39",
           929 => x"3d",
           930 => x"96",
           931 => x"51",
           932 => x"9c",
           933 => x"72",
           934 => x"71",
           935 => x"81",
           936 => x"72",
           937 => x"71",
           938 => x"81",
           939 => x"72",
           940 => x"71",
           941 => x"81",
           942 => x"72",
           943 => x"71",
           944 => x"53",
           945 => x"3d",
           946 => x"83",
           947 => x"51",
           948 => x"3d",
           949 => x"83",
           950 => x"51",
           951 => x"06",
           952 => x"39",
           953 => x"9c",
           954 => x"b7",
           955 => x"51",
           956 => x"c2",
           957 => x"d3",
           958 => x"9b",
           959 => x"06",
           960 => x"38",
           961 => x"3f",
           962 => x"80",
           963 => x"70",
           964 => x"fe",
           965 => x"9a",
           966 => x"ef",
           967 => x"84",
           968 => x"80",
           969 => x"81",
           970 => x"51",
           971 => x"3f",
           972 => x"52",
           973 => x"bd",
           974 => x"d3",
           975 => x"9a",
           976 => x"06",
           977 => x"38",
           978 => x"70",
           979 => x"0c",
           980 => x"fb",
           981 => x"06",
           982 => x"84",
           983 => x"b8",
           984 => x"51",
           985 => x"53",
           986 => x"0b",
           987 => x"ff",
           988 => x"f1",
           989 => x"78",
           990 => x"83",
           991 => x"80",
           992 => x"7b",
           993 => x"81",
           994 => x"2e",
           995 => x"be",
           996 => x"05",
           997 => x"84",
           998 => x"54",
           999 => x"da",
          1000 => x"84",
          1001 => x"80",
          1002 => x"5d",
          1003 => x"3d",
          1004 => x"38",
          1005 => x"3f",
          1006 => x"e4",
          1007 => x"b8",
          1008 => x"05",
          1009 => x"08",
          1010 => x"2e",
          1011 => x"51",
          1012 => x"8f",
          1013 => x"3d",
          1014 => x"38",
          1015 => x"81",
          1016 => x"53",
          1017 => x"dd",
          1018 => x"94",
          1019 => x"90",
          1020 => x"7c",
          1021 => x"08",
          1022 => x"70",
          1023 => x"42",
          1024 => x"81",
          1025 => x"2e",
          1026 => x"06",
          1027 => x"81",
          1028 => x"81",
          1029 => x"38",
          1030 => x"d5",
          1031 => x"80",
          1032 => x"bc",
          1033 => x"70",
          1034 => x"91",
          1035 => x"84",
          1036 => x"84",
          1037 => x"0b",
          1038 => x"cf",
          1039 => x"82",
          1040 => x"80",
          1041 => x"51",
          1042 => x"d8",
          1043 => x"7d",
          1044 => x"38",
          1045 => x"a1",
          1046 => x"ed",
          1047 => x"f8",
          1048 => x"70",
          1049 => x"39",
          1050 => x"59",
          1051 => x"78",
          1052 => x"79",
          1053 => x"52",
          1054 => x"7e",
          1055 => x"f3",
          1056 => x"09",
          1057 => x"9a",
          1058 => x"83",
          1059 => x"51",
          1060 => x"83",
          1061 => x"ac",
          1062 => x"7c",
          1063 => x"81",
          1064 => x"dd",
          1065 => x"51",
          1066 => x"8d",
          1067 => x"c0",
          1068 => x"04",
          1069 => x"d0",
          1070 => x"ff",
          1071 => x"ec",
          1072 => x"2e",
          1073 => x"f0",
          1074 => x"2d",
          1075 => x"a4",
          1076 => x"d6",
          1077 => x"39",
          1078 => x"80",
          1079 => x"e4",
          1080 => x"52",
          1081 => x"68",
          1082 => x"11",
          1083 => x"3f",
          1084 => x"dc",
          1085 => x"ff",
          1086 => x"b8",
          1087 => x"78",
          1088 => x"51",
          1089 => x"53",
          1090 => x"3f",
          1091 => x"2e",
          1092 => x"d3",
          1093 => x"cf",
          1094 => x"ff",
          1095 => x"b8",
          1096 => x"b8",
          1097 => x"05",
          1098 => x"08",
          1099 => x"53",
          1100 => x"a5",
          1101 => x"f8",
          1102 => x"48",
          1103 => x"c4",
          1104 => x"64",
          1105 => x"b8",
          1106 => x"05",
          1107 => x"08",
          1108 => x"fe",
          1109 => x"e9",
          1110 => x"2e",
          1111 => x"11",
          1112 => x"3f",
          1113 => x"f4",
          1114 => x"3f",
          1115 => x"83",
          1116 => x"5f",
          1117 => x"7a",
          1118 => x"52",
          1119 => x"66",
          1120 => x"47",
          1121 => x"11",
          1122 => x"3f",
          1123 => x"a4",
          1124 => x"ff",
          1125 => x"b8",
          1126 => x"b8",
          1127 => x"05",
          1128 => x"08",
          1129 => x"8c",
          1130 => x"67",
          1131 => x"70",
          1132 => x"81",
          1133 => x"84",
          1134 => x"93",
          1135 => x"f6",
          1136 => x"53",
          1137 => x"84",
          1138 => x"33",
          1139 => x"ed",
          1140 => x"f8",
          1141 => x"48",
          1142 => x"8c",
          1143 => x"68",
          1144 => x"02",
          1145 => x"81",
          1146 => x"53",
          1147 => x"84",
          1148 => x"38",
          1149 => x"79",
          1150 => x"fe",
          1151 => x"e7",
          1152 => x"bd",
          1153 => x"84",
          1154 => x"f3",
          1155 => x"f5",
          1156 => x"53",
          1157 => x"84",
          1158 => x"38",
          1159 => x"80",
          1160 => x"e4",
          1161 => x"46",
          1162 => x"68",
          1163 => x"38",
          1164 => x"5b",
          1165 => x"51",
          1166 => x"3d",
          1167 => x"84",
          1168 => x"05",
          1169 => x"84",
          1170 => x"83",
          1171 => x"f4",
          1172 => x"e7",
          1173 => x"ff",
          1174 => x"e5",
          1175 => x"38",
          1176 => x"2e",
          1177 => x"49",
          1178 => x"80",
          1179 => x"e4",
          1180 => x"5a",
          1181 => x"f1",
          1182 => x"11",
          1183 => x"3f",
          1184 => x"38",
          1185 => x"83",
          1186 => x"30",
          1187 => x"5c",
          1188 => x"7a",
          1189 => x"d7",
          1190 => x"68",
          1191 => x"eb",
          1192 => x"b0",
          1193 => x"0c",
          1194 => x"fe",
          1195 => x"e2",
          1196 => x"2e",
          1197 => x"59",
          1198 => x"f0",
          1199 => x"87",
          1200 => x"f2",
          1201 => x"05",
          1202 => x"7d",
          1203 => x"ff",
          1204 => x"b8",
          1205 => x"64",
          1206 => x"70",
          1207 => x"3d",
          1208 => x"51",
          1209 => x"ff",
          1210 => x"fe",
          1211 => x"e3",
          1212 => x"2e",
          1213 => x"db",
          1214 => x"49",
          1215 => x"11",
          1216 => x"3f",
          1217 => x"98",
          1218 => x"84",
          1219 => x"7a",
          1220 => x"38",
          1221 => x"53",
          1222 => x"f5",
          1223 => x"51",
          1224 => x"d7",
          1225 => x"39",
          1226 => x"80",
          1227 => x"e4",
          1228 => x"02",
          1229 => x"05",
          1230 => x"83",
          1231 => x"80",
          1232 => x"fc",
          1233 => x"7b",
          1234 => x"08",
          1235 => x"51",
          1236 => x"39",
          1237 => x"64",
          1238 => x"33",
          1239 => x"f1",
          1240 => x"d8",
          1241 => x"39",
          1242 => x"2e",
          1243 => x"fc",
          1244 => x"7d",
          1245 => x"08",
          1246 => x"33",
          1247 => x"f1",
          1248 => x"f1",
          1249 => x"38",
          1250 => x"39",
          1251 => x"2e",
          1252 => x"fb",
          1253 => x"80",
          1254 => x"d0",
          1255 => x"f3",
          1256 => x"34",
          1257 => x"57",
          1258 => x"d2",
          1259 => x"77",
          1260 => x"75",
          1261 => x"e4",
          1262 => x"9c",
          1263 => x"52",
          1264 => x"e4",
          1265 => x"87",
          1266 => x"3f",
          1267 => x"0c",
          1268 => x"84",
          1269 => x"94",
          1270 => x"c7",
          1271 => x"05",
          1272 => x"89",
          1273 => x"0c",
          1274 => x"3f",
          1275 => x"8d",
          1276 => x"52",
          1277 => x"83",
          1278 => x"87",
          1279 => x"b8",
          1280 => x"c0",
          1281 => x"ed",
          1282 => x"77",
          1283 => x"53",
          1284 => x"33",
          1285 => x"a0",
          1286 => x"15",
          1287 => x"53",
          1288 => x"81",
          1289 => x"82",
          1290 => x"e7",
          1291 => x"06",
          1292 => x"38",
          1293 => x"73",
          1294 => x"e1",
          1295 => x"54",
          1296 => x"38",
          1297 => x"70",
          1298 => x"72",
          1299 => x"81",
          1300 => x"51",
          1301 => x"0d",
          1302 => x"80",
          1303 => x"80",
          1304 => x"54",
          1305 => x"54",
          1306 => x"53",
          1307 => x"fe",
          1308 => x"76",
          1309 => x"84",
          1310 => x"86",
          1311 => x"87",
          1312 => x"e5",
          1313 => x"3d",
          1314 => x"11",
          1315 => x"70",
          1316 => x"33",
          1317 => x"26",
          1318 => x"83",
          1319 => x"85",
          1320 => x"26",
          1321 => x"85",
          1322 => x"88",
          1323 => x"e7",
          1324 => x"54",
          1325 => x"cc",
          1326 => x"0c",
          1327 => x"82",
          1328 => x"83",
          1329 => x"84",
          1330 => x"85",
          1331 => x"86",
          1332 => x"74",
          1333 => x"c0",
          1334 => x"98",
          1335 => x"e4",
          1336 => x"0d",
          1337 => x"81",
          1338 => x"5e",
          1339 => x"08",
          1340 => x"98",
          1341 => x"87",
          1342 => x"1c",
          1343 => x"79",
          1344 => x"08",
          1345 => x"98",
          1346 => x"87",
          1347 => x"1c",
          1348 => x"ff",
          1349 => x"58",
          1350 => x"56",
          1351 => x"54",
          1352 => x"ff",
          1353 => x"bf",
          1354 => x"3d",
          1355 => x"81",
          1356 => x"b0",
          1357 => x"70",
          1358 => x"09",
          1359 => x"e3",
          1360 => x"3d",
          1361 => x"3f",
          1362 => x"98",
          1363 => x"81",
          1364 => x"f0",
          1365 => x"70",
          1366 => x"d2",
          1367 => x"70",
          1368 => x"51",
          1369 => x"08",
          1370 => x"71",
          1371 => x"81",
          1372 => x"38",
          1373 => x"0d",
          1374 => x"33",
          1375 => x"06",
          1376 => x"f4",
          1377 => x"96",
          1378 => x"70",
          1379 => x"70",
          1380 => x"72",
          1381 => x"2e",
          1382 => x"52",
          1383 => x"51",
          1384 => x"2e",
          1385 => x"74",
          1386 => x"86",
          1387 => x"81",
          1388 => x"81",
          1389 => x"cb",
          1390 => x"71",
          1391 => x"84",
          1392 => x"53",
          1393 => x"ff",
          1394 => x"30",
          1395 => x"83",
          1396 => x"fa",
          1397 => x"70",
          1398 => x"e7",
          1399 => x"70",
          1400 => x"80",
          1401 => x"94",
          1402 => x"53",
          1403 => x"71",
          1404 => x"70",
          1405 => x"53",
          1406 => x"2a",
          1407 => x"81",
          1408 => x"52",
          1409 => x"94",
          1410 => x"75",
          1411 => x"76",
          1412 => x"04",
          1413 => x"51",
          1414 => x"06",
          1415 => x"93",
          1416 => x"ff",
          1417 => x"70",
          1418 => x"52",
          1419 => x"0d",
          1420 => x"2a",
          1421 => x"84",
          1422 => x"83",
          1423 => x"08",
          1424 => x"94",
          1425 => x"9e",
          1426 => x"c0",
          1427 => x"87",
          1428 => x"0c",
          1429 => x"b8",
          1430 => x"f1",
          1431 => x"83",
          1432 => x"08",
          1433 => x"bc",
          1434 => x"9e",
          1435 => x"c0",
          1436 => x"87",
          1437 => x"f1",
          1438 => x"83",
          1439 => x"08",
          1440 => x"8c",
          1441 => x"83",
          1442 => x"9e",
          1443 => x"51",
          1444 => x"83",
          1445 => x"9e",
          1446 => x"51",
          1447 => x"81",
          1448 => x"0b",
          1449 => x"80",
          1450 => x"2e",
          1451 => x"e7",
          1452 => x"08",
          1453 => x"52",
          1454 => x"71",
          1455 => x"c0",
          1456 => x"06",
          1457 => x"38",
          1458 => x"80",
          1459 => x"90",
          1460 => x"80",
          1461 => x"f1",
          1462 => x"90",
          1463 => x"52",
          1464 => x"52",
          1465 => x"87",
          1466 => x"80",
          1467 => x"83",
          1468 => x"34",
          1469 => x"70",
          1470 => x"70",
          1471 => x"83",
          1472 => x"9e",
          1473 => x"51",
          1474 => x"81",
          1475 => x"0b",
          1476 => x"80",
          1477 => x"83",
          1478 => x"34",
          1479 => x"06",
          1480 => x"f1",
          1481 => x"90",
          1482 => x"52",
          1483 => x"71",
          1484 => x"90",
          1485 => x"53",
          1486 => x"0b",
          1487 => x"06",
          1488 => x"38",
          1489 => x"87",
          1490 => x"70",
          1491 => x"04",
          1492 => x"0d",
          1493 => x"3f",
          1494 => x"aa",
          1495 => x"3f",
          1496 => x"fa",
          1497 => x"85",
          1498 => x"75",
          1499 => x"55",
          1500 => x"33",
          1501 => x"ef",
          1502 => x"f1",
          1503 => x"83",
          1504 => x"38",
          1505 => x"cf",
          1506 => x"83",
          1507 => x"74",
          1508 => x"56",
          1509 => x"33",
          1510 => x"cc",
          1511 => x"08",
          1512 => x"c5",
          1513 => x"d9",
          1514 => x"f1",
          1515 => x"ff",
          1516 => x"c2",
          1517 => x"83",
          1518 => x"83",
          1519 => x"52",
          1520 => x"e4",
          1521 => x"31",
          1522 => x"83",
          1523 => x"83",
          1524 => x"38",
          1525 => x"38",
          1526 => x"0d",
          1527 => x"84",
          1528 => x"84",
          1529 => x"76",
          1530 => x"08",
          1531 => x"ad",
          1532 => x"3d",
          1533 => x"bd",
          1534 => x"3f",
          1535 => x"29",
          1536 => x"e4",
          1537 => x"b3",
          1538 => x"74",
          1539 => x"39",
          1540 => x"83",
          1541 => x"f1",
          1542 => x"ff",
          1543 => x"52",
          1544 => x"3f",
          1545 => x"a8",
          1546 => x"d0",
          1547 => x"22",
          1548 => x"a5",
          1549 => x"84",
          1550 => x"84",
          1551 => x"76",
          1552 => x"08",
          1553 => x"fd",
          1554 => x"80",
          1555 => x"83",
          1556 => x"83",
          1557 => x"fd",
          1558 => x"94",
          1559 => x"ed",
          1560 => x"38",
          1561 => x"bf",
          1562 => x"74",
          1563 => x"83",
          1564 => x"83",
          1565 => x"fc",
          1566 => x"33",
          1567 => x"8d",
          1568 => x"80",
          1569 => x"f1",
          1570 => x"ff",
          1571 => x"55",
          1572 => x"39",
          1573 => x"80",
          1574 => x"f3",
          1575 => x"38",
          1576 => x"f1",
          1577 => x"a0",
          1578 => x"ef",
          1579 => x"38",
          1580 => x"f1",
          1581 => x"bc",
          1582 => x"ea",
          1583 => x"38",
          1584 => x"f1",
          1585 => x"d8",
          1586 => x"e9",
          1587 => x"38",
          1588 => x"f1",
          1589 => x"f4",
          1590 => x"e8",
          1591 => x"38",
          1592 => x"f1",
          1593 => x"90",
          1594 => x"eb",
          1595 => x"38",
          1596 => x"b0",
          1597 => x"bd",
          1598 => x"74",
          1599 => x"ff",
          1600 => x"71",
          1601 => x"83",
          1602 => x"83",
          1603 => x"83",
          1604 => x"ff",
          1605 => x"83",
          1606 => x"83",
          1607 => x"ff",
          1608 => x"83",
          1609 => x"83",
          1610 => x"ff",
          1611 => x"71",
          1612 => x"c0",
          1613 => x"08",
          1614 => x"3d",
          1615 => x"5a",
          1616 => x"83",
          1617 => x"3f",
          1618 => x"8b",
          1619 => x"08",
          1620 => x"82",
          1621 => x"80",
          1622 => x"3f",
          1623 => x"55",
          1624 => x"8e",
          1625 => x"70",
          1626 => x"09",
          1627 => x"51",
          1628 => x"73",
          1629 => x"8c",
          1630 => x"3f",
          1631 => x"76",
          1632 => x"0c",
          1633 => x"51",
          1634 => x"09",
          1635 => x"51",
          1636 => x"3f",
          1637 => x"08",
          1638 => x"51",
          1639 => x"b8",
          1640 => x"3d",
          1641 => x"71",
          1642 => x"57",
          1643 => x"0b",
          1644 => x"10",
          1645 => x"54",
          1646 => x"08",
          1647 => x"9a",
          1648 => x"84",
          1649 => x"88",
          1650 => x"16",
          1651 => x"76",
          1652 => x"b8",
          1653 => x"1a",
          1654 => x"ff",
          1655 => x"b8",
          1656 => x"1b",
          1657 => x"3f",
          1658 => x"54",
          1659 => x"70",
          1660 => x"27",
          1661 => x"33",
          1662 => x"e6",
          1663 => x"55",
          1664 => x"fe",
          1665 => x"80",
          1666 => x"39",
          1667 => x"f2",
          1668 => x"3f",
          1669 => x"83",
          1670 => x"77",
          1671 => x"e4",
          1672 => x"ff",
          1673 => x"55",
          1674 => x"9d",
          1675 => x"70",
          1676 => x"53",
          1677 => x"52",
          1678 => x"2e",
          1679 => x"0b",
          1680 => x"04",
          1681 => x"3d",
          1682 => x"80",
          1683 => x"33",
          1684 => x"9e",
          1685 => x"56",
          1686 => x"80",
          1687 => x"06",
          1688 => x"80",
          1689 => x"3d",
          1690 => x"84",
          1691 => x"2c",
          1692 => x"79",
          1693 => x"70",
          1694 => x"9c",
          1695 => x"71",
          1696 => x"dd",
          1697 => x"52",
          1698 => x"5c",
          1699 => x"cd",
          1700 => x"75",
          1701 => x"05",
          1702 => x"24",
          1703 => x"82",
          1704 => x"f0",
          1705 => x"91",
          1706 => x"70",
          1707 => x"95",
          1708 => x"84",
          1709 => x"2e",
          1710 => x"2b",
          1711 => x"70",
          1712 => x"2c",
          1713 => x"11",
          1714 => x"57",
          1715 => x"76",
          1716 => x"81",
          1717 => x"80",
          1718 => x"98",
          1719 => x"41",
          1720 => x"10",
          1721 => x"0b",
          1722 => x"77",
          1723 => x"15",
          1724 => x"61",
          1725 => x"ff",
          1726 => x"76",
          1727 => x"39",
          1728 => x"76",
          1729 => x"34",
          1730 => x"34",
          1731 => x"26",
          1732 => x"c3",
          1733 => x"dd",
          1734 => x"84",
          1735 => x"9c",
          1736 => x"56",
          1737 => x"d4",
          1738 => x"9b",
          1739 => x"57",
          1740 => x"39",
          1741 => x"06",
          1742 => x"75",
          1743 => x"c8",
          1744 => x"d0",
          1745 => x"55",
          1746 => x"7c",
          1747 => x"10",
          1748 => x"59",
          1749 => x"a4",
          1750 => x"33",
          1751 => x"80",
          1752 => x"52",
          1753 => x"d4",
          1754 => x"9b",
          1755 => x"51",
          1756 => x"33",
          1757 => x"34",
          1758 => x"38",
          1759 => x"84",
          1760 => x"8a",
          1761 => x"8d",
          1762 => x"fc",
          1763 => x"8e",
          1764 => x"2e",
          1765 => x"fd",
          1766 => x"a4",
          1767 => x"06",
          1768 => x"ff",
          1769 => x"84",
          1770 => x"2e",
          1771 => x"52",
          1772 => x"d4",
          1773 => x"83",
          1774 => x"51",
          1775 => x"33",
          1776 => x"34",
          1777 => x"84",
          1778 => x"84",
          1779 => x"79",
          1780 => x"08",
          1781 => x"a8",
          1782 => x"ff",
          1783 => x"70",
          1784 => x"5a",
          1785 => x"38",
          1786 => x"57",
          1787 => x"70",
          1788 => x"84",
          1789 => x"84",
          1790 => x"76",
          1791 => x"84",
          1792 => x"56",
          1793 => x"ff",
          1794 => x"75",
          1795 => x"ff",
          1796 => x"80",
          1797 => x"a0",
          1798 => x"a8",
          1799 => x"84",
          1800 => x"74",
          1801 => x"c8",
          1802 => x"3f",
          1803 => x"0a",
          1804 => x"33",
          1805 => x"e2",
          1806 => x"51",
          1807 => x"0a",
          1808 => x"2c",
          1809 => x"7a",
          1810 => x"39",
          1811 => x"34",
          1812 => x"51",
          1813 => x"0a",
          1814 => x"2c",
          1815 => x"75",
          1816 => x"58",
          1817 => x"c8",
          1818 => x"9b",
          1819 => x"80",
          1820 => x"a4",
          1821 => x"ff",
          1822 => x"a8",
          1823 => x"38",
          1824 => x"ff",
          1825 => x"ff",
          1826 => x"76",
          1827 => x"d0",
          1828 => x"34",
          1829 => x"ff",
          1830 => x"7b",
          1831 => x"08",
          1832 => x"38",
          1833 => x"2e",
          1834 => x"70",
          1835 => x"08",
          1836 => x"75",
          1837 => x"fc",
          1838 => x"80",
          1839 => x"7b",
          1840 => x"10",
          1841 => x"41",
          1842 => x"d0",
          1843 => x"83",
          1844 => x"8b",
          1845 => x"34",
          1846 => x"84",
          1847 => x"84",
          1848 => x"b6",
          1849 => x"51",
          1850 => x"08",
          1851 => x"84",
          1852 => x"af",
          1853 => x"05",
          1854 => x"81",
          1855 => x"d1",
          1856 => x"0b",
          1857 => x"d0",
          1858 => x"34",
          1859 => x"a8",
          1860 => x"84",
          1861 => x"ae",
          1862 => x"a0",
          1863 => x"c8",
          1864 => x"3f",
          1865 => x"7c",
          1866 => x"06",
          1867 => x"51",
          1868 => x"d0",
          1869 => x"34",
          1870 => x"0d",
          1871 => x"ff",
          1872 => x"ca",
          1873 => x"59",
          1874 => x"58",
          1875 => x"c8",
          1876 => x"3f",
          1877 => x"70",
          1878 => x"52",
          1879 => x"38",
          1880 => x"ff",
          1881 => x"70",
          1882 => x"a4",
          1883 => x"24",
          1884 => x"52",
          1885 => x"81",
          1886 => x"70",
          1887 => x"51",
          1888 => x"84",
          1889 => x"ac",
          1890 => x"81",
          1891 => x"d0",
          1892 => x"25",
          1893 => x"16",
          1894 => x"d4",
          1895 => x"ac",
          1896 => x"81",
          1897 => x"d0",
          1898 => x"25",
          1899 => x"17",
          1900 => x"52",
          1901 => x"75",
          1902 => x"05",
          1903 => x"43",
          1904 => x"38",
          1905 => x"70",
          1906 => x"2e",
          1907 => x"55",
          1908 => x"2b",
          1909 => x"24",
          1910 => x"81",
          1911 => x"81",
          1912 => x"d0",
          1913 => x"25",
          1914 => x"d0",
          1915 => x"05",
          1916 => x"d0",
          1917 => x"38",
          1918 => x"34",
          1919 => x"81",
          1920 => x"70",
          1921 => x"58",
          1922 => x"38",
          1923 => x"81",
          1924 => x"25",
          1925 => x"52",
          1926 => x"81",
          1927 => x"70",
          1928 => x"57",
          1929 => x"84",
          1930 => x"aa",
          1931 => x"81",
          1932 => x"d0",
          1933 => x"24",
          1934 => x"f1",
          1935 => x"9d",
          1936 => x"84",
          1937 => x"84",
          1938 => x"05",
          1939 => x"cf",
          1940 => x"a8",
          1941 => x"c8",
          1942 => x"51",
          1943 => x"08",
          1944 => x"84",
          1945 => x"a9",
          1946 => x"05",
          1947 => x"81",
          1948 => x"80",
          1949 => x"83",
          1950 => x"85",
          1951 => x"77",
          1952 => x"d4",
          1953 => x"52",
          1954 => x"80",
          1955 => x"98",
          1956 => x"57",
          1957 => x"a8",
          1958 => x"79",
          1959 => x"75",
          1960 => x"39",
          1961 => x"fc",
          1962 => x"76",
          1963 => x"84",
          1964 => x"38",
          1965 => x"f2",
          1966 => x"d4",
          1967 => x"83",
          1968 => x"3f",
          1969 => x"3d",
          1970 => x"74",
          1971 => x"0c",
          1972 => x"80",
          1973 => x"75",
          1974 => x"e4",
          1975 => x"e4",
          1976 => x"75",
          1977 => x"93",
          1978 => x"a8",
          1979 => x"f2",
          1980 => x"88",
          1981 => x"c8",
          1982 => x"3f",
          1983 => x"ff",
          1984 => x"ff",
          1985 => x"79",
          1986 => x"7c",
          1987 => x"80",
          1988 => x"b8",
          1989 => x"51",
          1990 => x"08",
          1991 => x"08",
          1992 => x"52",
          1993 => x"1d",
          1994 => x"33",
          1995 => x"56",
          1996 => x"d4",
          1997 => x"83",
          1998 => x"51",
          1999 => x"08",
          2000 => x"84",
          2001 => x"84",
          2002 => x"55",
          2003 => x"3f",
          2004 => x"34",
          2005 => x"81",
          2006 => x"a9",
          2007 => x"06",
          2008 => x"33",
          2009 => x"f0",
          2010 => x"88",
          2011 => x"c8",
          2012 => x"3f",
          2013 => x"ff",
          2014 => x"ff",
          2015 => x"60",
          2016 => x"51",
          2017 => x"33",
          2018 => x"f1",
          2019 => x"5c",
          2020 => x"e4",
          2021 => x"70",
          2022 => x"08",
          2023 => x"d5",
          2024 => x"ff",
          2025 => x"81",
          2026 => x"93",
          2027 => x"f2",
          2028 => x"fe",
          2029 => x"75",
          2030 => x"d0",
          2031 => x"3f",
          2032 => x"f3",
          2033 => x"80",
          2034 => x"b8",
          2035 => x"53",
          2036 => x"81",
          2037 => x"82",
          2038 => x"3d",
          2039 => x"80",
          2040 => x"3f",
          2041 => x"e4",
          2042 => x"ee",
          2043 => x"a6",
          2044 => x"80",
          2045 => x"e3",
          2046 => x"70",
          2047 => x"81",
          2048 => x"10",
          2049 => x"58",
          2050 => x"76",
          2051 => x"fc",
          2052 => x"80",
          2053 => x"75",
          2054 => x"10",
          2055 => x"40",
          2056 => x"81",
          2057 => x"83",
          2058 => x"81",
          2059 => x"38",
          2060 => x"74",
          2061 => x"d4",
          2062 => x"5b",
          2063 => x"80",
          2064 => x"39",
          2065 => x"f2",
          2066 => x"06",
          2067 => x"54",
          2068 => x"84",
          2069 => x"d4",
          2070 => x"05",
          2071 => x"2e",
          2072 => x"83",
          2073 => x"83",
          2074 => x"e0",
          2075 => x"e7",
          2076 => x"0d",
          2077 => x"05",
          2078 => x"83",
          2079 => x"81",
          2080 => x"38",
          2081 => x"a7",
          2082 => x"70",
          2083 => x"79",
          2084 => x"94",
          2085 => x"83",
          2086 => x"70",
          2087 => x"88",
          2088 => x"56",
          2089 => x"80",
          2090 => x"73",
          2091 => x"26",
          2092 => x"83",
          2093 => x"79",
          2094 => x"e0",
          2095 => x"05",
          2096 => x"38",
          2097 => x"80",
          2098 => x"10",
          2099 => x"29",
          2100 => x"59",
          2101 => x"d8",
          2102 => x"d7",
          2103 => x"92",
          2104 => x"75",
          2105 => x"5b",
          2106 => x"74",
          2107 => x"06",
          2108 => x"06",
          2109 => x"ff",
          2110 => x"57",
          2111 => x"38",
          2112 => x"05",
          2113 => x"83",
          2114 => x"38",
          2115 => x"fe",
          2116 => x"55",
          2117 => x"81",
          2118 => x"a0",
          2119 => x"84",
          2120 => x"84",
          2121 => x"83",
          2122 => x"5b",
          2123 => x"78",
          2124 => x"06",
          2125 => x"18",
          2126 => x"bb",
          2127 => x"80",
          2128 => x"90",
          2129 => x"07",
          2130 => x"7f",
          2131 => x"fd",
          2132 => x"e6",
          2133 => x"ff",
          2134 => x"95",
          2135 => x"a0",
          2136 => x"5f",
          2137 => x"b6",
          2138 => x"b6",
          2139 => x"f8",
          2140 => x"7c",
          2141 => x"5f",
          2142 => x"26",
          2143 => x"7d",
          2144 => x"06",
          2145 => x"7d",
          2146 => x"06",
          2147 => x"5d",
          2148 => x"75",
          2149 => x"83",
          2150 => x"76",
          2151 => x"fb",
          2152 => x"56",
          2153 => x"ee",
          2154 => x"87",
          2155 => x"34",
          2156 => x"75",
          2157 => x"80",
          2158 => x"34",
          2159 => x"34",
          2160 => x"81",
          2161 => x"a0",
          2162 => x"f8",
          2163 => x"06",
          2164 => x"73",
          2165 => x"07",
          2166 => x"87",
          2167 => x"51",
          2168 => x"73",
          2169 => x"72",
          2170 => x"d8",
          2171 => x"87",
          2172 => x"84",
          2173 => x"02",
          2174 => x"05",
          2175 => x"56",
          2176 => x"38",
          2177 => x"33",
          2178 => x"12",
          2179 => x"92",
          2180 => x"29",
          2181 => x"f6",
          2182 => x"81",
          2183 => x"22",
          2184 => x"23",
          2185 => x"81",
          2186 => x"5b",
          2187 => x"ff",
          2188 => x"83",
          2189 => x"06",
          2190 => x"79",
          2191 => x"d8",
          2192 => x"54",
          2193 => x"97",
          2194 => x"13",
          2195 => x"81",
          2196 => x"57",
          2197 => x"73",
          2198 => x"a1",
          2199 => x"b6",
          2200 => x"14",
          2201 => x"34",
          2202 => x"eb",
          2203 => x"56",
          2204 => x"78",
          2205 => x"06",
          2206 => x"38",
          2207 => x"d8",
          2208 => x"75",
          2209 => x"a7",
          2210 => x"81",
          2211 => x"5c",
          2212 => x"84",
          2213 => x"33",
          2214 => x"70",
          2215 => x"05",
          2216 => x"34",
          2217 => x"b6",
          2218 => x"5c",
          2219 => x"80",
          2220 => x"3d",
          2221 => x"83",
          2222 => x"06",
          2223 => x"73",
          2224 => x"2e",
          2225 => x"ff",
          2226 => x"72",
          2227 => x"38",
          2228 => x"d8",
          2229 => x"11",
          2230 => x"fe",
          2231 => x"97",
          2232 => x"56",
          2233 => x"75",
          2234 => x"53",
          2235 => x"0b",
          2236 => x"81",
          2237 => x"d8",
          2238 => x"b6",
          2239 => x"83",
          2240 => x"e0",
          2241 => x"33",
          2242 => x"76",
          2243 => x"51",
          2244 => x"10",
          2245 => x"04",
          2246 => x"27",
          2247 => x"80",
          2248 => x"0d",
          2249 => x"83",
          2250 => x"54",
          2251 => x"12",
          2252 => x"0b",
          2253 => x"04",
          2254 => x"70",
          2255 => x"55",
          2256 => x"de",
          2257 => x"84",
          2258 => x"51",
          2259 => x"72",
          2260 => x"b8",
          2261 => x"f8",
          2262 => x"70",
          2263 => x"55",
          2264 => x"84",
          2265 => x"83",
          2266 => x"d8",
          2267 => x"74",
          2268 => x"f8",
          2269 => x"0c",
          2270 => x"f8",
          2271 => x"b6",
          2272 => x"75",
          2273 => x"70",
          2274 => x"ff",
          2275 => x"70",
          2276 => x"83",
          2277 => x"83",
          2278 => x"71",
          2279 => x"84",
          2280 => x"80",
          2281 => x"80",
          2282 => x"0b",
          2283 => x"04",
          2284 => x"90",
          2285 => x"80",
          2286 => x"0d",
          2287 => x"07",
          2288 => x"39",
          2289 => x"86",
          2290 => x"d7",
          2291 => x"34",
          2292 => x"3d",
          2293 => x"fc",
          2294 => x"90",
          2295 => x"33",
          2296 => x"34",
          2297 => x"81",
          2298 => x"f8",
          2299 => x"90",
          2300 => x"70",
          2301 => x"83",
          2302 => x"07",
          2303 => x"ef",
          2304 => x"06",
          2305 => x"df",
          2306 => x"06",
          2307 => x"90",
          2308 => x"33",
          2309 => x"83",
          2310 => x"f8",
          2311 => x"07",
          2312 => x"a7",
          2313 => x"06",
          2314 => x"90",
          2315 => x"33",
          2316 => x"83",
          2317 => x"f8",
          2318 => x"83",
          2319 => x"f8",
          2320 => x"51",
          2321 => x"39",
          2322 => x"02",
          2323 => x"f8",
          2324 => x"f8",
          2325 => x"41",
          2326 => x"82",
          2327 => x"78",
          2328 => x"b6",
          2329 => x"34",
          2330 => x"f8",
          2331 => x"8f",
          2332 => x"81",
          2333 => x"da",
          2334 => x"82",
          2335 => x"83",
          2336 => x"92",
          2337 => x"57",
          2338 => x"d6",
          2339 => x"52",
          2340 => x"3f",
          2341 => x"84",
          2342 => x"34",
          2343 => x"f8",
          2344 => x"0b",
          2345 => x"b6",
          2346 => x"34",
          2347 => x"0b",
          2348 => x"33",
          2349 => x"b7",
          2350 => x"7c",
          2351 => x"ff",
          2352 => x"e5",
          2353 => x"38",
          2354 => x"22",
          2355 => x"80",
          2356 => x"06",
          2357 => x"78",
          2358 => x"51",
          2359 => x"da",
          2360 => x"7a",
          2361 => x"92",
          2362 => x"3d",
          2363 => x"34",
          2364 => x"0b",
          2365 => x"f8",
          2366 => x"23",
          2367 => x"3f",
          2368 => x"90",
          2369 => x"83",
          2370 => x"78",
          2371 => x"38",
          2372 => x"e3",
          2373 => x"19",
          2374 => x"39",
          2375 => x"a7",
          2376 => x"f8",
          2377 => x"71",
          2378 => x"83",
          2379 => x"71",
          2380 => x"06",
          2381 => x"55",
          2382 => x"38",
          2383 => x"89",
          2384 => x"83",
          2385 => x"38",
          2386 => x"33",
          2387 => x"05",
          2388 => x"33",
          2389 => x"b6",
          2390 => x"f8",
          2391 => x"5a",
          2392 => x"34",
          2393 => x"16",
          2394 => x"a7",
          2395 => x"33",
          2396 => x"22",
          2397 => x"11",
          2398 => x"90",
          2399 => x"18",
          2400 => x"78",
          2401 => x"33",
          2402 => x"53",
          2403 => x"db",
          2404 => x"84",
          2405 => x"80",
          2406 => x"0c",
          2407 => x"97",
          2408 => x"75",
          2409 => x"38",
          2410 => x"80",
          2411 => x"39",
          2412 => x"b6",
          2413 => x"2e",
          2414 => x"53",
          2415 => x"81",
          2416 => x"72",
          2417 => x"a0",
          2418 => x"81",
          2419 => x"d8",
          2420 => x"95",
          2421 => x"51",
          2422 => x"e4",
          2423 => x"ff",
          2424 => x"83",
          2425 => x"55",
          2426 => x"53",
          2427 => x"a0",
          2428 => x"33",
          2429 => x"53",
          2430 => x"83",
          2431 => x"0b",
          2432 => x"51",
          2433 => x"52",
          2434 => x"39",
          2435 => x"33",
          2436 => x"81",
          2437 => x"83",
          2438 => x"38",
          2439 => x"88",
          2440 => x"88",
          2441 => x"f8",
          2442 => x"72",
          2443 => x"e0",
          2444 => x"34",
          2445 => x"33",
          2446 => x"12",
          2447 => x"96",
          2448 => x"71",
          2449 => x"90",
          2450 => x"34",
          2451 => x"06",
          2452 => x"33",
          2453 => x"58",
          2454 => x"b6",
          2455 => x"06",
          2456 => x"38",
          2457 => x"f1",
          2458 => x"95",
          2459 => x"9c",
          2460 => x"8a",
          2461 => x"78",
          2462 => x"db",
          2463 => x"b7",
          2464 => x"f8",
          2465 => x"72",
          2466 => x"e0",
          2467 => x"34",
          2468 => x"33",
          2469 => x"12",
          2470 => x"96",
          2471 => x"71",
          2472 => x"33",
          2473 => x"b6",
          2474 => x"f8",
          2475 => x"72",
          2476 => x"83",
          2477 => x"05",
          2478 => x"06",
          2479 => x"77",
          2480 => x"b8",
          2481 => x"9b",
          2482 => x"83",
          2483 => x"06",
          2484 => x"95",
          2485 => x"9c",
          2486 => x"aa",
          2487 => x"84",
          2488 => x"11",
          2489 => x"78",
          2490 => x"ff",
          2491 => x"1a",
          2492 => x"9c",
          2493 => x"e9",
          2494 => x"84",
          2495 => x"83",
          2496 => x"5e",
          2497 => x"86",
          2498 => x"d8",
          2499 => x"92",
          2500 => x"59",
          2501 => x"83",
          2502 => x"5b",
          2503 => x"b0",
          2504 => x"70",
          2505 => x"83",
          2506 => x"44",
          2507 => x"33",
          2508 => x"1f",
          2509 => x"51",
          2510 => x"95",
          2511 => x"33",
          2512 => x"06",
          2513 => x"12",
          2514 => x"92",
          2515 => x"05",
          2516 => x"ea",
          2517 => x"81",
          2518 => x"06",
          2519 => x"38",
          2520 => x"fc",
          2521 => x"34",
          2522 => x"0b",
          2523 => x"b7",
          2524 => x"0c",
          2525 => x"3d",
          2526 => x"b8",
          2527 => x"b8",
          2528 => x"b8",
          2529 => x"0c",
          2530 => x"3d",
          2531 => x"81",
          2532 => x"33",
          2533 => x"06",
          2534 => x"06",
          2535 => x"80",
          2536 => x"72",
          2537 => x"06",
          2538 => x"5c",
          2539 => x"fe",
          2540 => x"58",
          2541 => x"83",
          2542 => x"7a",
          2543 => x"72",
          2544 => x"b7",
          2545 => x"34",
          2546 => x"33",
          2547 => x"12",
          2548 => x"f8",
          2549 => x"60",
          2550 => x"f8",
          2551 => x"34",
          2552 => x"06",
          2553 => x"33",
          2554 => x"5e",
          2555 => x"97",
          2556 => x"ff",
          2557 => x"ea",
          2558 => x"96",
          2559 => x"f8",
          2560 => x"81",
          2561 => x"ac",
          2562 => x"78",
          2563 => x"2e",
          2564 => x"5f",
          2565 => x"56",
          2566 => x"10",
          2567 => x"08",
          2568 => x"80",
          2569 => x"0b",
          2570 => x"04",
          2571 => x"33",
          2572 => x"33",
          2573 => x"11",
          2574 => x"92",
          2575 => x"70",
          2576 => x"33",
          2577 => x"7f",
          2578 => x"7a",
          2579 => x"7a",
          2580 => x"5c",
          2581 => x"a7",
          2582 => x"33",
          2583 => x"22",
          2584 => x"56",
          2585 => x"83",
          2586 => x"5a",
          2587 => x"b0",
          2588 => x"70",
          2589 => x"83",
          2590 => x"5b",
          2591 => x"33",
          2592 => x"05",
          2593 => x"7a",
          2594 => x"33",
          2595 => x"56",
          2596 => x"70",
          2597 => x"26",
          2598 => x"84",
          2599 => x"72",
          2600 => x"72",
          2601 => x"54",
          2602 => x"80",
          2603 => x"84",
          2604 => x"83",
          2605 => x"5e",
          2606 => x"96",
          2607 => x"71",
          2608 => x"33",
          2609 => x"b6",
          2610 => x"f8",
          2611 => x"72",
          2612 => x"83",
          2613 => x"34",
          2614 => x"5b",
          2615 => x"77",
          2616 => x"82",
          2617 => x"84",
          2618 => x"83",
          2619 => x"e0",
          2620 => x"33",
          2621 => x"56",
          2622 => x"e6",
          2623 => x"9c",
          2624 => x"33",
          2625 => x"34",
          2626 => x"33",
          2627 => x"80",
          2628 => x"42",
          2629 => x"51",
          2630 => x"08",
          2631 => x"e5",
          2632 => x"b7",
          2633 => x"41",
          2634 => x"b8",
          2635 => x"f8",
          2636 => x"1c",
          2637 => x"84",
          2638 => x"5b",
          2639 => x"d8",
          2640 => x"95",
          2641 => x"5b",
          2642 => x"a7",
          2643 => x"33",
          2644 => x"22",
          2645 => x"56",
          2646 => x"f8",
          2647 => x"5e",
          2648 => x"b0",
          2649 => x"70",
          2650 => x"83",
          2651 => x"41",
          2652 => x"33",
          2653 => x"70",
          2654 => x"26",
          2655 => x"58",
          2656 => x"75",
          2657 => x"b7",
          2658 => x"7f",
          2659 => x"dc",
          2660 => x"52",
          2661 => x"84",
          2662 => x"84",
          2663 => x"84",
          2664 => x"84",
          2665 => x"92",
          2666 => x"33",
          2667 => x"33",
          2668 => x"33",
          2669 => x"84",
          2670 => x"ff",
          2671 => x"7c",
          2672 => x"38",
          2673 => x"83",
          2674 => x"53",
          2675 => x"52",
          2676 => x"fe",
          2677 => x"81",
          2678 => x"76",
          2679 => x"38",
          2680 => x"fd",
          2681 => x"84",
          2682 => x"ff",
          2683 => x"38",
          2684 => x"11",
          2685 => x"a5",
          2686 => x"05",
          2687 => x"33",
          2688 => x"83",
          2689 => x"71",
          2690 => x"72",
          2691 => x"83",
          2692 => x"b7",
          2693 => x"e7",
          2694 => x"70",
          2695 => x"5d",
          2696 => x"38",
          2697 => x"39",
          2698 => x"f8",
          2699 => x"57",
          2700 => x"17",
          2701 => x"9c",
          2702 => x"83",
          2703 => x"ff",
          2704 => x"84",
          2705 => x"94",
          2706 => x"33",
          2707 => x"83",
          2708 => x"71",
          2709 => x"72",
          2710 => x"83",
          2711 => x"b7",
          2712 => x"c4",
          2713 => x"99",
          2714 => x"84",
          2715 => x"83",
          2716 => x"86",
          2717 => x"22",
          2718 => x"05",
          2719 => x"e8",
          2720 => x"5a",
          2721 => x"92",
          2722 => x"34",
          2723 => x"5a",
          2724 => x"b8",
          2725 => x"81",
          2726 => x"f6",
          2727 => x"e5",
          2728 => x"38",
          2729 => x"33",
          2730 => x"ff",
          2731 => x"83",
          2732 => x"34",
          2733 => x"57",
          2734 => x"b8",
          2735 => x"61",
          2736 => x"59",
          2737 => x"75",
          2738 => x"f4",
          2739 => x"ed",
          2740 => x"57",
          2741 => x"76",
          2742 => x"53",
          2743 => x"cd",
          2744 => x"84",
          2745 => x"39",
          2746 => x"57",
          2747 => x"b8",
          2748 => x"75",
          2749 => x"51",
          2750 => x"b7",
          2751 => x"b7",
          2752 => x"70",
          2753 => x"ff",
          2754 => x"d7",
          2755 => x"40",
          2756 => x"7e",
          2757 => x"f8",
          2758 => x"18",
          2759 => x"77",
          2760 => x"b6",
          2761 => x"60",
          2762 => x"83",
          2763 => x"b7",
          2764 => x"ef",
          2765 => x"d7",
          2766 => x"94",
          2767 => x"d8",
          2768 => x"95",
          2769 => x"a0",
          2770 => x"40",
          2771 => x"ff",
          2772 => x"59",
          2773 => x"f0",
          2774 => x"7c",
          2775 => x"fe",
          2776 => x"76",
          2777 => x"75",
          2778 => x"06",
          2779 => x"24",
          2780 => x"56",
          2781 => x"16",
          2782 => x"81",
          2783 => x"57",
          2784 => x"75",
          2785 => x"06",
          2786 => x"58",
          2787 => x"b0",
          2788 => x"ff",
          2789 => x"42",
          2790 => x"84",
          2791 => x"33",
          2792 => x"70",
          2793 => x"05",
          2794 => x"34",
          2795 => x"b6",
          2796 => x"40",
          2797 => x"38",
          2798 => x"e0",
          2799 => x"34",
          2800 => x"70",
          2801 => x"b6",
          2802 => x"71",
          2803 => x"78",
          2804 => x"84",
          2805 => x"87",
          2806 => x"33",
          2807 => x"80",
          2808 => x"84",
          2809 => x"79",
          2810 => x"22",
          2811 => x"8b",
          2812 => x"76",
          2813 => x"79",
          2814 => x"ed",
          2815 => x"60",
          2816 => x"06",
          2817 => x"7b",
          2818 => x"76",
          2819 => x"70",
          2820 => x"80",
          2821 => x"b0",
          2822 => x"5d",
          2823 => x"57",
          2824 => x"33",
          2825 => x"71",
          2826 => x"59",
          2827 => x"38",
          2828 => x"7d",
          2829 => x"77",
          2830 => x"84",
          2831 => x"ff",
          2832 => x"92",
          2833 => x"59",
          2834 => x"76",
          2835 => x"05",
          2836 => x"76",
          2837 => x"90",
          2838 => x"a0",
          2839 => x"70",
          2840 => x"76",
          2841 => x"e0",
          2842 => x"05",
          2843 => x"27",
          2844 => x"70",
          2845 => x"39",
          2846 => x"06",
          2847 => x"84",
          2848 => x"f0",
          2849 => x"f2",
          2850 => x"70",
          2851 => x"39",
          2852 => x"b6",
          2853 => x"94",
          2854 => x"92",
          2855 => x"5f",
          2856 => x"33",
          2857 => x"34",
          2858 => x"56",
          2859 => x"81",
          2860 => x"f8",
          2861 => x"33",
          2862 => x"83",
          2863 => x"90",
          2864 => x"75",
          2865 => x"f8",
          2866 => x"56",
          2867 => x"39",
          2868 => x"81",
          2869 => x"f4",
          2870 => x"8f",
          2871 => x"ff",
          2872 => x"9f",
          2873 => x"90",
          2874 => x"33",
          2875 => x"75",
          2876 => x"83",
          2877 => x"c0",
          2878 => x"fe",
          2879 => x"af",
          2880 => x"90",
          2881 => x"33",
          2882 => x"83",
          2883 => x"f8",
          2884 => x"56",
          2885 => x"39",
          2886 => x"82",
          2887 => x"fe",
          2888 => x"f8",
          2889 => x"fd",
          2890 => x"f0",
          2891 => x"fd",
          2892 => x"f0",
          2893 => x"fd",
          2894 => x"df",
          2895 => x"f8",
          2896 => x"90",
          2897 => x"75",
          2898 => x"80",
          2899 => x"81",
          2900 => x"84",
          2901 => x"84",
          2902 => x"84",
          2903 => x"92",
          2904 => x"e8",
          2905 => x"34",
          2906 => x"3d",
          2907 => x"83",
          2908 => x"58",
          2909 => x"b7",
          2910 => x"d8",
          2911 => x"b8",
          2912 => x"08",
          2913 => x"b7",
          2914 => x"0c",
          2915 => x"95",
          2916 => x"33",
          2917 => x"e5",
          2918 => x"02",
          2919 => x"1e",
          2920 => x"ca",
          2921 => x"80",
          2922 => x"f8",
          2923 => x"ff",
          2924 => x"83",
          2925 => x"d0",
          2926 => x"fe",
          2927 => x"f8",
          2928 => x"9f",
          2929 => x"a6",
          2930 => x"84",
          2931 => x"ee",
          2932 => x"ee",
          2933 => x"05",
          2934 => x"58",
          2935 => x"94",
          2936 => x"ff",
          2937 => x"f3",
          2938 => x"84",
          2939 => x"58",
          2940 => x"83",
          2941 => x"70",
          2942 => x"71",
          2943 => x"05",
          2944 => x"7e",
          2945 => x"83",
          2946 => x"5f",
          2947 => x"79",
          2948 => x"57",
          2949 => x"b6",
          2950 => x"98",
          2951 => x"92",
          2952 => x"57",
          2953 => x"84",
          2954 => x"82",
          2955 => x"f8",
          2956 => x"f8",
          2957 => x"76",
          2958 => x"05",
          2959 => x"5c",
          2960 => x"80",
          2961 => x"ff",
          2962 => x"29",
          2963 => x"27",
          2964 => x"57",
          2965 => x"e0",
          2966 => x"34",
          2967 => x"70",
          2968 => x"b6",
          2969 => x"71",
          2970 => x"76",
          2971 => x"33",
          2972 => x"70",
          2973 => x"05",
          2974 => x"34",
          2975 => x"b6",
          2976 => x"41",
          2977 => x"38",
          2978 => x"33",
          2979 => x"34",
          2980 => x"33",
          2981 => x"33",
          2982 => x"76",
          2983 => x"70",
          2984 => x"58",
          2985 => x"79",
          2986 => x"06",
          2987 => x"83",
          2988 => x"34",
          2989 => x"06",
          2990 => x"27",
          2991 => x"f8",
          2992 => x"95",
          2993 => x"ff",
          2994 => x"ef",
          2995 => x"75",
          2996 => x"38",
          2997 => x"06",
          2998 => x"5d",
          2999 => x"f4",
          3000 => x"56",
          3001 => x"39",
          3002 => x"23",
          3003 => x"75",
          3004 => x"77",
          3005 => x"8d",
          3006 => x"34",
          3007 => x"05",
          3008 => x"38",
          3009 => x"83",
          3010 => x"59",
          3011 => x"d3",
          3012 => x"f8",
          3013 => x"83",
          3014 => x"83",
          3015 => x"0b",
          3016 => x"80",
          3017 => x"39",
          3018 => x"b6",
          3019 => x"83",
          3020 => x"3d",
          3021 => x"da",
          3022 => x"38",
          3023 => x"84",
          3024 => x"76",
          3025 => x"0b",
          3026 => x"04",
          3027 => x"5c",
          3028 => x"81",
          3029 => x"58",
          3030 => x"d6",
          3031 => x"e8",
          3032 => x"0c",
          3033 => x"08",
          3034 => x"38",
          3035 => x"70",
          3036 => x"58",
          3037 => x"80",
          3038 => x"83",
          3039 => x"30",
          3040 => x"5d",
          3041 => x"b6",
          3042 => x"f8",
          3043 => x"a7",
          3044 => x"5b",
          3045 => x"83",
          3046 => x"58",
          3047 => x"8c",
          3048 => x"80",
          3049 => x"88",
          3050 => x"75",
          3051 => x"84",
          3052 => x"34",
          3053 => x"55",
          3054 => x"54",
          3055 => x"ff",
          3056 => x"54",
          3057 => x"72",
          3058 => x"83",
          3059 => x"06",
          3060 => x"38",
          3061 => x"f6",
          3062 => x"34",
          3063 => x"5e",
          3064 => x"f6",
          3065 => x"25",
          3066 => x"34",
          3067 => x"81",
          3068 => x"72",
          3069 => x"83",
          3070 => x"53",
          3071 => x"0b",
          3072 => x"f6",
          3073 => x"f6",
          3074 => x"83",
          3075 => x"5c",
          3076 => x"55",
          3077 => x"f6",
          3078 => x"82",
          3079 => x"53",
          3080 => x"f6",
          3081 => x"38",
          3082 => x"ff",
          3083 => x"33",
          3084 => x"74",
          3085 => x"2e",
          3086 => x"33",
          3087 => x"83",
          3088 => x"c0",
          3089 => x"27",
          3090 => x"98",
          3091 => x"81",
          3092 => x"89",
          3093 => x"f6",
          3094 => x"fe",
          3095 => x"8b",
          3096 => x"05",
          3097 => x"08",
          3098 => x"f4",
          3099 => x"5e",
          3100 => x"0b",
          3101 => x"81",
          3102 => x"f6",
          3103 => x"83",
          3104 => x"58",
          3105 => x"96",
          3106 => x"33",
          3107 => x"39",
          3108 => x"2e",
          3109 => x"f4",
          3110 => x"54",
          3111 => x"39",
          3112 => x"81",
          3113 => x"81",
          3114 => x"80",
          3115 => x"38",
          3116 => x"27",
          3117 => x"25",
          3118 => x"81",
          3119 => x"81",
          3120 => x"2b",
          3121 => x"24",
          3122 => x"10",
          3123 => x"83",
          3124 => x"54",
          3125 => x"f6",
          3126 => x"59",
          3127 => x"81",
          3128 => x"59",
          3129 => x"9f",
          3130 => x"54",
          3131 => x"7b",
          3132 => x"76",
          3133 => x"7b",
          3134 => x"38",
          3135 => x"53",
          3136 => x"05",
          3137 => x"83",
          3138 => x"06",
          3139 => x"84",
          3140 => x"f9",
          3141 => x"74",
          3142 => x"52",
          3143 => x"b8",
          3144 => x"76",
          3145 => x"72",
          3146 => x"ac",
          3147 => x"f6",
          3148 => x"0b",
          3149 => x"83",
          3150 => x"f6",
          3151 => x"81",
          3152 => x"fc",
          3153 => x"55",
          3154 => x"81",
          3155 => x"81",
          3156 => x"08",
          3157 => x"08",
          3158 => x"38",
          3159 => x"b8",
          3160 => x"d7",
          3161 => x"34",
          3162 => x"34",
          3163 => x"9e",
          3164 => x"0b",
          3165 => x"08",
          3166 => x"c0",
          3167 => x"42",
          3168 => x"79",
          3169 => x"38",
          3170 => x"38",
          3171 => x"c0",
          3172 => x"81",
          3173 => x"84",
          3174 => x"38",
          3175 => x"ff",
          3176 => x"b6",
          3177 => x"81",
          3178 => x"59",
          3179 => x"c4",
          3180 => x"0b",
          3181 => x"84",
          3182 => x"ff",
          3183 => x"83",
          3184 => x"23",
          3185 => x"53",
          3186 => x"73",
          3187 => x"33",
          3188 => x"53",
          3189 => x"72",
          3190 => x"b7",
          3191 => x"a5",
          3192 => x"54",
          3193 => x"83",
          3194 => x"81",
          3195 => x"c8",
          3196 => x"0d",
          3197 => x"0d",
          3198 => x"f2",
          3199 => x"33",
          3200 => x"51",
          3201 => x"f2",
          3202 => x"15",
          3203 => x"34",
          3204 => x"f0",
          3205 => x"87",
          3206 => x"98",
          3207 => x"38",
          3208 => x"08",
          3209 => x"71",
          3210 => x"98",
          3211 => x"27",
          3212 => x"2e",
          3213 => x"08",
          3214 => x"98",
          3215 => x"08",
          3216 => x"14",
          3217 => x"52",
          3218 => x"ff",
          3219 => x"08",
          3220 => x"52",
          3221 => x"06",
          3222 => x"74",
          3223 => x"38",
          3224 => x"b8",
          3225 => x"0b",
          3226 => x"04",
          3227 => x"a3",
          3228 => x"f2",
          3229 => x"80",
          3230 => x"51",
          3231 => x"72",
          3232 => x"71",
          3233 => x"72",
          3234 => x"52",
          3235 => x"08",
          3236 => x"83",
          3237 => x"81",
          3238 => x"e8",
          3239 => x"f2",
          3240 => x"53",
          3241 => x"c0",
          3242 => x"f6",
          3243 => x"9c",
          3244 => x"38",
          3245 => x"c0",
          3246 => x"73",
          3247 => x"ff",
          3248 => x"9c",
          3249 => x"c0",
          3250 => x"9c",
          3251 => x"81",
          3252 => x"52",
          3253 => x"81",
          3254 => x"a4",
          3255 => x"ff",
          3256 => x"ff",
          3257 => x"c7",
          3258 => x"fe",
          3259 => x"06",
          3260 => x"7b",
          3261 => x"73",
          3262 => x"53",
          3263 => x"72",
          3264 => x"e4",
          3265 => x"84",
          3266 => x"ff",
          3267 => x"02",
          3268 => x"80",
          3269 => x"2b",
          3270 => x"98",
          3271 => x"83",
          3272 => x"84",
          3273 => x"85",
          3274 => x"83",
          3275 => x"80",
          3276 => x"27",
          3277 => x"33",
          3278 => x"71",
          3279 => x"54",
          3280 => x"08",
          3281 => x"83",
          3282 => x"81",
          3283 => x"e8",
          3284 => x"f2",
          3285 => x"53",
          3286 => x"c0",
          3287 => x"f6",
          3288 => x"9c",
          3289 => x"38",
          3290 => x"c0",
          3291 => x"73",
          3292 => x"ff",
          3293 => x"9c",
          3294 => x"c0",
          3295 => x"9c",
          3296 => x"81",
          3297 => x"52",
          3298 => x"81",
          3299 => x"a4",
          3300 => x"ff",
          3301 => x"ff",
          3302 => x"38",
          3303 => x"d5",
          3304 => x"54",
          3305 => x"76",
          3306 => x"04",
          3307 => x"83",
          3308 => x"34",
          3309 => x"56",
          3310 => x"86",
          3311 => x"9c",
          3312 => x"ce",
          3313 => x"08",
          3314 => x"72",
          3315 => x"87",
          3316 => x"74",
          3317 => x"db",
          3318 => x"ff",
          3319 => x"71",
          3320 => x"87",
          3321 => x"05",
          3322 => x"87",
          3323 => x"2e",
          3324 => x"98",
          3325 => x"87",
          3326 => x"87",
          3327 => x"26",
          3328 => x"16",
          3329 => x"80",
          3330 => x"54",
          3331 => x"3d",
          3332 => x"d0",
          3333 => x"0d",
          3334 => x"83",
          3335 => x"83",
          3336 => x"33",
          3337 => x"77",
          3338 => x"98",
          3339 => x"41",
          3340 => x"57",
          3341 => x"72",
          3342 => x"71",
          3343 => x"05",
          3344 => x"2b",
          3345 => x"52",
          3346 => x"9e",
          3347 => x"71",
          3348 => x"05",
          3349 => x"74",
          3350 => x"54",
          3351 => x"08",
          3352 => x"33",
          3353 => x"5c",
          3354 => x"34",
          3355 => x"08",
          3356 => x"80",
          3357 => x"08",
          3358 => x"14",
          3359 => x"33",
          3360 => x"82",
          3361 => x"58",
          3362 => x"13",
          3363 => x"33",
          3364 => x"83",
          3365 => x"85",
          3366 => x"88",
          3367 => x"58",
          3368 => x"34",
          3369 => x"11",
          3370 => x"71",
          3371 => x"72",
          3372 => x"71",
          3373 => x"55",
          3374 => x"87",
          3375 => x"70",
          3376 => x"07",
          3377 => x"5a",
          3378 => x"81",
          3379 => x"17",
          3380 => x"2b",
          3381 => x"33",
          3382 => x"70",
          3383 => x"05",
          3384 => x"5c",
          3385 => x"34",
          3386 => x"08",
          3387 => x"71",
          3388 => x"05",
          3389 => x"2b",
          3390 => x"2a",
          3391 => x"52",
          3392 => x"84",
          3393 => x"33",
          3394 => x"83",
          3395 => x"12",
          3396 => x"07",
          3397 => x"53",
          3398 => x"33",
          3399 => x"82",
          3400 => x"59",
          3401 => x"34",
          3402 => x"33",
          3403 => x"83",
          3404 => x"83",
          3405 => x"88",
          3406 => x"52",
          3407 => x"15",
          3408 => x"0d",
          3409 => x"76",
          3410 => x"86",
          3411 => x"3d",
          3412 => x"b8",
          3413 => x"d0",
          3414 => x"84",
          3415 => x"84",
          3416 => x"81",
          3417 => x"08",
          3418 => x"85",
          3419 => x"76",
          3420 => x"34",
          3421 => x"22",
          3422 => x"83",
          3423 => x"51",
          3424 => x"89",
          3425 => x"10",
          3426 => x"f8",
          3427 => x"81",
          3428 => x"f7",
          3429 => x"51",
          3430 => x"83",
          3431 => x"06",
          3432 => x"84",
          3433 => x"12",
          3434 => x"59",
          3435 => x"75",
          3436 => x"10",
          3437 => x"71",
          3438 => x"06",
          3439 => x"70",
          3440 => x"52",
          3441 => x"2e",
          3442 => x"12",
          3443 => x"07",
          3444 => x"ff",
          3445 => x"56",
          3446 => x"33",
          3447 => x"70",
          3448 => x"56",
          3449 => x"81",
          3450 => x"8d",
          3451 => x"85",
          3452 => x"74",
          3453 => x"82",
          3454 => x"5c",
          3455 => x"81",
          3456 => x"76",
          3457 => x"34",
          3458 => x"08",
          3459 => x"71",
          3460 => x"ff",
          3461 => x"ff",
          3462 => x"57",
          3463 => x"72",
          3464 => x"34",
          3465 => x"74",
          3466 => x"d4",
          3467 => x"12",
          3468 => x"07",
          3469 => x"75",
          3470 => x"84",
          3471 => x"05",
          3472 => x"88",
          3473 => x"58",
          3474 => x"15",
          3475 => x"84",
          3476 => x"2b",
          3477 => x"5a",
          3478 => x"72",
          3479 => x"70",
          3480 => x"85",
          3481 => x"88",
          3482 => x"15",
          3483 => x"d4",
          3484 => x"b8",
          3485 => x"14",
          3486 => x"71",
          3487 => x"33",
          3488 => x"70",
          3489 => x"52",
          3490 => x"34",
          3491 => x"11",
          3492 => x"71",
          3493 => x"33",
          3494 => x"70",
          3495 => x"5b",
          3496 => x"87",
          3497 => x"70",
          3498 => x"07",
          3499 => x"59",
          3500 => x"81",
          3501 => x"84",
          3502 => x"0d",
          3503 => x"76",
          3504 => x"8a",
          3505 => x"3d",
          3506 => x"84",
          3507 => x"89",
          3508 => x"84",
          3509 => x"b8",
          3510 => x"52",
          3511 => x"3f",
          3512 => x"34",
          3513 => x"d4",
          3514 => x"0b",
          3515 => x"56",
          3516 => x"17",
          3517 => x"d0",
          3518 => x"70",
          3519 => x"58",
          3520 => x"73",
          3521 => x"70",
          3522 => x"05",
          3523 => x"34",
          3524 => x"77",
          3525 => x"39",
          3526 => x"80",
          3527 => x"41",
          3528 => x"80",
          3529 => x"88",
          3530 => x"8f",
          3531 => x"05",
          3532 => x"73",
          3533 => x"83",
          3534 => x"83",
          3535 => x"33",
          3536 => x"70",
          3537 => x"10",
          3538 => x"70",
          3539 => x"07",
          3540 => x"42",
          3541 => x"5c",
          3542 => x"7a",
          3543 => x"83",
          3544 => x"10",
          3545 => x"33",
          3546 => x"53",
          3547 => x"24",
          3548 => x"f6",
          3549 => x"87",
          3550 => x"38",
          3551 => x"be",
          3552 => x"92",
          3553 => x"12",
          3554 => x"07",
          3555 => x"71",
          3556 => x"43",
          3557 => x"60",
          3558 => x"11",
          3559 => x"71",
          3560 => x"33",
          3561 => x"83",
          3562 => x"85",
          3563 => x"88",
          3564 => x"58",
          3565 => x"34",
          3566 => x"08",
          3567 => x"33",
          3568 => x"74",
          3569 => x"71",
          3570 => x"42",
          3571 => x"86",
          3572 => x"b8",
          3573 => x"33",
          3574 => x"06",
          3575 => x"76",
          3576 => x"b8",
          3577 => x"83",
          3578 => x"2b",
          3579 => x"33",
          3580 => x"41",
          3581 => x"79",
          3582 => x"b8",
          3583 => x"12",
          3584 => x"07",
          3585 => x"33",
          3586 => x"41",
          3587 => x"79",
          3588 => x"84",
          3589 => x"33",
          3590 => x"66",
          3591 => x"52",
          3592 => x"fe",
          3593 => x"1e",
          3594 => x"83",
          3595 => x"62",
          3596 => x"84",
          3597 => x"84",
          3598 => x"a0",
          3599 => x"80",
          3600 => x"51",
          3601 => x"08",
          3602 => x"1f",
          3603 => x"84",
          3604 => x"84",
          3605 => x"34",
          3606 => x"d4",
          3607 => x"fe",
          3608 => x"06",
          3609 => x"78",
          3610 => x"84",
          3611 => x"84",
          3612 => x"56",
          3613 => x"15",
          3614 => x"fa",
          3615 => x"38",
          3616 => x"38",
          3617 => x"e4",
          3618 => x"0d",
          3619 => x"71",
          3620 => x"05",
          3621 => x"2b",
          3622 => x"2a",
          3623 => x"34",
          3624 => x"d4",
          3625 => x"75",
          3626 => x"84",
          3627 => x"81",
          3628 => x"83",
          3629 => x"64",
          3630 => x"4a",
          3631 => x"63",
          3632 => x"41",
          3633 => x"d4",
          3634 => x"81",
          3635 => x"05",
          3636 => x"54",
          3637 => x"83",
          3638 => x"39",
          3639 => x"70",
          3640 => x"83",
          3641 => x"10",
          3642 => x"33",
          3643 => x"53",
          3644 => x"73",
          3645 => x"39",
          3646 => x"7a",
          3647 => x"ff",
          3648 => x"38",
          3649 => x"84",
          3650 => x"b8",
          3651 => x"52",
          3652 => x"3f",
          3653 => x"34",
          3654 => x"d4",
          3655 => x"0b",
          3656 => x"58",
          3657 => x"19",
          3658 => x"d0",
          3659 => x"70",
          3660 => x"58",
          3661 => x"34",
          3662 => x"d0",
          3663 => x"d4",
          3664 => x"61",
          3665 => x"34",
          3666 => x"de",
          3667 => x"61",
          3668 => x"39",
          3669 => x"51",
          3670 => x"b8",
          3671 => x"1e",
          3672 => x"8b",
          3673 => x"86",
          3674 => x"2b",
          3675 => x"14",
          3676 => x"07",
          3677 => x"5b",
          3678 => x"64",
          3679 => x"34",
          3680 => x"11",
          3681 => x"71",
          3682 => x"33",
          3683 => x"70",
          3684 => x"59",
          3685 => x"7a",
          3686 => x"08",
          3687 => x"88",
          3688 => x"88",
          3689 => x"34",
          3690 => x"08",
          3691 => x"33",
          3692 => x"74",
          3693 => x"88",
          3694 => x"5e",
          3695 => x"34",
          3696 => x"08",
          3697 => x"71",
          3698 => x"05",
          3699 => x"88",
          3700 => x"40",
          3701 => x"18",
          3702 => x"d4",
          3703 => x"12",
          3704 => x"62",
          3705 => x"5d",
          3706 => x"ef",
          3707 => x"05",
          3708 => x"fc",
          3709 => x"b8",
          3710 => x"d0",
          3711 => x"84",
          3712 => x"84",
          3713 => x"81",
          3714 => x"08",
          3715 => x"85",
          3716 => x"7f",
          3717 => x"34",
          3718 => x"22",
          3719 => x"83",
          3720 => x"43",
          3721 => x"89",
          3722 => x"10",
          3723 => x"f8",
          3724 => x"81",
          3725 => x"bd",
          3726 => x"19",
          3727 => x"71",
          3728 => x"33",
          3729 => x"70",
          3730 => x"55",
          3731 => x"85",
          3732 => x"1e",
          3733 => x"8b",
          3734 => x"86",
          3735 => x"2b",
          3736 => x"48",
          3737 => x"05",
          3738 => x"b8",
          3739 => x"33",
          3740 => x"06",
          3741 => x"75",
          3742 => x"b8",
          3743 => x"12",
          3744 => x"07",
          3745 => x"71",
          3746 => x"ff",
          3747 => x"48",
          3748 => x"41",
          3749 => x"34",
          3750 => x"33",
          3751 => x"83",
          3752 => x"12",
          3753 => x"ff",
          3754 => x"5e",
          3755 => x"76",
          3756 => x"ff",
          3757 => x"33",
          3758 => x"83",
          3759 => x"85",
          3760 => x"88",
          3761 => x"78",
          3762 => x"84",
          3763 => x"33",
          3764 => x"83",
          3765 => x"87",
          3766 => x"88",
          3767 => x"55",
          3768 => x"60",
          3769 => x"18",
          3770 => x"2b",
          3771 => x"2a",
          3772 => x"78",
          3773 => x"70",
          3774 => x"8b",
          3775 => x"70",
          3776 => x"07",
          3777 => x"77",
          3778 => x"5f",
          3779 => x"17",
          3780 => x"d4",
          3781 => x"33",
          3782 => x"74",
          3783 => x"88",
          3784 => x"88",
          3785 => x"5d",
          3786 => x"34",
          3787 => x"11",
          3788 => x"71",
          3789 => x"33",
          3790 => x"83",
          3791 => x"85",
          3792 => x"88",
          3793 => x"59",
          3794 => x"1d",
          3795 => x"d4",
          3796 => x"12",
          3797 => x"07",
          3798 => x"33",
          3799 => x"5f",
          3800 => x"77",
          3801 => x"84",
          3802 => x"12",
          3803 => x"ff",
          3804 => x"59",
          3805 => x"84",
          3806 => x"33",
          3807 => x"83",
          3808 => x"15",
          3809 => x"2a",
          3810 => x"55",
          3811 => x"84",
          3812 => x"81",
          3813 => x"2b",
          3814 => x"15",
          3815 => x"2a",
          3816 => x"55",
          3817 => x"34",
          3818 => x"11",
          3819 => x"07",
          3820 => x"42",
          3821 => x"51",
          3822 => x"08",
          3823 => x"70",
          3824 => x"f1",
          3825 => x"33",
          3826 => x"79",
          3827 => x"71",
          3828 => x"48",
          3829 => x"05",
          3830 => x"b8",
          3831 => x"85",
          3832 => x"2b",
          3833 => x"15",
          3834 => x"2a",
          3835 => x"56",
          3836 => x"87",
          3837 => x"70",
          3838 => x"07",
          3839 => x"5c",
          3840 => x"81",
          3841 => x"1f",
          3842 => x"2b",
          3843 => x"33",
          3844 => x"70",
          3845 => x"05",
          3846 => x"58",
          3847 => x"34",
          3848 => x"08",
          3849 => x"71",
          3850 => x"05",
          3851 => x"2b",
          3852 => x"2a",
          3853 => x"5b",
          3854 => x"77",
          3855 => x"39",
          3856 => x"84",
          3857 => x"08",
          3858 => x"52",
          3859 => x"cf",
          3860 => x"5b",
          3861 => x"e9",
          3862 => x"84",
          3863 => x"2e",
          3864 => x"73",
          3865 => x"04",
          3866 => x"e4",
          3867 => x"2e",
          3868 => x"b8",
          3869 => x"73",
          3870 => x"04",
          3871 => x"0c",
          3872 => x"82",
          3873 => x"f4",
          3874 => x"d4",
          3875 => x"81",
          3876 => x"76",
          3877 => x"34",
          3878 => x"17",
          3879 => x"b8",
          3880 => x"05",
          3881 => x"ff",
          3882 => x"56",
          3883 => x"34",
          3884 => x"10",
          3885 => x"55",
          3886 => x"83",
          3887 => x"fe",
          3888 => x"0d",
          3889 => x"70",
          3890 => x"11",
          3891 => x"83",
          3892 => x"93",
          3893 => x"26",
          3894 => x"84",
          3895 => x"72",
          3896 => x"34",
          3897 => x"84",
          3898 => x"f7",
          3899 => x"05",
          3900 => x"81",
          3901 => x"b8",
          3902 => x"54",
          3903 => x"85",
          3904 => x"53",
          3905 => x"84",
          3906 => x"74",
          3907 => x"8c",
          3908 => x"26",
          3909 => x"54",
          3910 => x"73",
          3911 => x"3d",
          3912 => x"70",
          3913 => x"78",
          3914 => x"3d",
          3915 => x"af",
          3916 => x"54",
          3917 => x"e0",
          3918 => x"83",
          3919 => x"0b",
          3920 => x"75",
          3921 => x"b8",
          3922 => x"80",
          3923 => x"08",
          3924 => x"d6",
          3925 => x"73",
          3926 => x"55",
          3927 => x"0d",
          3928 => x"81",
          3929 => x"26",
          3930 => x"0d",
          3931 => x"02",
          3932 => x"55",
          3933 => x"84",
          3934 => x"06",
          3935 => x"0b",
          3936 => x"70",
          3937 => x"ad",
          3938 => x"53",
          3939 => x"0d",
          3940 => x"84",
          3941 => x"81",
          3942 => x"e4",
          3943 => x"2b",
          3944 => x"70",
          3945 => x"81",
          3946 => x"38",
          3947 => x"ea",
          3948 => x"70",
          3949 => x"92",
          3950 => x"54",
          3951 => x"08",
          3952 => x"90",
          3953 => x"0b",
          3954 => x"74",
          3955 => x"77",
          3956 => x"38",
          3957 => x"51",
          3958 => x"80",
          3959 => x"b8",
          3960 => x"54",
          3961 => x"53",
          3962 => x"3f",
          3963 => x"2e",
          3964 => x"e4",
          3965 => x"70",
          3966 => x"84",
          3967 => x"74",
          3968 => x"33",
          3969 => x"ff",
          3970 => x"79",
          3971 => x"3f",
          3972 => x"2e",
          3973 => x"18",
          3974 => x"06",
          3975 => x"80",
          3976 => x"05",
          3977 => x"38",
          3978 => x"ff",
          3979 => x"d2",
          3980 => x"34",
          3981 => x"c1",
          3982 => x"84",
          3983 => x"9d",
          3984 => x"19",
          3985 => x"34",
          3986 => x"19",
          3987 => x"a1",
          3988 => x"84",
          3989 => x"7a",
          3990 => x"5b",
          3991 => x"2a",
          3992 => x"90",
          3993 => x"7a",
          3994 => x"34",
          3995 => x"1a",
          3996 => x"52",
          3997 => x"76",
          3998 => x"81",
          3999 => x"b8",
          4000 => x"fd",
          4001 => x"70",
          4002 => x"88",
          4003 => x"38",
          4004 => x"8f",
          4005 => x"58",
          4006 => x"82",
          4007 => x"09",
          4008 => x"16",
          4009 => x"5a",
          4010 => x"2e",
          4011 => x"7b",
          4012 => x"81",
          4013 => x"17",
          4014 => x"e4",
          4015 => x"81",
          4016 => x"9a",
          4017 => x"11",
          4018 => x"1b",
          4019 => x"17",
          4020 => x"83",
          4021 => x"7d",
          4022 => x"81",
          4023 => x"17",
          4024 => x"e4",
          4025 => x"81",
          4026 => x"ca",
          4027 => x"11",
          4028 => x"81",
          4029 => x"59",
          4030 => x"ff",
          4031 => x"0d",
          4032 => x"05",
          4033 => x"38",
          4034 => x"5d",
          4035 => x"81",
          4036 => x"17",
          4037 => x"3f",
          4038 => x"38",
          4039 => x"0c",
          4040 => x"fe",
          4041 => x"33",
          4042 => x"b8",
          4043 => x"04",
          4044 => x"b8",
          4045 => x"05",
          4046 => x"38",
          4047 => x"5e",
          4048 => x"82",
          4049 => x"17",
          4050 => x"3f",
          4051 => x"38",
          4052 => x"0c",
          4053 => x"83",
          4054 => x"11",
          4055 => x"71",
          4056 => x"72",
          4057 => x"ff",
          4058 => x"e4",
          4059 => x"8f",
          4060 => x"08",
          4061 => x"33",
          4062 => x"84",
          4063 => x"06",
          4064 => x"83",
          4065 => x"08",
          4066 => x"7d",
          4067 => x"82",
          4068 => x"81",
          4069 => x"17",
          4070 => x"52",
          4071 => x"7a",
          4072 => x"17",
          4073 => x"18",
          4074 => x"b8",
          4075 => x"82",
          4076 => x"18",
          4077 => x"31",
          4078 => x"38",
          4079 => x"81",
          4080 => x"fb",
          4081 => x"53",
          4082 => x"52",
          4083 => x"b8",
          4084 => x"fd",
          4085 => x"18",
          4086 => x"31",
          4087 => x"a0",
          4088 => x"17",
          4089 => x"06",
          4090 => x"08",
          4091 => x"81",
          4092 => x"5a",
          4093 => x"08",
          4094 => x"33",
          4095 => x"84",
          4096 => x"06",
          4097 => x"83",
          4098 => x"08",
          4099 => x"74",
          4100 => x"82",
          4101 => x"81",
          4102 => x"17",
          4103 => x"52",
          4104 => x"7c",
          4105 => x"17",
          4106 => x"52",
          4107 => x"fa",
          4108 => x"38",
          4109 => x"62",
          4110 => x"76",
          4111 => x"27",
          4112 => x"2e",
          4113 => x"38",
          4114 => x"84",
          4115 => x"75",
          4116 => x"80",
          4117 => x"78",
          4118 => x"7c",
          4119 => x"06",
          4120 => x"b8",
          4121 => x"87",
          4122 => x"85",
          4123 => x"1a",
          4124 => x"75",
          4125 => x"83",
          4126 => x"1f",
          4127 => x"1f",
          4128 => x"84",
          4129 => x"74",
          4130 => x"38",
          4131 => x"58",
          4132 => x"76",
          4133 => x"33",
          4134 => x"81",
          4135 => x"53",
          4136 => x"f1",
          4137 => x"2e",
          4138 => x"b4",
          4139 => x"38",
          4140 => x"05",
          4141 => x"2b",
          4142 => x"07",
          4143 => x"7d",
          4144 => x"7d",
          4145 => x"7d",
          4146 => x"81",
          4147 => x"75",
          4148 => x"1b",
          4149 => x"5a",
          4150 => x"83",
          4151 => x"7d",
          4152 => x"81",
          4153 => x"19",
          4154 => x"e4",
          4155 => x"81",
          4156 => x"7b",
          4157 => x"19",
          4158 => x"5f",
          4159 => x"8f",
          4160 => x"77",
          4161 => x"74",
          4162 => x"7d",
          4163 => x"80",
          4164 => x"76",
          4165 => x"53",
          4166 => x"52",
          4167 => x"b8",
          4168 => x"80",
          4169 => x"1a",
          4170 => x"08",
          4171 => x"08",
          4172 => x"8b",
          4173 => x"2e",
          4174 => x"76",
          4175 => x"3f",
          4176 => x"38",
          4177 => x"0c",
          4178 => x"06",
          4179 => x"56",
          4180 => x"33",
          4181 => x"56",
          4182 => x"1a",
          4183 => x"53",
          4184 => x"52",
          4185 => x"b8",
          4186 => x"fc",
          4187 => x"1a",
          4188 => x"08",
          4189 => x"08",
          4190 => x"fb",
          4191 => x"82",
          4192 => x"81",
          4193 => x"19",
          4194 => x"fb",
          4195 => x"19",
          4196 => x"ee",
          4197 => x"08",
          4198 => x"38",
          4199 => x"b4",
          4200 => x"a0",
          4201 => x"40",
          4202 => x"38",
          4203 => x"09",
          4204 => x"7d",
          4205 => x"51",
          4206 => x"39",
          4207 => x"53",
          4208 => x"3f",
          4209 => x"2e",
          4210 => x"b8",
          4211 => x"08",
          4212 => x"08",
          4213 => x"5e",
          4214 => x"19",
          4215 => x"06",
          4216 => x"53",
          4217 => x"86",
          4218 => x"54",
          4219 => x"33",
          4220 => x"8b",
          4221 => x"7a",
          4222 => x"5f",
          4223 => x"2a",
          4224 => x"39",
          4225 => x"82",
          4226 => x"11",
          4227 => x"0a",
          4228 => x"58",
          4229 => x"88",
          4230 => x"90",
          4231 => x"98",
          4232 => x"cf",
          4233 => x"08",
          4234 => x"90",
          4235 => x"f4",
          4236 => x"ec",
          4237 => x"73",
          4238 => x"2e",
          4239 => x"56",
          4240 => x"82",
          4241 => x"75",
          4242 => x"b8",
          4243 => x"80",
          4244 => x"b1",
          4245 => x"30",
          4246 => x"07",
          4247 => x"38",
          4248 => x"b5",
          4249 => x"0c",
          4250 => x"91",
          4251 => x"39",
          4252 => x"81",
          4253 => x"db",
          4254 => x"b8",
          4255 => x"19",
          4256 => x"38",
          4257 => x"56",
          4258 => x"82",
          4259 => x"3f",
          4260 => x"2e",
          4261 => x"09",
          4262 => x"70",
          4263 => x"51",
          4264 => x"84",
          4265 => x"90",
          4266 => x"a3",
          4267 => x"9b",
          4268 => x"39",
          4269 => x"53",
          4270 => x"84",
          4271 => x"30",
          4272 => x"25",
          4273 => x"74",
          4274 => x"9c",
          4275 => x"56",
          4276 => x"15",
          4277 => x"07",
          4278 => x"74",
          4279 => x"04",
          4280 => x"3d",
          4281 => x"fe",
          4282 => x"38",
          4283 => x"8b",
          4284 => x"a7",
          4285 => x"e4",
          4286 => x"74",
          4287 => x"ff",
          4288 => x"71",
          4289 => x"0a",
          4290 => x"53",
          4291 => x"0c",
          4292 => x"38",
          4293 => x"cc",
          4294 => x"88",
          4295 => x"a9",
          4296 => x"74",
          4297 => x"82",
          4298 => x"89",
          4299 => x"ff",
          4300 => x"80",
          4301 => x"3d",
          4302 => x"0c",
          4303 => x"55",
          4304 => x"17",
          4305 => x"76",
          4306 => x"fe",
          4307 => x"75",
          4308 => x"76",
          4309 => x"53",
          4310 => x"74",
          4311 => x"b8",
          4312 => x"ff",
          4313 => x"e4",
          4314 => x"08",
          4315 => x"ff",
          4316 => x"76",
          4317 => x"0b",
          4318 => x"04",
          4319 => x"12",
          4320 => x"80",
          4321 => x"98",
          4322 => x"56",
          4323 => x"ff",
          4324 => x"94",
          4325 => x"79",
          4326 => x"74",
          4327 => x"18",
          4328 => x"b8",
          4329 => x"84",
          4330 => x"77",
          4331 => x"05",
          4332 => x"38",
          4333 => x"84",
          4334 => x"0b",
          4335 => x"81",
          4336 => x"c6",
          4337 => x"08",
          4338 => x"81",
          4339 => x"51",
          4340 => x"5d",
          4341 => x"2e",
          4342 => x"e4",
          4343 => x"56",
          4344 => x"86",
          4345 => x"33",
          4346 => x"18",
          4347 => x"80",
          4348 => x"19",
          4349 => x"05",
          4350 => x"19",
          4351 => x"76",
          4352 => x"55",
          4353 => x"22",
          4354 => x"81",
          4355 => x"19",
          4356 => x"e4",
          4357 => x"dd",
          4358 => x"84",
          4359 => x"75",
          4360 => x"70",
          4361 => x"86",
          4362 => x"38",
          4363 => x"b4",
          4364 => x"74",
          4365 => x"82",
          4366 => x"81",
          4367 => x"19",
          4368 => x"52",
          4369 => x"fe",
          4370 => x"83",
          4371 => x"09",
          4372 => x"0c",
          4373 => x"5e",
          4374 => x"85",
          4375 => x"b0",
          4376 => x"fc",
          4377 => x"0c",
          4378 => x"64",
          4379 => x"5b",
          4380 => x"5e",
          4381 => x"b8",
          4382 => x"19",
          4383 => x"19",
          4384 => x"09",
          4385 => x"75",
          4386 => x"51",
          4387 => x"80",
          4388 => x"79",
          4389 => x"90",
          4390 => x"58",
          4391 => x"18",
          4392 => x"5b",
          4393 => x"e5",
          4394 => x"30",
          4395 => x"54",
          4396 => x"74",
          4397 => x"2e",
          4398 => x"86",
          4399 => x"51",
          4400 => x"5b",
          4401 => x"98",
          4402 => x"7a",
          4403 => x"04",
          4404 => x"52",
          4405 => x"81",
          4406 => x"09",
          4407 => x"e4",
          4408 => x"a8",
          4409 => x"58",
          4410 => x"b5",
          4411 => x"2e",
          4412 => x"54",
          4413 => x"53",
          4414 => x"de",
          4415 => x"8f",
          4416 => x"76",
          4417 => x"2e",
          4418 => x"bf",
          4419 => x"05",
          4420 => x"ab",
          4421 => x"cc",
          4422 => x"81",
          4423 => x"5b",
          4424 => x"b8",
          4425 => x"5b",
          4426 => x"7d",
          4427 => x"8c",
          4428 => x"33",
          4429 => x"75",
          4430 => x"bf",
          4431 => x"81",
          4432 => x"33",
          4433 => x"71",
          4434 => x"80",
          4435 => x"26",
          4436 => x"76",
          4437 => x"5a",
          4438 => x"38",
          4439 => x"59",
          4440 => x"81",
          4441 => x"61",
          4442 => x"70",
          4443 => x"39",
          4444 => x"81",
          4445 => x"38",
          4446 => x"75",
          4447 => x"05",
          4448 => x"ff",
          4449 => x"e4",
          4450 => x"ff",
          4451 => x"e4",
          4452 => x"0d",
          4453 => x"7b",
          4454 => x"08",
          4455 => x"38",
          4456 => x"ac",
          4457 => x"08",
          4458 => x"2e",
          4459 => x"58",
          4460 => x"81",
          4461 => x"1b",
          4462 => x"3f",
          4463 => x"38",
          4464 => x"0c",
          4465 => x"1c",
          4466 => x"2e",
          4467 => x"06",
          4468 => x"86",
          4469 => x"f2",
          4470 => x"75",
          4471 => x"e2",
          4472 => x"7c",
          4473 => x"57",
          4474 => x"05",
          4475 => x"76",
          4476 => x"59",
          4477 => x"2e",
          4478 => x"06",
          4479 => x"1d",
          4480 => x"33",
          4481 => x"71",
          4482 => x"76",
          4483 => x"2e",
          4484 => x"ac",
          4485 => x"c8",
          4486 => x"b8",
          4487 => x"79",
          4488 => x"04",
          4489 => x"52",
          4490 => x"81",
          4491 => x"09",
          4492 => x"e4",
          4493 => x"a8",
          4494 => x"58",
          4495 => x"ea",
          4496 => x"2e",
          4497 => x"54",
          4498 => x"53",
          4499 => x"b6",
          4500 => x"5a",
          4501 => x"86",
          4502 => x"f2",
          4503 => x"79",
          4504 => x"77",
          4505 => x"7f",
          4506 => x"7d",
          4507 => x"5d",
          4508 => x"84",
          4509 => x"08",
          4510 => x"39",
          4511 => x"ff",
          4512 => x"a2",
          4513 => x"2e",
          4514 => x"08",
          4515 => x"88",
          4516 => x"b3",
          4517 => x"29",
          4518 => x"56",
          4519 => x"81",
          4520 => x"07",
          4521 => x"ed",
          4522 => x"38",
          4523 => x"b8",
          4524 => x"22",
          4525 => x"a0",
          4526 => x"2e",
          4527 => x"56",
          4528 => x"b0",
          4529 => x"06",
          4530 => x"74",
          4531 => x"05",
          4532 => x"38",
          4533 => x"5a",
          4534 => x"e4",
          4535 => x"ff",
          4536 => x"55",
          4537 => x"70",
          4538 => x"06",
          4539 => x"85",
          4540 => x"22",
          4541 => x"38",
          4542 => x"51",
          4543 => x"a0",
          4544 => x"58",
          4545 => x"77",
          4546 => x"55",
          4547 => x"33",
          4548 => x"2e",
          4549 => x"1f",
          4550 => x"8c",
          4551 => x"61",
          4552 => x"59",
          4553 => x"ff",
          4554 => x"27",
          4555 => x"57",
          4556 => x"1a",
          4557 => x"77",
          4558 => x"ff",
          4559 => x"44",
          4560 => x"38",
          4561 => x"18",
          4562 => x"22",
          4563 => x"05",
          4564 => x"07",
          4565 => x"38",
          4566 => x"16",
          4567 => x"56",
          4568 => x"fe",
          4569 => x"78",
          4570 => x"a0",
          4571 => x"78",
          4572 => x"33",
          4573 => x"06",
          4574 => x"77",
          4575 => x"05",
          4576 => x"59",
          4577 => x"87",
          4578 => x"84",
          4579 => x"5b",
          4580 => x"87",
          4581 => x"38",
          4582 => x"e4",
          4583 => x"d6",
          4584 => x"1f",
          4585 => x"db",
          4586 => x"81",
          4587 => x"90",
          4588 => x"8a",
          4589 => x"5b",
          4590 => x"84",
          4591 => x"08",
          4592 => x"b8",
          4593 => x"80",
          4594 => x"f3",
          4595 => x"2e",
          4596 => x"54",
          4597 => x"33",
          4598 => x"08",
          4599 => x"57",
          4600 => x"bc",
          4601 => x"42",
          4602 => x"74",
          4603 => x"5f",
          4604 => x"19",
          4605 => x"81",
          4606 => x"b8",
          4607 => x"80",
          4608 => x"84",
          4609 => x"81",
          4610 => x"f3",
          4611 => x"08",
          4612 => x"78",
          4613 => x"54",
          4614 => x"33",
          4615 => x"08",
          4616 => x"56",
          4617 => x"80",
          4618 => x"57",
          4619 => x"34",
          4620 => x"0b",
          4621 => x"75",
          4622 => x"81",
          4623 => x"ef",
          4624 => x"98",
          4625 => x"81",
          4626 => x"84",
          4627 => x"81",
          4628 => x"57",
          4629 => x"59",
          4630 => x"84",
          4631 => x"08",
          4632 => x"39",
          4633 => x"52",
          4634 => x"84",
          4635 => x"06",
          4636 => x"83",
          4637 => x"08",
          4638 => x"8b",
          4639 => x"2e",
          4640 => x"57",
          4641 => x"1f",
          4642 => x"e9",
          4643 => x"84",
          4644 => x"84",
          4645 => x"74",
          4646 => x"78",
          4647 => x"05",
          4648 => x"56",
          4649 => x"06",
          4650 => x"57",
          4651 => x"b2",
          4652 => x"2e",
          4653 => x"54",
          4654 => x"33",
          4655 => x"08",
          4656 => x"56",
          4657 => x"fe",
          4658 => x"08",
          4659 => x"60",
          4660 => x"34",
          4661 => x"34",
          4662 => x"f3",
          4663 => x"83",
          4664 => x"1f",
          4665 => x"83",
          4666 => x"76",
          4667 => x"88",
          4668 => x"38",
          4669 => x"8c",
          4670 => x"ff",
          4671 => x"70",
          4672 => x"a6",
          4673 => x"1d",
          4674 => x"3f",
          4675 => x"e4",
          4676 => x"40",
          4677 => x"81",
          4678 => x"70",
          4679 => x"96",
          4680 => x"fc",
          4681 => x"1d",
          4682 => x"31",
          4683 => x"a0",
          4684 => x"1c",
          4685 => x"06",
          4686 => x"08",
          4687 => x"81",
          4688 => x"56",
          4689 => x"70",
          4690 => x"2e",
          4691 => x"ff",
          4692 => x"2e",
          4693 => x"80",
          4694 => x"54",
          4695 => x"1c",
          4696 => x"e4",
          4697 => x"38",
          4698 => x"b4",
          4699 => x"74",
          4700 => x"1c",
          4701 => x"84",
          4702 => x"75",
          4703 => x"fa",
          4704 => x"57",
          4705 => x"75",
          4706 => x"39",
          4707 => x"08",
          4708 => x"51",
          4709 => x"54",
          4710 => x"53",
          4711 => x"96",
          4712 => x"7f",
          4713 => x"0b",
          4714 => x"2e",
          4715 => x"2e",
          4716 => x"8c",
          4717 => x"5c",
          4718 => x"54",
          4719 => x"55",
          4720 => x"80",
          4721 => x"5a",
          4722 => x"73",
          4723 => x"58",
          4724 => x"70",
          4725 => x"5c",
          4726 => x"0b",
          4727 => x"59",
          4728 => x"33",
          4729 => x"2e",
          4730 => x"38",
          4731 => x"07",
          4732 => x"26",
          4733 => x"ae",
          4734 => x"18",
          4735 => x"34",
          4736 => x"ba",
          4737 => x"0b",
          4738 => x"72",
          4739 => x"0b",
          4740 => x"94",
          4741 => x"9c",
          4742 => x"73",
          4743 => x"1c",
          4744 => x"34",
          4745 => x"33",
          4746 => x"88",
          4747 => x"07",
          4748 => x"0c",
          4749 => x"71",
          4750 => x"5a",
          4751 => x"99",
          4752 => x"2b",
          4753 => x"8f",
          4754 => x"c0",
          4755 => x"7a",
          4756 => x"7a",
          4757 => x"89",
          4758 => x"ff",
          4759 => x"38",
          4760 => x"88",
          4761 => x"18",
          4762 => x"8c",
          4763 => x"11",
          4764 => x"90",
          4765 => x"30",
          4766 => x"25",
          4767 => x"38",
          4768 => x"80",
          4769 => x"39",
          4770 => x"57",
          4771 => x"96",
          4772 => x"33",
          4773 => x"26",
          4774 => x"33",
          4775 => x"72",
          4776 => x"7d",
          4777 => x"83",
          4778 => x"70",
          4779 => x"16",
          4780 => x"57",
          4781 => x"fd",
          4782 => x"39",
          4783 => x"30",
          4784 => x"a9",
          4785 => x"70",
          4786 => x"57",
          4787 => x"81",
          4788 => x"38",
          4789 => x"16",
          4790 => x"3d",
          4791 => x"27",
          4792 => x"08",
          4793 => x"05",
          4794 => x"38",
          4795 => x"ec",
          4796 => x"38",
          4797 => x"81",
          4798 => x"70",
          4799 => x"71",
          4800 => x"73",
          4801 => x"82",
          4802 => x"38",
          4803 => x"33",
          4804 => x"73",
          4805 => x"2e",
          4806 => x"81",
          4807 => x"38",
          4808 => x"84",
          4809 => x"38",
          4810 => x"81",
          4811 => x"33",
          4812 => x"f0",
          4813 => x"dc",
          4814 => x"07",
          4815 => x"a1",
          4816 => x"74",
          4817 => x"38",
          4818 => x"80",
          4819 => x"e1",
          4820 => x"96",
          4821 => x"9f",
          4822 => x"b5",
          4823 => x"84",
          4824 => x"54",
          4825 => x"84",
          4826 => x"83",
          4827 => x"5c",
          4828 => x"e4",
          4829 => x"80",
          4830 => x"b8",
          4831 => x"3d",
          4832 => x"70",
          4833 => x"55",
          4834 => x"81",
          4835 => x"55",
          4836 => x"80",
          4837 => x"78",
          4838 => x"73",
          4839 => x"5a",
          4840 => x"82",
          4841 => x"76",
          4842 => x"11",
          4843 => x"70",
          4844 => x"5f",
          4845 => x"72",
          4846 => x"38",
          4847 => x"23",
          4848 => x"78",
          4849 => x"58",
          4850 => x"e6",
          4851 => x"72",
          4852 => x"2e",
          4853 => x"22",
          4854 => x"76",
          4855 => x"57",
          4856 => x"70",
          4857 => x"81",
          4858 => x"55",
          4859 => x"34",
          4860 => x"73",
          4861 => x"81",
          4862 => x"2e",
          4863 => x"d0",
          4864 => x"80",
          4865 => x"85",
          4866 => x"59",
          4867 => x"75",
          4868 => x"80",
          4869 => x"54",
          4870 => x"8b",
          4871 => x"8a",
          4872 => x"26",
          4873 => x"7e",
          4874 => x"57",
          4875 => x"18",
          4876 => x"a0",
          4877 => x"83",
          4878 => x"38",
          4879 => x"82",
          4880 => x"83",
          4881 => x"81",
          4882 => x"06",
          4883 => x"90",
          4884 => x"5e",
          4885 => x"07",
          4886 => x"e4",
          4887 => x"1d",
          4888 => x"80",
          4889 => x"08",
          4890 => x"38",
          4891 => x"80",
          4892 => x"81",
          4893 => x"08",
          4894 => x"08",
          4895 => x"16",
          4896 => x"40",
          4897 => x"75",
          4898 => x"07",
          4899 => x"56",
          4900 => x"ac",
          4901 => x"09",
          4902 => x"18",
          4903 => x"1d",
          4904 => x"83",
          4905 => x"05",
          4906 => x"27",
          4907 => x"ab",
          4908 => x"84",
          4909 => x"54",
          4910 => x"74",
          4911 => x"ce",
          4912 => x"81",
          4913 => x"cd",
          4914 => x"60",
          4915 => x"12",
          4916 => x"41",
          4917 => x"d8",
          4918 => x"65",
          4919 => x"55",
          4920 => x"17",
          4921 => x"39",
          4922 => x"fd",
          4923 => x"06",
          4924 => x"2e",
          4925 => x"82",
          4926 => x"a0",
          4927 => x"06",
          4928 => x"0b",
          4929 => x"e4",
          4930 => x"ff",
          4931 => x"80",
          4932 => x"26",
          4933 => x"77",
          4934 => x"79",
          4935 => x"51",
          4936 => x"08",
          4937 => x"81",
          4938 => x"38",
          4939 => x"11",
          4940 => x"ff",
          4941 => x"38",
          4942 => x"33",
          4943 => x"73",
          4944 => x"2e",
          4945 => x"81",
          4946 => x"38",
          4947 => x"d4",
          4948 => x"26",
          4949 => x"ff",
          4950 => x"78",
          4951 => x"70",
          4952 => x"ff",
          4953 => x"1b",
          4954 => x"1b",
          4955 => x"80",
          4956 => x"33",
          4957 => x"80",
          4958 => x"83",
          4959 => x"55",
          4960 => x"39",
          4961 => x"33",
          4962 => x"77",
          4963 => x"95",
          4964 => x"2a",
          4965 => x"7c",
          4966 => x"34",
          4967 => x"83",
          4968 => x"81",
          4969 => x"38",
          4970 => x"06",
          4971 => x"84",
          4972 => x"eb",
          4973 => x"80",
          4974 => x"61",
          4975 => x"42",
          4976 => x"70",
          4977 => x"56",
          4978 => x"74",
          4979 => x"38",
          4980 => x"24",
          4981 => x"d0",
          4982 => x"58",
          4983 => x"61",
          4984 => x"5d",
          4985 => x"17",
          4986 => x"b8",
          4987 => x"06",
          4988 => x"38",
          4989 => x"b8",
          4990 => x"52",
          4991 => x"3f",
          4992 => x"70",
          4993 => x"84",
          4994 => x"75",
          4995 => x"60",
          4996 => x"18",
          4997 => x"7b",
          4998 => x"17",
          4999 => x"ff",
          5000 => x"7b",
          5001 => x"74",
          5002 => x"38",
          5003 => x"33",
          5004 => x"56",
          5005 => x"38",
          5006 => x"d9",
          5007 => x"81",
          5008 => x"8d",
          5009 => x"80",
          5010 => x"71",
          5011 => x"80",
          5012 => x"80",
          5013 => x"71",
          5014 => x"38",
          5015 => x"12",
          5016 => x"07",
          5017 => x"2b",
          5018 => x"43",
          5019 => x"80",
          5020 => x"c8",
          5021 => x"06",
          5022 => x"26",
          5023 => x"76",
          5024 => x"5f",
          5025 => x"77",
          5026 => x"78",
          5027 => x"ca",
          5028 => x"88",
          5029 => x"23",
          5030 => x"58",
          5031 => x"33",
          5032 => x"07",
          5033 => x"17",
          5034 => x"90",
          5035 => x"33",
          5036 => x"71",
          5037 => x"42",
          5038 => x"33",
          5039 => x"58",
          5040 => x"1c",
          5041 => x"26",
          5042 => x"31",
          5043 => x"e4",
          5044 => x"2e",
          5045 => x"80",
          5046 => x"83",
          5047 => x"38",
          5048 => x"eb",
          5049 => x"19",
          5050 => x"70",
          5051 => x"0c",
          5052 => x"38",
          5053 => x"80",
          5054 => x"18",
          5055 => x"8d",
          5056 => x"7a",
          5057 => x"15",
          5058 => x"18",
          5059 => x"18",
          5060 => x"80",
          5061 => x"86",
          5062 => x"bc",
          5063 => x"bc",
          5064 => x"c4",
          5065 => x"18",
          5066 => x"0c",
          5067 => x"b8",
          5068 => x"33",
          5069 => x"57",
          5070 => x"17",
          5071 => x"59",
          5072 => x"7e",
          5073 => x"7c",
          5074 => x"05",
          5075 => x"33",
          5076 => x"99",
          5077 => x"ff",
          5078 => x"77",
          5079 => x"81",
          5080 => x"9f",
          5081 => x"81",
          5082 => x"78",
          5083 => x"9f",
          5084 => x"80",
          5085 => x"1e",
          5086 => x"38",
          5087 => x"2e",
          5088 => x"06",
          5089 => x"80",
          5090 => x"57",
          5091 => x"06",
          5092 => x"32",
          5093 => x"5a",
          5094 => x"81",
          5095 => x"77",
          5096 => x"33",
          5097 => x"38",
          5098 => x"33",
          5099 => x"83",
          5100 => x"2b",
          5101 => x"59",
          5102 => x"84",
          5103 => x"57",
          5104 => x"84",
          5105 => x"9f",
          5106 => x"10",
          5107 => x"44",
          5108 => x"5b",
          5109 => x"38",
          5110 => x"b4",
          5111 => x"ff",
          5112 => x"b8",
          5113 => x"b4",
          5114 => x"2e",
          5115 => x"b4",
          5116 => x"81",
          5117 => x"07",
          5118 => x"d5",
          5119 => x"0b",
          5120 => x"e9",
          5121 => x"32",
          5122 => x"42",
          5123 => x"e8",
          5124 => x"ff",
          5125 => x"1e",
          5126 => x"81",
          5127 => x"27",
          5128 => x"b7",
          5129 => x"83",
          5130 => x"39",
          5131 => x"94",
          5132 => x"5d",
          5133 => x"71",
          5134 => x"56",
          5135 => x"80",
          5136 => x"18",
          5137 => x"70",
          5138 => x"05",
          5139 => x"5b",
          5140 => x"8e",
          5141 => x"58",
          5142 => x"93",
          5143 => x"3d",
          5144 => x"fe",
          5145 => x"83",
          5146 => x"39",
          5147 => x"3d",
          5148 => x"83",
          5149 => x"81",
          5150 => x"5c",
          5151 => x"57",
          5152 => x"38",
          5153 => x"81",
          5154 => x"58",
          5155 => x"70",
          5156 => x"ff",
          5157 => x"2e",
          5158 => x"38",
          5159 => x"fc",
          5160 => x"80",
          5161 => x"71",
          5162 => x"2e",
          5163 => x"1b",
          5164 => x"2e",
          5165 => x"7a",
          5166 => x"81",
          5167 => x"17",
          5168 => x"b8",
          5169 => x"58",
          5170 => x"f9",
          5171 => x"b7",
          5172 => x"88",
          5173 => x"d5",
          5174 => x"b8",
          5175 => x"71",
          5176 => x"14",
          5177 => x"33",
          5178 => x"5c",
          5179 => x"2e",
          5180 => x"9c",
          5181 => x"71",
          5182 => x"14",
          5183 => x"33",
          5184 => x"5a",
          5185 => x"2e",
          5186 => x"a0",
          5187 => x"71",
          5188 => x"14",
          5189 => x"33",
          5190 => x"a4",
          5191 => x"71",
          5192 => x"14",
          5193 => x"33",
          5194 => x"44",
          5195 => x"56",
          5196 => x"22",
          5197 => x"23",
          5198 => x"0b",
          5199 => x"0c",
          5200 => x"f0",
          5201 => x"95",
          5202 => x"b8",
          5203 => x"59",
          5204 => x"08",
          5205 => x"38",
          5206 => x"b4",
          5207 => x"7f",
          5208 => x"17",
          5209 => x"38",
          5210 => x"39",
          5211 => x"38",
          5212 => x"98",
          5213 => x"e3",
          5214 => x"88",
          5215 => x"f6",
          5216 => x"f6",
          5217 => x"33",
          5218 => x"88",
          5219 => x"07",
          5220 => x"1e",
          5221 => x"44",
          5222 => x"58",
          5223 => x"58",
          5224 => x"a8",
          5225 => x"59",
          5226 => x"da",
          5227 => x"17",
          5228 => x"52",
          5229 => x"3f",
          5230 => x"80",
          5231 => x"3d",
          5232 => x"75",
          5233 => x"81",
          5234 => x"55",
          5235 => x"ed",
          5236 => x"84",
          5237 => x"80",
          5238 => x"ac",
          5239 => x"2e",
          5240 => x"73",
          5241 => x"62",
          5242 => x"80",
          5243 => x"70",
          5244 => x"84",
          5245 => x"e4",
          5246 => x"84",
          5247 => x"75",
          5248 => x"56",
          5249 => x"82",
          5250 => x"5c",
          5251 => x"80",
          5252 => x"5b",
          5253 => x"81",
          5254 => x"5a",
          5255 => x"76",
          5256 => x"81",
          5257 => x"57",
          5258 => x"70",
          5259 => x"70",
          5260 => x"09",
          5261 => x"38",
          5262 => x"07",
          5263 => x"79",
          5264 => x"1d",
          5265 => x"38",
          5266 => x"24",
          5267 => x"fe",
          5268 => x"84",
          5269 => x"89",
          5270 => x"bf",
          5271 => x"53",
          5272 => x"9f",
          5273 => x"b8",
          5274 => x"79",
          5275 => x"0c",
          5276 => x"52",
          5277 => x"3f",
          5278 => x"e4",
          5279 => x"9c",
          5280 => x"38",
          5281 => x"84",
          5282 => x"58",
          5283 => x"81",
          5284 => x"38",
          5285 => x"71",
          5286 => x"58",
          5287 => x"e9",
          5288 => x"0b",
          5289 => x"34",
          5290 => x"56",
          5291 => x"57",
          5292 => x"0b",
          5293 => x"83",
          5294 => x"0b",
          5295 => x"34",
          5296 => x"9f",
          5297 => x"16",
          5298 => x"7e",
          5299 => x"57",
          5300 => x"9c",
          5301 => x"82",
          5302 => x"02",
          5303 => x"5d",
          5304 => x"86",
          5305 => x"b8",
          5306 => x"c2",
          5307 => x"5d",
          5308 => x"2a",
          5309 => x"38",
          5310 => x"38",
          5311 => x"80",
          5312 => x"58",
          5313 => x"67",
          5314 => x"9a",
          5315 => x"33",
          5316 => x"2e",
          5317 => x"9c",
          5318 => x"71",
          5319 => x"14",
          5320 => x"33",
          5321 => x"60",
          5322 => x"5d",
          5323 => x"77",
          5324 => x"34",
          5325 => x"2a",
          5326 => x"ac",
          5327 => x"75",
          5328 => x"89",
          5329 => x"70",
          5330 => x"76",
          5331 => x"06",
          5332 => x"38",
          5333 => x"3f",
          5334 => x"e4",
          5335 => x"84",
          5336 => x"38",
          5337 => x"80",
          5338 => x"95",
          5339 => x"74",
          5340 => x"80",
          5341 => x"80",
          5342 => x"80",
          5343 => x"cd",
          5344 => x"88",
          5345 => x"fc",
          5346 => x"57",
          5347 => x"17",
          5348 => x"07",
          5349 => x"39",
          5350 => x"38",
          5351 => x"3f",
          5352 => x"e4",
          5353 => x"b8",
          5354 => x"84",
          5355 => x"38",
          5356 => x"b2",
          5357 => x"90",
          5358 => x"19",
          5359 => x"ff",
          5360 => x"84",
          5361 => x"18",
          5362 => x"a0",
          5363 => x"17",
          5364 => x"cc",
          5365 => x"71",
          5366 => x"07",
          5367 => x"34",
          5368 => x"90",
          5369 => x"34",
          5370 => x"7e",
          5371 => x"34",
          5372 => x"5d",
          5373 => x"84",
          5374 => x"72",
          5375 => x"7e",
          5376 => x"79",
          5377 => x"81",
          5378 => x"16",
          5379 => x"b8",
          5380 => x"57",
          5381 => x"56",
          5382 => x"7a",
          5383 => x"0c",
          5384 => x"08",
          5385 => x"33",
          5386 => x"b8",
          5387 => x"81",
          5388 => x"17",
          5389 => x"31",
          5390 => x"a0",
          5391 => x"16",
          5392 => x"06",
          5393 => x"08",
          5394 => x"81",
          5395 => x"7c",
          5396 => x"0c",
          5397 => x"1a",
          5398 => x"ff",
          5399 => x"38",
          5400 => x"05",
          5401 => x"df",
          5402 => x"b0",
          5403 => x"2e",
          5404 => x"9c",
          5405 => x"75",
          5406 => x"39",
          5407 => x"39",
          5408 => x"0c",
          5409 => x"fe",
          5410 => x"67",
          5411 => x"0c",
          5412 => x"79",
          5413 => x"75",
          5414 => x"86",
          5415 => x"78",
          5416 => x"74",
          5417 => x"91",
          5418 => x"90",
          5419 => x"76",
          5420 => x"08",
          5421 => x"7b",
          5422 => x"2e",
          5423 => x"ff",
          5424 => x"19",
          5425 => x"5b",
          5426 => x"88",
          5427 => x"85",
          5428 => x"74",
          5429 => x"08",
          5430 => x"41",
          5431 => x"8a",
          5432 => x"08",
          5433 => x"d5",
          5434 => x"57",
          5435 => x"1b",
          5436 => x"7b",
          5437 => x"52",
          5438 => x"3f",
          5439 => x"60",
          5440 => x"2e",
          5441 => x"56",
          5442 => x"76",
          5443 => x"55",
          5444 => x"70",
          5445 => x"74",
          5446 => x"78",
          5447 => x"1e",
          5448 => x"1d",
          5449 => x"80",
          5450 => x"3d",
          5451 => x"92",
          5452 => x"39",
          5453 => x"06",
          5454 => x"78",
          5455 => x"b4",
          5456 => x"0b",
          5457 => x"7f",
          5458 => x"38",
          5459 => x"81",
          5460 => x"84",
          5461 => x"ff",
          5462 => x"7a",
          5463 => x"83",
          5464 => x"b8",
          5465 => x"e6",
          5466 => x"77",
          5467 => x"56",
          5468 => x"70",
          5469 => x"05",
          5470 => x"38",
          5471 => x"08",
          5472 => x"33",
          5473 => x"5b",
          5474 => x"81",
          5475 => x"08",
          5476 => x"1a",
          5477 => x"55",
          5478 => x"38",
          5479 => x"09",
          5480 => x"b4",
          5481 => x"7f",
          5482 => x"fe",
          5483 => x"9c",
          5484 => x"84",
          5485 => x"ff",
          5486 => x"55",
          5487 => x"ff",
          5488 => x"81",
          5489 => x"7a",
          5490 => x"0b",
          5491 => x"e4",
          5492 => x"91",
          5493 => x"0c",
          5494 => x"62",
          5495 => x"80",
          5496 => x"9f",
          5497 => x"97",
          5498 => x"8f",
          5499 => x"59",
          5500 => x"80",
          5501 => x"c4",
          5502 => x"bc",
          5503 => x"81",
          5504 => x"2e",
          5505 => x"11",
          5506 => x"76",
          5507 => x"38",
          5508 => x"a2",
          5509 => x"78",
          5510 => x"38",
          5511 => x"55",
          5512 => x"81",
          5513 => x"86",
          5514 => x"1a",
          5515 => x"60",
          5516 => x"2e",
          5517 => x"05",
          5518 => x"77",
          5519 => x"22",
          5520 => x"56",
          5521 => x"78",
          5522 => x"80",
          5523 => x"76",
          5524 => x"58",
          5525 => x"16",
          5526 => x"b8",
          5527 => x"11",
          5528 => x"27",
          5529 => x"76",
          5530 => x"70",
          5531 => x"05",
          5532 => x"38",
          5533 => x"89",
          5534 => x"1a",
          5535 => x"1b",
          5536 => x"08",
          5537 => x"27",
          5538 => x"0c",
          5539 => x"58",
          5540 => x"1b",
          5541 => x"0c",
          5542 => x"e4",
          5543 => x"33",
          5544 => x"fe",
          5545 => x"56",
          5546 => x"31",
          5547 => x"7a",
          5548 => x"2e",
          5549 => x"71",
          5550 => x"81",
          5551 => x"53",
          5552 => x"ff",
          5553 => x"80",
          5554 => x"76",
          5555 => x"60",
          5556 => x"7a",
          5557 => x"78",
          5558 => x"05",
          5559 => x"34",
          5560 => x"58",
          5561 => x"39",
          5562 => x"16",
          5563 => x"ff",
          5564 => x"e4",
          5565 => x"ab",
          5566 => x"34",
          5567 => x"84",
          5568 => x"17",
          5569 => x"33",
          5570 => x"fe",
          5571 => x"a0",
          5572 => x"16",
          5573 => x"5c",
          5574 => x"8c",
          5575 => x"16",
          5576 => x"7c",
          5577 => x"56",
          5578 => x"f8",
          5579 => x"ff",
          5580 => x"55",
          5581 => x"90",
          5582 => x"52",
          5583 => x"b8",
          5584 => x"fb",
          5585 => x"16",
          5586 => x"17",
          5587 => x"84",
          5588 => x"b8",
          5589 => x"08",
          5590 => x"17",
          5591 => x"33",
          5592 => x"fc",
          5593 => x"a0",
          5594 => x"16",
          5595 => x"56",
          5596 => x"ff",
          5597 => x"81",
          5598 => x"7a",
          5599 => x"54",
          5600 => x"53",
          5601 => x"c6",
          5602 => x"38",
          5603 => x"b4",
          5604 => x"74",
          5605 => x"82",
          5606 => x"81",
          5607 => x"16",
          5608 => x"52",
          5609 => x"3f",
          5610 => x"08",
          5611 => x"91",
          5612 => x"0c",
          5613 => x"1b",
          5614 => x"92",
          5615 => x"58",
          5616 => x"77",
          5617 => x"75",
          5618 => x"86",
          5619 => x"78",
          5620 => x"74",
          5621 => x"90",
          5622 => x"5c",
          5623 => x"7b",
          5624 => x"08",
          5625 => x"5b",
          5626 => x"53",
          5627 => x"ff",
          5628 => x"80",
          5629 => x"78",
          5630 => x"a4",
          5631 => x"5a",
          5632 => x"88",
          5633 => x"5d",
          5634 => x"88",
          5635 => x"17",
          5636 => x"74",
          5637 => x"08",
          5638 => x"5b",
          5639 => x"56",
          5640 => x"59",
          5641 => x"80",
          5642 => x"18",
          5643 => x"80",
          5644 => x"18",
          5645 => x"34",
          5646 => x"b8",
          5647 => x"06",
          5648 => x"84",
          5649 => x"81",
          5650 => x"70",
          5651 => x"93",
          5652 => x"08",
          5653 => x"83",
          5654 => x"08",
          5655 => x"74",
          5656 => x"82",
          5657 => x"81",
          5658 => x"17",
          5659 => x"52",
          5660 => x"3f",
          5661 => x"2a",
          5662 => x"2a",
          5663 => x"08",
          5664 => x"5b",
          5665 => x"56",
          5666 => x"59",
          5667 => x"80",
          5668 => x"18",
          5669 => x"80",
          5670 => x"18",
          5671 => x"34",
          5672 => x"b8",
          5673 => x"06",
          5674 => x"ae",
          5675 => x"a5",
          5676 => x"55",
          5677 => x"56",
          5678 => x"79",
          5679 => x"b8",
          5680 => x"b1",
          5681 => x"38",
          5682 => x"38",
          5683 => x"38",
          5684 => x"52",
          5685 => x"71",
          5686 => x"75",
          5687 => x"3d",
          5688 => x"8f",
          5689 => x"06",
          5690 => x"53",
          5691 => x"7d",
          5692 => x"b2",
          5693 => x"70",
          5694 => x"ac",
          5695 => x"a4",
          5696 => x"71",
          5697 => x"34",
          5698 => x"3d",
          5699 => x"0c",
          5700 => x"11",
          5701 => x"70",
          5702 => x"81",
          5703 => x"76",
          5704 => x"e4",
          5705 => x"57",
          5706 => x"70",
          5707 => x"53",
          5708 => x"e0",
          5709 => x"ff",
          5710 => x"38",
          5711 => x"54",
          5712 => x"71",
          5713 => x"73",
          5714 => x"30",
          5715 => x"59",
          5716 => x"81",
          5717 => x"25",
          5718 => x"39",
          5719 => x"5e",
          5720 => x"80",
          5721 => x"3d",
          5722 => x"08",
          5723 => x"8a",
          5724 => x"3d",
          5725 => x"3d",
          5726 => x"b8",
          5727 => x"80",
          5728 => x"70",
          5729 => x"80",
          5730 => x"84",
          5731 => x"2e",
          5732 => x"9a",
          5733 => x"33",
          5734 => x"2e",
          5735 => x"84",
          5736 => x"84",
          5737 => x"06",
          5738 => x"e4",
          5739 => x"33",
          5740 => x"90",
          5741 => x"5b",
          5742 => x"0c",
          5743 => x"3d",
          5744 => x"e6",
          5745 => x"40",
          5746 => x"3d",
          5747 => x"51",
          5748 => x"59",
          5749 => x"60",
          5750 => x"11",
          5751 => x"db",
          5752 => x"82",
          5753 => x"40",
          5754 => x"aa",
          5755 => x"b8",
          5756 => x"df",
          5757 => x"77",
          5758 => x"83",
          5759 => x"38",
          5760 => x"81",
          5761 => x"84",
          5762 => x"ff",
          5763 => x"78",
          5764 => x"9b",
          5765 => x"2b",
          5766 => x"56",
          5767 => x"76",
          5768 => x"51",
          5769 => x"08",
          5770 => x"38",
          5771 => x"3f",
          5772 => x"e4",
          5773 => x"9b",
          5774 => x"2b",
          5775 => x"5e",
          5776 => x"76",
          5777 => x"08",
          5778 => x"84",
          5779 => x"08",
          5780 => x"2e",
          5781 => x"80",
          5782 => x"51",
          5783 => x"05",
          5784 => x"38",
          5785 => x"70",
          5786 => x"81",
          5787 => x"38",
          5788 => x"82",
          5789 => x"08",
          5790 => x"56",
          5791 => x"38",
          5792 => x"5f",
          5793 => x"08",
          5794 => x"2e",
          5795 => x"c0",
          5796 => x"05",
          5797 => x"5e",
          5798 => x"1a",
          5799 => x"74",
          5800 => x"26",
          5801 => x"94",
          5802 => x"70",
          5803 => x"79",
          5804 => x"81",
          5805 => x"81",
          5806 => x"7c",
          5807 => x"e4",
          5808 => x"17",
          5809 => x"07",
          5810 => x"39",
          5811 => x"98",
          5812 => x"80",
          5813 => x"7a",
          5814 => x"e4",
          5815 => x"2e",
          5816 => x"54",
          5817 => x"53",
          5818 => x"fe",
          5819 => x"fc",
          5820 => x"17",
          5821 => x"31",
          5822 => x"a0",
          5823 => x"16",
          5824 => x"06",
          5825 => x"08",
          5826 => x"81",
          5827 => x"7c",
          5828 => x"e6",
          5829 => x"34",
          5830 => x"10",
          5831 => x"70",
          5832 => x"7a",
          5833 => x"fd",
          5834 => x"81",
          5835 => x"81",
          5836 => x"8e",
          5837 => x"19",
          5838 => x"05",
          5839 => x"fd",
          5840 => x"78",
          5841 => x"0d",
          5842 => x"55",
          5843 => x"74",
          5844 => x"73",
          5845 => x"86",
          5846 => x"78",
          5847 => x"72",
          5848 => x"91",
          5849 => x"8c",
          5850 => x"b9",
          5851 => x"76",
          5852 => x"11",
          5853 => x"73",
          5854 => x"ff",
          5855 => x"b8",
          5856 => x"53",
          5857 => x"b8",
          5858 => x"75",
          5859 => x"77",
          5860 => x"59",
          5861 => x"77",
          5862 => x"94",
          5863 => x"16",
          5864 => x"5a",
          5865 => x"73",
          5866 => x"84",
          5867 => x"08",
          5868 => x"2e",
          5869 => x"38",
          5870 => x"82",
          5871 => x"ae",
          5872 => x"53",
          5873 => x"0d",
          5874 => x"81",
          5875 => x"75",
          5876 => x"76",
          5877 => x"38",
          5878 => x"54",
          5879 => x"16",
          5880 => x"57",
          5881 => x"06",
          5882 => x"15",
          5883 => x"16",
          5884 => x"8b",
          5885 => x"0c",
          5886 => x"80",
          5887 => x"80",
          5888 => x"84",
          5889 => x"17",
          5890 => x"56",
          5891 => x"15",
          5892 => x"56",
          5893 => x"16",
          5894 => x"05",
          5895 => x"78",
          5896 => x"08",
          5897 => x"51",
          5898 => x"08",
          5899 => x"51",
          5900 => x"08",
          5901 => x"72",
          5902 => x"73",
          5903 => x"84",
          5904 => x"08",
          5905 => x"08",
          5906 => x"e4",
          5907 => x"0c",
          5908 => x"34",
          5909 => x"3d",
          5910 => x"89",
          5911 => x"53",
          5912 => x"84",
          5913 => x"e4",
          5914 => x"2e",
          5915 => x"73",
          5916 => x"04",
          5917 => x"ff",
          5918 => x"55",
          5919 => x"ab",
          5920 => x"80",
          5921 => x"70",
          5922 => x"80",
          5923 => x"9b",
          5924 => x"2b",
          5925 => x"55",
          5926 => x"88",
          5927 => x"84",
          5928 => x"99",
          5929 => x"74",
          5930 => x"ff",
          5931 => x"39",
          5932 => x"39",
          5933 => x"98",
          5934 => x"88",
          5935 => x"fa",
          5936 => x"80",
          5937 => x"80",
          5938 => x"80",
          5939 => x"16",
          5940 => x"38",
          5941 => x"73",
          5942 => x"88",
          5943 => x"fe",
          5944 => x"81",
          5945 => x"08",
          5946 => x"7a",
          5947 => x"2e",
          5948 => x"2e",
          5949 => x"2e",
          5950 => x"22",
          5951 => x"38",
          5952 => x"80",
          5953 => x"38",
          5954 => x"3f",
          5955 => x"e4",
          5956 => x"e4",
          5957 => x"ff",
          5958 => x"ff",
          5959 => x"84",
          5960 => x"2c",
          5961 => x"54",
          5962 => x"0d",
          5963 => x"ff",
          5964 => x"ff",
          5965 => x"84",
          5966 => x"2c",
          5967 => x"54",
          5968 => x"96",
          5969 => x"b8",
          5970 => x"14",
          5971 => x"b8",
          5972 => x"d8",
          5973 => x"d2",
          5974 => x"53",
          5975 => x"56",
          5976 => x"55",
          5977 => x"38",
          5978 => x"0d",
          5979 => x"a9",
          5980 => x"b8",
          5981 => x"05",
          5982 => x"74",
          5983 => x"38",
          5984 => x"3f",
          5985 => x"0d",
          5986 => x"95",
          5987 => x"68",
          5988 => x"05",
          5989 => x"84",
          5990 => x"08",
          5991 => x"9c",
          5992 => x"59",
          5993 => x"38",
          5994 => x"0c",
          5995 => x"08",
          5996 => x"82",
          5997 => x"b8",
          5998 => x"c1",
          5999 => x"56",
          6000 => x"38",
          6001 => x"81",
          6002 => x"17",
          6003 => x"b7",
          6004 => x"85",
          6005 => x"18",
          6006 => x"cc",
          6007 => x"82",
          6008 => x"11",
          6009 => x"71",
          6010 => x"72",
          6011 => x"ff",
          6012 => x"70",
          6013 => x"83",
          6014 => x"43",
          6015 => x"56",
          6016 => x"7a",
          6017 => x"07",
          6018 => x"b8",
          6019 => x"54",
          6020 => x"53",
          6021 => x"a6",
          6022 => x"fe",
          6023 => x"18",
          6024 => x"31",
          6025 => x"a0",
          6026 => x"17",
          6027 => x"06",
          6028 => x"08",
          6029 => x"81",
          6030 => x"77",
          6031 => x"92",
          6032 => x"ff",
          6033 => x"ff",
          6034 => x"08",
          6035 => x"e4",
          6036 => x"07",
          6037 => x"5a",
          6038 => x"26",
          6039 => x"18",
          6040 => x"77",
          6041 => x"17",
          6042 => x"71",
          6043 => x"25",
          6044 => x"1f",
          6045 => x"78",
          6046 => x"5a",
          6047 => x"7a",
          6048 => x"17",
          6049 => x"34",
          6050 => x"e7",
          6051 => x"56",
          6052 => x"55",
          6053 => x"54",
          6054 => x"22",
          6055 => x"2e",
          6056 => x"75",
          6057 => x"75",
          6058 => x"81",
          6059 => x"73",
          6060 => x"08",
          6061 => x"38",
          6062 => x"77",
          6063 => x"38",
          6064 => x"82",
          6065 => x"17",
          6066 => x"07",
          6067 => x"2e",
          6068 => x"55",
          6069 => x"0d",
          6070 => x"ff",
          6071 => x"ca",
          6072 => x"b8",
          6073 => x"84",
          6074 => x"38",
          6075 => x"e5",
          6076 => x"ff",
          6077 => x"82",
          6078 => x"94",
          6079 => x"27",
          6080 => x"0c",
          6081 => x"84",
          6082 => x"ff",
          6083 => x"51",
          6084 => x"08",
          6085 => x"73",
          6086 => x"80",
          6087 => x"56",
          6088 => x"39",
          6089 => x"fd",
          6090 => x"2e",
          6091 => x"81",
          6092 => x"38",
          6093 => x"19",
          6094 => x"e4",
          6095 => x"56",
          6096 => x"27",
          6097 => x"9c",
          6098 => x"80",
          6099 => x"75",
          6100 => x"e4",
          6101 => x"e3",
          6102 => x"d2",
          6103 => x"b8",
          6104 => x"84",
          6105 => x"38",
          6106 => x"fe",
          6107 => x"ff",
          6108 => x"80",
          6109 => x"94",
          6110 => x"27",
          6111 => x"84",
          6112 => x"17",
          6113 => x"a1",
          6114 => x"33",
          6115 => x"bb",
          6116 => x"56",
          6117 => x"82",
          6118 => x"86",
          6119 => x"33",
          6120 => x"90",
          6121 => x"84",
          6122 => x"56",
          6123 => x"53",
          6124 => x"3d",
          6125 => x"e4",
          6126 => x"2e",
          6127 => x"a7",
          6128 => x"08",
          6129 => x"ab",
          6130 => x"84",
          6131 => x"93",
          6132 => x"59",
          6133 => x"98",
          6134 => x"02",
          6135 => x"5d",
          6136 => x"7d",
          6137 => x"12",
          6138 => x"41",
          6139 => x"80",
          6140 => x"57",
          6141 => x"56",
          6142 => x"38",
          6143 => x"08",
          6144 => x"8b",
          6145 => x"84",
          6146 => x"b8",
          6147 => x"b4",
          6148 => x"b8",
          6149 => x"b8",
          6150 => x"16",
          6151 => x"71",
          6152 => x"5d",
          6153 => x"84",
          6154 => x"fe",
          6155 => x"08",
          6156 => x"d3",
          6157 => x"92",
          6158 => x"b8",
          6159 => x"30",
          6160 => x"7a",
          6161 => x"95",
          6162 => x"7b",
          6163 => x"26",
          6164 => x"d2",
          6165 => x"84",
          6166 => x"a7",
          6167 => x"19",
          6168 => x"76",
          6169 => x"7a",
          6170 => x"06",
          6171 => x"b8",
          6172 => x"f1",
          6173 => x"2e",
          6174 => x"b4",
          6175 => x"9c",
          6176 => x"0b",
          6177 => x"27",
          6178 => x"ff",
          6179 => x"56",
          6180 => x"96",
          6181 => x"fe",
          6182 => x"81",
          6183 => x"81",
          6184 => x"81",
          6185 => x"09",
          6186 => x"e4",
          6187 => x"a8",
          6188 => x"59",
          6189 => x"eb",
          6190 => x"2e",
          6191 => x"54",
          6192 => x"53",
          6193 => x"f1",
          6194 => x"79",
          6195 => x"74",
          6196 => x"84",
          6197 => x"08",
          6198 => x"e4",
          6199 => x"b8",
          6200 => x"80",
          6201 => x"9b",
          6202 => x"9c",
          6203 => x"58",
          6204 => x"38",
          6205 => x"33",
          6206 => x"79",
          6207 => x"80",
          6208 => x"f7",
          6209 => x"95",
          6210 => x"3d",
          6211 => x"05",
          6212 => x"3f",
          6213 => x"e4",
          6214 => x"b8",
          6215 => x"43",
          6216 => x"ff",
          6217 => x"56",
          6218 => x"0b",
          6219 => x"04",
          6220 => x"81",
          6221 => x"33",
          6222 => x"86",
          6223 => x"74",
          6224 => x"83",
          6225 => x"57",
          6226 => x"87",
          6227 => x"80",
          6228 => x"2e",
          6229 => x"7d",
          6230 => x"5d",
          6231 => x"19",
          6232 => x"80",
          6233 => x"17",
          6234 => x"05",
          6235 => x"17",
          6236 => x"76",
          6237 => x"55",
          6238 => x"22",
          6239 => x"81",
          6240 => x"17",
          6241 => x"b8",
          6242 => x"58",
          6243 => x"81",
          6244 => x"70",
          6245 => x"ee",
          6246 => x"08",
          6247 => x"18",
          6248 => x"31",
          6249 => x"ee",
          6250 => x"2e",
          6251 => x"54",
          6252 => x"53",
          6253 => x"ed",
          6254 => x"7b",
          6255 => x"fd",
          6256 => x"fd",
          6257 => x"f2",
          6258 => x"84",
          6259 => x"38",
          6260 => x"8d",
          6261 => x"fd",
          6262 => x"51",
          6263 => x"08",
          6264 => x"11",
          6265 => x"7b",
          6266 => x"0c",
          6267 => x"84",
          6268 => x"ff",
          6269 => x"9f",
          6270 => x"74",
          6271 => x"76",
          6272 => x"38",
          6273 => x"75",
          6274 => x"56",
          6275 => x"b8",
          6276 => x"c3",
          6277 => x"1a",
          6278 => x"0b",
          6279 => x"80",
          6280 => x"ff",
          6281 => x"34",
          6282 => x"17",
          6283 => x"81",
          6284 => x"d8",
          6285 => x"70",
          6286 => x"05",
          6287 => x"38",
          6288 => x"34",
          6289 => x"5b",
          6290 => x"78",
          6291 => x"34",
          6292 => x"f0",
          6293 => x"34",
          6294 => x"b8",
          6295 => x"fd",
          6296 => x"08",
          6297 => x"97",
          6298 => x"80",
          6299 => x"58",
          6300 => x"2a",
          6301 => x"5a",
          6302 => x"55",
          6303 => x"81",
          6304 => x"ed",
          6305 => x"75",
          6306 => x"04",
          6307 => x"17",
          6308 => x"ed",
          6309 => x"2a",
          6310 => x"88",
          6311 => x"7d",
          6312 => x"1b",
          6313 => x"90",
          6314 => x"88",
          6315 => x"55",
          6316 => x"81",
          6317 => x"ec",
          6318 => x"ff",
          6319 => x"b4",
          6320 => x"80",
          6321 => x"5b",
          6322 => x"ba",
          6323 => x"75",
          6324 => x"b1",
          6325 => x"51",
          6326 => x"08",
          6327 => x"8a",
          6328 => x"3d",
          6329 => x"3d",
          6330 => x"ff",
          6331 => x"56",
          6332 => x"81",
          6333 => x"86",
          6334 => x"3d",
          6335 => x"70",
          6336 => x"05",
          6337 => x"38",
          6338 => x"58",
          6339 => x"77",
          6340 => x"55",
          6341 => x"77",
          6342 => x"e4",
          6343 => x"d8",
          6344 => x"cb",
          6345 => x"b1",
          6346 => x"70",
          6347 => x"89",
          6348 => x"ff",
          6349 => x"2e",
          6350 => x"e4",
          6351 => x"5f",
          6352 => x"79",
          6353 => x"12",
          6354 => x"38",
          6355 => x"55",
          6356 => x"89",
          6357 => x"58",
          6358 => x"55",
          6359 => x"38",
          6360 => x"70",
          6361 => x"07",
          6362 => x"38",
          6363 => x"83",
          6364 => x"5a",
          6365 => x"fd",
          6366 => x"b1",
          6367 => x"51",
          6368 => x"08",
          6369 => x"38",
          6370 => x"2e",
          6371 => x"51",
          6372 => x"08",
          6373 => x"38",
          6374 => x"88",
          6375 => x"75",
          6376 => x"81",
          6377 => x"ef",
          6378 => x"19",
          6379 => x"81",
          6380 => x"a0",
          6381 => x"5d",
          6382 => x"33",
          6383 => x"75",
          6384 => x"08",
          6385 => x"19",
          6386 => x"07",
          6387 => x"83",
          6388 => x"18",
          6389 => x"27",
          6390 => x"71",
          6391 => x"75",
          6392 => x"5d",
          6393 => x"38",
          6394 => x"38",
          6395 => x"81",
          6396 => x"84",
          6397 => x"ff",
          6398 => x"7f",
          6399 => x"7b",
          6400 => x"79",
          6401 => x"6a",
          6402 => x"7b",
          6403 => x"58",
          6404 => x"5b",
          6405 => x"38",
          6406 => x"18",
          6407 => x"ed",
          6408 => x"18",
          6409 => x"3d",
          6410 => x"95",
          6411 => x"a2",
          6412 => x"b8",
          6413 => x"5c",
          6414 => x"16",
          6415 => x"33",
          6416 => x"81",
          6417 => x"53",
          6418 => x"fe",
          6419 => x"80",
          6420 => x"76",
          6421 => x"38",
          6422 => x"81",
          6423 => x"7b",
          6424 => x"fe",
          6425 => x"55",
          6426 => x"98",
          6427 => x"e1",
          6428 => x"7f",
          6429 => x"e4",
          6430 => x"0d",
          6431 => x"b1",
          6432 => x"19",
          6433 => x"07",
          6434 => x"39",
          6435 => x"fe",
          6436 => x"fe",
          6437 => x"b1",
          6438 => x"08",
          6439 => x"fe",
          6440 => x"e4",
          6441 => x"db",
          6442 => x"34",
          6443 => x"84",
          6444 => x"17",
          6445 => x"33",
          6446 => x"fe",
          6447 => x"a0",
          6448 => x"16",
          6449 => x"58",
          6450 => x"08",
          6451 => x"33",
          6452 => x"5c",
          6453 => x"84",
          6454 => x"17",
          6455 => x"e4",
          6456 => x"27",
          6457 => x"7c",
          6458 => x"38",
          6459 => x"08",
          6460 => x"51",
          6461 => x"e8",
          6462 => x"05",
          6463 => x"33",
          6464 => x"05",
          6465 => x"3f",
          6466 => x"e4",
          6467 => x"b8",
          6468 => x"5a",
          6469 => x"ff",
          6470 => x"56",
          6471 => x"80",
          6472 => x"86",
          6473 => x"61",
          6474 => x"7a",
          6475 => x"73",
          6476 => x"83",
          6477 => x"3f",
          6478 => x"0c",
          6479 => x"67",
          6480 => x"52",
          6481 => x"84",
          6482 => x"08",
          6483 => x"e4",
          6484 => x"66",
          6485 => x"95",
          6486 => x"84",
          6487 => x"cf",
          6488 => x"55",
          6489 => x"86",
          6490 => x"59",
          6491 => x"2a",
          6492 => x"2a",
          6493 => x"2a",
          6494 => x"81",
          6495 => x"e1",
          6496 => x"b8",
          6497 => x"3d",
          6498 => x"9a",
          6499 => x"ff",
          6500 => x"84",
          6501 => x"e4",
          6502 => x"7a",
          6503 => x"06",
          6504 => x"30",
          6505 => x"7b",
          6506 => x"76",
          6507 => x"80",
          6508 => x"80",
          6509 => x"f6",
          6510 => x"74",
          6511 => x"38",
          6512 => x"81",
          6513 => x"84",
          6514 => x"ff",
          6515 => x"78",
          6516 => x"56",
          6517 => x"8b",
          6518 => x"83",
          6519 => x"83",
          6520 => x"2b",
          6521 => x"70",
          6522 => x"07",
          6523 => x"56",
          6524 => x"0d",
          6525 => x"8e",
          6526 => x"3f",
          6527 => x"e4",
          6528 => x"84",
          6529 => x"80",
          6530 => x"77",
          6531 => x"70",
          6532 => x"dc",
          6533 => x"08",
          6534 => x"38",
          6535 => x"b4",
          6536 => x"b8",
          6537 => x"08",
          6538 => x"55",
          6539 => x"a0",
          6540 => x"17",
          6541 => x"33",
          6542 => x"81",
          6543 => x"16",
          6544 => x"b8",
          6545 => x"fe",
          6546 => x"f8",
          6547 => x"84",
          6548 => x"b8",
          6549 => x"5c",
          6550 => x"1b",
          6551 => x"81",
          6552 => x"8b",
          6553 => x"77",
          6554 => x"7b",
          6555 => x"a0",
          6556 => x"57",
          6557 => x"53",
          6558 => x"3d",
          6559 => x"e4",
          6560 => x"a6",
          6561 => x"55",
          6562 => x"ff",
          6563 => x"3d",
          6564 => x"5b",
          6565 => x"b7",
          6566 => x"75",
          6567 => x"74",
          6568 => x"83",
          6569 => x"51",
          6570 => x"b8",
          6571 => x"b8",
          6572 => x"76",
          6573 => x"f4",
          6574 => x"ff",
          6575 => x"81",
          6576 => x"99",
          6577 => x"ff",
          6578 => x"89",
          6579 => x"e9",
          6580 => x"81",
          6581 => x"f8",
          6582 => x"81",
          6583 => x"2a",
          6584 => x"34",
          6585 => x"05",
          6586 => x"70",
          6587 => x"58",
          6588 => x"8f",
          6589 => x"e5",
          6590 => x"38",
          6591 => x"33",
          6592 => x"06",
          6593 => x"38",
          6594 => x"3d",
          6595 => x"84",
          6596 => x"08",
          6597 => x"84",
          6598 => x"83",
          6599 => x"84",
          6600 => x"55",
          6601 => x"84",
          6602 => x"83",
          6603 => x"81",
          6604 => x"84",
          6605 => x"08",
          6606 => x"c4",
          6607 => x"76",
          6608 => x"81",
          6609 => x"ef",
          6610 => x"34",
          6611 => x"b8",
          6612 => x"39",
          6613 => x"56",
          6614 => x"84",
          6615 => x"80",
          6616 => x"75",
          6617 => x"ee",
          6618 => x"84",
          6619 => x"06",
          6620 => x"b8",
          6621 => x"80",
          6622 => x"38",
          6623 => x"09",
          6624 => x"76",
          6625 => x"51",
          6626 => x"08",
          6627 => x"59",
          6628 => x"be",
          6629 => x"57",
          6630 => x"9e",
          6631 => x"07",
          6632 => x"38",
          6633 => x"38",
          6634 => x"3f",
          6635 => x"e4",
          6636 => x"55",
          6637 => x"55",
          6638 => x"55",
          6639 => x"ff",
          6640 => x"88",
          6641 => x"59",
          6642 => x"33",
          6643 => x"15",
          6644 => x"76",
          6645 => x"81",
          6646 => x"da",
          6647 => x"7a",
          6648 => x"34",
          6649 => x"b8",
          6650 => x"57",
          6651 => x"08",
          6652 => x"fe",
          6653 => x"79",
          6654 => x"84",
          6655 => x"18",
          6656 => x"a0",
          6657 => x"33",
          6658 => x"b8",
          6659 => x"5a",
          6660 => x"3f",
          6661 => x"e4",
          6662 => x"ae",
          6663 => x"2e",
          6664 => x"54",
          6665 => x"53",
          6666 => x"d3",
          6667 => x"0d",
          6668 => x"05",
          6669 => x"80",
          6670 => x"80",
          6671 => x"80",
          6672 => x"18",
          6673 => x"c2",
          6674 => x"a5",
          6675 => x"9d",
          6676 => x"8c",
          6677 => x"33",
          6678 => x"74",
          6679 => x"11",
          6680 => x"54",
          6681 => x"ff",
          6682 => x"07",
          6683 => x"90",
          6684 => x"58",
          6685 => x"08",
          6686 => x"78",
          6687 => x"51",
          6688 => x"55",
          6689 => x"38",
          6690 => x"2e",
          6691 => x"ff",
          6692 => x"08",
          6693 => x"7d",
          6694 => x"81",
          6695 => x"73",
          6696 => x"04",
          6697 => x"3d",
          6698 => x"d0",
          6699 => x"06",
          6700 => x"08",
          6701 => x"2e",
          6702 => x"7c",
          6703 => x"74",
          6704 => x"77",
          6705 => x"84",
          6706 => x"08",
          6707 => x"17",
          6708 => x"7e",
          6709 => x"ff",
          6710 => x"8c",
          6711 => x"07",
          6712 => x"08",
          6713 => x"76",
          6714 => x"31",
          6715 => x"07",
          6716 => x"fe",
          6717 => x"74",
          6718 => x"54",
          6719 => x"39",
          6720 => x"b8",
          6721 => x"08",
          6722 => x"87",
          6723 => x"a2",
          6724 => x"80",
          6725 => x"05",
          6726 => x"75",
          6727 => x"38",
          6728 => x"d0",
          6729 => x"e5",
          6730 => x"05",
          6731 => x"84",
          6732 => x"b8",
          6733 => x"33",
          6734 => x"fe",
          6735 => x"81",
          6736 => x"83",
          6737 => x"2a",
          6738 => x"9f",
          6739 => x"52",
          6740 => x"b8",
          6741 => x"74",
          6742 => x"80",
          6743 => x"75",
          6744 => x"80",
          6745 => x"83",
          6746 => x"83",
          6747 => x"74",
          6748 => x"3d",
          6749 => x"59",
          6750 => x"ab",
          6751 => x"07",
          6752 => x"38",
          6753 => x"54",
          6754 => x"cd",
          6755 => x"08",
          6756 => x"33",
          6757 => x"2b",
          6758 => x"d4",
          6759 => x"38",
          6760 => x"11",
          6761 => x"e7",
          6762 => x"82",
          6763 => x"2b",
          6764 => x"88",
          6765 => x"1f",
          6766 => x"90",
          6767 => x"33",
          6768 => x"71",
          6769 => x"3d",
          6770 => x"45",
          6771 => x"8e",
          6772 => x"38",
          6773 => x"87",
          6774 => x"45",
          6775 => x"61",
          6776 => x"38",
          6777 => x"38",
          6778 => x"7a",
          6779 => x"7a",
          6780 => x"0b",
          6781 => x"80",
          6782 => x"38",
          6783 => x"17",
          6784 => x"2e",
          6785 => x"77",
          6786 => x"84",
          6787 => x"84",
          6788 => x"38",
          6789 => x"84",
          6790 => x"2a",
          6791 => x"15",
          6792 => x"7b",
          6793 => x"ff",
          6794 => x"4e",
          6795 => x"38",
          6796 => x"70",
          6797 => x"82",
          6798 => x"78",
          6799 => x"80",
          6800 => x"62",
          6801 => x"2e",
          6802 => x"ff",
          6803 => x"82",
          6804 => x"18",
          6805 => x"38",
          6806 => x"76",
          6807 => x"84",
          6808 => x"fe",
          6809 => x"9f",
          6810 => x"7c",
          6811 => x"57",
          6812 => x"82",
          6813 => x"5d",
          6814 => x"80",
          6815 => x"08",
          6816 => x"5c",
          6817 => x"ff",
          6818 => x"26",
          6819 => x"06",
          6820 => x"99",
          6821 => x"ff",
          6822 => x"2a",
          6823 => x"06",
          6824 => x"7a",
          6825 => x"2a",
          6826 => x"2e",
          6827 => x"5f",
          6828 => x"7f",
          6829 => x"05",
          6830 => x"dd",
          6831 => x"fe",
          6832 => x"84",
          6833 => x"38",
          6834 => x"75",
          6835 => x"59",
          6836 => x"39",
          6837 => x"7a",
          6838 => x"61",
          6839 => x"2e",
          6840 => x"4a",
          6841 => x"e4",
          6842 => x"8b",
          6843 => x"27",
          6844 => x"b8",
          6845 => x"f0",
          6846 => x"86",
          6847 => x"38",
          6848 => x"fd",
          6849 => x"80",
          6850 => x"15",
          6851 => x"e4",
          6852 => x"05",
          6853 => x"34",
          6854 => x"8b",
          6855 => x"8c",
          6856 => x"7b",
          6857 => x"8e",
          6858 => x"61",
          6859 => x"34",
          6860 => x"80",
          6861 => x"82",
          6862 => x"6c",
          6863 => x"ad",
          6864 => x"74",
          6865 => x"4c",
          6866 => x"95",
          6867 => x"80",
          6868 => x"05",
          6869 => x"61",
          6870 => x"67",
          6871 => x"4c",
          6872 => x"2a",
          6873 => x"08",
          6874 => x"85",
          6875 => x"80",
          6876 => x"05",
          6877 => x"7c",
          6878 => x"96",
          6879 => x"61",
          6880 => x"05",
          6881 => x"61",
          6882 => x"55",
          6883 => x"70",
          6884 => x"74",
          6885 => x"80",
          6886 => x"4b",
          6887 => x"53",
          6888 => x"3f",
          6889 => x"e7",
          6890 => x"87",
          6891 => x"76",
          6892 => x"55",
          6893 => x"62",
          6894 => x"ff",
          6895 => x"f8",
          6896 => x"7c",
          6897 => x"46",
          6898 => x"70",
          6899 => x"56",
          6900 => x"76",
          6901 => x"54",
          6902 => x"c5",
          6903 => x"e6",
          6904 => x"76",
          6905 => x"55",
          6906 => x"31",
          6907 => x"05",
          6908 => x"77",
          6909 => x"56",
          6910 => x"75",
          6911 => x"79",
          6912 => x"e4",
          6913 => x"76",
          6914 => x"58",
          6915 => x"6c",
          6916 => x"58",
          6917 => x"7d",
          6918 => x"06",
          6919 => x"61",
          6920 => x"57",
          6921 => x"80",
          6922 => x"60",
          6923 => x"81",
          6924 => x"05",
          6925 => x"67",
          6926 => x"c1",
          6927 => x"3f",
          6928 => x"e4",
          6929 => x"67",
          6930 => x"67",
          6931 => x"05",
          6932 => x"6b",
          6933 => x"f0",
          6934 => x"61",
          6935 => x"45",
          6936 => x"90",
          6937 => x"34",
          6938 => x"cd",
          6939 => x"52",
          6940 => x"57",
          6941 => x"80",
          6942 => x"dd",
          6943 => x"f7",
          6944 => x"b8",
          6945 => x"f0",
          6946 => x"74",
          6947 => x"39",
          6948 => x"81",
          6949 => x"74",
          6950 => x"98",
          6951 => x"82",
          6952 => x"80",
          6953 => x"38",
          6954 => x"3f",
          6955 => x"87",
          6956 => x"5c",
          6957 => x"80",
          6958 => x"0a",
          6959 => x"f8",
          6960 => x"ff",
          6961 => x"d3",
          6962 => x"bf",
          6963 => x"81",
          6964 => x"38",
          6965 => x"a0",
          6966 => x"61",
          6967 => x"7a",
          6968 => x"57",
          6969 => x"39",
          6970 => x"61",
          6971 => x"c5",
          6972 => x"05",
          6973 => x"88",
          6974 => x"7c",
          6975 => x"34",
          6976 => x"05",
          6977 => x"61",
          6978 => x"34",
          6979 => x"b0",
          6980 => x"86",
          6981 => x"05",
          6982 => x"34",
          6983 => x"61",
          6984 => x"57",
          6985 => x"76",
          6986 => x"55",
          6987 => x"70",
          6988 => x"05",
          6989 => x"38",
          6990 => x"60",
          6991 => x"81",
          6992 => x"38",
          6993 => x"62",
          6994 => x"b8",
          6995 => x"fe",
          6996 => x"0b",
          6997 => x"84",
          6998 => x"7b",
          6999 => x"34",
          7000 => x"ff",
          7001 => x"ff",
          7002 => x"05",
          7003 => x"61",
          7004 => x"34",
          7005 => x"34",
          7006 => x"86",
          7007 => x"be",
          7008 => x"80",
          7009 => x"17",
          7010 => x"d2",
          7011 => x"55",
          7012 => x"34",
          7013 => x"34",
          7014 => x"83",
          7015 => x"e5",
          7016 => x"05",
          7017 => x"34",
          7018 => x"e8",
          7019 => x"61",
          7020 => x"56",
          7021 => x"98",
          7022 => x"34",
          7023 => x"61",
          7024 => x"ee",
          7025 => x"34",
          7026 => x"34",
          7027 => x"79",
          7028 => x"81",
          7029 => x"bd",
          7030 => x"a6",
          7031 => x"5b",
          7032 => x"57",
          7033 => x"59",
          7034 => x"78",
          7035 => x"7b",
          7036 => x"8d",
          7037 => x"38",
          7038 => x"81",
          7039 => x"77",
          7040 => x"7a",
          7041 => x"84",
          7042 => x"f7",
          7043 => x"05",
          7044 => x"d5",
          7045 => x"24",
          7046 => x"8c",
          7047 => x"16",
          7048 => x"84",
          7049 => x"8b",
          7050 => x"54",
          7051 => x"51",
          7052 => x"70",
          7053 => x"30",
          7054 => x"0c",
          7055 => x"76",
          7056 => x"e3",
          7057 => x"8d",
          7058 => x"55",
          7059 => x"ff",
          7060 => x"08",
          7061 => x"38",
          7062 => x"38",
          7063 => x"77",
          7064 => x"24",
          7065 => x"19",
          7066 => x"24",
          7067 => x"55",
          7068 => x"51",
          7069 => x"08",
          7070 => x"ff",
          7071 => x"0d",
          7072 => x"75",
          7073 => x"ff",
          7074 => x"30",
          7075 => x"52",
          7076 => x"52",
          7077 => x"39",
          7078 => x"0d",
          7079 => x"05",
          7080 => x"72",
          7081 => x"ff",
          7082 => x"0c",
          7083 => x"73",
          7084 => x"81",
          7085 => x"38",
          7086 => x"2e",
          7087 => x"ff",
          7088 => x"8d",
          7089 => x"70",
          7090 => x"12",
          7091 => x"0c",
          7092 => x"0d",
          7093 => x"96",
          7094 => x"80",
          7095 => x"84",
          7096 => x"71",
          7097 => x"38",
          7098 => x"10",
          7099 => x"b8",
          7100 => x"fb",
          7101 => x"ff",
          7102 => x"ff",
          7103 => x"9f",
          7104 => x"82",
          7105 => x"80",
          7106 => x"53",
          7107 => x"05",
          7108 => x"56",
          7109 => x"70",
          7110 => x"73",
          7111 => x"22",
          7112 => x"79",
          7113 => x"2e",
          7114 => x"e4",
          7115 => x"9c",
          7116 => x"ea",
          7117 => x"05",
          7118 => x"70",
          7119 => x"51",
          7120 => x"ff",
          7121 => x"16",
          7122 => x"e6",
          7123 => x"06",
          7124 => x"83",
          7125 => x"e0",
          7126 => x"51",
          7127 => x"ff",
          7128 => x"73",
          7129 => x"83",
          7130 => x"a6",
          7131 => x"70",
          7132 => x"00",
          7133 => x"ff",
          7134 => x"ff",
          7135 => x"19",
          7136 => x"19",
          7137 => x"19",
          7138 => x"19",
          7139 => x"19",
          7140 => x"19",
          7141 => x"18",
          7142 => x"18",
          7143 => x"18",
          7144 => x"18",
          7145 => x"1f",
          7146 => x"1f",
          7147 => x"1f",
          7148 => x"1f",
          7149 => x"1f",
          7150 => x"1f",
          7151 => x"1f",
          7152 => x"1f",
          7153 => x"1f",
          7154 => x"1f",
          7155 => x"1f",
          7156 => x"1f",
          7157 => x"1f",
          7158 => x"1f",
          7159 => x"1f",
          7160 => x"1f",
          7161 => x"1f",
          7162 => x"1f",
          7163 => x"1f",
          7164 => x"1f",
          7165 => x"1f",
          7166 => x"24",
          7167 => x"1f",
          7168 => x"1f",
          7169 => x"1f",
          7170 => x"1f",
          7171 => x"1f",
          7172 => x"1f",
          7173 => x"1f",
          7174 => x"1f",
          7175 => x"23",
          7176 => x"22",
          7177 => x"23",
          7178 => x"21",
          7179 => x"1f",
          7180 => x"1f",
          7181 => x"1f",
          7182 => x"1f",
          7183 => x"1f",
          7184 => x"1f",
          7185 => x"1f",
          7186 => x"1f",
          7187 => x"1f",
          7188 => x"1f",
          7189 => x"1f",
          7190 => x"1f",
          7191 => x"1f",
          7192 => x"1f",
          7193 => x"1f",
          7194 => x"1f",
          7195 => x"1f",
          7196 => x"1f",
          7197 => x"1f",
          7198 => x"1f",
          7199 => x"1f",
          7200 => x"1f",
          7201 => x"1f",
          7202 => x"1f",
          7203 => x"1f",
          7204 => x"1f",
          7205 => x"21",
          7206 => x"1f",
          7207 => x"1f",
          7208 => x"1f",
          7209 => x"1f",
          7210 => x"21",
          7211 => x"21",
          7212 => x"21",
          7213 => x"21",
          7214 => x"32",
          7215 => x"32",
          7216 => x"32",
          7217 => x"3a",
          7218 => x"36",
          7219 => x"34",
          7220 => x"36",
          7221 => x"36",
          7222 => x"39",
          7223 => x"38",
          7224 => x"37",
          7225 => x"34",
          7226 => x"36",
          7227 => x"36",
          7228 => x"46",
          7229 => x"46",
          7230 => x"46",
          7231 => x"47",
          7232 => x"47",
          7233 => x"47",
          7234 => x"47",
          7235 => x"47",
          7236 => x"47",
          7237 => x"47",
          7238 => x"47",
          7239 => x"47",
          7240 => x"47",
          7241 => x"47",
          7242 => x"47",
          7243 => x"47",
          7244 => x"47",
          7245 => x"47",
          7246 => x"48",
          7247 => x"48",
          7248 => x"47",
          7249 => x"48",
          7250 => x"47",
          7251 => x"47",
          7252 => x"47",
          7253 => x"47",
          7254 => x"47",
          7255 => x"47",
          7256 => x"53",
          7257 => x"55",
          7258 => x"54",
          7259 => x"54",
          7260 => x"52",
          7261 => x"57",
          7262 => x"52",
          7263 => x"52",
          7264 => x"52",
          7265 => x"57",
          7266 => x"52",
          7267 => x"52",
          7268 => x"52",
          7269 => x"52",
          7270 => x"52",
          7271 => x"52",
          7272 => x"52",
          7273 => x"52",
          7274 => x"52",
          7275 => x"52",
          7276 => x"52",
          7277 => x"52",
          7278 => x"53",
          7279 => x"52",
          7280 => x"52",
          7281 => x"53",
          7282 => x"53",
          7283 => x"59",
          7284 => x"59",
          7285 => x"59",
          7286 => x"58",
          7287 => x"59",
          7288 => x"59",
          7289 => x"59",
          7290 => x"59",
          7291 => x"59",
          7292 => x"59",
          7293 => x"59",
          7294 => x"59",
          7295 => x"59",
          7296 => x"59",
          7297 => x"59",
          7298 => x"59",
          7299 => x"59",
          7300 => x"5a",
          7301 => x"5a",
          7302 => x"5a",
          7303 => x"5a",
          7304 => x"5a",
          7305 => x"59",
          7306 => x"59",
          7307 => x"59",
          7308 => x"61",
          7309 => x"61",
          7310 => x"61",
          7311 => x"61",
          7312 => x"61",
          7313 => x"61",
          7314 => x"61",
          7315 => x"61",
          7316 => x"61",
          7317 => x"61",
          7318 => x"63",
          7319 => x"61",
          7320 => x"61",
          7321 => x"5e",
          7322 => x"de",
          7323 => x"de",
          7324 => x"de",
          7325 => x"de",
          7326 => x"de",
          7327 => x"0b",
          7328 => x"0f",
          7329 => x"0b",
          7330 => x"0b",
          7331 => x"0b",
          7332 => x"0d",
          7333 => x"0f",
          7334 => x"0b",
          7335 => x"0b",
          7336 => x"0b",
          7337 => x"0b",
          7338 => x"0b",
          7339 => x"0b",
          7340 => x"0b",
          7341 => x"0b",
          7342 => x"0b",
          7343 => x"0b",
          7344 => x"0b",
          7345 => x"0b",
          7346 => x"0b",
          7347 => x"0b",
          7348 => x"0b",
          7349 => x"0b",
          7350 => x"0b",
          7351 => x"0b",
          7352 => x"0f",
          7353 => x"0b",
          7354 => x"0b",
          7355 => x"0b",
          7356 => x"0b",
          7357 => x"0b",
          7358 => x"0b",
          7359 => x"0b",
          7360 => x"0e",
          7361 => x"0e",
          7362 => x"0e",
          7363 => x"0e",
          7364 => x"0b",
          7365 => x"0b",
          7366 => x"0c",
          7367 => x"0b",
          7368 => x"0f",
          7369 => x"0c",
          7370 => x"0b",
          7371 => x"6e",
          7372 => x"6f",
          7373 => x"6e",
          7374 => x"6f",
          7375 => x"78",
          7376 => x"6c",
          7377 => x"6f",
          7378 => x"69",
          7379 => x"75",
          7380 => x"62",
          7381 => x"77",
          7382 => x"65",
          7383 => x"65",
          7384 => x"00",
          7385 => x"73",
          7386 => x"73",
          7387 => x"66",
          7388 => x"73",
          7389 => x"73",
          7390 => x"61",
          7391 => x"61",
          7392 => x"6c",
          7393 => x"00",
          7394 => x"6e",
          7395 => x"00",
          7396 => x"74",
          7397 => x"6f",
          7398 => x"00",
          7399 => x"6e",
          7400 => x"66",
          7401 => x"00",
          7402 => x"69",
          7403 => x"65",
          7404 => x"00",
          7405 => x"73",
          7406 => x"2e",
          7407 => x"74",
          7408 => x"74",
          7409 => x"63",
          7410 => x"00",
          7411 => x"20",
          7412 => x"2e",
          7413 => x"70",
          7414 => x"66",
          7415 => x"65",
          7416 => x"20",
          7417 => x"2e",
          7418 => x"6f",
          7419 => x"65",
          7420 => x"69",
          7421 => x"65",
          7422 => x"76",
          7423 => x"00",
          7424 => x"77",
          7425 => x"6f",
          7426 => x"00",
          7427 => x"61",
          7428 => x"76",
          7429 => x"00",
          7430 => x"6c",
          7431 => x"78",
          7432 => x"00",
          7433 => x"20",
          7434 => x"00",
          7435 => x"64",
          7436 => x"6d",
          7437 => x"20",
          7438 => x"75",
          7439 => x"20",
          7440 => x"75",
          7441 => x"73",
          7442 => x"65",
          7443 => x"74",
          7444 => x"72",
          7445 => x"73",
          7446 => x"00",
          7447 => x"73",
          7448 => x"6c",
          7449 => x"20",
          7450 => x"6c",
          7451 => x"2f",
          7452 => x"00",
          7453 => x"00",
          7454 => x"00",
          7455 => x"32",
          7456 => x"00",
          7457 => x"00",
          7458 => x"00",
          7459 => x"20",
          7460 => x"53",
          7461 => x"28",
          7462 => x"32",
          7463 => x"2e",
          7464 => x"50",
          7465 => x"25",
          7466 => x"20",
          7467 => x"00",
          7468 => x"74",
          7469 => x"48",
          7470 => x"00",
          7471 => x"54",
          7472 => x"72",
          7473 => x"52",
          7474 => x"6e",
          7475 => x"00",
          7476 => x"54",
          7477 => x"72",
          7478 => x"52",
          7479 => x"6e",
          7480 => x"00",
          7481 => x"57",
          7482 => x"72",
          7483 => x"43",
          7484 => x"6e",
          7485 => x"00",
          7486 => x"74",
          7487 => x"00",
          7488 => x"69",
          7489 => x"74",
          7490 => x"67",
          7491 => x"65",
          7492 => x"61",
          7493 => x"69",
          7494 => x"00",
          7495 => x"65",
          7496 => x"00",
          7497 => x"75",
          7498 => x"69",
          7499 => x"69",
          7500 => x"73",
          7501 => x"72",
          7502 => x"65",
          7503 => x"74",
          7504 => x"6c",
          7505 => x"00",
          7506 => x"00",
          7507 => x"64",
          7508 => x"64",
          7509 => x"55",
          7510 => x"3a",
          7511 => x"25",
          7512 => x"6c",
          7513 => x"74",
          7514 => x"00",
          7515 => x"74",
          7516 => x"6c",
          7517 => x"2e",
          7518 => x"6c",
          7519 => x"64",
          7520 => x"6c",
          7521 => x"00",
          7522 => x"65",
          7523 => x"63",
          7524 => x"29",
          7525 => x"65",
          7526 => x"63",
          7527 => x"30",
          7528 => x"0a",
          7529 => x"25",
          7530 => x"00",
          7531 => x"25",
          7532 => x"6d",
          7533 => x"2e",
          7534 => x"38",
          7535 => x"29",
          7536 => x"28",
          7537 => x"00",
          7538 => x"67",
          7539 => x"38",
          7540 => x"2d",
          7541 => x"6e",
          7542 => x"00",
          7543 => x"65",
          7544 => x"6f",
          7545 => x"00",
          7546 => x"5c",
          7547 => x"6d",
          7548 => x"61",
          7549 => x"63",
          7550 => x"72",
          7551 => x"6f",
          7552 => x"00",
          7553 => x"2f",
          7554 => x"64",
          7555 => x"25",
          7556 => x"43",
          7557 => x"75",
          7558 => x"00",
          7559 => x"63",
          7560 => x"65",
          7561 => x"00",
          7562 => x"73",
          7563 => x"20",
          7564 => x"73",
          7565 => x"6f",
          7566 => x"73",
          7567 => x"58",
          7568 => x"20",
          7569 => x"6d",
          7570 => x"72",
          7571 => x"73",
          7572 => x"58",
          7573 => x"20",
          7574 => x"53",
          7575 => x"64",
          7576 => x"20",
          7577 => x"58",
          7578 => x"73",
          7579 => x"20",
          7580 => x"20",
          7581 => x"20",
          7582 => x"20",
          7583 => x"58",
          7584 => x"20",
          7585 => x"20",
          7586 => x"72",
          7587 => x"20",
          7588 => x"25",
          7589 => x"00",
          7590 => x"73",
          7591 => x"44",
          7592 => x"63",
          7593 => x"20",
          7594 => x"4d",
          7595 => x"20",
          7596 => x"43",
          7597 => x"65",
          7598 => x"20",
          7599 => x"25",
          7600 => x"00",
          7601 => x"49",
          7602 => x"32",
          7603 => x"43",
          7604 => x"20",
          7605 => x"00",
          7606 => x"53",
          7607 => x"55",
          7608 => x"20",
          7609 => x"54",
          7610 => x"6e",
          7611 => x"32",
          7612 => x"20",
          7613 => x"20",
          7614 => x"65",
          7615 => x"32",
          7616 => x"20",
          7617 => x"44",
          7618 => x"69",
          7619 => x"32",
          7620 => x"20",
          7621 => x"20",
          7622 => x"58",
          7623 => x"0a",
          7624 => x"41",
          7625 => x"28",
          7626 => x"38",
          7627 => x"20",
          7628 => x"52",
          7629 => x"58",
          7630 => x"0a",
          7631 => x"52",
          7632 => x"28",
          7633 => x"38",
          7634 => x"20",
          7635 => x"41",
          7636 => x"58",
          7637 => x"0a",
          7638 => x"20",
          7639 => x"66",
          7640 => x"6b",
          7641 => x"4f",
          7642 => x"61",
          7643 => x"64",
          7644 => x"65",
          7645 => x"4f",
          7646 => x"00",
          7647 => x"f0",
          7648 => x"00",
          7649 => x"00",
          7650 => x"f0",
          7651 => x"00",
          7652 => x"00",
          7653 => x"f0",
          7654 => x"00",
          7655 => x"00",
          7656 => x"f0",
          7657 => x"00",
          7658 => x"00",
          7659 => x"f0",
          7660 => x"00",
          7661 => x"00",
          7662 => x"f0",
          7663 => x"00",
          7664 => x"00",
          7665 => x"f0",
          7666 => x"00",
          7667 => x"00",
          7668 => x"f0",
          7669 => x"00",
          7670 => x"00",
          7671 => x"f0",
          7672 => x"00",
          7673 => x"00",
          7674 => x"ef",
          7675 => x"00",
          7676 => x"00",
          7677 => x"ef",
          7678 => x"00",
          7679 => x"43",
          7680 => x"41",
          7681 => x"35",
          7682 => x"46",
          7683 => x"32",
          7684 => x"00",
          7685 => x"00",
          7686 => x"00",
          7687 => x"00",
          7688 => x"00",
          7689 => x"00",
          7690 => x"20",
          7691 => x"65",
          7692 => x"74",
          7693 => x"65",
          7694 => x"6c",
          7695 => x"73",
          7696 => x"73",
          7697 => x"00",
          7698 => x"20",
          7699 => x"69",
          7700 => x"72",
          7701 => x"65",
          7702 => x"79",
          7703 => x"6f",
          7704 => x"00",
          7705 => x"00",
          7706 => x"00",
          7707 => x"42",
          7708 => x"44",
          7709 => x"00",
          7710 => x"00",
          7711 => x"00",
          7712 => x"00",
          7713 => x"00",
          7714 => x"00",
          7715 => x"00",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"00",
          7721 => x"35",
          7722 => x"36",
          7723 => x"25",
          7724 => x"2c",
          7725 => x"64",
          7726 => x"00",
          7727 => x"64",
          7728 => x"25",
          7729 => x"3a",
          7730 => x"25",
          7731 => x"32",
          7732 => x"5b",
          7733 => x"00",
          7734 => x"20",
          7735 => x"00",
          7736 => x"78",
          7737 => x"00",
          7738 => x"78",
          7739 => x"00",
          7740 => x"78",
          7741 => x"20",
          7742 => x"66",
          7743 => x"00",
          7744 => x"3a",
          7745 => x"00",
          7746 => x"00",
          7747 => x"54",
          7748 => x"90",
          7749 => x"30",
          7750 => x"45",
          7751 => x"20",
          7752 => x"20",
          7753 => x"20",
          7754 => x"20",
          7755 => x"00",
          7756 => x"00",
          7757 => x"10",
          7758 => x"00",
          7759 => x"8f",
          7760 => x"8e",
          7761 => x"55",
          7762 => x"9e",
          7763 => x"a6",
          7764 => x"ae",
          7765 => x"b6",
          7766 => x"be",
          7767 => x"c6",
          7768 => x"ce",
          7769 => x"d6",
          7770 => x"de",
          7771 => x"e6",
          7772 => x"ee",
          7773 => x"f6",
          7774 => x"fe",
          7775 => x"5d",
          7776 => x"3f",
          7777 => x"00",
          7778 => x"02",
          7779 => x"00",
          7780 => x"00",
          7781 => x"00",
          7782 => x"00",
          7783 => x"00",
          7784 => x"00",
          7785 => x"00",
          7786 => x"00",
          7787 => x"00",
          7788 => x"00",
          7789 => x"00",
          7790 => x"00",
          7791 => x"23",
          7792 => x"00",
          7793 => x"25",
          7794 => x"25",
          7795 => x"25",
          7796 => x"25",
          7797 => x"25",
          7798 => x"25",
          7799 => x"25",
          7800 => x"25",
          7801 => x"25",
          7802 => x"25",
          7803 => x"25",
          7804 => x"25",
          7805 => x"00",
          7806 => x"03",
          7807 => x"03",
          7808 => x"03",
          7809 => x"00",
          7810 => x"23",
          7811 => x"22",
          7812 => x"00",
          7813 => x"03",
          7814 => x"03",
          7815 => x"01",
          7816 => x"01",
          7817 => x"01",
          7818 => x"02",
          7819 => x"01",
          7820 => x"01",
          7821 => x"01",
          7822 => x"01",
          7823 => x"01",
          7824 => x"01",
          7825 => x"01",
          7826 => x"01",
          7827 => x"01",
          7828 => x"01",
          7829 => x"01",
          7830 => x"01",
          7831 => x"01",
          7832 => x"01",
          7833 => x"01",
          7834 => x"01",
          7835 => x"01",
          7836 => x"01",
          7837 => x"01",
          7838 => x"00",
          7839 => x"01",
          7840 => x"01",
          7841 => x"01",
          7842 => x"02",
          7843 => x"02",
          7844 => x"02",
          7845 => x"01",
          7846 => x"01",
          7847 => x"01",
          7848 => x"02",
          7849 => x"01",
          7850 => x"02",
          7851 => x"2c",
          7852 => x"01",
          7853 => x"02",
          7854 => x"02",
          7855 => x"02",
          7856 => x"02",
          7857 => x"01",
          7858 => x"02",
          7859 => x"01",
          7860 => x"02",
          7861 => x"03",
          7862 => x"03",
          7863 => x"03",
          7864 => x"03",
          7865 => x"03",
          7866 => x"00",
          7867 => x"03",
          7868 => x"03",
          7869 => x"03",
          7870 => x"03",
          7871 => x"04",
          7872 => x"04",
          7873 => x"04",
          7874 => x"01",
          7875 => x"00",
          7876 => x"1e",
          7877 => x"1f",
          7878 => x"1f",
          7879 => x"1f",
          7880 => x"1f",
          7881 => x"1f",
          7882 => x"06",
          7883 => x"1f",
          7884 => x"1f",
          7885 => x"1f",
          7886 => x"1f",
          7887 => x"06",
          7888 => x"00",
          7889 => x"1f",
          7890 => x"1f",
          7891 => x"1f",
          7892 => x"00",
          7893 => x"21",
          7894 => x"00",
          7895 => x"2c",
          7896 => x"2c",
          7897 => x"2c",
          7898 => x"ff",
          7899 => x"00",
          7900 => x"01",
          7901 => x"00",
          7902 => x"01",
          7903 => x"00",
          7904 => x"03",
          7905 => x"00",
          7906 => x"03",
          7907 => x"00",
          7908 => x"03",
          7909 => x"00",
          7910 => x"04",
          7911 => x"00",
          7912 => x"04",
          7913 => x"00",
          7914 => x"04",
          7915 => x"00",
          7916 => x"04",
          7917 => x"00",
          7918 => x"04",
          7919 => x"00",
          7920 => x"04",
          7921 => x"00",
          7922 => x"04",
          7923 => x"00",
          7924 => x"05",
          7925 => x"00",
          7926 => x"05",
          7927 => x"00",
          7928 => x"05",
          7929 => x"00",
          7930 => x"05",
          7931 => x"00",
          7932 => x"07",
          7933 => x"00",
          7934 => x"07",
          7935 => x"00",
          7936 => x"08",
          7937 => x"00",
          7938 => x"08",
          7939 => x"00",
          7940 => x"08",
          7941 => x"00",
          7942 => x"08",
          7943 => x"00",
          7944 => x"08",
          7945 => x"00",
          7946 => x"08",
          7947 => x"00",
          7948 => x"09",
          7949 => x"00",
          7950 => x"09",
          7951 => x"00",
          7952 => x"09",
          7953 => x"00",
          7954 => x"09",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"00",
          7959 => x"00",
          7960 => x"00",
          7961 => x"00",
          7962 => x"78",
          7963 => x"e1",
          7964 => x"e1",
          7965 => x"01",
          7966 => x"10",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"f0",
          7980 => x"f0",
          7981 => x"f0",
          7982 => x"fd",
          7983 => x"3a",
          7984 => x"f0",
          7985 => x"77",
          7986 => x"6f",
          7987 => x"67",
          7988 => x"37",
          7989 => x"2c",
          7990 => x"3f",
          7991 => x"f0",
          7992 => x"f0",
          7993 => x"3b",
          7994 => x"f0",
          7995 => x"57",
          7996 => x"4f",
          7997 => x"47",
          7998 => x"37",
          7999 => x"2c",
          8000 => x"3f",
          8001 => x"f0",
          8002 => x"f0",
          8003 => x"2a",
          8004 => x"f0",
          8005 => x"57",
          8006 => x"4f",
          8007 => x"47",
          8008 => x"27",
          8009 => x"3c",
          8010 => x"3f",
          8011 => x"f0",
          8012 => x"f0",
          8013 => x"f0",
          8014 => x"f0",
          8015 => x"17",
          8016 => x"0f",
          8017 => x"07",
          8018 => x"f0",
          8019 => x"f0",
          8020 => x"f0",
          8021 => x"f0",
          8022 => x"f0",
          8023 => x"4d",
          8024 => x"f0",
          8025 => x"78",
          8026 => x"d5",
          8027 => x"4c",
          8028 => x"5f",
          8029 => x"d0",
          8030 => x"bb",
          8031 => x"f0",
          8032 => x"f0",
          8033 => x"00",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"00",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"01",
          9068 => x"f2",
          9069 => x"fa",
          9070 => x"c2",
          9071 => x"e5",
          9072 => x"62",
          9073 => x"6b",
          9074 => x"22",
          9075 => x"4f",
          9076 => x"02",
          9077 => x"0a",
          9078 => x"12",
          9079 => x"1a",
          9080 => x"82",
          9081 => x"8a",
          9082 => x"92",
          9083 => x"9a",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"93",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"2d",
             6 => x"00",
             7 => x"00",
             8 => x"fd",
             9 => x"05",
            10 => x"ff",
            11 => x"00",
            12 => x"fd",
            13 => x"06",
            14 => x"2b",
            15 => x"0b",
            16 => x"09",
            17 => x"06",
            18 => x"0a",
            19 => x"00",
            20 => x"72",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"73",
            25 => x"81",
            26 => x"10",
            27 => x"51",
            28 => x"72",
            29 => x"04",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"0a",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"72",
            45 => x"0b",
            46 => x"00",
            47 => x"00",
            48 => x"72",
            49 => x"74",
            50 => x"07",
            51 => x"00",
            52 => x"71",
            53 => x"09",
            54 => x"2b",
            55 => x"04",
            56 => x"09",
            57 => x"05",
            58 => x"04",
            59 => x"00",
            60 => x"09",
            61 => x"05",
            62 => x"51",
            63 => x"00",
            64 => x"09",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"72",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"09",
            73 => x"53",
            74 => x"00",
            75 => x"00",
            76 => x"fc",
            77 => x"05",
            78 => x"ff",
            79 => x"00",
            80 => x"fc",
            81 => x"73",
            82 => x"0b",
            83 => x"00",
            84 => x"08",
            85 => x"0b",
            86 => x"08",
            87 => x"51",
            88 => x"08",
            89 => x"0b",
            90 => x"08",
            91 => x"51",
            92 => x"09",
            93 => x"06",
            94 => x"09",
            95 => x"51",
            96 => x"09",
            97 => x"81",
            98 => x"73",
            99 => x"07",
           100 => x"ff",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"81",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"84",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"0d",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"8c",
           134 => x"04",
           135 => x"0b",
           136 => x"8c",
           137 => x"04",
           138 => x"0b",
           139 => x"8d",
           140 => x"04",
           141 => x"0b",
           142 => x"8d",
           143 => x"04",
           144 => x"0b",
           145 => x"8e",
           146 => x"04",
           147 => x"0b",
           148 => x"8e",
           149 => x"04",
           150 => x"0b",
           151 => x"8f",
           152 => x"04",
           153 => x"0b",
           154 => x"8f",
           155 => x"04",
           156 => x"0b",
           157 => x"90",
           158 => x"04",
           159 => x"0b",
           160 => x"90",
           161 => x"04",
           162 => x"0b",
           163 => x"91",
           164 => x"04",
           165 => x"0b",
           166 => x"91",
           167 => x"04",
           168 => x"0b",
           169 => x"92",
           170 => x"04",
           171 => x"0b",
           172 => x"92",
           173 => x"04",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"00",
           193 => x"80",
           194 => x"80",
           195 => x"0c",
           196 => x"80",
           197 => x"0c",
           198 => x"80",
           199 => x"0c",
           200 => x"80",
           201 => x"0c",
           202 => x"80",
           203 => x"0c",
           204 => x"80",
           205 => x"0c",
           206 => x"80",
           207 => x"0c",
           208 => x"80",
           209 => x"0c",
           210 => x"80",
           211 => x"0c",
           212 => x"80",
           213 => x"0c",
           214 => x"80",
           215 => x"0c",
           216 => x"80",
           217 => x"0c",
           218 => x"08",
           219 => x"f0",
           220 => x"f0",
           221 => x"b8",
           222 => x"b8",
           223 => x"84",
           224 => x"84",
           225 => x"04",
           226 => x"2d",
           227 => x"90",
           228 => x"ef",
           229 => x"80",
           230 => x"d2",
           231 => x"c0",
           232 => x"82",
           233 => x"80",
           234 => x"0c",
           235 => x"08",
           236 => x"f0",
           237 => x"f0",
           238 => x"b8",
           239 => x"b8",
           240 => x"84",
           241 => x"84",
           242 => x"04",
           243 => x"2d",
           244 => x"90",
           245 => x"cf",
           246 => x"80",
           247 => x"84",
           248 => x"c0",
           249 => x"82",
           250 => x"80",
           251 => x"0c",
           252 => x"08",
           253 => x"f0",
           254 => x"f0",
           255 => x"b8",
           256 => x"b8",
           257 => x"84",
           258 => x"84",
           259 => x"04",
           260 => x"2d",
           261 => x"90",
           262 => x"d6",
           263 => x"80",
           264 => x"e6",
           265 => x"c0",
           266 => x"82",
           267 => x"80",
           268 => x"0c",
           269 => x"08",
           270 => x"f0",
           271 => x"f0",
           272 => x"b8",
           273 => x"b8",
           274 => x"84",
           275 => x"84",
           276 => x"04",
           277 => x"2d",
           278 => x"90",
           279 => x"82",
           280 => x"80",
           281 => x"b7",
           282 => x"c0",
           283 => x"81",
           284 => x"80",
           285 => x"0c",
           286 => x"08",
           287 => x"f0",
           288 => x"f0",
           289 => x"b8",
           290 => x"b8",
           291 => x"84",
           292 => x"84",
           293 => x"04",
           294 => x"2d",
           295 => x"90",
           296 => x"2d",
           297 => x"90",
           298 => x"f0",
           299 => x"80",
           300 => x"dc",
           301 => x"c0",
           302 => x"81",
           303 => x"80",
           304 => x"0c",
           305 => x"08",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"51",
           311 => x"73",
           312 => x"10",
           313 => x"0c",
           314 => x"81",
           315 => x"71",
           316 => x"72",
           317 => x"84",
           318 => x"8e",
           319 => x"0c",
           320 => x"81",
           321 => x"3d",
           322 => x"52",
           323 => x"c8",
           324 => x"0d",
           325 => x"85",
           326 => x"73",
           327 => x"52",
           328 => x"d3",
           329 => x"70",
           330 => x"55",
           331 => x"38",
           332 => x"8e",
           333 => x"84",
           334 => x"84",
           335 => x"57",
           336 => x"30",
           337 => x"54",
           338 => x"75",
           339 => x"0c",
           340 => x"b8",
           341 => x"3d",
           342 => x"99",
           343 => x"8e",
           344 => x"3d",
           345 => x"54",
           346 => x"fd",
           347 => x"76",
           348 => x"0d",
           349 => x"42",
           350 => x"85",
           351 => x"81",
           352 => x"7b",
           353 => x"7b",
           354 => x"38",
           355 => x"72",
           356 => x"5f",
           357 => x"b0",
           358 => x"54",
           359 => x"a9",
           360 => x"81",
           361 => x"38",
           362 => x"57",
           363 => x"54",
           364 => x"0d",
           365 => x"10",
           366 => x"70",
           367 => x"29",
           368 => x"5a",
           369 => x"86",
           370 => x"bd",
           371 => x"fe",
           372 => x"2e",
           373 => x"74",
           374 => x"5a",
           375 => x"7c",
           376 => x"33",
           377 => x"39",
           378 => x"55",
           379 => x"40",
           380 => x"72",
           381 => x"10",
           382 => x"04",
           383 => x"73",
           384 => x"8a",
           385 => x"76",
           386 => x"ff",
           387 => x"60",
           388 => x"cf",
           389 => x"f4",
           390 => x"3f",
           391 => x"84",
           392 => x"53",
           393 => x"e4",
           394 => x"81",
           395 => x"90",
           396 => x"84",
           397 => x"b8",
           398 => x"40",
           399 => x"84",
           400 => x"70",
           401 => x"70",
           402 => x"9e",
           403 => x"80",
           404 => x"38",
           405 => x"80",
           406 => x"83",
           407 => x"80",
           408 => x"81",
           409 => x"86",
           410 => x"70",
           411 => x"5b",
           412 => x"85",
           413 => x"70",
           414 => x"59",
           415 => x"7a",
           416 => x"eb",
           417 => x"73",
           418 => x"06",
           419 => x"06",
           420 => x"2a",
           421 => x"38",
           422 => x"80",
           423 => x"54",
           424 => x"b0",
           425 => x"80",
           426 => x"90",
           427 => x"e5",
           428 => x"2e",
           429 => x"29",
           430 => x"5b",
           431 => x"7c",
           432 => x"79",
           433 => x"05",
           434 => x"80",
           435 => x"81",
           436 => x"b9",
           437 => x"38",
           438 => x"76",
           439 => x"84",
           440 => x"ff",
           441 => x"3f",
           442 => x"06",
           443 => x"80",
           444 => x"80",
           445 => x"90",
           446 => x"fc",
           447 => x"f4",
           448 => x"7a",
           449 => x"fa",
           450 => x"c0",
           451 => x"61",
           452 => x"cf",
           453 => x"fd",
           454 => x"80",
           455 => x"2b",
           456 => x"fc",
           457 => x"52",
           458 => x"2a",
           459 => x"c9",
           460 => x"fc",
           461 => x"54",
           462 => x"7c",
           463 => x"39",
           464 => x"5b",
           465 => x"ca",
           466 => x"57",
           467 => x"ff",
           468 => x"54",
           469 => x"38",
           470 => x"33",
           471 => x"fc",
           472 => x"84",
           473 => x"70",
           474 => x"7b",
           475 => x"57",
           476 => x"7f",
           477 => x"40",
           478 => x"38",
           479 => x"b8",
           480 => x"07",
           481 => x"38",
           482 => x"80",
           483 => x"38",
           484 => x"71",
           485 => x"5f",
           486 => x"f6",
           487 => x"ff",
           488 => x"5a",
           489 => x"7a",
           490 => x"76",
           491 => x"60",
           492 => x"5d",
           493 => x"75",
           494 => x"08",
           495 => x"90",
           496 => x"80",
           497 => x"88",
           498 => x"80",
           499 => x"90",
           500 => x"fa",
           501 => x"c4",
           502 => x"83",
           503 => x"06",
           504 => x"83",
           505 => x"5f",
           506 => x"d8",
           507 => x"90",
           508 => x"06",
           509 => x"38",
           510 => x"82",
           511 => x"80",
           512 => x"7c",
           513 => x"3f",
           514 => x"f7",
           515 => x"31",
           516 => x"f9",
           517 => x"c4",
           518 => x"82",
           519 => x"75",
           520 => x"08",
           521 => x"90",
           522 => x"82",
           523 => x"06",
           524 => x"3d",
           525 => x"52",
           526 => x"0d",
           527 => x"0b",
           528 => x"70",
           529 => x"51",
           530 => x"77",
           531 => x"74",
           532 => x"77",
           533 => x"52",
           534 => x"2d",
           535 => x"38",
           536 => x"33",
           537 => x"d4",
           538 => x"c8",
           539 => x"8a",
           540 => x"84",
           541 => x"ff",
           542 => x"0c",
           543 => x"78",
           544 => x"33",
           545 => x"06",
           546 => x"77",
           547 => x"70",
           548 => x"2e",
           549 => x"75",
           550 => x"04",
           551 => x"72",
           552 => x"51",
           553 => x"b8",
           554 => x"74",
           555 => x"72",
           556 => x"84",
           557 => x"3f",
           558 => x"78",
           559 => x"81",
           560 => x"ff",
           561 => x"81",
           562 => x"8c",
           563 => x"25",
           564 => x"34",
           565 => x"15",
           566 => x"76",
           567 => x"3d",
           568 => x"06",
           569 => x"ff",
           570 => x"8c",
           571 => x"76",
           572 => x"85",
           573 => x"81",
           574 => x"ff",
           575 => x"81",
           576 => x"2a",
           577 => x"c3",
           578 => x"71",
           579 => x"76",
           580 => x"17",
           581 => x"84",
           582 => x"74",
           583 => x"34",
           584 => x"0c",
           585 => x"87",
           586 => x"08",
           587 => x"52",
           588 => x"b9",
           589 => x"54",
           590 => x"85",
           591 => x"17",
           592 => x"0c",
           593 => x"53",
           594 => x"39",
           595 => x"54",
           596 => x"51",
           597 => x"70",
           598 => x"70",
           599 => x"73",
           600 => x"04",
           601 => x"55",
           602 => x"38",
           603 => x"2e",
           604 => x"33",
           605 => x"11",
           606 => x"e4",
           607 => x"55",
           608 => x"75",
           609 => x"53",
           610 => x"70",
           611 => x"13",
           612 => x"11",
           613 => x"3d",
           614 => x"81",
           615 => x"ff",
           616 => x"0c",
           617 => x"0d",
           618 => x"70",
           619 => x"70",
           620 => x"73",
           621 => x"04",
           622 => x"55",
           623 => x"38",
           624 => x"70",
           625 => x"70",
           626 => x"85",
           627 => x"78",
           628 => x"a1",
           629 => x"57",
           630 => x"81",
           631 => x"80",
           632 => x"e1",
           633 => x"0c",
           634 => x"f1",
           635 => x"80",
           636 => x"81",
           637 => x"72",
           638 => x"0d",
           639 => x"3d",
           640 => x"53",
           641 => x"b8",
           642 => x"05",
           643 => x"b8",
           644 => x"80",
           645 => x"15",
           646 => x"52",
           647 => x"3f",
           648 => x"b8",
           649 => x"3d",
           650 => x"53",
           651 => x"70",
           652 => x"2e",
           653 => x"2e",
           654 => x"70",
           655 => x"e4",
           656 => x"0d",
           657 => x"54",
           658 => x"70",
           659 => x"70",
           660 => x"85",
           661 => x"7a",
           662 => x"8b",
           663 => x"b8",
           664 => x"80",
           665 => x"3f",
           666 => x"80",
           667 => x"73",
           668 => x"81",
           669 => x"76",
           670 => x"56",
           671 => x"74",
           672 => x"78",
           673 => x"81",
           674 => x"ff",
           675 => x"55",
           676 => x"07",
           677 => x"3d",
           678 => x"fc",
           679 => x"07",
           680 => x"31",
           681 => x"06",
           682 => x"88",
           683 => x"f0",
           684 => x"2b",
           685 => x"53",
           686 => x"30",
           687 => x"77",
           688 => x"70",
           689 => x"06",
           690 => x"51",
           691 => x"53",
           692 => x"56",
           693 => x"0d",
           694 => x"54",
           695 => x"84",
           696 => x"31",
           697 => x"0d",
           698 => x"54",
           699 => x"76",
           700 => x"08",
           701 => x"8d",
           702 => x"84",
           703 => x"71",
           704 => x"71",
           705 => x"71",
           706 => x"57",
           707 => x"2e",
           708 => x"07",
           709 => x"ff",
           710 => x"72",
           711 => x"56",
           712 => x"da",
           713 => x"3d",
           714 => x"2c",
           715 => x"32",
           716 => x"32",
           717 => x"56",
           718 => x"3f",
           719 => x"31",
           720 => x"04",
           721 => x"80",
           722 => x"56",
           723 => x"06",
           724 => x"70",
           725 => x"38",
           726 => x"b0",
           727 => x"80",
           728 => x"8a",
           729 => x"c4",
           730 => x"e0",
           731 => x"d0",
           732 => x"90",
           733 => x"81",
           734 => x"81",
           735 => x"38",
           736 => x"79",
           737 => x"a0",
           738 => x"84",
           739 => x"81",
           740 => x"3d",
           741 => x"0c",
           742 => x"2e",
           743 => x"15",
           744 => x"73",
           745 => x"73",
           746 => x"a0",
           747 => x"80",
           748 => x"e1",
           749 => x"3d",
           750 => x"78",
           751 => x"fe",
           752 => x"0c",
           753 => x"7b",
           754 => x"77",
           755 => x"a0",
           756 => x"15",
           757 => x"73",
           758 => x"80",
           759 => x"38",
           760 => x"26",
           761 => x"a0",
           762 => x"74",
           763 => x"ff",
           764 => x"ff",
           765 => x"38",
           766 => x"54",
           767 => x"78",
           768 => x"13",
           769 => x"56",
           770 => x"38",
           771 => x"56",
           772 => x"b8",
           773 => x"70",
           774 => x"56",
           775 => x"fe",
           776 => x"70",
           777 => x"a6",
           778 => x"a0",
           779 => x"38",
           780 => x"89",
           781 => x"b8",
           782 => x"58",
           783 => x"55",
           784 => x"0b",
           785 => x"04",
           786 => x"08",
           787 => x"04",
           788 => x"26",
           789 => x"f4",
           790 => x"8c",
           791 => x"04",
           792 => x"83",
           793 => x"ef",
           794 => x"ce",
           795 => x"0d",
           796 => x"3f",
           797 => x"51",
           798 => x"83",
           799 => x"3d",
           800 => x"f1",
           801 => x"cc",
           802 => x"04",
           803 => x"83",
           804 => x"ee",
           805 => x"d0",
           806 => x"0d",
           807 => x"3f",
           808 => x"51",
           809 => x"83",
           810 => x"3d",
           811 => x"99",
           812 => x"f8",
           813 => x"04",
           814 => x"83",
           815 => x"ed",
           816 => x"d1",
           817 => x"0d",
           818 => x"3f",
           819 => x"66",
           820 => x"5b",
           821 => x"07",
           822 => x"57",
           823 => x"57",
           824 => x"51",
           825 => x"81",
           826 => x"58",
           827 => x"08",
           828 => x"80",
           829 => x"3f",
           830 => x"7b",
           831 => x"57",
           832 => x"87",
           833 => x"e7",
           834 => x"87",
           835 => x"b8",
           836 => x"78",
           837 => x"3f",
           838 => x"0d",
           839 => x"98",
           840 => x"96",
           841 => x"75",
           842 => x"84",
           843 => x"08",
           844 => x"2e",
           845 => x"57",
           846 => x"51",
           847 => x"52",
           848 => x"e4",
           849 => x"52",
           850 => x"ff",
           851 => x"84",
           852 => x"58",
           853 => x"ec",
           854 => x"76",
           855 => x"8a",
           856 => x"3d",
           857 => x"56",
           858 => x"53",
           859 => x"b8",
           860 => x"3d",
           861 => x"63",
           862 => x"73",
           863 => x"5f",
           864 => x"38",
           865 => x"fe",
           866 => x"3f",
           867 => x"7c",
           868 => x"2e",
           869 => x"7a",
           870 => x"83",
           871 => x"14",
           872 => x"51",
           873 => x"38",
           874 => x"80",
           875 => x"75",
           876 => x"72",
           877 => x"53",
           878 => x"74",
           879 => x"57",
           880 => x"74",
           881 => x"08",
           882 => x"16",
           883 => x"d2",
           884 => x"79",
           885 => x"3f",
           886 => x"98",
           887 => x"ee",
           888 => x"7b",
           889 => x"38",
           890 => x"3d",
           891 => x"ae",
           892 => x"53",
           893 => x"74",
           894 => x"83",
           895 => x"14",
           896 => x"51",
           897 => x"c0",
           898 => x"df",
           899 => x"51",
           900 => x"c8",
           901 => x"3f",
           902 => x"39",
           903 => x"84",
           904 => x"a0",
           905 => x"fd",
           906 => x"27",
           907 => x"ec",
           908 => x"d4",
           909 => x"84",
           910 => x"d8",
           911 => x"51",
           912 => x"91",
           913 => x"e4",
           914 => x"72",
           915 => x"72",
           916 => x"e0",
           917 => x"51",
           918 => x"98",
           919 => x"70",
           920 => x"72",
           921 => x"58",
           922 => x"fd",
           923 => x"84",
           924 => x"2c",
           925 => x"32",
           926 => x"07",
           927 => x"53",
           928 => x"b9",
           929 => x"8f",
           930 => x"c0",
           931 => x"81",
           932 => x"51",
           933 => x"3f",
           934 => x"52",
           935 => x"70",
           936 => x"38",
           937 => x"52",
           938 => x"70",
           939 => x"38",
           940 => x"52",
           941 => x"70",
           942 => x"38",
           943 => x"52",
           944 => x"06",
           945 => x"84",
           946 => x"3f",
           947 => x"80",
           948 => x"84",
           949 => x"3f",
           950 => x"80",
           951 => x"81",
           952 => x"cb",
           953 => x"d3",
           954 => x"9b",
           955 => x"06",
           956 => x"38",
           957 => x"83",
           958 => x"51",
           959 => x"81",
           960 => x"f0",
           961 => x"80",
           962 => x"3f",
           963 => x"2a",
           964 => x"2e",
           965 => x"51",
           966 => x"9a",
           967 => x"72",
           968 => x"71",
           969 => x"39",
           970 => x"ec",
           971 => x"b0",
           972 => x"51",
           973 => x"ff",
           974 => x"83",
           975 => x"51",
           976 => x"81",
           977 => x"b8",
           978 => x"80",
           979 => x"f0",
           980 => x"b5",
           981 => x"ff",
           982 => x"2e",
           983 => x"e3",
           984 => x"88",
           985 => x"f8",
           986 => x"3f",
           987 => x"81",
           988 => x"82",
           989 => x"38",
           990 => x"2e",
           991 => x"79",
           992 => x"5c",
           993 => x"38",
           994 => x"a0",
           995 => x"26",
           996 => x"dc",
           997 => x"3f",
           998 => x"08",
           999 => x"e8",
          1000 => x"38",
          1001 => x"83",
          1002 => x"06",
          1003 => x"9a",
          1004 => x"dd",
          1005 => x"92",
          1006 => x"b8",
          1007 => x"84",
          1008 => x"80",
          1009 => x"e4",
          1010 => x"80",
          1011 => x"08",
          1012 => x"08",
          1013 => x"a5",
          1014 => x"85",
          1015 => x"7a",
          1016 => x"80",
          1017 => x"d5",
          1018 => x"b9",
          1019 => x"54",
          1020 => x"52",
          1021 => x"e4",
          1022 => x"30",
          1023 => x"5b",
          1024 => x"38",
          1025 => x"80",
          1026 => x"ff",
          1027 => x"7f",
          1028 => x"7c",
          1029 => x"e8",
          1030 => x"83",
          1031 => x"48",
          1032 => x"e8",
          1033 => x"33",
          1034 => x"fd",
          1035 => x"52",
          1036 => x"3f",
          1037 => x"81",
          1038 => x"84",
          1039 => x"51",
          1040 => x"08",
          1041 => x"08",
          1042 => x"ed",
          1043 => x"59",
          1044 => x"d3",
          1045 => x"82",
          1046 => x"83",
          1047 => x"80",
          1048 => x"67",
          1049 => x"90",
          1050 => x"33",
          1051 => x"38",
          1052 => x"5a",
          1053 => x"94",
          1054 => x"53",
          1055 => x"84",
          1056 => x"2e",
          1057 => x"70",
          1058 => x"39",
          1059 => x"7d",
          1060 => x"39",
          1061 => x"d5",
          1062 => x"52",
          1063 => x"39",
          1064 => x"9a",
          1065 => x"83",
          1066 => x"81",
          1067 => x"d5",
          1068 => x"78",
          1069 => x"3f",
          1070 => x"3d",
          1071 => x"51",
          1072 => x"80",
          1073 => x"d5",
          1074 => x"79",
          1075 => x"fa",
          1076 => x"83",
          1077 => x"95",
          1078 => x"ff",
          1079 => x"b8",
          1080 => x"68",
          1081 => x"3f",
          1082 => x"f4",
          1083 => x"a8",
          1084 => x"f9",
          1085 => x"53",
          1086 => x"84",
          1087 => x"59",
          1088 => x"c4",
          1089 => x"08",
          1090 => x"91",
          1091 => x"ae",
          1092 => x"87",
          1093 => x"59",
          1094 => x"53",
          1095 => x"84",
          1096 => x"38",
          1097 => x"80",
          1098 => x"e4",
          1099 => x"22",
          1100 => x"cf",
          1101 => x"80",
          1102 => x"7e",
          1103 => x"f8",
          1104 => x"38",
          1105 => x"39",
          1106 => x"80",
          1107 => x"e4",
          1108 => x"3d",
          1109 => x"51",
          1110 => x"80",
          1111 => x"f8",
          1112 => x"c4",
          1113 => x"f7",
          1114 => x"b6",
          1115 => x"27",
          1116 => x"33",
          1117 => x"38",
          1118 => x"78",
          1119 => x"3f",
          1120 => x"1b",
          1121 => x"84",
          1122 => x"f4",
          1123 => x"f7",
          1124 => x"53",
          1125 => x"84",
          1126 => x"38",
          1127 => x"80",
          1128 => x"e4",
          1129 => x"d7",
          1130 => x"79",
          1131 => x"79",
          1132 => x"65",
          1133 => x"ff",
          1134 => x"e8",
          1135 => x"2e",
          1136 => x"11",
          1137 => x"3f",
          1138 => x"70",
          1139 => x"cc",
          1140 => x"80",
          1141 => x"7e",
          1142 => x"f6",
          1143 => x"38",
          1144 => x"59",
          1145 => x"68",
          1146 => x"11",
          1147 => x"3f",
          1148 => x"dd",
          1149 => x"33",
          1150 => x"3d",
          1151 => x"51",
          1152 => x"ff",
          1153 => x"ff",
          1154 => x"e6",
          1155 => x"2e",
          1156 => x"11",
          1157 => x"3f",
          1158 => x"8d",
          1159 => x"ff",
          1160 => x"b8",
          1161 => x"08",
          1162 => x"3f",
          1163 => x"8f",
          1164 => x"05",
          1165 => x"8a",
          1166 => x"b8",
          1167 => x"3f",
          1168 => x"80",
          1169 => x"53",
          1170 => x"ea",
          1171 => x"2e",
          1172 => x"51",
          1173 => x"3d",
          1174 => x"51",
          1175 => x"91",
          1176 => x"80",
          1177 => x"08",
          1178 => x"ff",
          1179 => x"b8",
          1180 => x"33",
          1181 => x"83",
          1182 => x"f8",
          1183 => x"8c",
          1184 => x"a5",
          1185 => x"2e",
          1186 => x"70",
          1187 => x"06",
          1188 => x"38",
          1189 => x"83",
          1190 => x"55",
          1191 => x"51",
          1192 => x"d6",
          1193 => x"71",
          1194 => x"3d",
          1195 => x"51",
          1196 => x"80",
          1197 => x"0c",
          1198 => x"fe",
          1199 => x"e2",
          1200 => x"38",
          1201 => x"ce",
          1202 => x"23",
          1203 => x"53",
          1204 => x"84",
          1205 => x"38",
          1206 => x"7e",
          1207 => x"b8",
          1208 => x"05",
          1209 => x"08",
          1210 => x"3d",
          1211 => x"51",
          1212 => x"80",
          1213 => x"80",
          1214 => x"05",
          1215 => x"f0",
          1216 => x"80",
          1217 => x"81",
          1218 => x"64",
          1219 => x"39",
          1220 => x"9d",
          1221 => x"80",
          1222 => x"c8",
          1223 => x"7c",
          1224 => x"83",
          1225 => x"f5",
          1226 => x"ff",
          1227 => x"b8",
          1228 => x"59",
          1229 => x"82",
          1230 => x"39",
          1231 => x"2e",
          1232 => x"47",
          1233 => x"5c",
          1234 => x"a8",
          1235 => x"84",
          1236 => x"b6",
          1237 => x"3f",
          1238 => x"ea",
          1239 => x"83",
          1240 => x"83",
          1241 => x"c6",
          1242 => x"80",
          1243 => x"47",
          1244 => x"5e",
          1245 => x"b8",
          1246 => x"eb",
          1247 => x"83",
          1248 => x"83",
          1249 => x"9b",
          1250 => x"b9",
          1251 => x"80",
          1252 => x"47",
          1253 => x"fc",
          1254 => x"f1",
          1255 => x"39",
          1256 => x"94",
          1257 => x"56",
          1258 => x"da",
          1259 => x"2b",
          1260 => x"52",
          1261 => x"b8",
          1262 => x"94",
          1263 => x"80",
          1264 => x"b8",
          1265 => x"55",
          1266 => x"93",
          1267 => x"77",
          1268 => x"94",
          1269 => x"c0",
          1270 => x"81",
          1271 => x"a1",
          1272 => x"0b",
          1273 => x"72",
          1274 => x"f4",
          1275 => x"ba",
          1276 => x"a0",
          1277 => x"3f",
          1278 => x"94",
          1279 => x"d2",
          1280 => x"d2",
          1281 => x"3f",
          1282 => x"0d",
          1283 => x"52",
          1284 => x"74",
          1285 => x"70",
          1286 => x"81",
          1287 => x"53",
          1288 => x"71",
          1289 => x"81",
          1290 => x"80",
          1291 => x"ff",
          1292 => x"83",
          1293 => x"38",
          1294 => x"52",
          1295 => x"52",
          1296 => x"83",
          1297 => x"30",
          1298 => x"53",
          1299 => x"70",
          1300 => x"74",
          1301 => x"3d",
          1302 => x"73",
          1303 => x"52",
          1304 => x"53",
          1305 => x"81",
          1306 => x"75",
          1307 => x"06",
          1308 => x"0d",
          1309 => x"0b",
          1310 => x"04",
          1311 => x"db",
          1312 => x"2e",
          1313 => x"86",
          1314 => x"82",
          1315 => x"52",
          1316 => x"13",
          1317 => x"9e",
          1318 => x"51",
          1319 => x"38",
          1320 => x"bb",
          1321 => x"55",
          1322 => x"38",
          1323 => x"87",
          1324 => x"22",
          1325 => x"80",
          1326 => x"9c",
          1327 => x"0c",
          1328 => x"0c",
          1329 => x"0c",
          1330 => x"0c",
          1331 => x"0c",
          1332 => x"0c",
          1333 => x"87",
          1334 => x"c0",
          1335 => x"b8",
          1336 => x"3d",
          1337 => x"5d",
          1338 => x"08",
          1339 => x"b8",
          1340 => x"c0",
          1341 => x"34",
          1342 => x"84",
          1343 => x"5a",
          1344 => x"a8",
          1345 => x"c0",
          1346 => x"23",
          1347 => x"8a",
          1348 => x"ff",
          1349 => x"06",
          1350 => x"33",
          1351 => x"33",
          1352 => x"ff",
          1353 => x"ff",
          1354 => x"fe",
          1355 => x"72",
          1356 => x"e8",
          1357 => x"2b",
          1358 => x"2e",
          1359 => x"2e",
          1360 => x"84",
          1361 => x"89",
          1362 => x"70",
          1363 => x"09",
          1364 => x"e7",
          1365 => x"2b",
          1366 => x"2e",
          1367 => x"80",
          1368 => x"81",
          1369 => x"e4",
          1370 => x"52",
          1371 => x"07",
          1372 => x"db",
          1373 => x"3d",
          1374 => x"05",
          1375 => x"ff",
          1376 => x"80",
          1377 => x"70",
          1378 => x"52",
          1379 => x"2a",
          1380 => x"38",
          1381 => x"80",
          1382 => x"06",
          1383 => x"06",
          1384 => x"80",
          1385 => x"52",
          1386 => x"0c",
          1387 => x"70",
          1388 => x"72",
          1389 => x"2e",
          1390 => x"52",
          1391 => x"94",
          1392 => x"06",
          1393 => x"39",
          1394 => x"70",
          1395 => x"70",
          1396 => x"04",
          1397 => x"33",
          1398 => x"80",
          1399 => x"33",
          1400 => x"71",
          1401 => x"94",
          1402 => x"06",
          1403 => x"38",
          1404 => x"51",
          1405 => x"06",
          1406 => x"93",
          1407 => x"75",
          1408 => x"80",
          1409 => x"c0",
          1410 => x"17",
          1411 => x"38",
          1412 => x"0d",
          1413 => x"51",
          1414 => x"81",
          1415 => x"71",
          1416 => x"2e",
          1417 => x"08",
          1418 => x"54",
          1419 => x"3d",
          1420 => x"9c",
          1421 => x"2e",
          1422 => x"08",
          1423 => x"a8",
          1424 => x"9e",
          1425 => x"c0",
          1426 => x"87",
          1427 => x"0c",
          1428 => x"b4",
          1429 => x"f1",
          1430 => x"83",
          1431 => x"08",
          1432 => x"b8",
          1433 => x"9e",
          1434 => x"c0",
          1435 => x"87",
          1436 => x"0c",
          1437 => x"83",
          1438 => x"08",
          1439 => x"88",
          1440 => x"9e",
          1441 => x"0b",
          1442 => x"c0",
          1443 => x"06",
          1444 => x"71",
          1445 => x"c0",
          1446 => x"06",
          1447 => x"38",
          1448 => x"80",
          1449 => x"90",
          1450 => x"80",
          1451 => x"f1",
          1452 => x"90",
          1453 => x"52",
          1454 => x"52",
          1455 => x"87",
          1456 => x"80",
          1457 => x"83",
          1458 => x"34",
          1459 => x"70",
          1460 => x"70",
          1461 => x"83",
          1462 => x"9e",
          1463 => x"51",
          1464 => x"81",
          1465 => x"0b",
          1466 => x"80",
          1467 => x"2e",
          1468 => x"ec",
          1469 => x"08",
          1470 => x"52",
          1471 => x"71",
          1472 => x"c0",
          1473 => x"06",
          1474 => x"38",
          1475 => x"80",
          1476 => x"a0",
          1477 => x"2e",
          1478 => x"ef",
          1479 => x"80",
          1480 => x"83",
          1481 => x"9e",
          1482 => x"52",
          1483 => x"52",
          1484 => x"9e",
          1485 => x"2a",
          1486 => x"80",
          1487 => x"88",
          1488 => x"83",
          1489 => x"34",
          1490 => x"51",
          1491 => x"0d",
          1492 => x"3d",
          1493 => x"de",
          1494 => x"86",
          1495 => x"b9",
          1496 => x"85",
          1497 => x"73",
          1498 => x"56",
          1499 => x"33",
          1500 => x"ea",
          1501 => x"f1",
          1502 => x"83",
          1503 => x"38",
          1504 => x"ed",
          1505 => x"83",
          1506 => x"73",
          1507 => x"55",
          1508 => x"33",
          1509 => x"ee",
          1510 => x"d8",
          1511 => x"c8",
          1512 => x"b5",
          1513 => x"83",
          1514 => x"83",
          1515 => x"51",
          1516 => x"51",
          1517 => x"52",
          1518 => x"3f",
          1519 => x"c0",
          1520 => x"b8",
          1521 => x"71",
          1522 => x"52",
          1523 => x"3f",
          1524 => x"c3",
          1525 => x"8a",
          1526 => x"3d",
          1527 => x"bd",
          1528 => x"3f",
          1529 => x"29",
          1530 => x"e4",
          1531 => x"b4",
          1532 => x"87",
          1533 => x"56",
          1534 => x"b3",
          1535 => x"c0",
          1536 => x"b8",
          1537 => x"ff",
          1538 => x"55",
          1539 => x"9a",
          1540 => x"3f",
          1541 => x"83",
          1542 => x"51",
          1543 => x"08",
          1544 => x"c6",
          1545 => x"d9",
          1546 => x"d9",
          1547 => x"d4",
          1548 => x"b3",
          1549 => x"bd",
          1550 => x"3f",
          1551 => x"29",
          1552 => x"e4",
          1553 => x"b2",
          1554 => x"74",
          1555 => x"39",
          1556 => x"3f",
          1557 => x"2e",
          1558 => x"db",
          1559 => x"f1",
          1560 => x"e5",
          1561 => x"ff",
          1562 => x"55",
          1563 => x"39",
          1564 => x"3f",
          1565 => x"2e",
          1566 => x"f2",
          1567 => x"b2",
          1568 => x"75",
          1569 => x"83",
          1570 => x"51",
          1571 => x"33",
          1572 => x"cd",
          1573 => x"dc",
          1574 => x"f1",
          1575 => x"c0",
          1576 => x"83",
          1577 => x"dc",
          1578 => x"f1",
          1579 => x"97",
          1580 => x"83",
          1581 => x"dc",
          1582 => x"f1",
          1583 => x"ee",
          1584 => x"83",
          1585 => x"dc",
          1586 => x"f1",
          1587 => x"c5",
          1588 => x"83",
          1589 => x"dc",
          1590 => x"f1",
          1591 => x"9c",
          1592 => x"83",
          1593 => x"dd",
          1594 => x"f1",
          1595 => x"f3",
          1596 => x"ff",
          1597 => x"ff",
          1598 => x"55",
          1599 => x"39",
          1600 => x"52",
          1601 => x"10",
          1602 => x"04",
          1603 => x"3f",
          1604 => x"51",
          1605 => x"04",
          1606 => x"3f",
          1607 => x"51",
          1608 => x"04",
          1609 => x"3f",
          1610 => x"51",
          1611 => x"04",
          1612 => x"87",
          1613 => x"f8",
          1614 => x"d9",
          1615 => x"08",
          1616 => x"52",
          1617 => x"82",
          1618 => x"38",
          1619 => x"d0",
          1620 => x"51",
          1621 => x"08",
          1622 => x"f6",
          1623 => x"57",
          1624 => x"25",
          1625 => x"05",
          1626 => x"74",
          1627 => x"2a",
          1628 => x"38",
          1629 => x"08",
          1630 => x"9a",
          1631 => x"78",
          1632 => x"e4",
          1633 => x"98",
          1634 => x"2e",
          1635 => x"79",
          1636 => x"86",
          1637 => x"e4",
          1638 => x"c4",
          1639 => x"84",
          1640 => x"d8",
          1641 => x"08",
          1642 => x"5a",
          1643 => x"80",
          1644 => x"10",
          1645 => x"52",
          1646 => x"e4",
          1647 => x"c0",
          1648 => x"38",
          1649 => x"81",
          1650 => x"81",
          1651 => x"82",
          1652 => x"84",
          1653 => x"81",
          1654 => x"53",
          1655 => x"84",
          1656 => x"ff",
          1657 => x"a7",
          1658 => x"06",
          1659 => x"16",
          1660 => x"76",
          1661 => x"78",
          1662 => x"fe",
          1663 => x"33",
          1664 => x"06",
          1665 => x"38",
          1666 => x"cd",
          1667 => x"83",
          1668 => x"ea",
          1669 => x"38",
          1670 => x"52",
          1671 => x"b8",
          1672 => x"51",
          1673 => x"08",
          1674 => x"25",
          1675 => x"05",
          1676 => x"77",
          1677 => x"8c",
          1678 => x"ff",
          1679 => x"81",
          1680 => x"0d",
          1681 => x"b7",
          1682 => x"5c",
          1683 => x"d4",
          1684 => x"74",
          1685 => x"56",
          1686 => x"77",
          1687 => x"77",
          1688 => x"77",
          1689 => x"b4",
          1690 => x"3f",
          1691 => x"98",
          1692 => x"38",
          1693 => x"33",
          1694 => x"d0",
          1695 => x"2c",
          1696 => x"83",
          1697 => x"33",
          1698 => x"58",
          1699 => x"80",
          1700 => x"38",
          1701 => x"0a",
          1702 => x"76",
          1703 => x"70",
          1704 => x"dd",
          1705 => x"25",
          1706 => x"18",
          1707 => x"81",
          1708 => x"75",
          1709 => x"80",
          1710 => x"98",
          1711 => x"33",
          1712 => x"98",
          1713 => x"f0",
          1714 => x"5d",
          1715 => x"38",
          1716 => x"39",
          1717 => x"81",
          1718 => x"70",
          1719 => x"57",
          1720 => x"75",
          1721 => x"80",
          1722 => x"57",
          1723 => x"ec",
          1724 => x"78",
          1725 => x"2e",
          1726 => x"57",
          1727 => x"e7",
          1728 => x"57",
          1729 => x"a0",
          1730 => x"7e",
          1731 => x"95",
          1732 => x"83",
          1733 => x"83",
          1734 => x"0b",
          1735 => x"d0",
          1736 => x"33",
          1737 => x"84",
          1738 => x"b6",
          1739 => x"05",
          1740 => x"eb",
          1741 => x"ff",
          1742 => x"55",
          1743 => x"d4",
          1744 => x"84",
          1745 => x"52",
          1746 => x"39",
          1747 => x"10",
          1748 => x"57",
          1749 => x"d0",
          1750 => x"a4",
          1751 => x"74",
          1752 => x"08",
          1753 => x"84",
          1754 => x"b5",
          1755 => x"88",
          1756 => x"a8",
          1757 => x"a8",
          1758 => x"cc",
          1759 => x"75",
          1760 => x"7c",
          1761 => x"75",
          1762 => x"f1",
          1763 => x"75",
          1764 => x"80",
          1765 => x"b7",
          1766 => x"d0",
          1767 => x"ff",
          1768 => x"51",
          1769 => x"33",
          1770 => x"80",
          1771 => x"08",
          1772 => x"84",
          1773 => x"b4",
          1774 => x"88",
          1775 => x"a8",
          1776 => x"a8",
          1777 => x"39",
          1778 => x"06",
          1779 => x"75",
          1780 => x"c8",
          1781 => x"d0",
          1782 => x"55",
          1783 => x"33",
          1784 => x"33",
          1785 => x"83",
          1786 => x"15",
          1787 => x"16",
          1788 => x"3f",
          1789 => x"06",
          1790 => x"77",
          1791 => x"39",
          1792 => x"33",
          1793 => x"38",
          1794 => x"34",
          1795 => x"81",
          1796 => x"24",
          1797 => x"52",
          1798 => x"d0",
          1799 => x"2c",
          1800 => x"41",
          1801 => x"d4",
          1802 => x"9c",
          1803 => x"80",
          1804 => x"a4",
          1805 => x"f8",
          1806 => x"88",
          1807 => x"80",
          1808 => x"98",
          1809 => x"5a",
          1810 => x"bb",
          1811 => x"78",
          1812 => x"33",
          1813 => x"80",
          1814 => x"98",
          1815 => x"55",
          1816 => x"16",
          1817 => x"d4",
          1818 => x"b1",
          1819 => x"81",
          1820 => x"d0",
          1821 => x"24",
          1822 => x"d0",
          1823 => x"d3",
          1824 => x"51",
          1825 => x"33",
          1826 => x"34",
          1827 => x"84",
          1828 => x"7f",
          1829 => x"51",
          1830 => x"52",
          1831 => x"e4",
          1832 => x"cf",
          1833 => x"80",
          1834 => x"33",
          1835 => x"70",
          1836 => x"38",
          1837 => x"f1",
          1838 => x"5b",
          1839 => x"08",
          1840 => x"10",
          1841 => x"57",
          1842 => x"f2",
          1843 => x"38",
          1844 => x"2e",
          1845 => x"a8",
          1846 => x"7b",
          1847 => x"04",
          1848 => x"2e",
          1849 => x"88",
          1850 => x"c8",
          1851 => x"3f",
          1852 => x"ff",
          1853 => x"ff",
          1854 => x"75",
          1855 => x"83",
          1856 => x"80",
          1857 => x"84",
          1858 => x"7c",
          1859 => x"d0",
          1860 => x"38",
          1861 => x"ff",
          1862 => x"52",
          1863 => x"d4",
          1864 => x"ac",
          1865 => x"5d",
          1866 => x"ff",
          1867 => x"e0",
          1868 => x"84",
          1869 => x"a4",
          1870 => x"3d",
          1871 => x"81",
          1872 => x"f4",
          1873 => x"05",
          1874 => x"16",
          1875 => x"d4",
          1876 => x"cc",
          1877 => x"2b",
          1878 => x"5a",
          1879 => x"ef",
          1880 => x"51",
          1881 => x"33",
          1882 => x"d0",
          1883 => x"7a",
          1884 => x"08",
          1885 => x"74",
          1886 => x"05",
          1887 => x"5b",
          1888 => x"38",
          1889 => x"ff",
          1890 => x"29",
          1891 => x"84",
          1892 => x"75",
          1893 => x"7b",
          1894 => x"84",
          1895 => x"ff",
          1896 => x"29",
          1897 => x"84",
          1898 => x"61",
          1899 => x"81",
          1900 => x"08",
          1901 => x"3f",
          1902 => x"0a",
          1903 => x"33",
          1904 => x"a7",
          1905 => x"33",
          1906 => x"60",
          1907 => x"33",
          1908 => x"98",
          1909 => x"76",
          1910 => x"33",
          1911 => x"29",
          1912 => x"84",
          1913 => x"78",
          1914 => x"84",
          1915 => x"7c",
          1916 => x"84",
          1917 => x"8b",
          1918 => x"a4",
          1919 => x"70",
          1920 => x"05",
          1921 => x"44",
          1922 => x"ef",
          1923 => x"78",
          1924 => x"7a",
          1925 => x"08",
          1926 => x"75",
          1927 => x"05",
          1928 => x"57",
          1929 => x"38",
          1930 => x"ff",
          1931 => x"29",
          1932 => x"84",
          1933 => x"76",
          1934 => x"83",
          1935 => x"f4",
          1936 => x"3f",
          1937 => x"34",
          1938 => x"81",
          1939 => x"ad",
          1940 => x"d0",
          1941 => x"f4",
          1942 => x"88",
          1943 => x"c8",
          1944 => x"3f",
          1945 => x"ff",
          1946 => x"ff",
          1947 => x"7a",
          1948 => x"51",
          1949 => x"08",
          1950 => x"08",
          1951 => x"34",
          1952 => x"84",
          1953 => x"33",
          1954 => x"81",
          1955 => x"70",
          1956 => x"57",
          1957 => x"d0",
          1958 => x"2c",
          1959 => x"58",
          1960 => x"e4",
          1961 => x"ee",
          1962 => x"56",
          1963 => x"16",
          1964 => x"f0",
          1965 => x"83",
          1966 => x"ee",
          1967 => x"3f",
          1968 => x"fe",
          1969 => x"93",
          1970 => x"39",
          1971 => x"77",
          1972 => x"75",
          1973 => x"39",
          1974 => x"b8",
          1975 => x"b8",
          1976 => x"53",
          1977 => x"3f",
          1978 => x"d0",
          1979 => x"2e",
          1980 => x"52",
          1981 => x"d4",
          1982 => x"fc",
          1983 => x"51",
          1984 => x"33",
          1985 => x"34",
          1986 => x"80",
          1987 => x"34",
          1988 => x"84",
          1989 => x"75",
          1990 => x"e4",
          1991 => x"e4",
          1992 => x"75",
          1993 => x"81",
          1994 => x"a4",
          1995 => x"5e",
          1996 => x"84",
          1997 => x"a6",
          1998 => x"a0",
          1999 => x"c8",
          2000 => x"3f",
          2001 => x"76",
          2002 => x"06",
          2003 => x"8e",
          2004 => x"a4",
          2005 => x"06",
          2006 => x"ff",
          2007 => x"ff",
          2008 => x"a8",
          2009 => x"2e",
          2010 => x"52",
          2011 => x"d4",
          2012 => x"8c",
          2013 => x"51",
          2014 => x"33",
          2015 => x"34",
          2016 => x"74",
          2017 => x"d4",
          2018 => x"83",
          2019 => x"52",
          2020 => x"b8",
          2021 => x"33",
          2022 => x"70",
          2023 => x"f4",
          2024 => x"51",
          2025 => x"33",
          2026 => x"56",
          2027 => x"83",
          2028 => x"3d",
          2029 => x"52",
          2030 => x"f2",
          2031 => x"88",
          2032 => x"df",
          2033 => x"34",
          2034 => x"84",
          2035 => x"93",
          2036 => x"51",
          2037 => x"08",
          2038 => x"96",
          2039 => x"53",
          2040 => x"f2",
          2041 => x"b8",
          2042 => x"e9",
          2043 => x"ff",
          2044 => x"56",
          2045 => x"80",
          2046 => x"05",
          2047 => x"75",
          2048 => x"70",
          2049 => x"08",
          2050 => x"38",
          2051 => x"f1",
          2052 => x"55",
          2053 => x"08",
          2054 => x"10",
          2055 => x"57",
          2056 => x"70",
          2057 => x"27",
          2058 => x"09",
          2059 => x"ed",
          2060 => x"52",
          2061 => x"f2",
          2062 => x"06",
          2063 => x"38",
          2064 => x"bd",
          2065 => x"83",
          2066 => x"fc",
          2067 => x"70",
          2068 => x"3f",
          2069 => x"f2",
          2070 => x"fc",
          2071 => x"80",
          2072 => x"76",
          2073 => x"75",
          2074 => x"83",
          2075 => x"77",
          2076 => x"3d",
          2077 => x"84",
          2078 => x"72",
          2079 => x"2e",
          2080 => x"9e",
          2081 => x"86",
          2082 => x"80",
          2083 => x"58",
          2084 => x"f8",
          2085 => x"75",
          2086 => x"33",
          2087 => x"71",
          2088 => x"56",
          2089 => x"38",
          2090 => x"74",
          2091 => x"74",
          2092 => x"38",
          2093 => x"17",
          2094 => x"0b",
          2095 => x"81",
          2096 => x"ee",
          2097 => x"a0",
          2098 => x"10",
          2099 => x"90",
          2100 => x"40",
          2101 => x"b6",
          2102 => x"b6",
          2103 => x"f8",
          2104 => x"70",
          2105 => x"57",
          2106 => x"72",
          2107 => x"ff",
          2108 => x"ff",
          2109 => x"81",
          2110 => x"42",
          2111 => x"8f",
          2112 => x"31",
          2113 => x"76",
          2114 => x"9c",
          2115 => x"26",
          2116 => x"05",
          2117 => x"70",
          2118 => x"a7",
          2119 => x"70",
          2120 => x"06",
          2121 => x"06",
          2122 => x"5d",
          2123 => x"74",
          2124 => x"ff",
          2125 => x"29",
          2126 => x"fd",
          2127 => x"34",
          2128 => x"f8",
          2129 => x"2b",
          2130 => x"7a",
          2131 => x"26",
          2132 => x"fc",
          2133 => x"81",
          2134 => x"f8",
          2135 => x"a7",
          2136 => x"56",
          2137 => x"84",
          2138 => x"84",
          2139 => x"83",
          2140 => x"06",
          2141 => x"41",
          2142 => x"73",
          2143 => x"70",
          2144 => x"ff",
          2145 => x"29",
          2146 => x"ff",
          2147 => x"5c",
          2148 => x"77",
          2149 => x"79",
          2150 => x"38",
          2151 => x"38",
          2152 => x"29",
          2153 => x"86",
          2154 => x"34",
          2155 => x"73",
          2156 => x"f4",
          2157 => x"ee",
          2158 => x"76",
          2159 => x"74",
          2160 => x"34",
          2161 => x"86",
          2162 => x"81",
          2163 => x"77",
          2164 => x"34",
          2165 => x"c0",
          2166 => x"a0",
          2167 => x"07",
          2168 => x"34",
          2169 => x"53",
          2170 => x"b6",
          2171 => x"0c",
          2172 => x"33",
          2173 => x"0d",
          2174 => x"b3",
          2175 => x"59",
          2176 => x"da",
          2177 => x"95",
          2178 => x"29",
          2179 => x"f8",
          2180 => x"7c",
          2181 => x"83",
          2182 => x"72",
          2183 => x"92",
          2184 => x"92",
          2185 => x"70",
          2186 => x"55",
          2187 => x"38",
          2188 => x"34",
          2189 => x"ff",
          2190 => x"57",
          2191 => x"b6",
          2192 => x"80",
          2193 => x"84",
          2194 => x"e0",
          2195 => x"70",
          2196 => x"05",
          2197 => x"d5",
          2198 => x"26",
          2199 => x"97",
          2200 => x"e0",
          2201 => x"55",
          2202 => x"27",
          2203 => x"05",
          2204 => x"57",
          2205 => x"ff",
          2206 => x"fd",
          2207 => x"b6",
          2208 => x"57",
          2209 => x"86",
          2210 => x"75",
          2211 => x"5c",
          2212 => x"38",
          2213 => x"14",
          2214 => x"78",
          2215 => x"81",
          2216 => x"59",
          2217 => x"84",
          2218 => x"56",
          2219 => x"38",
          2220 => x"8b",
          2221 => x"34",
          2222 => x"ff",
          2223 => x"57",
          2224 => x"80",
          2225 => x"06",
          2226 => x"53",
          2227 => x"c8",
          2228 => x"b6",
          2229 => x"29",
          2230 => x"27",
          2231 => x"84",
          2232 => x"56",
          2233 => x"75",
          2234 => x"13",
          2235 => x"a0",
          2236 => x"70",
          2237 => x"72",
          2238 => x"84",
          2239 => x"39",
          2240 => x"b6",
          2241 => x"d7",
          2242 => x"0d",
          2243 => x"53",
          2244 => x"10",
          2245 => x"08",
          2246 => x"71",
          2247 => x"34",
          2248 => x"3d",
          2249 => x"34",
          2250 => x"06",
          2251 => x"ff",
          2252 => x"80",
          2253 => x"0d",
          2254 => x"31",
          2255 => x"54",
          2256 => x"34",
          2257 => x"05",
          2258 => x"56",
          2259 => x"53",
          2260 => x"84",
          2261 => x"83",
          2262 => x"09",
          2263 => x"53",
          2264 => x"0b",
          2265 => x"04",
          2266 => x"b6",
          2267 => x"70",
          2268 => x"83",
          2269 => x"e4",
          2270 => x"83",
          2271 => x"84",
          2272 => x"71",
          2273 => x"51",
          2274 => x"39",
          2275 => x"51",
          2276 => x"10",
          2277 => x"04",
          2278 => x"06",
          2279 => x"72",
          2280 => x"71",
          2281 => x"38",
          2282 => x"80",
          2283 => x"0d",
          2284 => x"06",
          2285 => x"34",
          2286 => x"3d",
          2287 => x"f0",
          2288 => x"e8",
          2289 => x"06",
          2290 => x"34",
          2291 => x"90",
          2292 => x"83",
          2293 => x"81",
          2294 => x"f8",
          2295 => x"90",
          2296 => x"90",
          2297 => x"33",
          2298 => x"83",
          2299 => x"f8",
          2300 => x"51",
          2301 => x"39",
          2302 => x"81",
          2303 => x"fe",
          2304 => x"f8",
          2305 => x"fe",
          2306 => x"df",
          2307 => x"f8",
          2308 => x"90",
          2309 => x"70",
          2310 => x"83",
          2311 => x"e0",
          2312 => x"fe",
          2313 => x"cf",
          2314 => x"f8",
          2315 => x"90",
          2316 => x"70",
          2317 => x"83",
          2318 => x"70",
          2319 => x"83",
          2320 => x"07",
          2321 => x"e0",
          2322 => x"33",
          2323 => x"83",
          2324 => x"83",
          2325 => x"43",
          2326 => x"2e",
          2327 => x"38",
          2328 => x"84",
          2329 => x"dc",
          2330 => x"83",
          2331 => x"34",
          2332 => x"09",
          2333 => x"b6",
          2334 => x"34",
          2335 => x"0b",
          2336 => x"f8",
          2337 => x"33",
          2338 => x"b6",
          2339 => x"7a",
          2340 => x"e6",
          2341 => x"0b",
          2342 => x"94",
          2343 => x"83",
          2344 => x"80",
          2345 => x"84",
          2346 => x"94",
          2347 => x"80",
          2348 => x"e7",
          2349 => x"84",
          2350 => x"54",
          2351 => x"51",
          2352 => x"b7",
          2353 => x"a5",
          2354 => x"70",
          2355 => x"ff",
          2356 => x"ff",
          2357 => x"59",
          2358 => x"94",
          2359 => x"b6",
          2360 => x"34",
          2361 => x"f8",
          2362 => x"8f",
          2363 => x"da",
          2364 => x"81",
          2365 => x"83",
          2366 => x"92",
          2367 => x"ae",
          2368 => x"e3",
          2369 => x"59",
          2370 => x"3f",
          2371 => x"a6",
          2372 => x"83",
          2373 => x"81",
          2374 => x"d8",
          2375 => x"05",
          2376 => x"83",
          2377 => x"72",
          2378 => x"11",
          2379 => x"5c",
          2380 => x"ff",
          2381 => x"51",
          2382 => x"e9",
          2383 => x"75",
          2384 => x"2e",
          2385 => x"d5",
          2386 => x"94",
          2387 => x"29",
          2388 => x"16",
          2389 => x"84",
          2390 => x"83",
          2391 => x"5a",
          2392 => x"18",
          2393 => x"29",
          2394 => x"86",
          2395 => x"d8",
          2396 => x"92",
          2397 => x"29",
          2398 => x"f8",
          2399 => x"81",
          2400 => x"73",
          2401 => x"d9",
          2402 => x"17",
          2403 => x"b6",
          2404 => x"38",
          2405 => x"2e",
          2406 => x"e4",
          2407 => x"2e",
          2408 => x"38",
          2409 => x"c1",
          2410 => x"3f",
          2411 => x"be",
          2412 => x"84",
          2413 => x"89",
          2414 => x"80",
          2415 => x"3f",
          2416 => x"54",
          2417 => x"52",
          2418 => x"70",
          2419 => x"27",
          2420 => x"f8",
          2421 => x"83",
          2422 => x"b8",
          2423 => x"80",
          2424 => x"38",
          2425 => x"06",
          2426 => x"73",
          2427 => x"52",
          2428 => x"95",
          2429 => x"05",
          2430 => x"72",
          2431 => x"80",
          2432 => x"81",
          2433 => x"80",
          2434 => x"86",
          2435 => x"05",
          2436 => x"75",
          2437 => x"2e",
          2438 => x"b5",
          2439 => x"78",
          2440 => x"2e",
          2441 => x"83",
          2442 => x"72",
          2443 => x"b6",
          2444 => x"17",
          2445 => x"95",
          2446 => x"29",
          2447 => x"f8",
          2448 => x"60",
          2449 => x"f8",
          2450 => x"05",
          2451 => x"ff",
          2452 => x"95",
          2453 => x"5d",
          2454 => x"97",
          2455 => x"ff",
          2456 => x"b8",
          2457 => x"86",
          2458 => x"f8",
          2459 => x"0c",
          2460 => x"84",
          2461 => x"38",
          2462 => x"80",
          2463 => x"84",
          2464 => x"83",
          2465 => x"72",
          2466 => x"b6",
          2467 => x"1d",
          2468 => x"95",
          2469 => x"29",
          2470 => x"f8",
          2471 => x"76",
          2472 => x"90",
          2473 => x"84",
          2474 => x"83",
          2475 => x"72",
          2476 => x"59",
          2477 => x"b6",
          2478 => x"ff",
          2479 => x"38",
          2480 => x"84",
          2481 => x"78",
          2482 => x"24",
          2483 => x"81",
          2484 => x"f8",
          2485 => x"0c",
          2486 => x"82",
          2487 => x"26",
          2488 => x"81",
          2489 => x"34",
          2490 => x"81",
          2491 => x"e8",
          2492 => x"0c",
          2493 => x"fd",
          2494 => x"0c",
          2495 => x"33",
          2496 => x"05",
          2497 => x"33",
          2498 => x"b6",
          2499 => x"f8",
          2500 => x"5f",
          2501 => x"34",
          2502 => x"19",
          2503 => x"a7",
          2504 => x"33",
          2505 => x"22",
          2506 => x"11",
          2507 => x"90",
          2508 => x"81",
          2509 => x"81",
          2510 => x"f8",
          2511 => x"d8",
          2512 => x"ff",
          2513 => x"29",
          2514 => x"f8",
          2515 => x"29",
          2516 => x"f6",
          2517 => x"75",
          2518 => x"ff",
          2519 => x"95",
          2520 => x"34",
          2521 => x"e4",
          2522 => x"80",
          2523 => x"84",
          2524 => x"e0",
          2525 => x"9c",
          2526 => x"84",
          2527 => x"84",
          2528 => x"84",
          2529 => x"e0",
          2530 => x"9c",
          2531 => x"09",
          2532 => x"94",
          2533 => x"ff",
          2534 => x"ff",
          2535 => x"a0",
          2536 => x"40",
          2537 => x"ff",
          2538 => x"43",
          2539 => x"85",
          2540 => x"1a",
          2541 => x"76",
          2542 => x"06",
          2543 => x"06",
          2544 => x"84",
          2545 => x"1e",
          2546 => x"95",
          2547 => x"29",
          2548 => x"83",
          2549 => x"33",
          2550 => x"83",
          2551 => x"1a",
          2552 => x"ff",
          2553 => x"95",
          2554 => x"5a",
          2555 => x"84",
          2556 => x"81",
          2557 => x"95",
          2558 => x"79",
          2559 => x"83",
          2560 => x"70",
          2561 => x"fd",
          2562 => x"38",
          2563 => x"bf",
          2564 => x"33",
          2565 => x"19",
          2566 => x"75",
          2567 => x"77",
          2568 => x"34",
          2569 => x"80",
          2570 => x"0d",
          2571 => x"d8",
          2572 => x"95",
          2573 => x"29",
          2574 => x"f8",
          2575 => x"05",
          2576 => x"ea",
          2577 => x"5b",
          2578 => x"5c",
          2579 => x"06",
          2580 => x"05",
          2581 => x"86",
          2582 => x"d8",
          2583 => x"92",
          2584 => x"5e",
          2585 => x"34",
          2586 => x"1e",
          2587 => x"a7",
          2588 => x"33",
          2589 => x"22",
          2590 => x"11",
          2591 => x"90",
          2592 => x"81",
          2593 => x"7e",
          2594 => x"d9",
          2595 => x"19",
          2596 => x"1c",
          2597 => x"83",
          2598 => x"33",
          2599 => x"33",
          2600 => x"06",
          2601 => x"05",
          2602 => x"b7",
          2603 => x"34",
          2604 => x"33",
          2605 => x"12",
          2606 => x"f8",
          2607 => x"76",
          2608 => x"90",
          2609 => x"84",
          2610 => x"83",
          2611 => x"72",
          2612 => x"59",
          2613 => x"18",
          2614 => x"06",
          2615 => x"38",
          2616 => x"39",
          2617 => x"0b",
          2618 => x"04",
          2619 => x"b6",
          2620 => x"95",
          2621 => x"05",
          2622 => x"b7",
          2623 => x"0c",
          2624 => x"17",
          2625 => x"7c",
          2626 => x"d8",
          2627 => x"5b",
          2628 => x"e8",
          2629 => x"05",
          2630 => x"e4",
          2631 => x"b7",
          2632 => x"84",
          2633 => x"06",
          2634 => x"84",
          2635 => x"83",
          2636 => x"e0",
          2637 => x"33",
          2638 => x"33",
          2639 => x"b6",
          2640 => x"f8",
          2641 => x"5d",
          2642 => x"86",
          2643 => x"d8",
          2644 => x"92",
          2645 => x"5b",
          2646 => x"83",
          2647 => x"41",
          2648 => x"a7",
          2649 => x"33",
          2650 => x"22",
          2651 => x"11",
          2652 => x"90",
          2653 => x"1c",
          2654 => x"7b",
          2655 => x"33",
          2656 => x"56",
          2657 => x"84",
          2658 => x"40",
          2659 => x"b6",
          2660 => x"78",
          2661 => x"0b",
          2662 => x"04",
          2663 => x"34",
          2664 => x"34",
          2665 => x"f8",
          2666 => x"94",
          2667 => x"95",
          2668 => x"93",
          2669 => x"39",
          2670 => x"2e",
          2671 => x"5d",
          2672 => x"85",
          2673 => x"55",
          2674 => x"9b",
          2675 => x"70",
          2676 => x"51",
          2677 => x"08",
          2678 => x"57",
          2679 => x"cd",
          2680 => x"fe",
          2681 => x"0b",
          2682 => x"81",
          2683 => x"ad",
          2684 => x"81",
          2685 => x"8a",
          2686 => x"94",
          2687 => x"e5",
          2688 => x"38",
          2689 => x"33",
          2690 => x"2c",
          2691 => x"75",
          2692 => x"84",
          2693 => x"8e",
          2694 => x"05",
          2695 => x"33",
          2696 => x"c5",
          2697 => x"bd",
          2698 => x"83",
          2699 => x"5d",
          2700 => x"ff",
          2701 => x"fd",
          2702 => x"34",
          2703 => x"33",
          2704 => x"fd",
          2705 => x"f8",
          2706 => x"e5",
          2707 => x"38",
          2708 => x"33",
          2709 => x"2c",
          2710 => x"75",
          2711 => x"84",
          2712 => x"fc",
          2713 => x"60",
          2714 => x"38",
          2715 => x"33",
          2716 => x"12",
          2717 => x"92",
          2718 => x"29",
          2719 => x"f6",
          2720 => x"42",
          2721 => x"2e",
          2722 => x"e9",
          2723 => x"33",
          2724 => x"84",
          2725 => x"09",
          2726 => x"83",
          2727 => x"b7",
          2728 => x"be",
          2729 => x"95",
          2730 => x"33",
          2731 => x"25",
          2732 => x"95",
          2733 => x"33",
          2734 => x"84",
          2735 => x"42",
          2736 => x"11",
          2737 => x"38",
          2738 => x"fa",
          2739 => x"e8",
          2740 => x"33",
          2741 => x"38",
          2742 => x"22",
          2743 => x"e8",
          2744 => x"06",
          2745 => x"da",
          2746 => x"5f",
          2747 => x"b8",
          2748 => x"38",
          2749 => x"06",
          2750 => x"84",
          2751 => x"8e",
          2752 => x"05",
          2753 => x"33",
          2754 => x"b6",
          2755 => x"11",
          2756 => x"77",
          2757 => x"83",
          2758 => x"ff",
          2759 => x"38",
          2760 => x"84",
          2761 => x"7a",
          2762 => x"75",
          2763 => x"84",
          2764 => x"8a",
          2765 => x"b6",
          2766 => x"f9",
          2767 => x"b6",
          2768 => x"f8",
          2769 => x"a7",
          2770 => x"5f",
          2771 => x"ff",
          2772 => x"52",
          2773 => x"84",
          2774 => x"70",
          2775 => x"8e",
          2776 => x"76",
          2777 => x"56",
          2778 => x"ff",
          2779 => x"60",
          2780 => x"33",
          2781 => x"ff",
          2782 => x"7e",
          2783 => x"57",
          2784 => x"38",
          2785 => x"ff",
          2786 => x"79",
          2787 => x"a7",
          2788 => x"81",
          2789 => x"58",
          2790 => x"38",
          2791 => x"17",
          2792 => x"7b",
          2793 => x"81",
          2794 => x"5e",
          2795 => x"84",
          2796 => x"43",
          2797 => x"9d",
          2798 => x"b6",
          2799 => x"5d",
          2800 => x"7c",
          2801 => x"84",
          2802 => x"71",
          2803 => x"7f",
          2804 => x"39",
          2805 => x"2e",
          2806 => x"b9",
          2807 => x"39",
          2808 => x"11",
          2809 => x"58",
          2810 => x"b8",
          2811 => x"06",
          2812 => x"58",
          2813 => x"33",
          2814 => x"81",
          2815 => x"7a",
          2816 => x"ff",
          2817 => x"38",
          2818 => x"57",
          2819 => x"1b",
          2820 => x"a0",
          2821 => x"a7",
          2822 => x"51",
          2823 => x"06",
          2824 => x"90",
          2825 => x"07",
          2826 => x"7f",
          2827 => x"9e",
          2828 => x"0c",
          2829 => x"79",
          2830 => x"33",
          2831 => x"81",
          2832 => x"f8",
          2833 => x"59",
          2834 => x"38",
          2835 => x"62",
          2836 => x"57",
          2837 => x"f8",
          2838 => x"5a",
          2839 => x"78",
          2840 => x"57",
          2841 => x"0b",
          2842 => x"81",
          2843 => x"77",
          2844 => x"1f",
          2845 => x"8a",
          2846 => x"f0",
          2847 => x"71",
          2848 => x"80",
          2849 => x"80",
          2850 => x"18",
          2851 => x"b6",
          2852 => x"84",
          2853 => x"f8",
          2854 => x"f8",
          2855 => x"5c",
          2856 => x"90",
          2857 => x"90",
          2858 => x"59",
          2859 => x"33",
          2860 => x"83",
          2861 => x"90",
          2862 => x"75",
          2863 => x"f8",
          2864 => x"56",
          2865 => x"83",
          2866 => x"07",
          2867 => x"b1",
          2868 => x"34",
          2869 => x"56",
          2870 => x"81",
          2871 => x"34",
          2872 => x"81",
          2873 => x"f8",
          2874 => x"90",
          2875 => x"56",
          2876 => x"39",
          2877 => x"80",
          2878 => x"34",
          2879 => x"81",
          2880 => x"f8",
          2881 => x"90",
          2882 => x"75",
          2883 => x"83",
          2884 => x"07",
          2885 => x"a1",
          2886 => x"06",
          2887 => x"34",
          2888 => x"81",
          2889 => x"34",
          2890 => x"80",
          2891 => x"34",
          2892 => x"80",
          2893 => x"34",
          2894 => x"81",
          2895 => x"83",
          2896 => x"f8",
          2897 => x"56",
          2898 => x"39",
          2899 => x"52",
          2900 => x"39",
          2901 => x"34",
          2902 => x"34",
          2903 => x"f8",
          2904 => x"0c",
          2905 => x"e7",
          2906 => x"9c",
          2907 => x"34",
          2908 => x"06",
          2909 => x"84",
          2910 => x"53",
          2911 => x"84",
          2912 => x"e4",
          2913 => x"84",
          2914 => x"e4",
          2915 => x"f8",
          2916 => x"e5",
          2917 => x"b7",
          2918 => x"5d",
          2919 => x"b8",
          2920 => x"34",
          2921 => x"34",
          2922 => x"83",
          2923 => x"58",
          2924 => x"0b",
          2925 => x"51",
          2926 => x"51",
          2927 => x"83",
          2928 => x"70",
          2929 => x"f2",
          2930 => x"39",
          2931 => x"27",
          2932 => x"34",
          2933 => x"ff",
          2934 => x"06",
          2935 => x"f8",
          2936 => x"33",
          2937 => x"25",
          2938 => x"39",
          2939 => x"06",
          2940 => x"38",
          2941 => x"33",
          2942 => x"33",
          2943 => x"80",
          2944 => x"71",
          2945 => x"06",
          2946 => x"42",
          2947 => x"38",
          2948 => x"5c",
          2949 => x"84",
          2950 => x"83",
          2951 => x"f8",
          2952 => x"11",
          2953 => x"38",
          2954 => x"27",
          2955 => x"83",
          2956 => x"83",
          2957 => x"76",
          2958 => x"81",
          2959 => x"29",
          2960 => x"a0",
          2961 => x"81",
          2962 => x"71",
          2963 => x"7e",
          2964 => x"1a",
          2965 => x"b6",
          2966 => x"5d",
          2967 => x"7d",
          2968 => x"84",
          2969 => x"71",
          2970 => x"77",
          2971 => x"17",
          2972 => x"7b",
          2973 => x"81",
          2974 => x"5f",
          2975 => x"84",
          2976 => x"59",
          2977 => x"99",
          2978 => x"17",
          2979 => x"7b",
          2980 => x"d8",
          2981 => x"d7",
          2982 => x"39",
          2983 => x"33",
          2984 => x"42",
          2985 => x"5a",
          2986 => x"ff",
          2987 => x"27",
          2988 => x"94",
          2989 => x"ff",
          2990 => x"78",
          2991 => x"83",
          2992 => x"f8",
          2993 => x"33",
          2994 => x"25",
          2995 => x"39",
          2996 => x"c0",
          2997 => x"ff",
          2998 => x"5d",
          2999 => x"06",
          3000 => x"1d",
          3001 => x"93",
          3002 => x"92",
          3003 => x"56",
          3004 => x"39",
          3005 => x"f5",
          3006 => x"58",
          3007 => x"81",
          3008 => x"ec",
          3009 => x"34",
          3010 => x"05",
          3011 => x"f4",
          3012 => x"83",
          3013 => x"0b",
          3014 => x"7e",
          3015 => x"80",
          3016 => x"39",
          3017 => x"a7",
          3018 => x"84",
          3019 => x"0b",
          3020 => x"fd",
          3021 => x"b6",
          3022 => x"90",
          3023 => x"0b",
          3024 => x"04",
          3025 => x"80",
          3026 => x"0d",
          3027 => x"33",
          3028 => x"70",
          3029 => x"33",
          3030 => x"80",
          3031 => x"f6",
          3032 => x"e4",
          3033 => x"c4",
          3034 => x"91",
          3035 => x"07",
          3036 => x"5e",
          3037 => x"59",
          3038 => x"06",
          3039 => x"70",
          3040 => x"5c",
          3041 => x"84",
          3042 => x"83",
          3043 => x"86",
          3044 => x"22",
          3045 => x"70",
          3046 => x"33",
          3047 => x"83",
          3048 => x"ee",
          3049 => x"98",
          3050 => x"56",
          3051 => x"80",
          3052 => x"15",
          3053 => x"55",
          3054 => x"80",
          3055 => x"81",
          3056 => x"58",
          3057 => x"38",
          3058 => x"74",
          3059 => x"ff",
          3060 => x"cd",
          3061 => x"83",
          3062 => x"15",
          3063 => x"55",
          3064 => x"83",
          3065 => x"80",
          3066 => x"bc",
          3067 => x"2a",
          3068 => x"58",
          3069 => x"0b",
          3070 => x"06",
          3071 => x"81",
          3072 => x"83",
          3073 => x"83",
          3074 => x"33",
          3075 => x"5e",
          3076 => x"33",
          3077 => x"83",
          3078 => x"2e",
          3079 => x"33",
          3080 => x"83",
          3081 => x"ec",
          3082 => x"81",
          3083 => x"16",
          3084 => x"38",
          3085 => x"ff",
          3086 => x"16",
          3087 => x"38",
          3088 => x"87",
          3089 => x"73",
          3090 => x"c0",
          3091 => x"58",
          3092 => x"54",
          3093 => x"83",
          3094 => x"34",
          3095 => x"82",
          3096 => x"dc",
          3097 => x"ec",
          3098 => x"83",
          3099 => x"5e",
          3100 => x"80",
          3101 => x"72",
          3102 => x"83",
          3103 => x"08",
          3104 => x"06",
          3105 => x"f8",
          3106 => x"14",
          3107 => x"a5",
          3108 => x"80",
          3109 => x"83",
          3110 => x"f0",
          3111 => x"e0",
          3112 => x"7c",
          3113 => x"09",
          3114 => x"2e",
          3115 => x"d7",
          3116 => x"77",
          3117 => x"80",
          3118 => x"38",
          3119 => x"10",
          3120 => x"98",
          3121 => x"73",
          3122 => x"79",
          3123 => x"05",
          3124 => x"56",
          3125 => x"83",
          3126 => x"80",
          3127 => x"79",
          3128 => x"82",
          3129 => x"fa",
          3130 => x"33",
          3131 => x"38",
          3132 => x"25",
          3133 => x"38",
          3134 => x"cc",
          3135 => x"80",
          3136 => x"f0",
          3137 => x"2e",
          3138 => x"ff",
          3139 => x"38",
          3140 => x"2e",
          3141 => x"55",
          3142 => x"06",
          3143 => x"84",
          3144 => x"be",
          3145 => x"39",
          3146 => x"f6",
          3147 => x"83",
          3148 => x"80",
          3149 => x"0b",
          3150 => x"83",
          3151 => x"74",
          3152 => x"2e",
          3153 => x"33",
          3154 => x"77",
          3155 => x"09",
          3156 => x"b8",
          3157 => x"9c",
          3158 => x"e8",
          3159 => x"f6",
          3160 => x"fb",
          3161 => x"15",
          3162 => x"bd",
          3163 => x"fa",
          3164 => x"80",
          3165 => x"c4",
          3166 => x"f6",
          3167 => x"5d",
          3168 => x"39",
          3169 => x"cb",
          3170 => x"ce",
          3171 => x"fc",
          3172 => x"34",
          3173 => x"0b",
          3174 => x"83",
          3175 => x"34",
          3176 => x"84",
          3177 => x"38",
          3178 => x"ff",
          3179 => x"f6",
          3180 => x"84",
          3181 => x"39",
          3182 => x"06",
          3183 => x"27",
          3184 => x"92",
          3185 => x"55",
          3186 => x"54",
          3187 => x"d8",
          3188 => x"05",
          3189 => x"53",
          3190 => x"f6",
          3191 => x"ba",
          3192 => x"72",
          3193 => x"52",
          3194 => x"3f",
          3195 => x"f6",
          3196 => x"3d",
          3197 => x"3d",
          3198 => x"83",
          3199 => x"05",
          3200 => x"08",
          3201 => x"83",
          3202 => x"81",
          3203 => x"e8",
          3204 => x"f2",
          3205 => x"53",
          3206 => x"c0",
          3207 => x"f6",
          3208 => x"9c",
          3209 => x"38",
          3210 => x"c0",
          3211 => x"73",
          3212 => x"ff",
          3213 => x"9c",
          3214 => x"c0",
          3215 => x"9c",
          3216 => x"81",
          3217 => x"52",
          3218 => x"81",
          3219 => x"a4",
          3220 => x"ff",
          3221 => x"ff",
          3222 => x"38",
          3223 => x"d5",
          3224 => x"84",
          3225 => x"81",
          3226 => x"0d",
          3227 => x"05",
          3228 => x"83",
          3229 => x"fc",
          3230 => x"07",
          3231 => x"34",
          3232 => x"34",
          3233 => x"34",
          3234 => x"08",
          3235 => x"f0",
          3236 => x"0b",
          3237 => x"0b",
          3238 => x"80",
          3239 => x"83",
          3240 => x"05",
          3241 => x"87",
          3242 => x"2e",
          3243 => x"98",
          3244 => x"87",
          3245 => x"87",
          3246 => x"70",
          3247 => x"71",
          3248 => x"98",
          3249 => x"87",
          3250 => x"98",
          3251 => x"38",
          3252 => x"08",
          3253 => x"71",
          3254 => x"98",
          3255 => x"38",
          3256 => x"81",
          3257 => x"80",
          3258 => x"71",
          3259 => x"ff",
          3260 => x"14",
          3261 => x"70",
          3262 => x"05",
          3263 => x"34",
          3264 => x"b8",
          3265 => x"0b",
          3266 => x"04",
          3267 => x"79",
          3268 => x"56",
          3269 => x"88",
          3270 => x"79",
          3271 => x"75",
          3272 => x"70",
          3273 => x"71",
          3274 => x"7a",
          3275 => x"84",
          3276 => x"73",
          3277 => x"52",
          3278 => x"72",
          3279 => x"08",
          3280 => x"f0",
          3281 => x"0b",
          3282 => x"0b",
          3283 => x"80",
          3284 => x"83",
          3285 => x"05",
          3286 => x"87",
          3287 => x"2e",
          3288 => x"98",
          3289 => x"87",
          3290 => x"87",
          3291 => x"70",
          3292 => x"71",
          3293 => x"98",
          3294 => x"87",
          3295 => x"98",
          3296 => x"38",
          3297 => x"08",
          3298 => x"71",
          3299 => x"98",
          3300 => x"38",
          3301 => x"81",
          3302 => x"a1",
          3303 => x"fe",
          3304 => x"06",
          3305 => x"57",
          3306 => x"0d",
          3307 => x"0d",
          3308 => x"71",
          3309 => x"56",
          3310 => x"0b",
          3311 => x"98",
          3312 => x"80",
          3313 => x"9c",
          3314 => x"53",
          3315 => x"33",
          3316 => x"70",
          3317 => x"2e",
          3318 => x"51",
          3319 => x"38",
          3320 => x"38",
          3321 => x"90",
          3322 => x"52",
          3323 => x"72",
          3324 => x"c0",
          3325 => x"27",
          3326 => x"38",
          3327 => x"71",
          3328 => x"ff",
          3329 => x"75",
          3330 => x"06",
          3331 => x"80",
          3332 => x"d0",
          3333 => x"3d",
          3334 => x"31",
          3335 => x"70",
          3336 => x"12",
          3337 => x"07",
          3338 => x"71",
          3339 => x"54",
          3340 => x"56",
          3341 => x"38",
          3342 => x"33",
          3343 => x"76",
          3344 => x"98",
          3345 => x"5c",
          3346 => x"83",
          3347 => x"33",
          3348 => x"75",
          3349 => x"57",
          3350 => x"06",
          3351 => x"d4",
          3352 => x"13",
          3353 => x"2a",
          3354 => x"14",
          3355 => x"d4",
          3356 => x"34",
          3357 => x"d4",
          3358 => x"85",
          3359 => x"70",
          3360 => x"07",
          3361 => x"58",
          3362 => x"81",
          3363 => x"12",
          3364 => x"71",
          3365 => x"33",
          3366 => x"70",
          3367 => x"58",
          3368 => x"12",
          3369 => x"84",
          3370 => x"2b",
          3371 => x"52",
          3372 => x"33",
          3373 => x"52",
          3374 => x"72",
          3375 => x"15",
          3376 => x"2b",
          3377 => x"2a",
          3378 => x"77",
          3379 => x"70",
          3380 => x"8b",
          3381 => x"70",
          3382 => x"07",
          3383 => x"77",
          3384 => x"54",
          3385 => x"14",
          3386 => x"d4",
          3387 => x"33",
          3388 => x"74",
          3389 => x"88",
          3390 => x"88",
          3391 => x"54",
          3392 => x"34",
          3393 => x"11",
          3394 => x"71",
          3395 => x"81",
          3396 => x"2b",
          3397 => x"53",
          3398 => x"71",
          3399 => x"07",
          3400 => x"59",
          3401 => x"16",
          3402 => x"70",
          3403 => x"71",
          3404 => x"33",
          3405 => x"70",
          3406 => x"56",
          3407 => x"83",
          3408 => x"3d",
          3409 => x"58",
          3410 => x"2e",
          3411 => x"89",
          3412 => x"84",
          3413 => x"b8",
          3414 => x"52",
          3415 => x"3f",
          3416 => x"34",
          3417 => x"d4",
          3418 => x"0b",
          3419 => x"56",
          3420 => x"17",
          3421 => x"d0",
          3422 => x"70",
          3423 => x"58",
          3424 => x"73",
          3425 => x"70",
          3426 => x"05",
          3427 => x"34",
          3428 => x"39",
          3429 => x"81",
          3430 => x"12",
          3431 => x"ff",
          3432 => x"06",
          3433 => x"85",
          3434 => x"52",
          3435 => x"54",
          3436 => x"10",
          3437 => x"33",
          3438 => x"ff",
          3439 => x"06",
          3440 => x"54",
          3441 => x"80",
          3442 => x"84",
          3443 => x"2b",
          3444 => x"81",
          3445 => x"54",
          3446 => x"70",
          3447 => x"07",
          3448 => x"5d",
          3449 => x"38",
          3450 => x"82",
          3451 => x"82",
          3452 => x"38",
          3453 => x"74",
          3454 => x"5b",
          3455 => x"78",
          3456 => x"15",
          3457 => x"14",
          3458 => x"d4",
          3459 => x"33",
          3460 => x"8f",
          3461 => x"ff",
          3462 => x"53",
          3463 => x"34",
          3464 => x"12",
          3465 => x"75",
          3466 => x"b8",
          3467 => x"87",
          3468 => x"2b",
          3469 => x"57",
          3470 => x"34",
          3471 => x"78",
          3472 => x"71",
          3473 => x"54",
          3474 => x"87",
          3475 => x"19",
          3476 => x"8b",
          3477 => x"58",
          3478 => x"34",
          3479 => x"08",
          3480 => x"33",
          3481 => x"70",
          3482 => x"84",
          3483 => x"b8",
          3484 => x"84",
          3485 => x"86",
          3486 => x"2b",
          3487 => x"17",
          3488 => x"07",
          3489 => x"54",
          3490 => x"12",
          3491 => x"84",
          3492 => x"2b",
          3493 => x"14",
          3494 => x"07",
          3495 => x"56",
          3496 => x"76",
          3497 => x"18",
          3498 => x"2b",
          3499 => x"2a",
          3500 => x"74",
          3501 => x"18",
          3502 => x"3d",
          3503 => x"58",
          3504 => x"77",
          3505 => x"89",
          3506 => x"3f",
          3507 => x"0c",
          3508 => x"0b",
          3509 => x"84",
          3510 => x"76",
          3511 => x"c5",
          3512 => x"75",
          3513 => x"b8",
          3514 => x"81",
          3515 => x"08",
          3516 => x"87",
          3517 => x"b8",
          3518 => x"07",
          3519 => x"2a",
          3520 => x"34",
          3521 => x"22",
          3522 => x"08",
          3523 => x"15",
          3524 => x"54",
          3525 => x"e3",
          3526 => x"5f",
          3527 => x"45",
          3528 => x"7e",
          3529 => x"2e",
          3530 => x"27",
          3531 => x"82",
          3532 => x"58",
          3533 => x"31",
          3534 => x"70",
          3535 => x"12",
          3536 => x"31",
          3537 => x"10",
          3538 => x"11",
          3539 => x"2b",
          3540 => x"53",
          3541 => x"44",
          3542 => x"80",
          3543 => x"33",
          3544 => x"70",
          3545 => x"12",
          3546 => x"07",
          3547 => x"74",
          3548 => x"82",
          3549 => x"2e",
          3550 => x"f9",
          3551 => x"87",
          3552 => x"24",
          3553 => x"81",
          3554 => x"2b",
          3555 => x"33",
          3556 => x"47",
          3557 => x"80",
          3558 => x"82",
          3559 => x"2b",
          3560 => x"11",
          3561 => x"71",
          3562 => x"33",
          3563 => x"70",
          3564 => x"41",
          3565 => x"1d",
          3566 => x"d4",
          3567 => x"12",
          3568 => x"07",
          3569 => x"33",
          3570 => x"5f",
          3571 => x"77",
          3572 => x"84",
          3573 => x"12",
          3574 => x"ff",
          3575 => x"59",
          3576 => x"84",
          3577 => x"33",
          3578 => x"83",
          3579 => x"15",
          3580 => x"2a",
          3581 => x"55",
          3582 => x"84",
          3583 => x"81",
          3584 => x"2b",
          3585 => x"15",
          3586 => x"2a",
          3587 => x"55",
          3588 => x"34",
          3589 => x"11",
          3590 => x"07",
          3591 => x"42",
          3592 => x"51",
          3593 => x"08",
          3594 => x"70",
          3595 => x"7a",
          3596 => x"73",
          3597 => x"04",
          3598 => x"0c",
          3599 => x"82",
          3600 => x"f4",
          3601 => x"d4",
          3602 => x"81",
          3603 => x"60",
          3604 => x"34",
          3605 => x"1d",
          3606 => x"b8",
          3607 => x"05",
          3608 => x"ff",
          3609 => x"57",
          3610 => x"34",
          3611 => x"10",
          3612 => x"55",
          3613 => x"83",
          3614 => x"7e",
          3615 => x"8c",
          3616 => x"df",
          3617 => x"b8",
          3618 => x"3d",
          3619 => x"08",
          3620 => x"7f",
          3621 => x"88",
          3622 => x"88",
          3623 => x"7b",
          3624 => x"b8",
          3625 => x"58",
          3626 => x"34",
          3627 => x"33",
          3628 => x"70",
          3629 => x"05",
          3630 => x"2a",
          3631 => x"63",
          3632 => x"06",
          3633 => x"b8",
          3634 => x"60",
          3635 => x"08",
          3636 => x"7e",
          3637 => x"70",
          3638 => x"ac",
          3639 => x"31",
          3640 => x"33",
          3641 => x"70",
          3642 => x"12",
          3643 => x"07",
          3644 => x"54",
          3645 => x"bc",
          3646 => x"80",
          3647 => x"ff",
          3648 => x"dd",
          3649 => x"0b",
          3650 => x"84",
          3651 => x"7e",
          3652 => x"dd",
          3653 => x"7a",
          3654 => x"b8",
          3655 => x"81",
          3656 => x"08",
          3657 => x"87",
          3658 => x"b8",
          3659 => x"07",
          3660 => x"2a",
          3661 => x"05",
          3662 => x"b8",
          3663 => x"b8",
          3664 => x"7e",
          3665 => x"05",
          3666 => x"83",
          3667 => x"5b",
          3668 => x"f2",
          3669 => x"7e",
          3670 => x"84",
          3671 => x"76",
          3672 => x"71",
          3673 => x"11",
          3674 => x"8b",
          3675 => x"84",
          3676 => x"2b",
          3677 => x"56",
          3678 => x"78",
          3679 => x"05",
          3680 => x"84",
          3681 => x"2b",
          3682 => x"14",
          3683 => x"07",
          3684 => x"5d",
          3685 => x"34",
          3686 => x"d4",
          3687 => x"71",
          3688 => x"70",
          3689 => x"7d",
          3690 => x"d4",
          3691 => x"12",
          3692 => x"07",
          3693 => x"71",
          3694 => x"5c",
          3695 => x"7c",
          3696 => x"d4",
          3697 => x"33",
          3698 => x"74",
          3699 => x"71",
          3700 => x"47",
          3701 => x"82",
          3702 => x"b8",
          3703 => x"83",
          3704 => x"57",
          3705 => x"58",
          3706 => x"bd",
          3707 => x"84",
          3708 => x"5f",
          3709 => x"84",
          3710 => x"b8",
          3711 => x"52",
          3712 => x"3f",
          3713 => x"34",
          3714 => x"d4",
          3715 => x"0b",
          3716 => x"54",
          3717 => x"15",
          3718 => x"d0",
          3719 => x"70",
          3720 => x"45",
          3721 => x"60",
          3722 => x"70",
          3723 => x"05",
          3724 => x"34",
          3725 => x"e7",
          3726 => x"86",
          3727 => x"2b",
          3728 => x"1c",
          3729 => x"07",
          3730 => x"59",
          3731 => x"61",
          3732 => x"70",
          3733 => x"71",
          3734 => x"05",
          3735 => x"88",
          3736 => x"48",
          3737 => x"86",
          3738 => x"84",
          3739 => x"12",
          3740 => x"ff",
          3741 => x"58",
          3742 => x"84",
          3743 => x"81",
          3744 => x"2b",
          3745 => x"33",
          3746 => x"8f",
          3747 => x"2a",
          3748 => x"44",
          3749 => x"17",
          3750 => x"70",
          3751 => x"71",
          3752 => x"81",
          3753 => x"ff",
          3754 => x"5e",
          3755 => x"34",
          3756 => x"ff",
          3757 => x"15",
          3758 => x"71",
          3759 => x"33",
          3760 => x"70",
          3761 => x"5d",
          3762 => x"34",
          3763 => x"11",
          3764 => x"71",
          3765 => x"33",
          3766 => x"70",
          3767 => x"42",
          3768 => x"75",
          3769 => x"08",
          3770 => x"88",
          3771 => x"88",
          3772 => x"34",
          3773 => x"08",
          3774 => x"71",
          3775 => x"05",
          3776 => x"2b",
          3777 => x"06",
          3778 => x"5f",
          3779 => x"82",
          3780 => x"b8",
          3781 => x"12",
          3782 => x"07",
          3783 => x"71",
          3784 => x"70",
          3785 => x"59",
          3786 => x"1d",
          3787 => x"82",
          3788 => x"2b",
          3789 => x"11",
          3790 => x"71",
          3791 => x"33",
          3792 => x"70",
          3793 => x"42",
          3794 => x"84",
          3795 => x"b8",
          3796 => x"85",
          3797 => x"2b",
          3798 => x"15",
          3799 => x"2a",
          3800 => x"57",
          3801 => x"34",
          3802 => x"81",
          3803 => x"ff",
          3804 => x"5e",
          3805 => x"34",
          3806 => x"11",
          3807 => x"71",
          3808 => x"81",
          3809 => x"88",
          3810 => x"55",
          3811 => x"34",
          3812 => x"33",
          3813 => x"83",
          3814 => x"83",
          3815 => x"88",
          3816 => x"55",
          3817 => x"1a",
          3818 => x"82",
          3819 => x"2b",
          3820 => x"2b",
          3821 => x"05",
          3822 => x"d4",
          3823 => x"1c",
          3824 => x"5f",
          3825 => x"1a",
          3826 => x"07",
          3827 => x"33",
          3828 => x"40",
          3829 => x"84",
          3830 => x"84",
          3831 => x"33",
          3832 => x"83",
          3833 => x"87",
          3834 => x"88",
          3835 => x"41",
          3836 => x"64",
          3837 => x"1d",
          3838 => x"2b",
          3839 => x"2a",
          3840 => x"7c",
          3841 => x"70",
          3842 => x"8b",
          3843 => x"70",
          3844 => x"07",
          3845 => x"77",
          3846 => x"49",
          3847 => x"1e",
          3848 => x"d4",
          3849 => x"33",
          3850 => x"74",
          3851 => x"88",
          3852 => x"88",
          3853 => x"5e",
          3854 => x"34",
          3855 => x"83",
          3856 => x"3f",
          3857 => x"e4",
          3858 => x"73",
          3859 => x"b5",
          3860 => x"61",
          3861 => x"f0",
          3862 => x"29",
          3863 => x"80",
          3864 => x"38",
          3865 => x"0d",
          3866 => x"b8",
          3867 => x"80",
          3868 => x"84",
          3869 => x"3f",
          3870 => x"0d",
          3871 => x"d4",
          3872 => x"23",
          3873 => x"ff",
          3874 => x"b8",
          3875 => x"0b",
          3876 => x"54",
          3877 => x"15",
          3878 => x"86",
          3879 => x"84",
          3880 => x"ff",
          3881 => x"ff",
          3882 => x"55",
          3883 => x"17",
          3884 => x"10",
          3885 => x"05",
          3886 => x"0b",
          3887 => x"2e",
          3888 => x"3d",
          3889 => x"52",
          3890 => x"e0",
          3891 => x"0c",
          3892 => x"02",
          3893 => x"81",
          3894 => x"3f",
          3895 => x"53",
          3896 => x"13",
          3897 => x"72",
          3898 => x"04",
          3899 => x"8c",
          3900 => x"59",
          3901 => x"84",
          3902 => x"06",
          3903 => x"58",
          3904 => x"78",
          3905 => x"3f",
          3906 => x"55",
          3907 => x"98",
          3908 => x"78",
          3909 => x"06",
          3910 => x"54",
          3911 => x"8b",
          3912 => x"19",
          3913 => x"79",
          3914 => x"f7",
          3915 => x"05",
          3916 => x"81",
          3917 => x"b8",
          3918 => x"54",
          3919 => x"85",
          3920 => x"53",
          3921 => x"84",
          3922 => x"74",
          3923 => x"8c",
          3924 => x"26",
          3925 => x"54",
          3926 => x"73",
          3927 => x"3d",
          3928 => x"70",
          3929 => x"78",
          3930 => x"3d",
          3931 => x"33",
          3932 => x"53",
          3933 => x"38",
          3934 => x"81",
          3935 => x"85",
          3936 => x"53",
          3937 => x"25",
          3938 => x"84",
          3939 => x"3d",
          3940 => x"73",
          3941 => x"04",
          3942 => x"b8",
          3943 => x"84",
          3944 => x"54",
          3945 => x"2a",
          3946 => x"8a",
          3947 => x"74",
          3948 => x"51",
          3949 => x"c0",
          3950 => x"06",
          3951 => x"71",
          3952 => x"ff",
          3953 => x"80",
          3954 => x"57",
          3955 => x"38",
          3956 => x"87",
          3957 => x"33",
          3958 => x"08",
          3959 => x"84",
          3960 => x"81",
          3961 => x"70",
          3962 => x"ff",
          3963 => x"77",
          3964 => x"b8",
          3965 => x"08",
          3966 => x"08",
          3967 => x"5b",
          3968 => x"18",
          3969 => x"06",
          3970 => x"53",
          3971 => x"b7",
          3972 => x"83",
          3973 => x"84",
          3974 => x"81",
          3975 => x"84",
          3976 => x"81",
          3977 => x"f4",
          3978 => x"34",
          3979 => x"80",
          3980 => x"19",
          3981 => x"80",
          3982 => x"0b",
          3983 => x"84",
          3984 => x"9e",
          3985 => x"19",
          3986 => x"a0",
          3987 => x"84",
          3988 => x"75",
          3989 => x"5b",
          3990 => x"08",
          3991 => x"88",
          3992 => x"7a",
          3993 => x"34",
          3994 => x"19",
          3995 => x"b4",
          3996 => x"79",
          3997 => x"3f",
          3998 => x"52",
          3999 => x"84",
          4000 => x"38",
          4001 => x"60",
          4002 => x"27",
          4003 => x"8c",
          4004 => x"0c",
          4005 => x"56",
          4006 => x"74",
          4007 => x"2e",
          4008 => x"2a",
          4009 => x"05",
          4010 => x"79",
          4011 => x"7b",
          4012 => x"38",
          4013 => x"81",
          4014 => x"b8",
          4015 => x"59",
          4016 => x"ff",
          4017 => x"b8",
          4018 => x"a8",
          4019 => x"b4",
          4020 => x"0b",
          4021 => x"74",
          4022 => x"38",
          4023 => x"81",
          4024 => x"b8",
          4025 => x"59",
          4026 => x"fe",
          4027 => x"b8",
          4028 => x"78",
          4029 => x"59",
          4030 => x"9f",
          4031 => x"3d",
          4032 => x"08",
          4033 => x"b5",
          4034 => x"5c",
          4035 => x"06",
          4036 => x"b8",
          4037 => x"a8",
          4038 => x"85",
          4039 => x"18",
          4040 => x"83",
          4041 => x"11",
          4042 => x"84",
          4043 => x"0d",
          4044 => x"fd",
          4045 => x"08",
          4046 => x"b5",
          4047 => x"5c",
          4048 => x"06",
          4049 => x"b8",
          4050 => x"c0",
          4051 => x"85",
          4052 => x"18",
          4053 => x"2b",
          4054 => x"83",
          4055 => x"2b",
          4056 => x"70",
          4057 => x"80",
          4058 => x"b8",
          4059 => x"56",
          4060 => x"17",
          4061 => x"18",
          4062 => x"5a",
          4063 => x"81",
          4064 => x"08",
          4065 => x"18",
          4066 => x"5e",
          4067 => x"38",
          4068 => x"09",
          4069 => x"b4",
          4070 => x"7b",
          4071 => x"3f",
          4072 => x"b4",
          4073 => x"81",
          4074 => x"84",
          4075 => x"06",
          4076 => x"83",
          4077 => x"08",
          4078 => x"8b",
          4079 => x"2e",
          4080 => x"5b",
          4081 => x"08",
          4082 => x"33",
          4083 => x"84",
          4084 => x"06",
          4085 => x"83",
          4086 => x"08",
          4087 => x"7d",
          4088 => x"82",
          4089 => x"81",
          4090 => x"17",
          4091 => x"52",
          4092 => x"7a",
          4093 => x"17",
          4094 => x"18",
          4095 => x"5a",
          4096 => x"81",
          4097 => x"08",
          4098 => x"18",
          4099 => x"55",
          4100 => x"38",
          4101 => x"09",
          4102 => x"b4",
          4103 => x"7d",
          4104 => x"3f",
          4105 => x"b4",
          4106 => x"7b",
          4107 => x"3f",
          4108 => x"bb",
          4109 => x"60",
          4110 => x"81",
          4111 => x"08",
          4112 => x"78",
          4113 => x"80",
          4114 => x"77",
          4115 => x"04",
          4116 => x"58",
          4117 => x"76",
          4118 => x"33",
          4119 => x"81",
          4120 => x"53",
          4121 => x"f2",
          4122 => x"2e",
          4123 => x"b4",
          4124 => x"38",
          4125 => x"7b",
          4126 => x"b8",
          4127 => x"b9",
          4128 => x"77",
          4129 => x"04",
          4130 => x"ff",
          4131 => x"05",
          4132 => x"5c",
          4133 => x"19",
          4134 => x"09",
          4135 => x"77",
          4136 => x"51",
          4137 => x"80",
          4138 => x"77",
          4139 => x"b7",
          4140 => x"79",
          4141 => x"98",
          4142 => x"06",
          4143 => x"34",
          4144 => x"34",
          4145 => x"34",
          4146 => x"34",
          4147 => x"39",
          4148 => x"a8",
          4149 => x"59",
          4150 => x"0b",
          4151 => x"74",
          4152 => x"38",
          4153 => x"81",
          4154 => x"b8",
          4155 => x"58",
          4156 => x"58",
          4157 => x"06",
          4158 => x"06",
          4159 => x"2e",
          4160 => x"06",
          4161 => x"5a",
          4162 => x"34",
          4163 => x"56",
          4164 => x"74",
          4165 => x"74",
          4166 => x"33",
          4167 => x"84",
          4168 => x"06",
          4169 => x"83",
          4170 => x"1b",
          4171 => x"e4",
          4172 => x"27",
          4173 => x"82",
          4174 => x"53",
          4175 => x"d8",
          4176 => x"85",
          4177 => x"1a",
          4178 => x"ff",
          4179 => x"56",
          4180 => x"76",
          4181 => x"07",
          4182 => x"83",
          4183 => x"76",
          4184 => x"33",
          4185 => x"84",
          4186 => x"06",
          4187 => x"83",
          4188 => x"1b",
          4189 => x"e4",
          4190 => x"27",
          4191 => x"74",
          4192 => x"38",
          4193 => x"81",
          4194 => x"5a",
          4195 => x"b8",
          4196 => x"57",
          4197 => x"e4",
          4198 => x"ae",
          4199 => x"34",
          4200 => x"31",
          4201 => x"5f",
          4202 => x"f0",
          4203 => x"2e",
          4204 => x"54",
          4205 => x"33",
          4206 => x"d0",
          4207 => x"70",
          4208 => x"cf",
          4209 => x"7c",
          4210 => x"84",
          4211 => x"19",
          4212 => x"1b",
          4213 => x"40",
          4214 => x"82",
          4215 => x"81",
          4216 => x"1e",
          4217 => x"ed",
          4218 => x"81",
          4219 => x"19",
          4220 => x"fd",
          4221 => x"06",
          4222 => x"59",
          4223 => x"88",
          4224 => x"fa",
          4225 => x"76",
          4226 => x"b8",
          4227 => x"8f",
          4228 => x"42",
          4229 => x"7d",
          4230 => x"7d",
          4231 => x"7d",
          4232 => x"fa",
          4233 => x"71",
          4234 => x"38",
          4235 => x"80",
          4236 => x"80",
          4237 => x"54",
          4238 => x"7b",
          4239 => x"16",
          4240 => x"38",
          4241 => x"38",
          4242 => x"84",
          4243 => x"38",
          4244 => x"2e",
          4245 => x"70",
          4246 => x"7b",
          4247 => x"aa",
          4248 => x"ff",
          4249 => x"e4",
          4250 => x"ff",
          4251 => x"ca",
          4252 => x"3f",
          4253 => x"27",
          4254 => x"84",
          4255 => x"9c",
          4256 => x"c4",
          4257 => x"1b",
          4258 => x"38",
          4259 => x"eb",
          4260 => x"81",
          4261 => x"08",
          4262 => x"25",
          4263 => x"54",
          4264 => x"38",
          4265 => x"38",
          4266 => x"fe",
          4267 => x"fe",
          4268 => x"96",
          4269 => x"ff",
          4270 => x"3f",
          4271 => x"08",
          4272 => x"80",
          4273 => x"38",
          4274 => x"0c",
          4275 => x"08",
          4276 => x"ff",
          4277 => x"81",
          4278 => x"55",
          4279 => x"0d",
          4280 => x"8c",
          4281 => x"58",
          4282 => x"b8",
          4283 => x"f5",
          4284 => x"ff",
          4285 => x"b8",
          4286 => x"56",
          4287 => x"55",
          4288 => x"7c",
          4289 => x"80",
          4290 => x"06",
          4291 => x"19",
          4292 => x"df",
          4293 => x"80",
          4294 => x"0b",
          4295 => x"27",
          4296 => x"0c",
          4297 => x"53",
          4298 => x"73",
          4299 => x"83",
          4300 => x"0c",
          4301 => x"8a",
          4302 => x"e4",
          4303 => x"08",
          4304 => x"8a",
          4305 => x"73",
          4306 => x"53",
          4307 => x"59",
          4308 => x"22",
          4309 => x"5a",
          4310 => x"39",
          4311 => x"84",
          4312 => x"08",
          4313 => x"b8",
          4314 => x"17",
          4315 => x"27",
          4316 => x"73",
          4317 => x"81",
          4318 => x"0d",
          4319 => x"90",
          4320 => x"f0",
          4321 => x"0b",
          4322 => x"84",
          4323 => x"83",
          4324 => x"15",
          4325 => x"38",
          4326 => x"55",
          4327 => x"98",
          4328 => x"1b",
          4329 => x"75",
          4330 => x"04",
          4331 => x"ff",
          4332 => x"da",
          4333 => x"3f",
          4334 => x"81",
          4335 => x"38",
          4336 => x"2e",
          4337 => x"e4",
          4338 => x"2e",
          4339 => x"76",
          4340 => x"08",
          4341 => x"80",
          4342 => x"b8",
          4343 => x"81",
          4344 => x"ff",
          4345 => x"1a",
          4346 => x"fe",
          4347 => x"56",
          4348 => x"8a",
          4349 => x"08",
          4350 => x"b8",
          4351 => x"80",
          4352 => x"15",
          4353 => x"19",
          4354 => x"38",
          4355 => x"81",
          4356 => x"b8",
          4357 => x"56",
          4358 => x"0b",
          4359 => x"04",
          4360 => x"19",
          4361 => x"e4",
          4362 => x"f3",
          4363 => x"34",
          4364 => x"55",
          4365 => x"38",
          4366 => x"09",
          4367 => x"b4",
          4368 => x"75",
          4369 => x"3f",
          4370 => x"74",
          4371 => x"2e",
          4372 => x"18",
          4373 => x"05",
          4374 => x"fd",
          4375 => x"29",
          4376 => x"5c",
          4377 => x"e4",
          4378 => x"0d",
          4379 => x"5a",
          4380 => x"58",
          4381 => x"38",
          4382 => x"b4",
          4383 => x"83",
          4384 => x"2e",
          4385 => x"54",
          4386 => x"33",
          4387 => x"08",
          4388 => x"57",
          4389 => x"82",
          4390 => x"58",
          4391 => x"8b",
          4392 => x"06",
          4393 => x"81",
          4394 => x"70",
          4395 => x"07",
          4396 => x"38",
          4397 => x"88",
          4398 => x"81",
          4399 => x"7b",
          4400 => x"08",
          4401 => x"38",
          4402 => x"38",
          4403 => x"0d",
          4404 => x"7e",
          4405 => x"3f",
          4406 => x"2e",
          4407 => x"b8",
          4408 => x"08",
          4409 => x"08",
          4410 => x"fe",
          4411 => x"82",
          4412 => x"81",
          4413 => x"05",
          4414 => x"e0",
          4415 => x"79",
          4416 => x"38",
          4417 => x"80",
          4418 => x"81",
          4419 => x"ac",
          4420 => x"2e",
          4421 => x"fe",
          4422 => x"09",
          4423 => x"84",
          4424 => x"84",
          4425 => x"77",
          4426 => x"57",
          4427 => x"38",
          4428 => x"1a",
          4429 => x"41",
          4430 => x"81",
          4431 => x"5a",
          4432 => x"17",
          4433 => x"33",
          4434 => x"7a",
          4435 => x"fe",
          4436 => x"05",
          4437 => x"1a",
          4438 => x"cc",
          4439 => x"06",
          4440 => x"79",
          4441 => x"10",
          4442 => x"1d",
          4443 => x"9d",
          4444 => x"38",
          4445 => x"a8",
          4446 => x"2a",
          4447 => x"81",
          4448 => x"81",
          4449 => x"76",
          4450 => x"38",
          4451 => x"b8",
          4452 => x"3d",
          4453 => x"52",
          4454 => x"e4",
          4455 => x"80",
          4456 => x"0b",
          4457 => x"1c",
          4458 => x"76",
          4459 => x"78",
          4460 => x"06",
          4461 => x"b8",
          4462 => x"e0",
          4463 => x"85",
          4464 => x"1c",
          4465 => x"9c",
          4466 => x"80",
          4467 => x"bf",
          4468 => x"77",
          4469 => x"80",
          4470 => x"55",
          4471 => x"80",
          4472 => x"38",
          4473 => x"8b",
          4474 => x"29",
          4475 => x"57",
          4476 => x"19",
          4477 => x"7f",
          4478 => x"81",
          4479 => x"a0",
          4480 => x"5a",
          4481 => x"71",
          4482 => x"40",
          4483 => x"80",
          4484 => x"0b",
          4485 => x"f5",
          4486 => x"84",
          4487 => x"38",
          4488 => x"0d",
          4489 => x"7d",
          4490 => x"3f",
          4491 => x"2e",
          4492 => x"b8",
          4493 => x"08",
          4494 => x"08",
          4495 => x"fd",
          4496 => x"82",
          4497 => x"81",
          4498 => x"05",
          4499 => x"db",
          4500 => x"77",
          4501 => x"70",
          4502 => x"fe",
          4503 => x"5a",
          4504 => x"33",
          4505 => x"08",
          4506 => x"76",
          4507 => x"74",
          4508 => x"3f",
          4509 => x"e4",
          4510 => x"c8",
          4511 => x"81",
          4512 => x"fe",
          4513 => x"77",
          4514 => x"1b",
          4515 => x"71",
          4516 => x"ff",
          4517 => x"8d",
          4518 => x"59",
          4519 => x"05",
          4520 => x"2b",
          4521 => x"80",
          4522 => x"84",
          4523 => x"84",
          4524 => x"70",
          4525 => x"81",
          4526 => x"08",
          4527 => x"76",
          4528 => x"ff",
          4529 => x"81",
          4530 => x"38",
          4531 => x"60",
          4532 => x"b4",
          4533 => x"5e",
          4534 => x"b8",
          4535 => x"83",
          4536 => x"ff",
          4537 => x"68",
          4538 => x"a0",
          4539 => x"74",
          4540 => x"70",
          4541 => x"8e",
          4542 => x"22",
          4543 => x"3d",
          4544 => x"58",
          4545 => x"33",
          4546 => x"15",
          4547 => x"05",
          4548 => x"80",
          4549 => x"ab",
          4550 => x"5b",
          4551 => x"7a",
          4552 => x"05",
          4553 => x"34",
          4554 => x"7b",
          4555 => x"56",
          4556 => x"82",
          4557 => x"06",
          4558 => x"83",
          4559 => x"06",
          4560 => x"87",
          4561 => x"ff",
          4562 => x"78",
          4563 => x"84",
          4564 => x"b0",
          4565 => x"84",
          4566 => x"ff",
          4567 => x"59",
          4568 => x"80",
          4569 => x"80",
          4570 => x"74",
          4571 => x"75",
          4572 => x"70",
          4573 => x"81",
          4574 => x"55",
          4575 => x"78",
          4576 => x"57",
          4577 => x"27",
          4578 => x"3f",
          4579 => x"1b",
          4580 => x"38",
          4581 => x"e7",
          4582 => x"b8",
          4583 => x"82",
          4584 => x"ab",
          4585 => x"80",
          4586 => x"2a",
          4587 => x"2e",
          4588 => x"fe",
          4589 => x"1b",
          4590 => x"3f",
          4591 => x"e4",
          4592 => x"08",
          4593 => x"56",
          4594 => x"85",
          4595 => x"77",
          4596 => x"81",
          4597 => x"18",
          4598 => x"e4",
          4599 => x"81",
          4600 => x"76",
          4601 => x"56",
          4602 => x"38",
          4603 => x"56",
          4604 => x"81",
          4605 => x"38",
          4606 => x"84",
          4607 => x"08",
          4608 => x"75",
          4609 => x"75",
          4610 => x"81",
          4611 => x"1c",
          4612 => x"33",
          4613 => x"81",
          4614 => x"1c",
          4615 => x"e4",
          4616 => x"81",
          4617 => x"75",
          4618 => x"08",
          4619 => x"58",
          4620 => x"8b",
          4621 => x"55",
          4622 => x"70",
          4623 => x"74",
          4624 => x"33",
          4625 => x"34",
          4626 => x"75",
          4627 => x"04",
          4628 => x"07",
          4629 => x"74",
          4630 => x"3f",
          4631 => x"e4",
          4632 => x"bd",
          4633 => x"7c",
          4634 => x"3f",
          4635 => x"81",
          4636 => x"08",
          4637 => x"19",
          4638 => x"27",
          4639 => x"82",
          4640 => x"08",
          4641 => x"90",
          4642 => x"51",
          4643 => x"58",
          4644 => x"79",
          4645 => x"57",
          4646 => x"05",
          4647 => x"76",
          4648 => x"59",
          4649 => x"ff",
          4650 => x"08",
          4651 => x"2e",
          4652 => x"76",
          4653 => x"81",
          4654 => x"1c",
          4655 => x"e4",
          4656 => x"81",
          4657 => x"75",
          4658 => x"1f",
          4659 => x"5f",
          4660 => x"1c",
          4661 => x"1c",
          4662 => x"29",
          4663 => x"76",
          4664 => x"10",
          4665 => x"56",
          4666 => x"55",
          4667 => x"76",
          4668 => x"85",
          4669 => x"58",
          4670 => x"ff",
          4671 => x"1f",
          4672 => x"81",
          4673 => x"83",
          4674 => x"e1",
          4675 => x"b8",
          4676 => x"05",
          4677 => x"39",
          4678 => x"1c",
          4679 => x"d0",
          4680 => x"08",
          4681 => x"83",
          4682 => x"08",
          4683 => x"60",
          4684 => x"82",
          4685 => x"81",
          4686 => x"1c",
          4687 => x"52",
          4688 => x"77",
          4689 => x"08",
          4690 => x"e5",
          4691 => x"fb",
          4692 => x"80",
          4693 => x"7c",
          4694 => x"81",
          4695 => x"81",
          4696 => x"b8",
          4697 => x"bc",
          4698 => x"34",
          4699 => x"55",
          4700 => x"82",
          4701 => x"38",
          4702 => x"39",
          4703 => x"2e",
          4704 => x"1a",
          4705 => x"56",
          4706 => x"fd",
          4707 => x"1d",
          4708 => x"33",
          4709 => x"81",
          4710 => x"05",
          4711 => x"ce",
          4712 => x"0d",
          4713 => x"80",
          4714 => x"80",
          4715 => x"ff",
          4716 => x"60",
          4717 => x"5b",
          4718 => x"77",
          4719 => x"5b",
          4720 => x"d0",
          4721 => x"58",
          4722 => x"38",
          4723 => x"5d",
          4724 => x"30",
          4725 => x"5a",
          4726 => x"80",
          4727 => x"1f",
          4728 => x"70",
          4729 => x"a0",
          4730 => x"bc",
          4731 => x"72",
          4732 => x"8b",
          4733 => x"38",
          4734 => x"81",
          4735 => x"59",
          4736 => x"ff",
          4737 => x"80",
          4738 => x"53",
          4739 => x"bf",
          4740 => x"17",
          4741 => x"34",
          4742 => x"53",
          4743 => x"9c",
          4744 => x"1e",
          4745 => x"11",
          4746 => x"71",
          4747 => x"72",
          4748 => x"64",
          4749 => x"33",
          4750 => x"40",
          4751 => x"23",
          4752 => x"88",
          4753 => x"23",
          4754 => x"fe",
          4755 => x"ff",
          4756 => x"52",
          4757 => x"91",
          4758 => x"ff",
          4759 => x"ad",
          4760 => x"74",
          4761 => x"97",
          4762 => x"0b",
          4763 => x"75",
          4764 => x"fd",
          4765 => x"76",
          4766 => x"80",
          4767 => x"f9",
          4768 => x"58",
          4769 => x"cd",
          4770 => x"57",
          4771 => x"7c",
          4772 => x"14",
          4773 => x"99",
          4774 => x"11",
          4775 => x"38",
          4776 => x"5e",
          4777 => x"70",
          4778 => x"78",
          4779 => x"81",
          4780 => x"5e",
          4781 => x"38",
          4782 => x"cc",
          4783 => x"70",
          4784 => x"fc",
          4785 => x"08",
          4786 => x"33",
          4787 => x"38",
          4788 => x"df",
          4789 => x"98",
          4790 => x"96",
          4791 => x"75",
          4792 => x"16",
          4793 => x"81",
          4794 => x"df",
          4795 => x"81",
          4796 => x"8b",
          4797 => x"23",
          4798 => x"06",
          4799 => x"27",
          4800 => x"55",
          4801 => x"2e",
          4802 => x"b2",
          4803 => x"80",
          4804 => x"56",
          4805 => x"75",
          4806 => x"70",
          4807 => x"ee",
          4808 => x"81",
          4809 => x"fd",
          4810 => x"23",
          4811 => x"52",
          4812 => x"fe",
          4813 => x"80",
          4814 => x"73",
          4815 => x"2e",
          4816 => x"80",
          4817 => x"dd",
          4818 => x"70",
          4819 => x"72",
          4820 => x"33",
          4821 => x"74",
          4822 => x"83",
          4823 => x"3f",
          4824 => x"06",
          4825 => x"73",
          4826 => x"04",
          4827 => x"06",
          4828 => x"38",
          4829 => x"34",
          4830 => x"84",
          4831 => x"93",
          4832 => x"32",
          4833 => x"41",
          4834 => x"38",
          4835 => x"55",
          4836 => x"72",
          4837 => x"25",
          4838 => x"38",
          4839 => x"2b",
          4840 => x"76",
          4841 => x"59",
          4842 => x"78",
          4843 => x"32",
          4844 => x"56",
          4845 => x"38",
          4846 => x"dd",
          4847 => x"76",
          4848 => x"80",
          4849 => x"72",
          4850 => x"82",
          4851 => x"53",
          4852 => x"80",
          4853 => x"70",
          4854 => x"38",
          4855 => x"17",
          4856 => x"14",
          4857 => x"09",
          4858 => x"1d",
          4859 => x"56",
          4860 => x"72",
          4861 => x"22",
          4862 => x"80",
          4863 => x"83",
          4864 => x"70",
          4865 => x"2e",
          4866 => x"72",
          4867 => x"59",
          4868 => x"07",
          4869 => x"54",
          4870 => x"7c",
          4871 => x"2e",
          4872 => x"77",
          4873 => x"8b",
          4874 => x"18",
          4875 => x"81",
          4876 => x"38",
          4877 => x"2e",
          4878 => x"e3",
          4879 => x"2e",
          4880 => x"74",
          4881 => x"2a",
          4882 => x"81",
          4883 => x"79",
          4884 => x"06",
          4885 => x"88",
          4886 => x"51",
          4887 => x"ab",
          4888 => x"08",
          4889 => x"e4",
          4890 => x"f7",
          4891 => x"79",
          4892 => x"2a",
          4893 => x"7b",
          4894 => x"16",
          4895 => x"81",
          4896 => x"40",
          4897 => x"38",
          4898 => x"83",
          4899 => x"22",
          4900 => x"fc",
          4901 => x"2e",
          4902 => x"10",
          4903 => x"a0",
          4904 => x"26",
          4905 => x"81",
          4906 => x"73",
          4907 => x"77",
          4908 => x"3f",
          4909 => x"56",
          4910 => x"38",
          4911 => x"fa",
          4912 => x"2a",
          4913 => x"83",
          4914 => x"06",
          4915 => x"d2",
          4916 => x"33",
          4917 => x"82",
          4918 => x"08",
          4919 => x"22",
          4920 => x"76",
          4921 => x"ab",
          4922 => x"5a",
          4923 => x"fc",
          4924 => x"8c",
          4925 => x"79",
          4926 => x"0b",
          4927 => x"81",
          4928 => x"80",
          4929 => x"b8",
          4930 => x"80",
          4931 => x"27",
          4932 => x"7b",
          4933 => x"7d",
          4934 => x"39",
          4935 => x"74",
          4936 => x"e4",
          4937 => x"2a",
          4938 => x"c4",
          4939 => x"f4",
          4940 => x"26",
          4941 => x"85",
          4942 => x"8c",
          4943 => x"59",
          4944 => x"75",
          4945 => x"70",
          4946 => x"ee",
          4947 => x"80",
          4948 => x"99",
          4949 => x"81",
          4950 => x"59",
          4951 => x"07",
          4952 => x"83",
          4953 => x"7b",
          4954 => x"81",
          4955 => x"39",
          4956 => x"8c",
          4957 => x"78",
          4958 => x"7a",
          4959 => x"5b",
          4960 => x"d2",
          4961 => x"15",
          4962 => x"07",
          4963 => x"fd",
          4964 => x"88",
          4965 => x"1b",
          4966 => x"79",
          4967 => x"79",
          4968 => x"76",
          4969 => x"a3",
          4970 => x"81",
          4971 => x"0b",
          4972 => x"04",
          4973 => x"05",
          4974 => x"80",
          4975 => x"5b",
          4976 => x"79",
          4977 => x"26",
          4978 => x"38",
          4979 => x"c7",
          4980 => x"76",
          4981 => x"84",
          4982 => x"8c",
          4983 => x"76",
          4984 => x"33",
          4985 => x"81",
          4986 => x"84",
          4987 => x"81",
          4988 => x"96",
          4989 => x"84",
          4990 => x"81",
          4991 => x"a4",
          4992 => x"06",
          4993 => x"7f",
          4994 => x"38",
          4995 => x"58",
          4996 => x"83",
          4997 => x"7a",
          4998 => x"b8",
          4999 => x"58",
          5000 => x"08",
          5001 => x"59",
          5002 => x"99",
          5003 => x"18",
          5004 => x"83",
          5005 => x"a5",
          5006 => x"b8",
          5007 => x"38",
          5008 => x"38",
          5009 => x"38",
          5010 => x"33",
          5011 => x"84",
          5012 => x"38",
          5013 => x"33",
          5014 => x"a4",
          5015 => x"82",
          5016 => x"2b",
          5017 => x"88",
          5018 => x"45",
          5019 => x"0c",
          5020 => x"80",
          5021 => x"ff",
          5022 => x"81",
          5023 => x"06",
          5024 => x"5a",
          5025 => x"59",
          5026 => x"18",
          5027 => x"80",
          5028 => x"71",
          5029 => x"18",
          5030 => x"8d",
          5031 => x"17",
          5032 => x"2b",
          5033 => x"d8",
          5034 => x"71",
          5035 => x"14",
          5036 => x"33",
          5037 => x"42",
          5038 => x"18",
          5039 => x"8d",
          5040 => x"7d",
          5041 => x"75",
          5042 => x"7a",
          5043 => x"b8",
          5044 => x"80",
          5045 => x"08",
          5046 => x"38",
          5047 => x"83",
          5048 => x"85",
          5049 => x"9c",
          5050 => x"1d",
          5051 => x"1a",
          5052 => x"87",
          5053 => x"7b",
          5054 => x"ac",
          5055 => x"2e",
          5056 => x"2a",
          5057 => x"ff",
          5058 => x"a0",
          5059 => x"94",
          5060 => x"ff",
          5061 => x"2e",
          5062 => x"d0",
          5063 => x"d0",
          5064 => x"d0",
          5065 => x"98",
          5066 => x"e4",
          5067 => x"84",
          5068 => x"76",
          5069 => x"57",
          5070 => x"82",
          5071 => x"5d",
          5072 => x"80",
          5073 => x"5c",
          5074 => x"81",
          5075 => x"5b",
          5076 => x"77",
          5077 => x"81",
          5078 => x"58",
          5079 => x"70",
          5080 => x"70",
          5081 => x"09",
          5082 => x"38",
          5083 => x"07",
          5084 => x"7a",
          5085 => x"84",
          5086 => x"98",
          5087 => x"80",
          5088 => x"81",
          5089 => x"38",
          5090 => x"33",
          5091 => x"81",
          5092 => x"eb",
          5093 => x"07",
          5094 => x"75",
          5095 => x"3d",
          5096 => x"16",
          5097 => x"a5",
          5098 => x"17",
          5099 => x"07",
          5100 => x"88",
          5101 => x"52",
          5102 => x"70",
          5103 => x"17",
          5104 => x"38",
          5105 => x"70",
          5106 => x"71",
          5107 => x"1c",
          5108 => x"08",
          5109 => x"fb",
          5110 => x"0b",
          5111 => x"7a",
          5112 => x"53",
          5113 => x"ff",
          5114 => x"76",
          5115 => x"74",
          5116 => x"38",
          5117 => x"2b",
          5118 => x"d4",
          5119 => x"80",
          5120 => x"81",
          5121 => x"eb",
          5122 => x"07",
          5123 => x"81",
          5124 => x"81",
          5125 => x"d9",
          5126 => x"09",
          5127 => x"76",
          5128 => x"f8",
          5129 => x"5a",
          5130 => x"a8",
          5131 => x"e4",
          5132 => x"05",
          5133 => x"33",
          5134 => x"56",
          5135 => x"75",
          5136 => x"8a",
          5137 => x"7b",
          5138 => x"81",
          5139 => x"1b",
          5140 => x"85",
          5141 => x"82",
          5142 => x"fa",
          5143 => x"97",
          5144 => x"2e",
          5145 => x"18",
          5146 => x"b7",
          5147 => x"97",
          5148 => x"18",
          5149 => x"70",
          5150 => x"05",
          5151 => x"5b",
          5152 => x"d1",
          5153 => x"0b",
          5154 => x"5a",
          5155 => x"7a",
          5156 => x"31",
          5157 => x"80",
          5158 => x"e1",
          5159 => x"59",
          5160 => x"39",
          5161 => x"33",
          5162 => x"81",
          5163 => x"81",
          5164 => x"78",
          5165 => x"7a",
          5166 => x"38",
          5167 => x"81",
          5168 => x"84",
          5169 => x"ff",
          5170 => x"79",
          5171 => x"84",
          5172 => x"71",
          5173 => x"d4",
          5174 => x"38",
          5175 => x"33",
          5176 => x"81",
          5177 => x"75",
          5178 => x"42",
          5179 => x"d2",
          5180 => x"84",
          5181 => x"33",
          5182 => x"81",
          5183 => x"75",
          5184 => x"5c",
          5185 => x"f2",
          5186 => x"84",
          5187 => x"33",
          5188 => x"81",
          5189 => x"75",
          5190 => x"84",
          5191 => x"33",
          5192 => x"81",
          5193 => x"75",
          5194 => x"59",
          5195 => x"5b",
          5196 => x"bc",
          5197 => x"bc",
          5198 => x"c4",
          5199 => x"18",
          5200 => x"f8",
          5201 => x"f2",
          5202 => x"53",
          5203 => x"52",
          5204 => x"e4",
          5205 => x"a4",
          5206 => x"34",
          5207 => x"40",
          5208 => x"82",
          5209 => x"8d",
          5210 => x"a0",
          5211 => x"91",
          5212 => x"e4",
          5213 => x"80",
          5214 => x"71",
          5215 => x"7d",
          5216 => x"61",
          5217 => x"11",
          5218 => x"71",
          5219 => x"72",
          5220 => x"ac",
          5221 => x"43",
          5222 => x"75",
          5223 => x"82",
          5224 => x"f2",
          5225 => x"83",
          5226 => x"f5",
          5227 => x"b4",
          5228 => x"78",
          5229 => x"e7",
          5230 => x"02",
          5231 => x"93",
          5232 => x"40",
          5233 => x"70",
          5234 => x"55",
          5235 => x"73",
          5236 => x"38",
          5237 => x"24",
          5238 => x"d0",
          5239 => x"80",
          5240 => x"54",
          5241 => x"34",
          5242 => x"7c",
          5243 => x"3d",
          5244 => x"3f",
          5245 => x"b8",
          5246 => x"0b",
          5247 => x"04",
          5248 => x"06",
          5249 => x"38",
          5250 => x"05",
          5251 => x"38",
          5252 => x"5f",
          5253 => x"70",
          5254 => x"05",
          5255 => x"55",
          5256 => x"70",
          5257 => x"16",
          5258 => x"16",
          5259 => x"30",
          5260 => x"2e",
          5261 => x"be",
          5262 => x"72",
          5263 => x"54",
          5264 => x"84",
          5265 => x"99",
          5266 => x"83",
          5267 => x"54",
          5268 => x"02",
          5269 => x"59",
          5270 => x"74",
          5271 => x"05",
          5272 => x"ed",
          5273 => x"84",
          5274 => x"80",
          5275 => x"e4",
          5276 => x"6d",
          5277 => x"9a",
          5278 => x"b8",
          5279 => x"77",
          5280 => x"ca",
          5281 => x"76",
          5282 => x"07",
          5283 => x"2a",
          5284 => x"d1",
          5285 => x"33",
          5286 => x"42",
          5287 => x"84",
          5288 => x"80",
          5289 => x"17",
          5290 => x"66",
          5291 => x"67",
          5292 => x"80",
          5293 => x"7c",
          5294 => x"80",
          5295 => x"1c",
          5296 => x"0b",
          5297 => x"83",
          5298 => x"38",
          5299 => x"53",
          5300 => x"38",
          5301 => x"38",
          5302 => x"39",
          5303 => x"2b",
          5304 => x"38",
          5305 => x"fe",
          5306 => x"80",
          5307 => x"06",
          5308 => x"81",
          5309 => x"89",
          5310 => x"f6",
          5311 => x"75",
          5312 => x"07",
          5313 => x"0c",
          5314 => x"33",
          5315 => x"73",
          5316 => x"83",
          5317 => x"0c",
          5318 => x"33",
          5319 => x"81",
          5320 => x"75",
          5321 => x"0c",
          5322 => x"57",
          5323 => x"23",
          5324 => x"1a",
          5325 => x"85",
          5326 => x"84",
          5327 => x"38",
          5328 => x"70",
          5329 => x"30",
          5330 => x"79",
          5331 => x"76",
          5332 => x"86",
          5333 => x"db",
          5334 => x"b8",
          5335 => x"57",
          5336 => x"cb",
          5337 => x"02",
          5338 => x"7d",
          5339 => x"55",
          5340 => x"57",
          5341 => x"57",
          5342 => x"57",
          5343 => x"51",
          5344 => x"78",
          5345 => x"38",
          5346 => x"57",
          5347 => x"94",
          5348 => x"2b",
          5349 => x"fc",
          5350 => x"bd",
          5351 => x"cb",
          5352 => x"b8",
          5353 => x"84",
          5354 => x"38",
          5355 => x"99",
          5356 => x"ff",
          5357 => x"83",
          5358 => x"94",
          5359 => x"27",
          5360 => x"0c",
          5361 => x"84",
          5362 => x"ff",
          5363 => x"94",
          5364 => x"fb",
          5365 => x"33",
          5366 => x"7e",
          5367 => x"17",
          5368 => x"0b",
          5369 => x"17",
          5370 => x"34",
          5371 => x"17",
          5372 => x"33",
          5373 => x"fb",
          5374 => x"7f",
          5375 => x"08",
          5376 => x"5a",
          5377 => x"38",
          5378 => x"81",
          5379 => x"84",
          5380 => x"ff",
          5381 => x"7e",
          5382 => x"57",
          5383 => x"79",
          5384 => x"16",
          5385 => x"17",
          5386 => x"84",
          5387 => x"06",
          5388 => x"83",
          5389 => x"08",
          5390 => x"74",
          5391 => x"82",
          5392 => x"81",
          5393 => x"16",
          5394 => x"52",
          5395 => x"3f",
          5396 => x"1a",
          5397 => x"98",
          5398 => x"83",
          5399 => x"9a",
          5400 => x"fe",
          5401 => x"f9",
          5402 => x"29",
          5403 => x"80",
          5404 => x"15",
          5405 => x"39",
          5406 => x"e4",
          5407 => x"da",
          5408 => x"79",
          5409 => x"5b",
          5410 => x"65",
          5411 => x"7e",
          5412 => x"38",
          5413 => x"38",
          5414 => x"38",
          5415 => x"59",
          5416 => x"55",
          5417 => x"38",
          5418 => x"38",
          5419 => x"56",
          5420 => x"1a",
          5421 => x"56",
          5422 => x"80",
          5423 => x"83",
          5424 => x"8a",
          5425 => x"06",
          5426 => x"38",
          5427 => x"84",
          5428 => x"38",
          5429 => x"1a",
          5430 => x"05",
          5431 => x"38",
          5432 => x"1b",
          5433 => x"83",
          5434 => x"59",
          5435 => x"77",
          5436 => x"75",
          5437 => x"7c",
          5438 => x"e0",
          5439 => x"38",
          5440 => x"80",
          5441 => x"31",
          5442 => x"80",
          5443 => x"58",
          5444 => x"77",
          5445 => x"55",
          5446 => x"7b",
          5447 => x"78",
          5448 => x"94",
          5449 => x"38",
          5450 => x"92",
          5451 => x"0c",
          5452 => x"8e",
          5453 => x"ff",
          5454 => x"7b",
          5455 => x"56",
          5456 => x"80",
          5457 => x"5f",
          5458 => x"e4",
          5459 => x"52",
          5460 => x"3f",
          5461 => x"38",
          5462 => x"0c",
          5463 => x"08",
          5464 => x"58",
          5465 => x"fe",
          5466 => x"33",
          5467 => x"16",
          5468 => x"74",
          5469 => x"81",
          5470 => x"da",
          5471 => x"19",
          5472 => x"1a",
          5473 => x"81",
          5474 => x"09",
          5475 => x"e4",
          5476 => x"a8",
          5477 => x"5c",
          5478 => x"e1",
          5479 => x"2e",
          5480 => x"54",
          5481 => x"53",
          5482 => x"9d",
          5483 => x"76",
          5484 => x"fe",
          5485 => x"51",
          5486 => x"08",
          5487 => x"51",
          5488 => x"08",
          5489 => x"74",
          5490 => x"81",
          5491 => x"b8",
          5492 => x"0b",
          5493 => x"e4",
          5494 => x"0d",
          5495 => x"5a",
          5496 => x"2e",
          5497 => x"2e",
          5498 => x"2e",
          5499 => x"22",
          5500 => x"38",
          5501 => x"82",
          5502 => x"82",
          5503 => x"2a",
          5504 => x"80",
          5505 => x"7b",
          5506 => x"38",
          5507 => x"81",
          5508 => x"82",
          5509 => x"05",
          5510 => x"aa",
          5511 => x"08",
          5512 => x"74",
          5513 => x"2e",
          5514 => x"88",
          5515 => x"0c",
          5516 => x"08",
          5517 => x"fe",
          5518 => x"58",
          5519 => x"16",
          5520 => x"05",
          5521 => x"38",
          5522 => x"77",
          5523 => x"5f",
          5524 => x"31",
          5525 => x"81",
          5526 => x"84",
          5527 => x"b4",
          5528 => x"78",
          5529 => x"18",
          5530 => x"74",
          5531 => x"81",
          5532 => x"ef",
          5533 => x"77",
          5534 => x"08",
          5535 => x"08",
          5536 => x"1e",
          5537 => x"75",
          5538 => x"1b",
          5539 => x"33",
          5540 => x"90",
          5541 => x"e4",
          5542 => x"b8",
          5543 => x"16",
          5544 => x"56",
          5545 => x"59",
          5546 => x"71",
          5547 => x"38",
          5548 => x"78",
          5549 => x"33",
          5550 => x"09",
          5551 => x"77",
          5552 => x"51",
          5553 => x"08",
          5554 => x"5c",
          5555 => x"38",
          5556 => x"11",
          5557 => x"58",
          5558 => x"81",
          5559 => x"57",
          5560 => x"60",
          5561 => x"a3",
          5562 => x"b8",
          5563 => x"40",
          5564 => x"b8",
          5565 => x"ff",
          5566 => x"17",
          5567 => x"31",
          5568 => x"a0",
          5569 => x"16",
          5570 => x"06",
          5571 => x"08",
          5572 => x"81",
          5573 => x"7e",
          5574 => x"57",
          5575 => x"83",
          5576 => x"60",
          5577 => x"58",
          5578 => x"fd",
          5579 => x"51",
          5580 => x"08",
          5581 => x"38",
          5582 => x"76",
          5583 => x"84",
          5584 => x"08",
          5585 => x"b4",
          5586 => x"81",
          5587 => x"3f",
          5588 => x"84",
          5589 => x"16",
          5590 => x"a0",
          5591 => x"16",
          5592 => x"06",
          5593 => x"08",
          5594 => x"81",
          5595 => x"60",
          5596 => x"51",
          5597 => x"08",
          5598 => x"74",
          5599 => x"81",
          5600 => x"70",
          5601 => x"96",
          5602 => x"c6",
          5603 => x"34",
          5604 => x"55",
          5605 => x"38",
          5606 => x"09",
          5607 => x"b4",
          5608 => x"76",
          5609 => x"87",
          5610 => x"1b",
          5611 => x"0b",
          5612 => x"e4",
          5613 => x"91",
          5614 => x"0c",
          5615 => x"7d",
          5616 => x"38",
          5617 => x"38",
          5618 => x"38",
          5619 => x"59",
          5620 => x"55",
          5621 => x"38",
          5622 => x"06",
          5623 => x"38",
          5624 => x"17",
          5625 => x"33",
          5626 => x"78",
          5627 => x"51",
          5628 => x"08",
          5629 => x"56",
          5630 => x"38",
          5631 => x"07",
          5632 => x"08",
          5633 => x"06",
          5634 => x"7a",
          5635 => x"9c",
          5636 => x"5b",
          5637 => x"18",
          5638 => x"2a",
          5639 => x"2a",
          5640 => x"2a",
          5641 => x"34",
          5642 => x"98",
          5643 => x"34",
          5644 => x"93",
          5645 => x"1c",
          5646 => x"84",
          5647 => x"bf",
          5648 => x"75",
          5649 => x"04",
          5650 => x"17",
          5651 => x"ff",
          5652 => x"e4",
          5653 => x"08",
          5654 => x"18",
          5655 => x"55",
          5656 => x"38",
          5657 => x"09",
          5658 => x"b4",
          5659 => x"7a",
          5660 => x"ef",
          5661 => x"90",
          5662 => x"88",
          5663 => x"18",
          5664 => x"2a",
          5665 => x"2a",
          5666 => x"2a",
          5667 => x"34",
          5668 => x"98",
          5669 => x"34",
          5670 => x"93",
          5671 => x"1c",
          5672 => x"84",
          5673 => x"bf",
          5674 => x"fe",
          5675 => x"90",
          5676 => x"06",
          5677 => x"08",
          5678 => x"0d",
          5679 => x"84",
          5680 => x"08",
          5681 => x"9e",
          5682 => x"96",
          5683 => x"8e",
          5684 => x"58",
          5685 => x"52",
          5686 => x"75",
          5687 => x"89",
          5688 => x"ff",
          5689 => x"81",
          5690 => x"08",
          5691 => x"ff",
          5692 => x"2e",
          5693 => x"33",
          5694 => x"2e",
          5695 => x"2e",
          5696 => x"80",
          5697 => x"c0",
          5698 => x"8c",
          5699 => x"e4",
          5700 => x"d0",
          5701 => x"53",
          5702 => x"73",
          5703 => x"73",
          5704 => x"83",
          5705 => x"56",
          5706 => x"75",
          5707 => x"12",
          5708 => x"38",
          5709 => x"54",
          5710 => x"89",
          5711 => x"54",
          5712 => x"51",
          5713 => x"38",
          5714 => x"70",
          5715 => x"07",
          5716 => x"38",
          5717 => x"78",
          5718 => x"cf",
          5719 => x"76",
          5720 => x"0d",
          5721 => x"99",
          5722 => x"e4",
          5723 => x"2e",
          5724 => x"98",
          5725 => x"98",
          5726 => x"84",
          5727 => x"08",
          5728 => x"33",
          5729 => x"24",
          5730 => x"70",
          5731 => x"80",
          5732 => x"33",
          5733 => x"73",
          5734 => x"83",
          5735 => x"74",
          5736 => x"04",
          5737 => x"81",
          5738 => x"b8",
          5739 => x"16",
          5740 => x"71",
          5741 => x"0c",
          5742 => x"12",
          5743 => x"98",
          5744 => x"80",
          5745 => x"5d",
          5746 => x"e4",
          5747 => x"3d",
          5748 => x"08",
          5749 => x"38",
          5750 => x"98",
          5751 => x"80",
          5752 => x"2e",
          5753 => x"3d",
          5754 => x"a4",
          5755 => x"84",
          5756 => x"80",
          5757 => x"08",
          5758 => x"08",
          5759 => x"c7",
          5760 => x"52",
          5761 => x"3f",
          5762 => x"38",
          5763 => x"0c",
          5764 => x"08",
          5765 => x"88",
          5766 => x"59",
          5767 => x"38",
          5768 => x"7a",
          5769 => x"e4",
          5770 => x"9f",
          5771 => x"f5",
          5772 => x"b8",
          5773 => x"08",
          5774 => x"88",
          5775 => x"59",
          5776 => x"38",
          5777 => x"e4",
          5778 => x"3f",
          5779 => x"e4",
          5780 => x"84",
          5781 => x"38",
          5782 => x"7a",
          5783 => x"82",
          5784 => x"90",
          5785 => x"17",
          5786 => x"38",
          5787 => x"95",
          5788 => x"17",
          5789 => x"3d",
          5790 => x"59",
          5791 => x"eb",
          5792 => x"11",
          5793 => x"3d",
          5794 => x"60",
          5795 => x"d0",
          5796 => x"d4",
          5797 => x"59",
          5798 => x"81",
          5799 => x"5a",
          5800 => x"78",
          5801 => x"27",
          5802 => x"7c",
          5803 => x"57",
          5804 => x"70",
          5805 => x"09",
          5806 => x"80",
          5807 => x"80",
          5808 => x"94",
          5809 => x"2b",
          5810 => x"f0",
          5811 => x"71",
          5812 => x"07",
          5813 => x"52",
          5814 => x"b8",
          5815 => x"80",
          5816 => x"81",
          5817 => x"70",
          5818 => x"88",
          5819 => x"08",
          5820 => x"83",
          5821 => x"08",
          5822 => x"74",
          5823 => x"82",
          5824 => x"81",
          5825 => x"16",
          5826 => x"52",
          5827 => x"3f",
          5828 => x"80",
          5829 => x"7b",
          5830 => x"70",
          5831 => x"08",
          5832 => x"7e",
          5833 => x"38",
          5834 => x"18",
          5835 => x"70",
          5836 => x"fe",
          5837 => x"81",
          5838 => x"81",
          5839 => x"38",
          5840 => x"34",
          5841 => x"3d",
          5842 => x"58",
          5843 => x"38",
          5844 => x"38",
          5845 => x"38",
          5846 => x"59",
          5847 => x"53",
          5848 => x"38",
          5849 => x"38",
          5850 => x"81",
          5851 => x"58",
          5852 => x"8a",
          5853 => x"56",
          5854 => x"52",
          5855 => x"84",
          5856 => x"70",
          5857 => x"84",
          5858 => x"38",
          5859 => x"0c",
          5860 => x"58",
          5861 => x"75",
          5862 => x"31",
          5863 => x"90",
          5864 => x"51",
          5865 => x"38",
          5866 => x"3f",
          5867 => x"e4",
          5868 => x"ff",
          5869 => x"b4",
          5870 => x"27",
          5871 => x"ff",
          5872 => x"81",
          5873 => x"3d",
          5874 => x"2a",
          5875 => x"38",
          5876 => x"58",
          5877 => x"b6",
          5878 => x"08",
          5879 => x"8c",
          5880 => x"07",
          5881 => x"ff",
          5882 => x"9c",
          5883 => x"9c",
          5884 => x"0c",
          5885 => x"16",
          5886 => x"2e",
          5887 => x"73",
          5888 => x"39",
          5889 => x"08",
          5890 => x"06",
          5891 => x"fe",
          5892 => x"55",
          5893 => x"8a",
          5894 => x"08",
          5895 => x"53",
          5896 => x"15",
          5897 => x"74",
          5898 => x"e4",
          5899 => x"33",
          5900 => x"e4",
          5901 => x"38",
          5902 => x"39",
          5903 => x"3f",
          5904 => x"e4",
          5905 => x"e4",
          5906 => x"b8",
          5907 => x"16",
          5908 => x"16",
          5909 => x"8b",
          5910 => x"56",
          5911 => x"80",
          5912 => x"3d",
          5913 => x"b8",
          5914 => x"80",
          5915 => x"54",
          5916 => x"0d",
          5917 => x"51",
          5918 => x"08",
          5919 => x"38",
          5920 => x"59",
          5921 => x"33",
          5922 => x"79",
          5923 => x"08",
          5924 => x"88",
          5925 => x"5a",
          5926 => x"77",
          5927 => x"22",
          5928 => x"ff",
          5929 => x"55",
          5930 => x"2e",
          5931 => x"fe",
          5932 => x"f6",
          5933 => x"71",
          5934 => x"07",
          5935 => x"39",
          5936 => x"74",
          5937 => x"72",
          5938 => x"71",
          5939 => x"84",
          5940 => x"94",
          5941 => x"38",
          5942 => x"0c",
          5943 => x"51",
          5944 => x"08",
          5945 => x"75",
          5946 => x"0d",
          5947 => x"80",
          5948 => x"80",
          5949 => x"80",
          5950 => x"16",
          5951 => x"97",
          5952 => x"75",
          5953 => x"f3",
          5954 => x"bd",
          5955 => x"b8",
          5956 => x"b8",
          5957 => x"51",
          5958 => x"51",
          5959 => x"08",
          5960 => x"9f",
          5961 => x"57",
          5962 => x"3d",
          5963 => x"53",
          5964 => x"51",
          5965 => x"08",
          5966 => x"9f",
          5967 => x"57",
          5968 => x"ff",
          5969 => x"84",
          5970 => x"81",
          5971 => x"84",
          5972 => x"fe",
          5973 => x"fe",
          5974 => x"80",
          5975 => x"52",
          5976 => x"08",
          5977 => x"8a",
          5978 => x"3d",
          5979 => x"b5",
          5980 => x"84",
          5981 => x"cb",
          5982 => x"80",
          5983 => x"d1",
          5984 => x"bd",
          5985 => x"3d",
          5986 => x"0c",
          5987 => x"66",
          5988 => x"ec",
          5989 => x"3f",
          5990 => x"e4",
          5991 => x"08",
          5992 => x"08",
          5993 => x"8d",
          5994 => x"e4",
          5995 => x"e4",
          5996 => x"2e",
          5997 => x"84",
          5998 => x"80",
          5999 => x"5d",
          6000 => x"ef",
          6001 => x"7c",
          6002 => x"b8",
          6003 => x"fc",
          6004 => x"2e",
          6005 => x"b4",
          6006 => x"80",
          6007 => x"2e",
          6008 => x"83",
          6009 => x"2b",
          6010 => x"70",
          6011 => x"80",
          6012 => x"30",
          6013 => x"05",
          6014 => x"41",
          6015 => x"5e",
          6016 => x"0c",
          6017 => x"81",
          6018 => x"84",
          6019 => x"81",
          6020 => x"70",
          6021 => x"fc",
          6022 => x"08",
          6023 => x"83",
          6024 => x"08",
          6025 => x"74",
          6026 => x"82",
          6027 => x"81",
          6028 => x"17",
          6029 => x"52",
          6030 => x"3f",
          6031 => x"42",
          6032 => x"51",
          6033 => x"08",
          6034 => x"e4",
          6035 => x"b8",
          6036 => x"08",
          6037 => x"62",
          6038 => x"76",
          6039 => x"94",
          6040 => x"58",
          6041 => x"77",
          6042 => x"33",
          6043 => x"80",
          6044 => x"ff",
          6045 => x"55",
          6046 => x"77",
          6047 => x"5a",
          6048 => x"84",
          6049 => x"18",
          6050 => x"5a",
          6051 => x"89",
          6052 => x"08",
          6053 => x"33",
          6054 => x"15",
          6055 => x"78",
          6056 => x"5a",
          6057 => x"56",
          6058 => x"70",
          6059 => x"55",
          6060 => x"17",
          6061 => x"b7",
          6062 => x"08",
          6063 => x"88",
          6064 => x"38",
          6065 => x"94",
          6066 => x"c0",
          6067 => x"80",
          6068 => x"75",
          6069 => x"3d",
          6070 => x"80",
          6071 => x"fe",
          6072 => x"84",
          6073 => x"38",
          6074 => x"d8",
          6075 => x"82",
          6076 => x"51",
          6077 => x"08",
          6078 => x"11",
          6079 => x"74",
          6080 => x"17",
          6081 => x"73",
          6082 => x"26",
          6083 => x"33",
          6084 => x"e4",
          6085 => x"38",
          6086 => x"39",
          6087 => x"73",
          6088 => x"c7",
          6089 => x"fe",
          6090 => x"ff",
          6091 => x"08",
          6092 => x"ae",
          6093 => x"9c",
          6094 => x"b8",
          6095 => x"58",
          6096 => x"08",
          6097 => x"08",
          6098 => x"74",
          6099 => x"52",
          6100 => x"b8",
          6101 => x"80",
          6102 => x"fc",
          6103 => x"84",
          6104 => x"38",
          6105 => x"dc",
          6106 => x"80",
          6107 => x"51",
          6108 => x"08",
          6109 => x"11",
          6110 => x"74",
          6111 => x"0c",
          6112 => x"84",
          6113 => x"ff",
          6114 => x"17",
          6115 => x"fe",
          6116 => x"59",
          6117 => x"39",
          6118 => x"fe",
          6119 => x"18",
          6120 => x"0b",
          6121 => x"39",
          6122 => x"81",
          6123 => x"82",
          6124 => x"a8",
          6125 => x"b8",
          6126 => x"80",
          6127 => x"0c",
          6128 => x"3d",
          6129 => x"ff",
          6130 => x"56",
          6131 => x"81",
          6132 => x"06",
          6133 => x"76",
          6134 => x"38",
          6135 => x"06",
          6136 => x"38",
          6137 => x"9a",
          6138 => x"33",
          6139 => x"2e",
          6140 => x"06",
          6141 => x"87",
          6142 => x"83",
          6143 => x"e4",
          6144 => x"ff",
          6145 => x"56",
          6146 => x"84",
          6147 => x"91",
          6148 => x"84",
          6149 => x"84",
          6150 => x"95",
          6151 => x"2b",
          6152 => x"5d",
          6153 => x"08",
          6154 => x"08",
          6155 => x"3d",
          6156 => x"80",
          6157 => x"8b",
          6158 => x"84",
          6159 => x"75",
          6160 => x"5a",
          6161 => x"2e",
          6162 => x"81",
          6163 => x"7b",
          6164 => x"fd",
          6165 => x"3f",
          6166 => x"0c",
          6167 => x"98",
          6168 => x"08",
          6169 => x"33",
          6170 => x"81",
          6171 => x"53",
          6172 => x"fe",
          6173 => x"80",
          6174 => x"75",
          6175 => x"38",
          6176 => x"81",
          6177 => x"7c",
          6178 => x"51",
          6179 => x"08",
          6180 => x"ff",
          6181 => x"06",
          6182 => x"39",
          6183 => x"52",
          6184 => x"3f",
          6185 => x"2e",
          6186 => x"b8",
          6187 => x"08",
          6188 => x"08",
          6189 => x"fe",
          6190 => x"82",
          6191 => x"81",
          6192 => x"05",
          6193 => x"fe",
          6194 => x"39",
          6195 => x"38",
          6196 => x"3f",
          6197 => x"e4",
          6198 => x"b8",
          6199 => x"84",
          6200 => x"38",
          6201 => x"fd",
          6202 => x"38",
          6203 => x"08",
          6204 => x"b0",
          6205 => x"17",
          6206 => x"34",
          6207 => x"38",
          6208 => x"fd",
          6209 => x"fd",
          6210 => x"e3",
          6211 => x"bc",
          6212 => x"c0",
          6213 => x"b8",
          6214 => x"84",
          6215 => x"7d",
          6216 => x"5a",
          6217 => x"08",
          6218 => x"88",
          6219 => x"0d",
          6220 => x"09",
          6221 => x"05",
          6222 => x"58",
          6223 => x"5f",
          6224 => x"ff",
          6225 => x"75",
          6226 => x"38",
          6227 => x"2e",
          6228 => x"ff",
          6229 => x"38",
          6230 => x"33",
          6231 => x"fe",
          6232 => x"56",
          6233 => x"8a",
          6234 => x"08",
          6235 => x"b8",
          6236 => x"80",
          6237 => x"15",
          6238 => x"17",
          6239 => x"38",
          6240 => x"81",
          6241 => x"84",
          6242 => x"18",
          6243 => x"39",
          6244 => x"17",
          6245 => x"fe",
          6246 => x"e4",
          6247 => x"83",
          6248 => x"08",
          6249 => x"fe",
          6250 => x"82",
          6251 => x"75",
          6252 => x"05",
          6253 => x"fe",
          6254 => x"56",
          6255 => x"27",
          6256 => x"27",
          6257 => x"fe",
          6258 => x"5a",
          6259 => x"96",
          6260 => x"fd",
          6261 => x"2e",
          6262 => x"76",
          6263 => x"e4",
          6264 => x"fe",
          6265 => x"77",
          6266 => x"18",
          6267 => x"7b",
          6268 => x"26",
          6269 => x"0c",
          6270 => x"55",
          6271 => x"56",
          6272 => x"f0",
          6273 => x"a0",
          6274 => x"16",
          6275 => x"0b",
          6276 => x"80",
          6277 => x"ce",
          6278 => x"a1",
          6279 => x"0b",
          6280 => x"ff",
          6281 => x"17",
          6282 => x"d3",
          6283 => x"2e",
          6284 => x"80",
          6285 => x"74",
          6286 => x"81",
          6287 => x"ef",
          6288 => x"17",
          6289 => x"06",
          6290 => x"34",
          6291 => x"17",
          6292 => x"80",
          6293 => x"1c",
          6294 => x"84",
          6295 => x"08",
          6296 => x"e4",
          6297 => x"08",
          6298 => x"34",
          6299 => x"6a",
          6300 => x"88",
          6301 => x"33",
          6302 => x"69",
          6303 => x"57",
          6304 => x"fe",
          6305 => x"56",
          6306 => x"0d",
          6307 => x"ec",
          6308 => x"80",
          6309 => x"90",
          6310 => x"7a",
          6311 => x"34",
          6312 => x"b8",
          6313 => x"7b",
          6314 => x"77",
          6315 => x"69",
          6316 => x"57",
          6317 => x"fe",
          6318 => x"56",
          6319 => x"3d",
          6320 => x"79",
          6321 => x"05",
          6322 => x"75",
          6323 => x"38",
          6324 => x"53",
          6325 => x"3d",
          6326 => x"e4",
          6327 => x"2e",
          6328 => x"b1",
          6329 => x"b2",
          6330 => x"59",
          6331 => x"08",
          6332 => x"02",
          6333 => x"5d",
          6334 => x"92",
          6335 => x"75",
          6336 => x"81",
          6337 => x"ef",
          6338 => x"58",
          6339 => x"33",
          6340 => x"15",
          6341 => x"52",
          6342 => x"b8",
          6343 => x"85",
          6344 => x"81",
          6345 => x"0c",
          6346 => x"11",
          6347 => x"74",
          6348 => x"81",
          6349 => x"7a",
          6350 => x"83",
          6351 => x"5f",
          6352 => x"33",
          6353 => x"9f",
          6354 => x"89",
          6355 => x"57",
          6356 => x"26",
          6357 => x"06",
          6358 => x"59",
          6359 => x"85",
          6360 => x"32",
          6361 => x"7a",
          6362 => x"95",
          6363 => x"7b",
          6364 => x"7e",
          6365 => x"24",
          6366 => x"53",
          6367 => x"3d",
          6368 => x"e4",
          6369 => x"b2",
          6370 => x"08",
          6371 => x"77",
          6372 => x"e4",
          6373 => x"92",
          6374 => x"02",
          6375 => x"5a",
          6376 => x"70",
          6377 => x"79",
          6378 => x"8b",
          6379 => x"2a",
          6380 => x"75",
          6381 => x"7f",
          6382 => x"18",
          6383 => x"5c",
          6384 => x"3d",
          6385 => x"9b",
          6386 => x"2b",
          6387 => x"7d",
          6388 => x"9c",
          6389 => x"7d",
          6390 => x"76",
          6391 => x"5e",
          6392 => x"7a",
          6393 => x"aa",
          6394 => x"bc",
          6395 => x"52",
          6396 => x"3f",
          6397 => x"38",
          6398 => x"0c",
          6399 => x"56",
          6400 => x"5a",
          6401 => x"38",
          6402 => x"56",
          6403 => x"2a",
          6404 => x"33",
          6405 => x"93",
          6406 => x"ec",
          6407 => x"80",
          6408 => x"83",
          6409 => x"b2",
          6410 => x"2e",
          6411 => x"fb",
          6412 => x"84",
          6413 => x"16",
          6414 => x"b4",
          6415 => x"16",
          6416 => x"09",
          6417 => x"76",
          6418 => x"51",
          6419 => x"08",
          6420 => x"58",
          6421 => x"aa",
          6422 => x"34",
          6423 => x"08",
          6424 => x"51",
          6425 => x"08",
          6426 => x"ff",
          6427 => x"f9",
          6428 => x"38",
          6429 => x"b8",
          6430 => x"3d",
          6431 => x"0c",
          6432 => x"94",
          6433 => x"2b",
          6434 => x"8d",
          6435 => x"fb",
          6436 => x"2e",
          6437 => x"0c",
          6438 => x"16",
          6439 => x"51",
          6440 => x"b8",
          6441 => x"fe",
          6442 => x"17",
          6443 => x"31",
          6444 => x"a0",
          6445 => x"16",
          6446 => x"06",
          6447 => x"08",
          6448 => x"81",
          6449 => x"79",
          6450 => x"17",
          6451 => x"18",
          6452 => x"81",
          6453 => x"38",
          6454 => x"b4",
          6455 => x"b8",
          6456 => x"08",
          6457 => x"5d",
          6458 => x"81",
          6459 => x"18",
          6460 => x"33",
          6461 => x"fb",
          6462 => x"df",
          6463 => x"05",
          6464 => x"cc",
          6465 => x"d8",
          6466 => x"b8",
          6467 => x"84",
          6468 => x"78",
          6469 => x"51",
          6470 => x"08",
          6471 => x"02",
          6472 => x"54",
          6473 => x"06",
          6474 => x"06",
          6475 => x"55",
          6476 => x"0b",
          6477 => x"9a",
          6478 => x"e4",
          6479 => x"0d",
          6480 => x"05",
          6481 => x"3f",
          6482 => x"e4",
          6483 => x"b8",
          6484 => x"5a",
          6485 => x"ff",
          6486 => x"55",
          6487 => x"80",
          6488 => x"86",
          6489 => x"22",
          6490 => x"59",
          6491 => x"88",
          6492 => x"90",
          6493 => x"98",
          6494 => x"57",
          6495 => x"fe",
          6496 => x"84",
          6497 => x"e8",
          6498 => x"53",
          6499 => x"51",
          6500 => x"08",
          6501 => x"b8",
          6502 => x"57",
          6503 => x"76",
          6504 => x"76",
          6505 => x"5b",
          6506 => x"70",
          6507 => x"81",
          6508 => x"56",
          6509 => x"82",
          6510 => x"55",
          6511 => x"98",
          6512 => x"52",
          6513 => x"3f",
          6514 => x"38",
          6515 => x"0c",
          6516 => x"33",
          6517 => x"2e",
          6518 => x"2e",
          6519 => x"05",
          6520 => x"90",
          6521 => x"33",
          6522 => x"71",
          6523 => x"59",
          6524 => x"3d",
          6525 => x"52",
          6526 => x"8b",
          6527 => x"b8",
          6528 => x"76",
          6529 => x"38",
          6530 => x"39",
          6531 => x"16",
          6532 => x"fe",
          6533 => x"e4",
          6534 => x"e8",
          6535 => x"34",
          6536 => x"84",
          6537 => x"17",
          6538 => x"33",
          6539 => x"fe",
          6540 => x"a0",
          6541 => x"16",
          6542 => x"59",
          6543 => x"81",
          6544 => x"84",
          6545 => x"38",
          6546 => x"fe",
          6547 => x"57",
          6548 => x"84",
          6549 => x"66",
          6550 => x"7c",
          6551 => x"34",
          6552 => x"38",
          6553 => x"34",
          6554 => x"18",
          6555 => x"79",
          6556 => x"79",
          6557 => x"82",
          6558 => x"a2",
          6559 => x"b8",
          6560 => x"82",
          6561 => x"57",
          6562 => x"34",
          6563 => x"a3",
          6564 => x"06",
          6565 => x"81",
          6566 => x"5c",
          6567 => x"55",
          6568 => x"74",
          6569 => x"74",
          6570 => x"84",
          6571 => x"84",
          6572 => x"57",
          6573 => x"e5",
          6574 => x"81",
          6575 => x"2e",
          6576 => x"2e",
          6577 => x"81",
          6578 => x"2e",
          6579 => x"06",
          6580 => x"78",
          6581 => x"81",
          6582 => x"38",
          6583 => x"88",
          6584 => x"5d",
          6585 => x"81",
          6586 => x"08",
          6587 => x"58",
          6588 => x"38",
          6589 => x"81",
          6590 => x"99",
          6591 => x"70",
          6592 => x"81",
          6593 => x"ed",
          6594 => x"95",
          6595 => x"3f",
          6596 => x"e4",
          6597 => x"75",
          6598 => x"04",
          6599 => x"3f",
          6600 => x"06",
          6601 => x"75",
          6602 => x"04",
          6603 => x"39",
          6604 => x"3f",
          6605 => x"e4",
          6606 => x"82",
          6607 => x"55",
          6608 => x"70",
          6609 => x"74",
          6610 => x"1e",
          6611 => x"84",
          6612 => x"87",
          6613 => x"86",
          6614 => x"08",
          6615 => x"38",
          6616 => x"38",
          6617 => x"fe",
          6618 => x"57",
          6619 => x"81",
          6620 => x"08",
          6621 => x"57",
          6622 => x"b2",
          6623 => x"2e",
          6624 => x"54",
          6625 => x"33",
          6626 => x"e4",
          6627 => x"81",
          6628 => x"78",
          6629 => x"33",
          6630 => x"81",
          6631 => x"78",
          6632 => x"d7",
          6633 => x"a5",
          6634 => x"a1",
          6635 => x"b8",
          6636 => x"87",
          6637 => x"76",
          6638 => x"57",
          6639 => x"34",
          6640 => x"56",
          6641 => x"7e",
          6642 => x"58",
          6643 => x"ff",
          6644 => x"38",
          6645 => x"70",
          6646 => x"74",
          6647 => x"e5",
          6648 => x"1e",
          6649 => x"84",
          6650 => x"81",
          6651 => x"18",
          6652 => x"51",
          6653 => x"08",
          6654 => x"38",
          6655 => x"b4",
          6656 => x"7b",
          6657 => x"18",
          6658 => x"84",
          6659 => x"74",
          6660 => x"d1",
          6661 => x"b8",
          6662 => x"fe",
          6663 => x"80",
          6664 => x"81",
          6665 => x"05",
          6666 => x"fe",
          6667 => x"3d",
          6668 => x"cb",
          6669 => x"76",
          6670 => x"74",
          6671 => x"73",
          6672 => x"84",
          6673 => x"81",
          6674 => x"81",
          6675 => x"81",
          6676 => x"38",
          6677 => x"17",
          6678 => x"5d",
          6679 => x"8a",
          6680 => x"7c",
          6681 => x"3f",
          6682 => x"72",
          6683 => x"05",
          6684 => x"55",
          6685 => x"19",
          6686 => x"77",
          6687 => x"76",
          6688 => x"7f",
          6689 => x"83",
          6690 => x"81",
          6691 => x"08",
          6692 => x"e4",
          6693 => x"78",
          6694 => x"09",
          6695 => x"54",
          6696 => x"0d",
          6697 => x"90",
          6698 => x"fe",
          6699 => x"81",
          6700 => x"77",
          6701 => x"80",
          6702 => x"58",
          6703 => x"54",
          6704 => x"53",
          6705 => x"3f",
          6706 => x"e4",
          6707 => x"ff",
          6708 => x"7e",
          6709 => x"2e",
          6710 => x"79",
          6711 => x"c0",
          6712 => x"15",
          6713 => x"5a",
          6714 => x"7d",
          6715 => x"81",
          6716 => x"54",
          6717 => x"39",
          6718 => x"82",
          6719 => x"c0",
          6720 => x"84",
          6721 => x"3d",
          6722 => x"81",
          6723 => x"0b",
          6724 => x"79",
          6725 => x"81",
          6726 => x"56",
          6727 => x"ed",
          6728 => x"84",
          6729 => x"84",
          6730 => x"ac",
          6731 => x"2e",
          6732 => x"84",
          6733 => x"12",
          6734 => x"51",
          6735 => x"08",
          6736 => x"56",
          6737 => x"82",
          6738 => x"84",
          6739 => x"83",
          6740 => x"84",
          6741 => x"55",
          6742 => x"82",
          6743 => x"15",
          6744 => x"7e",
          6745 => x"26",
          6746 => x"26",
          6747 => x"55",
          6748 => x"a6",
          6749 => x"77",
          6750 => x"85",
          6751 => x"77",
          6752 => x"b0",
          6753 => x"81",
          6754 => x"fe",
          6755 => x"e4",
          6756 => x"05",
          6757 => x"88",
          6758 => x"82",
          6759 => x"f8",
          6760 => x"b2",
          6761 => x"82",
          6762 => x"33",
          6763 => x"88",
          6764 => x"07",
          6765 => x"ba",
          6766 => x"71",
          6767 => x"14",
          6768 => x"33",
          6769 => x"a3",
          6770 => x"54",
          6771 => x"4d",
          6772 => x"90",
          6773 => x"82",
          6774 => x"06",
          6775 => x"38",
          6776 => x"89",
          6777 => x"f4",
          6778 => x"43",
          6779 => x"38",
          6780 => x"81",
          6781 => x"74",
          6782 => x"98",
          6783 => x"82",
          6784 => x"80",
          6785 => x"38",
          6786 => x"3f",
          6787 => x"55",
          6788 => x"96",
          6789 => x"10",
          6790 => x"72",
          6791 => x"ff",
          6792 => x"47",
          6793 => x"11",
          6794 => x"58",
          6795 => x"b8",
          6796 => x"16",
          6797 => x"26",
          6798 => x"31",
          6799 => x"fd",
          6800 => x"40",
          6801 => x"82",
          6802 => x"83",
          6803 => x"27",
          6804 => x"77",
          6805 => x"ef",
          6806 => x"57",
          6807 => x"0d",
          6808 => x"fb",
          6809 => x"0c",
          6810 => x"04",
          6811 => x"06",
          6812 => x"38",
          6813 => x"05",
          6814 => x"38",
          6815 => x"7d",
          6816 => x"05",
          6817 => x"33",
          6818 => x"99",
          6819 => x"ff",
          6820 => x"64",
          6821 => x"81",
          6822 => x"9f",
          6823 => x"81",
          6824 => x"75",
          6825 => x"9f",
          6826 => x"80",
          6827 => x"1f",
          6828 => x"38",
          6829 => x"f8",
          6830 => x"ca",
          6831 => x"08",
          6832 => x"06",
          6833 => x"83",
          6834 => x"7e",
          6835 => x"31",
          6836 => x"d2",
          6837 => x"7b",
          6838 => x"39",
          6839 => x"80",
          6840 => x"30",
          6841 => x"b8",
          6842 => x"7a",
          6843 => x"7b",
          6844 => x"84",
          6845 => x"b8",
          6846 => x"2e",
          6847 => x"8b",
          6848 => x"7a",
          6849 => x"55",
          6850 => x"ff",
          6851 => x"83",
          6852 => x"81",
          6853 => x"58",
          6854 => x"60",
          6855 => x"61",
          6856 => x"34",
          6857 => x"61",
          6858 => x"7b",
          6859 => x"05",
          6860 => x"48",
          6861 => x"2a",
          6862 => x"34",
          6863 => x"86",
          6864 => x"55",
          6865 => x"2a",
          6866 => x"61",
          6867 => x"34",
          6868 => x"9a",
          6869 => x"7e",
          6870 => x"48",
          6871 => x"2a",
          6872 => x"98",
          6873 => x"f0",
          6874 => x"2e",
          6875 => x"34",
          6876 => x"a9",
          6877 => x"34",
          6878 => x"61",
          6879 => x"6a",
          6880 => x"a4",
          6881 => x"93",
          6882 => x"57",
          6883 => x"76",
          6884 => x"55",
          6885 => x"49",
          6886 => x"05",
          6887 => x"7e",
          6888 => x"8f",
          6889 => x"fa",
          6890 => x"2e",
          6891 => x"80",
          6892 => x"15",
          6893 => x"5b",
          6894 => x"ff",
          6895 => x"38",
          6896 => x"2a",
          6897 => x"05",
          6898 => x"64",
          6899 => x"2a",
          6900 => x"59",
          6901 => x"78",
          6902 => x"fe",
          6903 => x"85",
          6904 => x"80",
          6905 => x"15",
          6906 => x"7a",
          6907 => x"81",
          6908 => x"38",
          6909 => x"66",
          6910 => x"38",
          6911 => x"52",
          6912 => x"b8",
          6913 => x"76",
          6914 => x"8c",
          6915 => x"58",
          6916 => x"84",
          6917 => x"58",
          6918 => x"81",
          6919 => x"80",
          6920 => x"05",
          6921 => x"38",
          6922 => x"34",
          6923 => x"34",
          6924 => x"82",
          6925 => x"77",
          6926 => x"fd",
          6927 => x"ab",
          6928 => x"b8",
          6929 => x"76",
          6930 => x"08",
          6931 => x"c6",
          6932 => x"34",
          6933 => x"b8",
          6934 => x"62",
          6935 => x"2a",
          6936 => x"62",
          6937 => x"05",
          6938 => x"83",
          6939 => x"60",
          6940 => x"81",
          6941 => x"38",
          6942 => x"c3",
          6943 => x"08",
          6944 => x"84",
          6945 => x"b8",
          6946 => x"39",
          6947 => x"c4",
          6948 => x"57",
          6949 => x"58",
          6950 => x"26",
          6951 => x"10",
          6952 => x"74",
          6953 => x"ee",
          6954 => x"d3",
          6955 => x"84",
          6956 => x"a0",
          6957 => x"fc",
          6958 => x"f0",
          6959 => x"57",
          6960 => x"83",
          6961 => x"f8",
          6962 => x"f4",
          6963 => x"68",
          6964 => x"af",
          6965 => x"61",
          6966 => x"68",
          6967 => x"5b",
          6968 => x"2a",
          6969 => x"c6",
          6970 => x"80",
          6971 => x"80",
          6972 => x"c6",
          6973 => x"7c",
          6974 => x"34",
          6975 => x"05",
          6976 => x"a7",
          6977 => x"80",
          6978 => x"05",
          6979 => x"61",
          6980 => x"34",
          6981 => x"b3",
          6982 => x"05",
          6983 => x"93",
          6984 => x"59",
          6985 => x"33",
          6986 => x"15",
          6987 => x"76",
          6988 => x"81",
          6989 => x"da",
          6990 => x"53",
          6991 => x"3f",
          6992 => x"b0",
          6993 => x"77",
          6994 => x"84",
          6995 => x"51",
          6996 => x"81",
          6997 => x"0d",
          6998 => x"34",
          6999 => x"4c",
          7000 => x"34",
          7001 => x"34",
          7002 => x"86",
          7003 => x"ff",
          7004 => x"05",
          7005 => x"65",
          7006 => x"54",
          7007 => x"fe",
          7008 => x"57",
          7009 => x"ff",
          7010 => x"80",
          7011 => x"7b",
          7012 => x"57",
          7013 => x"57",
          7014 => x"61",
          7015 => x"83",
          7016 => x"e6",
          7017 => x"05",
          7018 => x"83",
          7019 => x"78",
          7020 => x"2a",
          7021 => x"7a",
          7022 => x"05",
          7023 => x"76",
          7024 => x"83",
          7025 => x"05",
          7026 => x"6b",
          7027 => x"52",
          7028 => x"54",
          7029 => x"fe",
          7030 => x"f7",
          7031 => x"5b",
          7032 => x"57",
          7033 => x"3d",
          7034 => x"53",
          7035 => x"3f",
          7036 => x"38",
          7037 => x"90",
          7038 => x"34",
          7039 => x"38",
          7040 => x"34",
          7041 => x"74",
          7042 => x"04",
          7043 => x"b3",
          7044 => x"80",
          7045 => x"76",
          7046 => x"17",
          7047 => x"81",
          7048 => x"74",
          7049 => x"0c",
          7050 => x"05",
          7051 => x"08",
          7052 => x"32",
          7053 => x"70",
          7054 => x"1b",
          7055 => x"52",
          7056 => x"39",
          7057 => x"33",
          7058 => x"57",
          7059 => x"34",
          7060 => x"3d",
          7061 => x"f7",
          7062 => x"c0",
          7063 => x"59",
          7064 => x"bb",
          7065 => x"81",
          7066 => x"75",
          7067 => x"11",
          7068 => x"08",
          7069 => x"e4",
          7070 => x"38",
          7071 => x"3d",
          7072 => x"55",
          7073 => x"51",
          7074 => x"70",
          7075 => x"30",
          7076 => x"8d",
          7077 => x"81",
          7078 => x"3d",
          7079 => x"84",
          7080 => x"52",
          7081 => x"83",
          7082 => x"e4",
          7083 => x"ff",
          7084 => x"09",
          7085 => x"e4",
          7086 => x"71",
          7087 => x"ff",
          7088 => x"26",
          7089 => x"05",
          7090 => x"80",
          7091 => x"e4",
          7092 => x"3d",
          7093 => x"05",
          7094 => x"70",
          7095 => x"72",
          7096 => x"04",
          7097 => x"ef",
          7098 => x"70",
          7099 => x"84",
          7100 => x"04",
          7101 => x"ff",
          7102 => x"ff",
          7103 => x"75",
          7104 => x"70",
          7105 => x"70",
          7106 => x"56",
          7107 => x"82",
          7108 => x"54",
          7109 => x"54",
          7110 => x"38",
          7111 => x"52",
          7112 => x"75",
          7113 => x"80",
          7114 => x"b8",
          7115 => x"ec",
          7116 => x"26",
          7117 => x"d0",
          7118 => x"16",
          7119 => x"75",
          7120 => x"83",
          7121 => x"88",
          7122 => x"51",
          7123 => x"ff",
          7124 => x"70",
          7125 => x"39",
          7126 => x"57",
          7127 => x"ff",
          7128 => x"75",
          7129 => x"70",
          7130 => x"ff",
          7131 => x"05",
          7132 => x"00",
          7133 => x"00",
          7134 => x"ff",
          7135 => x"00",
          7136 => x"00",
          7137 => x"00",
          7138 => x"00",
          7139 => x"00",
          7140 => x"00",
          7141 => x"00",
          7142 => x"00",
          7143 => x"00",
          7144 => x"00",
          7145 => x"00",
          7146 => x"00",
          7147 => x"00",
          7148 => x"00",
          7149 => x"00",
          7150 => x"00",
          7151 => x"00",
          7152 => x"00",
          7153 => x"00",
          7154 => x"00",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"69",
          7372 => x"69",
          7373 => x"69",
          7374 => x"6c",
          7375 => x"65",
          7376 => x"63",
          7377 => x"63",
          7378 => x"64",
          7379 => x"64",
          7380 => x"65",
          7381 => x"65",
          7382 => x"69",
          7383 => x"66",
          7384 => x"00",
          7385 => x"65",
          7386 => x"65",
          7387 => x"6e",
          7388 => x"65",
          7389 => x"6c",
          7390 => x"62",
          7391 => x"62",
          7392 => x"69",
          7393 => x"64",
          7394 => x"77",
          7395 => x"2e",
          7396 => x"65",
          7397 => x"63",
          7398 => x"00",
          7399 => x"61",
          7400 => x"20",
          7401 => x"00",
          7402 => x"66",
          7403 => x"6d",
          7404 => x"00",
          7405 => x"69",
          7406 => x"64",
          7407 => x"75",
          7408 => x"61",
          7409 => x"6e",
          7410 => x"00",
          7411 => x"74",
          7412 => x"64",
          7413 => x"6d",
          7414 => x"20",
          7415 => x"74",
          7416 => x"64",
          7417 => x"6b",
          7418 => x"6e",
          7419 => x"6c",
          7420 => x"72",
          7421 => x"62",
          7422 => x"6e",
          7423 => x"00",
          7424 => x"20",
          7425 => x"72",
          7426 => x"2e",
          7427 => x"68",
          7428 => x"6e",
          7429 => x"00",
          7430 => x"61",
          7431 => x"65",
          7432 => x"00",
          7433 => x"73",
          7434 => x"2e",
          7435 => x"69",
          7436 => x"61",
          7437 => x"6f",
          7438 => x"6f",
          7439 => x"6f",
          7440 => x"6f",
          7441 => x"69",
          7442 => x"72",
          7443 => x"6e",
          7444 => x"65",
          7445 => x"69",
          7446 => x"72",
          7447 => x"73",
          7448 => x"25",
          7449 => x"73",
          7450 => x"25",
          7451 => x"73",
          7452 => x"00",
          7453 => x"00",
          7454 => x"00",
          7455 => x"30",
          7456 => x"7c",
          7457 => x"20",
          7458 => x"00",
          7459 => x"20",
          7460 => x"4f",
          7461 => x"20",
          7462 => x"2f",
          7463 => x"31",
          7464 => x"5a",
          7465 => x"20",
          7466 => x"73",
          7467 => x"0a",
          7468 => x"6e",
          7469 => x"20",
          7470 => x"00",
          7471 => x"20",
          7472 => x"72",
          7473 => x"41",
          7474 => x"69",
          7475 => x"74",
          7476 => x"20",
          7477 => x"72",
          7478 => x"41",
          7479 => x"69",
          7480 => x"74",
          7481 => x"20",
          7482 => x"72",
          7483 => x"4f",
          7484 => x"69",
          7485 => x"74",
          7486 => x"6e",
          7487 => x"00",
          7488 => x"20",
          7489 => x"70",
          7490 => x"6e",
          7491 => x"6d",
          7492 => x"6e",
          7493 => x"74",
          7494 => x"00",
          7495 => x"78",
          7496 => x"00",
          7497 => x"70",
          7498 => x"61",
          7499 => x"20",
          7500 => x"69",
          7501 => x"61",
          7502 => x"6c",
          7503 => x"69",
          7504 => x"6c",
          7505 => x"20",
          7506 => x"73",
          7507 => x"61",
          7508 => x"6e",
          7509 => x"50",
          7510 => x"64",
          7511 => x"2e",
          7512 => x"6f",
          7513 => x"6f",
          7514 => x"00",
          7515 => x"72",
          7516 => x"70",
          7517 => x"6e",
          7518 => x"61",
          7519 => x"6f",
          7520 => x"38",
          7521 => x"00",
          7522 => x"72",
          7523 => x"20",
          7524 => x"64",
          7525 => x"78",
          7526 => x"20",
          7527 => x"25",
          7528 => x"2e",
          7529 => x"20",
          7530 => x"00",
          7531 => x"20",
          7532 => x"6f",
          7533 => x"2e",
          7534 => x"30",
          7535 => x"78",
          7536 => x"78",
          7537 => x"00",
          7538 => x"6e",
          7539 => x"30",
          7540 => x"58",
          7541 => x"69",
          7542 => x"00",
          7543 => x"4d",
          7544 => x"43",
          7545 => x"2e",
          7546 => x"73",
          7547 => x"65",
          7548 => x"68",
          7549 => x"20",
          7550 => x"70",
          7551 => x"63",
          7552 => x"00",
          7553 => x"64",
          7554 => x"25",
          7555 => x"2e",
          7556 => x"6f",
          7557 => x"67",
          7558 => x"00",
          7559 => x"69",
          7560 => x"6c",
          7561 => x"3a",
          7562 => x"73",
          7563 => x"20",
          7564 => x"65",
          7565 => x"74",
          7566 => x"65",
          7567 => x"38",
          7568 => x"20",
          7569 => x"65",
          7570 => x"61",
          7571 => x"65",
          7572 => x"38",
          7573 => x"20",
          7574 => x"20",
          7575 => x"64",
          7576 => x"20",
          7577 => x"38",
          7578 => x"69",
          7579 => x"20",
          7580 => x"64",
          7581 => x"20",
          7582 => x"20",
          7583 => x"34",
          7584 => x"20",
          7585 => x"6d",
          7586 => x"46",
          7587 => x"20",
          7588 => x"2e",
          7589 => x"0a",
          7590 => x"69",
          7591 => x"53",
          7592 => x"6f",
          7593 => x"3d",
          7594 => x"64",
          7595 => x"20",
          7596 => x"20",
          7597 => x"72",
          7598 => x"20",
          7599 => x"2e",
          7600 => x"0a",
          7601 => x"50",
          7602 => x"53",
          7603 => x"4f",
          7604 => x"20",
          7605 => x"43",
          7606 => x"49",
          7607 => x"42",
          7608 => x"20",
          7609 => x"43",
          7610 => x"61",
          7611 => x"30",
          7612 => x"20",
          7613 => x"31",
          7614 => x"6d",
          7615 => x"30",
          7616 => x"20",
          7617 => x"52",
          7618 => x"76",
          7619 => x"30",
          7620 => x"20",
          7621 => x"20",
          7622 => x"38",
          7623 => x"2e",
          7624 => x"52",
          7625 => x"20",
          7626 => x"30",
          7627 => x"20",
          7628 => x"42",
          7629 => x"38",
          7630 => x"2e",
          7631 => x"44",
          7632 => x"20",
          7633 => x"30",
          7634 => x"20",
          7635 => x"52",
          7636 => x"38",
          7637 => x"2e",
          7638 => x"6d",
          7639 => x"6e",
          7640 => x"6e",
          7641 => x"56",
          7642 => x"6d",
          7643 => x"65",
          7644 => x"6c",
          7645 => x"56",
          7646 => x"00",
          7647 => x"00",
          7648 => x"00",
          7649 => x"00",
          7650 => x"00",
          7651 => x"00",
          7652 => x"00",
          7653 => x"00",
          7654 => x"00",
          7655 => x"00",
          7656 => x"00",
          7657 => x"00",
          7658 => x"00",
          7659 => x"00",
          7660 => x"00",
          7661 => x"00",
          7662 => x"00",
          7663 => x"00",
          7664 => x"00",
          7665 => x"00",
          7666 => x"00",
          7667 => x"00",
          7668 => x"00",
          7669 => x"00",
          7670 => x"00",
          7671 => x"00",
          7672 => x"00",
          7673 => x"00",
          7674 => x"00",
          7675 => x"00",
          7676 => x"00",
          7677 => x"00",
          7678 => x"00",
          7679 => x"5b",
          7680 => x"5b",
          7681 => x"5b",
          7682 => x"30",
          7683 => x"5b",
          7684 => x"00",
          7685 => x"00",
          7686 => x"00",
          7687 => x"00",
          7688 => x"00",
          7689 => x"00",
          7690 => x"74",
          7691 => x"72",
          7692 => x"73",
          7693 => x"6c",
          7694 => x"62",
          7695 => x"69",
          7696 => x"69",
          7697 => x"00",
          7698 => x"20",
          7699 => x"61",
          7700 => x"20",
          7701 => x"68",
          7702 => x"72",
          7703 => x"74",
          7704 => x"00",
          7705 => x"00",
          7706 => x"00",
          7707 => x"5b",
          7708 => x"5b",
          7709 => x"00",
          7710 => x"00",
          7711 => x"00",
          7712 => x"00",
          7713 => x"00",
          7714 => x"00",
          7715 => x"00",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"00",
          7721 => x"5b",
          7722 => x"5b",
          7723 => x"3a",
          7724 => x"64",
          7725 => x"25",
          7726 => x"00",
          7727 => x"25",
          7728 => x"3a",
          7729 => x"64",
          7730 => x"3a",
          7731 => x"30",
          7732 => x"63",
          7733 => x"00",
          7734 => x"74",
          7735 => x"3a",
          7736 => x"32",
          7737 => x"00",
          7738 => x"32",
          7739 => x"00",
          7740 => x"32",
          7741 => x"6f",
          7742 => x"65",
          7743 => x"00",
          7744 => x"2a",
          7745 => x"00",
          7746 => x"5d",
          7747 => x"41",
          7748 => x"fe",
          7749 => x"2e",
          7750 => x"4d",
          7751 => x"54",
          7752 => x"4f",
          7753 => x"20",
          7754 => x"20",
          7755 => x"00",
          7756 => x"00",
          7757 => x"0e",
          7758 => x"00",
          7759 => x"41",
          7760 => x"49",
          7761 => x"4f",
          7762 => x"9d",
          7763 => x"a5",
          7764 => x"ad",
          7765 => x"b5",
          7766 => x"bd",
          7767 => x"c5",
          7768 => x"cd",
          7769 => x"d5",
          7770 => x"dd",
          7771 => x"e5",
          7772 => x"ed",
          7773 => x"f5",
          7774 => x"fd",
          7775 => x"5b",
          7776 => x"3e",
          7777 => x"01",
          7778 => x"00",
          7779 => x"01",
          7780 => x"10",
          7781 => x"c7",
          7782 => x"e4",
          7783 => x"ea",
          7784 => x"ee",
          7785 => x"c9",
          7786 => x"f6",
          7787 => x"ff",
          7788 => x"a3",
          7789 => x"e1",
          7790 => x"f1",
          7791 => x"bf",
          7792 => x"bc",
          7793 => x"91",
          7794 => x"24",
          7795 => x"55",
          7796 => x"5d",
          7797 => x"14",
          7798 => x"00",
          7799 => x"5a",
          7800 => x"60",
          7801 => x"68",
          7802 => x"58",
          7803 => x"6a",
          7804 => x"84",
          7805 => x"b1",
          7806 => x"a3",
          7807 => x"a6",
          7808 => x"1e",
          7809 => x"61",
          7810 => x"20",
          7811 => x"b0",
          7812 => x"7f",
          7813 => x"61",
          7814 => x"f8",
          7815 => x"78",
          7816 => x"06",
          7817 => x"2e",
          7818 => x"4d",
          7819 => x"82",
          7820 => x"87",
          7821 => x"8b",
          7822 => x"8f",
          7823 => x"93",
          7824 => x"97",
          7825 => x"9b",
          7826 => x"9f",
          7827 => x"a2",
          7828 => x"a7",
          7829 => x"ab",
          7830 => x"af",
          7831 => x"b3",
          7832 => x"b7",
          7833 => x"bb",
          7834 => x"f7",
          7835 => x"c3",
          7836 => x"c7",
          7837 => x"cb",
          7838 => x"dd",
          7839 => x"12",
          7840 => x"f4",
          7841 => x"22",
          7842 => x"65",
          7843 => x"66",
          7844 => x"41",
          7845 => x"40",
          7846 => x"89",
          7847 => x"5a",
          7848 => x"5e",
          7849 => x"62",
          7850 => x"66",
          7851 => x"6a",
          7852 => x"6e",
          7853 => x"9d",
          7854 => x"76",
          7855 => x"7a",
          7856 => x"7e",
          7857 => x"82",
          7858 => x"86",
          7859 => x"b1",
          7860 => x"8e",
          7861 => x"b7",
          7862 => x"fe",
          7863 => x"86",
          7864 => x"b1",
          7865 => x"a3",
          7866 => x"cc",
          7867 => x"8f",
          7868 => x"0a",
          7869 => x"f5",
          7870 => x"f9",
          7871 => x"20",
          7872 => x"22",
          7873 => x"0e",
          7874 => x"d0",
          7875 => x"00",
          7876 => x"63",
          7877 => x"5a",
          7878 => x"06",
          7879 => x"08",
          7880 => x"07",
          7881 => x"54",
          7882 => x"60",
          7883 => x"ba",
          7884 => x"ca",
          7885 => x"f8",
          7886 => x"fa",
          7887 => x"90",
          7888 => x"b0",
          7889 => x"b2",
          7890 => x"c3",
          7891 => x"02",
          7892 => x"f3",
          7893 => x"01",
          7894 => x"84",
          7895 => x"1a",
          7896 => x"02",
          7897 => x"02",
          7898 => x"26",
          7899 => x"00",
          7900 => x"02",
          7901 => x"00",
          7902 => x"04",
          7903 => x"00",
          7904 => x"14",
          7905 => x"00",
          7906 => x"2b",
          7907 => x"00",
          7908 => x"30",
          7909 => x"00",
          7910 => x"3c",
          7911 => x"00",
          7912 => x"3d",
          7913 => x"00",
          7914 => x"3f",
          7915 => x"00",
          7916 => x"40",
          7917 => x"00",
          7918 => x"41",
          7919 => x"00",
          7920 => x"42",
          7921 => x"00",
          7922 => x"43",
          7923 => x"00",
          7924 => x"50",
          7925 => x"00",
          7926 => x"51",
          7927 => x"00",
          7928 => x"54",
          7929 => x"00",
          7930 => x"55",
          7931 => x"00",
          7932 => x"79",
          7933 => x"00",
          7934 => x"78",
          7935 => x"00",
          7936 => x"82",
          7937 => x"00",
          7938 => x"83",
          7939 => x"00",
          7940 => x"85",
          7941 => x"00",
          7942 => x"87",
          7943 => x"00",
          7944 => x"88",
          7945 => x"00",
          7946 => x"89",
          7947 => x"00",
          7948 => x"8c",
          7949 => x"00",
          7950 => x"8d",
          7951 => x"00",
          7952 => x"8e",
          7953 => x"00",
          7954 => x"8f",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"01",
          7959 => x"01",
          7960 => x"00",
          7961 => x"00",
          7962 => x"00",
          7963 => x"f5",
          7964 => x"f5",
          7965 => x"01",
          7966 => x"01",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"01",
          7983 => x"3b",
          7984 => x"f0",
          7985 => x"76",
          7986 => x"6e",
          7987 => x"66",
          7988 => x"36",
          7989 => x"39",
          7990 => x"f2",
          7991 => x"f0",
          7992 => x"f0",
          7993 => x"3a",
          7994 => x"f0",
          7995 => x"56",
          7996 => x"4e",
          7997 => x"46",
          7998 => x"36",
          7999 => x"39",
          8000 => x"f2",
          8001 => x"f0",
          8002 => x"f0",
          8003 => x"2b",
          8004 => x"f0",
          8005 => x"56",
          8006 => x"4e",
          8007 => x"46",
          8008 => x"26",
          8009 => x"29",
          8010 => x"f8",
          8011 => x"f0",
          8012 => x"f0",
          8013 => x"f0",
          8014 => x"f0",
          8015 => x"16",
          8016 => x"0e",
          8017 => x"06",
          8018 => x"f0",
          8019 => x"1f",
          8020 => x"f0",
          8021 => x"f0",
          8022 => x"f0",
          8023 => x"b5",
          8024 => x"f0",
          8025 => x"a6",
          8026 => x"33",
          8027 => x"43",
          8028 => x"1e",
          8029 => x"a3",
          8030 => x"c4",
          8031 => x"f0",
          8032 => x"f0",
          8033 => x"00",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"00",
          8045 => x"01",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"e0",
          9069 => x"f9",
          9070 => x"c1",
          9071 => x"e4",
          9072 => x"61",
          9073 => x"69",
          9074 => x"21",
          9075 => x"29",
          9076 => x"01",
          9077 => x"09",
          9078 => x"11",
          9079 => x"19",
          9080 => x"81",
          9081 => x"89",
          9082 => x"91",
          9083 => x"99",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"02",
          9100 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"00",
             3 => x"00",
             4 => x"88",
             5 => x"08",
             6 => x"04",
             7 => x"00",
             8 => x"71",
             9 => x"81",
            10 => x"ff",
            11 => x"00",
            12 => x"71",
            13 => x"83",
            14 => x"2b",
            15 => x"0b",
            16 => x"72",
            17 => x"09",
            18 => x"07",
            19 => x"00",
            20 => x"72",
            21 => x"51",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"09",
            26 => x"0a",
            27 => x"51",
            28 => x"72",
            29 => x"51",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"72",
            45 => x"0b",
            46 => x"00",
            47 => x"00",
            48 => x"72",
            49 => x"09",
            50 => x"06",
            51 => x"00",
            52 => x"71",
            53 => x"06",
            54 => x"0b",
            55 => x"51",
            56 => x"72",
            57 => x"81",
            58 => x"51",
            59 => x"00",
            60 => x"72",
            61 => x"81",
            62 => x"53",
            63 => x"00",
            64 => x"71",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"72",
            69 => x"04",
            70 => x"00",
            71 => x"00",
            72 => x"72",
            73 => x"07",
            74 => x"00",
            75 => x"00",
            76 => x"71",
            77 => x"81",
            78 => x"81",
            79 => x"00",
            80 => x"71",
            81 => x"e4",
            82 => x"06",
            83 => x"00",
            84 => x"88",
            85 => x"0b",
            86 => x"88",
            87 => x"0c",
            88 => x"88",
            89 => x"0b",
            90 => x"88",
            91 => x"0c",
            92 => x"72",
            93 => x"81",
            94 => x"73",
            95 => x"07",
            96 => x"72",
            97 => x"09",
            98 => x"06",
            99 => x"06",
           100 => x"05",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"04",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"71",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"04",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"02",
           117 => x"04",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"02",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"0b",
           134 => x"96",
           135 => x"0b",
           136 => x"0b",
           137 => x"d6",
           138 => x"0b",
           139 => x"0b",
           140 => x"96",
           141 => x"0b",
           142 => x"0b",
           143 => x"d7",
           144 => x"0b",
           145 => x"0b",
           146 => x"9b",
           147 => x"0b",
           148 => x"0b",
           149 => x"df",
           150 => x"0b",
           151 => x"0b",
           152 => x"a3",
           153 => x"0b",
           154 => x"0b",
           155 => x"e7",
           156 => x"0b",
           157 => x"0b",
           158 => x"ab",
           159 => x"0b",
           160 => x"0b",
           161 => x"ef",
           162 => x"0b",
           163 => x"0b",
           164 => x"b3",
           165 => x"0b",
           166 => x"0b",
           167 => x"f7",
           168 => x"0b",
           169 => x"0b",
           170 => x"bb",
           171 => x"0b",
           172 => x"0b",
           173 => x"fe",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"04",
           193 => x"0c",
           194 => x"08",
           195 => x"f0",
           196 => x"08",
           197 => x"f0",
           198 => x"08",
           199 => x"f0",
           200 => x"08",
           201 => x"f0",
           202 => x"08",
           203 => x"f0",
           204 => x"08",
           205 => x"f0",
           206 => x"08",
           207 => x"f0",
           208 => x"08",
           209 => x"f0",
           210 => x"08",
           211 => x"f0",
           212 => x"08",
           213 => x"f0",
           214 => x"08",
           215 => x"f0",
           216 => x"08",
           217 => x"f0",
           218 => x"f0",
           219 => x"b8",
           220 => x"b8",
           221 => x"84",
           222 => x"84",
           223 => x"04",
           224 => x"2d",
           225 => x"90",
           226 => x"9d",
           227 => x"80",
           228 => x"e2",
           229 => x"c0",
           230 => x"82",
           231 => x"80",
           232 => x"0c",
           233 => x"08",
           234 => x"f0",
           235 => x"f0",
           236 => x"b8",
           237 => x"b8",
           238 => x"84",
           239 => x"84",
           240 => x"04",
           241 => x"2d",
           242 => x"90",
           243 => x"fa",
           244 => x"80",
           245 => x"f3",
           246 => x"c0",
           247 => x"83",
           248 => x"80",
           249 => x"0c",
           250 => x"08",
           251 => x"f0",
           252 => x"f0",
           253 => x"b8",
           254 => x"b8",
           255 => x"84",
           256 => x"84",
           257 => x"04",
           258 => x"2d",
           259 => x"90",
           260 => x"bf",
           261 => x"80",
           262 => x"e3",
           263 => x"c0",
           264 => x"82",
           265 => x"80",
           266 => x"0c",
           267 => x"08",
           268 => x"f0",
           269 => x"f0",
           270 => x"b8",
           271 => x"b8",
           272 => x"84",
           273 => x"84",
           274 => x"04",
           275 => x"2d",
           276 => x"90",
           277 => x"81",
           278 => x"80",
           279 => x"b9",
           280 => x"c0",
           281 => x"83",
           282 => x"80",
           283 => x"0c",
           284 => x"08",
           285 => x"f0",
           286 => x"f0",
           287 => x"b8",
           288 => x"b8",
           289 => x"84",
           290 => x"84",
           291 => x"04",
           292 => x"2d",
           293 => x"90",
           294 => x"8a",
           295 => x"80",
           296 => x"9a",
           297 => x"80",
           298 => x"da",
           299 => x"c0",
           300 => x"81",
           301 => x"80",
           302 => x"0c",
           303 => x"08",
           304 => x"f0",
           305 => x"f0",
           306 => x"04",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"53",
           311 => x"06",
           312 => x"05",
           313 => x"06",
           314 => x"72",
           315 => x"05",
           316 => x"53",
           317 => x"04",
           318 => x"27",
           319 => x"53",
           320 => x"8c",
           321 => x"fc",
           322 => x"05",
           323 => x"d4",
           324 => x"3d",
           325 => x"7c",
           326 => x"80",
           327 => x"80",
           328 => x"80",
           329 => x"32",
           330 => x"51",
           331 => x"b7",
           332 => x"51",
           333 => x"53",
           334 => x"38",
           335 => x"05",
           336 => x"70",
           337 => x"54",
           338 => x"80",
           339 => x"e4",
           340 => x"84",
           341 => x"f5",
           342 => x"05",
           343 => x"58",
           344 => x"8d",
           345 => x"19",
           346 => x"04",
           347 => x"53",
           348 => x"3d",
           349 => x"65",
           350 => x"0c",
           351 => x"32",
           352 => x"72",
           353 => x"38",
           354 => x"c5",
           355 => x"5c",
           356 => x"17",
           357 => x"76",
           358 => x"51",
           359 => x"2e",
           360 => x"32",
           361 => x"9e",
           362 => x"33",
           363 => x"08",
           364 => x"3d",
           365 => x"10",
           366 => x"2b",
           367 => x"0a",
           368 => x"52",
           369 => x"81",
           370 => x"ff",
           371 => x"76",
           372 => x"a5",
           373 => x"73",
           374 => x"58",
           375 => x"39",
           376 => x"7b",
           377 => x"8d",
           378 => x"54",
           379 => x"06",
           380 => x"53",
           381 => x"10",
           382 => x"08",
           383 => x"d8",
           384 => x"51",
           385 => x"5b",
           386 => x"80",
           387 => x"7f",
           388 => x"ff",
           389 => x"b8",
           390 => x"9a",
           391 => x"06",
           392 => x"56",
           393 => x"b8",
           394 => x"70",
           395 => x"51",
           396 => x"56",
           397 => x"84",
           398 => x"06",
           399 => x"77",
           400 => x"05",
           401 => x"2a",
           402 => x"2e",
           403 => x"f8",
           404 => x"8b",
           405 => x"80",
           406 => x"7a",
           407 => x"72",
           408 => x"70",
           409 => x"24",
           410 => x"06",
           411 => x"56",
           412 => x"2e",
           413 => x"2b",
           414 => x"56",
           415 => x"38",
           416 => x"85",
           417 => x"54",
           418 => x"81",
           419 => x"81",
           420 => x"88",
           421 => x"b2",
           422 => x"fc",
           423 => x"40",
           424 => x"52",
           425 => x"84",
           426 => x"70",
           427 => x"24",
           428 => x"80",
           429 => x"0a",
           430 => x"2c",
           431 => x"38",
           432 => x"78",
           433 => x"0a",
           434 => x"74",
           435 => x"70",
           436 => x"81",
           437 => x"d8",
           438 => x"38",
           439 => x"7d",
           440 => x"52",
           441 => x"a5",
           442 => x"81",
           443 => x"7a",
           444 => x"84",
           445 => x"70",
           446 => x"25",
           447 => x"86",
           448 => x"5b",
           449 => x"76",
           450 => x"80",
           451 => x"60",
           452 => x"ff",
           453 => x"fb",
           454 => x"fe",
           455 => x"98",
           456 => x"29",
           457 => x"5e",
           458 => x"87",
           459 => x"fe",
           460 => x"29",
           461 => x"5a",
           462 => x"38",
           463 => x"e2",
           464 => x"06",
           465 => x"fe",
           466 => x"05",
           467 => x"39",
           468 => x"5b",
           469 => x"ab",
           470 => x"57",
           471 => x"75",
           472 => x"78",
           473 => x"05",
           474 => x"e3",
           475 => x"56",
           476 => x"39",
           477 => x"53",
           478 => x"df",
           479 => x"84",
           480 => x"84",
           481 => x"89",
           482 => x"5b",
           483 => x"f9",
           484 => x"05",
           485 => x"41",
           486 => x"87",
           487 => x"ff",
           488 => x"54",
           489 => x"39",
           490 => x"5b",
           491 => x"7f",
           492 => x"06",
           493 => x"38",
           494 => x"e4",
           495 => x"31",
           496 => x"81",
           497 => x"f7",
           498 => x"84",
           499 => x"70",
           500 => x"25",
           501 => x"83",
           502 => x"51",
           503 => x"81",
           504 => x"51",
           505 => x"06",
           506 => x"fa",
           507 => x"31",
           508 => x"80",
           509 => x"90",
           510 => x"51",
           511 => x"73",
           512 => x"39",
           513 => x"e5",
           514 => x"2e",
           515 => x"74",
           516 => x"53",
           517 => x"82",
           518 => x"51",
           519 => x"52",
           520 => x"e4",
           521 => x"31",
           522 => x"7a",
           523 => x"bf",
           524 => x"fe",
           525 => x"75",
           526 => x"3d",
           527 => x"80",
           528 => x"33",
           529 => x"06",
           530 => x"72",
           531 => x"38",
           532 => x"72",
           533 => x"08",
           534 => x"72",
           535 => x"83",
           536 => x"56",
           537 => x"84",
           538 => x"d4",
           539 => x"52",
           540 => x"2d",
           541 => x"38",
           542 => x"e4",
           543 => x"0d",
           544 => x"16",
           545 => x"81",
           546 => x"72",
           547 => x"73",
           548 => x"77",
           549 => x"56",
           550 => x"0d",
           551 => x"53",
           552 => x"72",
           553 => x"84",
           554 => x"ff",
           555 => x"57",
           556 => x"0d",
           557 => x"85",
           558 => x"0d",
           559 => x"2a",
           560 => x"57",
           561 => x"2a",
           562 => x"38",
           563 => x"08",
           564 => x"76",
           565 => x"8c",
           566 => x"0c",
           567 => x"88",
           568 => x"ff",
           569 => x"2d",
           570 => x"38",
           571 => x"0c",
           572 => x"77",
           573 => x"70",
           574 => x"56",
           575 => x"2a",
           576 => x"82",
           577 => x"80",
           578 => x"53",
           579 => x"13",
           580 => x"8c",
           581 => x"73",
           582 => x"04",
           583 => x"17",
           584 => x"17",
           585 => x"0c",
           586 => x"16",
           587 => x"08",
           588 => x"ff",
           589 => x"07",
           590 => x"2e",
           591 => x"85",
           592 => x"e4",
           593 => x"07",
           594 => x"ec",
           595 => x"54",
           596 => x"33",
           597 => x"72",
           598 => x"72",
           599 => x"38",
           600 => x"0d",
           601 => x"7a",
           602 => x"9d",
           603 => x"80",
           604 => x"53",
           605 => x"ff",
           606 => x"b8",
           607 => x"12",
           608 => x"14",
           609 => x"53",
           610 => x"51",
           611 => x"ff",
           612 => x"ff",
           613 => x"fe",
           614 => x"70",
           615 => x"38",
           616 => x"e4",
           617 => x"3d",
           618 => x"72",
           619 => x"72",
           620 => x"38",
           621 => x"0d",
           622 => x"79",
           623 => x"93",
           624 => x"73",
           625 => x"51",
           626 => x"0c",
           627 => x"76",
           628 => x"2e",
           629 => x"05",
           630 => x"09",
           631 => x"71",
           632 => x"72",
           633 => x"e4",
           634 => x"2e",
           635 => x"72",
           636 => x"52",
           637 => x"72",
           638 => x"3d",
           639 => x"86",
           640 => x"79",
           641 => x"84",
           642 => x"81",
           643 => x"84",
           644 => x"08",
           645 => x"08",
           646 => x"75",
           647 => x"b1",
           648 => x"84",
           649 => x"fd",
           650 => x"55",
           651 => x"72",
           652 => x"80",
           653 => x"ff",
           654 => x"13",
           655 => x"b8",
           656 => x"3d",
           657 => x"54",
           658 => x"72",
           659 => x"51",
           660 => x"0c",
           661 => x"78",
           662 => x"2e",
           663 => x"84",
           664 => x"73",
           665 => x"e3",
           666 => x"53",
           667 => x"38",
           668 => x"38",
           669 => x"31",
           670 => x"80",
           671 => x"10",
           672 => x"07",
           673 => x"70",
           674 => x"31",
           675 => x"58",
           676 => x"76",
           677 => x"88",
           678 => x"70",
           679 => x"72",
           680 => x"71",
           681 => x"80",
           682 => x"2b",
           683 => x"81",
           684 => x"82",
           685 => x"55",
           686 => x"70",
           687 => x"31",
           688 => x"32",
           689 => x"31",
           690 => x"0c",
           691 => x"5a",
           692 => x"56",
           693 => x"3d",
           694 => x"70",
           695 => x"3f",
           696 => x"71",
           697 => x"3d",
           698 => x"58",
           699 => x"38",
           700 => x"e4",
           701 => x"2e",
           702 => x"72",
           703 => x"53",
           704 => x"53",
           705 => x"74",
           706 => x"2b",
           707 => x"76",
           708 => x"2a",
           709 => x"31",
           710 => x"7b",
           711 => x"5c",
           712 => x"74",
           713 => x"88",
           714 => x"9f",
           715 => x"7b",
           716 => x"73",
           717 => x"31",
           718 => x"b4",
           719 => x"75",
           720 => x"0d",
           721 => x"57",
           722 => x"33",
           723 => x"81",
           724 => x"0c",
           725 => x"f3",
           726 => x"73",
           727 => x"58",
           728 => x"38",
           729 => x"80",
           730 => x"38",
           731 => x"53",
           732 => x"53",
           733 => x"70",
           734 => x"27",
           735 => x"83",
           736 => x"70",
           737 => x"73",
           738 => x"2e",
           739 => x"0c",
           740 => x"8b",
           741 => x"79",
           742 => x"b0",
           743 => x"81",
           744 => x"55",
           745 => x"58",
           746 => x"56",
           747 => x"53",
           748 => x"fe",
           749 => x"8b",
           750 => x"70",
           751 => x"56",
           752 => x"e4",
           753 => x"0d",
           754 => x"0c",
           755 => x"73",
           756 => x"81",
           757 => x"55",
           758 => x"2e",
           759 => x"83",
           760 => x"89",
           761 => x"56",
           762 => x"e0",
           763 => x"81",
           764 => x"81",
           765 => x"8f",
           766 => x"54",
           767 => x"72",
           768 => x"29",
           769 => x"33",
           770 => x"be",
           771 => x"30",
           772 => x"84",
           773 => x"81",
           774 => x"56",
           775 => x"06",
           776 => x"0c",
           777 => x"2e",
           778 => x"2e",
           779 => x"c6",
           780 => x"58",
           781 => x"84",
           782 => x"82",
           783 => x"33",
           784 => x"80",
           785 => x"0d",
           786 => x"e4",
           787 => x"0c",
           788 => x"93",
           789 => x"bd",
           790 => x"ce",
           791 => x"0d",
           792 => x"3f",
           793 => x"51",
           794 => x"83",
           795 => x"3d",
           796 => x"92",
           797 => x"f4",
           798 => x"04",
           799 => x"83",
           800 => x"ee",
           801 => x"cf",
           802 => x"0d",
           803 => x"3f",
           804 => x"51",
           805 => x"83",
           806 => x"3d",
           807 => x"ba",
           808 => x"c4",
           809 => x"04",
           810 => x"83",
           811 => x"ee",
           812 => x"d0",
           813 => x"0d",
           814 => x"3f",
           815 => x"51",
           816 => x"83",
           817 => x"3d",
           818 => x"e2",
           819 => x"0d",
           820 => x"33",
           821 => x"7b",
           822 => x"78",
           823 => x"81",
           824 => x"06",
           825 => x"38",
           826 => x"52",
           827 => x"e4",
           828 => x"2e",
           829 => x"86",
           830 => x"25",
           831 => x"53",
           832 => x"38",
           833 => x"87",
           834 => x"78",
           835 => x"84",
           836 => x"53",
           837 => x"df",
           838 => x"3d",
           839 => x"c0",
           840 => x"59",
           841 => x"53",
           842 => x"3f",
           843 => x"e4",
           844 => x"80",
           845 => x"17",
           846 => x"74",
           847 => x"08",
           848 => x"b8",
           849 => x"78",
           850 => x"3f",
           851 => x"02",
           852 => x"ff",
           853 => x"fd",
           854 => x"38",
           855 => x"2e",
           856 => x"8a",
           857 => x"c4",
           858 => x"e4",
           859 => x"84",
           860 => x"8a",
           861 => x"61",
           862 => x"33",
           863 => x"5c",
           864 => x"82",
           865 => x"dd",
           866 => x"f7",
           867 => x"38",
           868 => x"a0",
           869 => x"72",
           870 => x"52",
           871 => x"81",
           872 => x"a0",
           873 => x"dc",
           874 => x"3f",
           875 => x"38",
           876 => x"55",
           877 => x"80",
           878 => x"53",
           879 => x"56",
           880 => x"fe",
           881 => x"c8",
           882 => x"81",
           883 => x"83",
           884 => x"18",
           885 => x"a8",
           886 => x"70",
           887 => x"81",
           888 => x"38",
           889 => x"b9",
           890 => x"8f",
           891 => x"dc",
           892 => x"08",
           893 => x"78",
           894 => x"39",
           895 => x"82",
           896 => x"a0",
           897 => x"fe",
           898 => x"27",
           899 => x"8c",
           900 => x"d4",
           901 => x"c5",
           902 => x"99",
           903 => x"3f",
           904 => x"54",
           905 => x"27",
           906 => x"7a",
           907 => x"d1",
           908 => x"84",
           909 => x"ea",
           910 => x"fd",
           911 => x"73",
           912 => x"fe",
           913 => x"b8",
           914 => x"59",
           915 => x"59",
           916 => x"fc",
           917 => x"80",
           918 => x"08",
           919 => x"32",
           920 => x"70",
           921 => x"55",
           922 => x"25",
           923 => x"3f",
           924 => x"98",
           925 => x"9b",
           926 => x"75",
           927 => x"58",
           928 => x"fd",
           929 => x"0c",
           930 => x"87",
           931 => x"3f",
           932 => x"dc",
           933 => x"e1",
           934 => x"51",
           935 => x"2a",
           936 => x"89",
           937 => x"51",
           938 => x"2a",
           939 => x"ad",
           940 => x"51",
           941 => x"2a",
           942 => x"d2",
           943 => x"51",
           944 => x"81",
           945 => x"3f",
           946 => x"f9",
           947 => x"3f",
           948 => x"3f",
           949 => x"e1",
           950 => x"3f",
           951 => x"2a",
           952 => x"38",
           953 => x"83",
           954 => x"51",
           955 => x"81",
           956 => x"9c",
           957 => x"3f",
           958 => x"80",
           959 => x"70",
           960 => x"fe",
           961 => x"9b",
           962 => x"91",
           963 => x"85",
           964 => x"80",
           965 => x"81",
           966 => x"51",
           967 => x"3f",
           968 => x"52",
           969 => x"bd",
           970 => x"d3",
           971 => x"9a",
           972 => x"06",
           973 => x"38",
           974 => x"3f",
           975 => x"80",
           976 => x"70",
           977 => x"fd",
           978 => x"0d",
           979 => x"cf",
           980 => x"81",
           981 => x"81",
           982 => x"61",
           983 => x"51",
           984 => x"d5",
           985 => x"80",
           986 => x"ae",
           987 => x"70",
           988 => x"2e",
           989 => x"88",
           990 => x"82",
           991 => x"5a",
           992 => x"33",
           993 => x"8c",
           994 => x"7b",
           995 => x"9b",
           996 => x"ed",
           997 => x"ff",
           998 => x"e4",
           999 => x"5d",
          1000 => x"8b",
          1001 => x"2e",
          1002 => x"ff",
          1003 => x"38",
          1004 => x"fe",
          1005 => x"e9",
          1006 => x"84",
          1007 => x"38",
          1008 => x"ff",
          1009 => x"b8",
          1010 => x"7a",
          1011 => x"e4",
          1012 => x"e4",
          1013 => x"0b",
          1014 => x"8d",
          1015 => x"38",
          1016 => x"54",
          1017 => x"51",
          1018 => x"84",
          1019 => x"80",
          1020 => x"0a",
          1021 => x"b8",
          1022 => x"70",
          1023 => x"5b",
          1024 => x"83",
          1025 => x"78",
          1026 => x"81",
          1027 => x"38",
          1028 => x"5d",
          1029 => x"81",
          1030 => x"3f",
          1031 => x"7e",
          1032 => x"51",
          1033 => x"d8",
          1034 => x"79",
          1035 => x"b4",
          1036 => x"bc",
          1037 => x"38",
          1038 => x"34",
          1039 => x"7e",
          1040 => x"e4",
          1041 => x"e4",
          1042 => x"83",
          1043 => x"5f",
          1044 => x"fc",
          1045 => x"51",
          1046 => x"0b",
          1047 => x"53",
          1048 => x"3f",
          1049 => x"38",
          1050 => x"1b",
          1051 => x"80",
          1052 => x"05",
          1053 => x"d5",
          1054 => x"60",
          1055 => x"82",
          1056 => x"61",
          1057 => x"81",
          1058 => x"ae",
          1059 => x"3f",
          1060 => x"90",
          1061 => x"83",
          1062 => x"b0",
          1063 => x"93",
          1064 => x"39",
          1065 => x"52",
          1066 => x"39",
          1067 => x"83",
          1068 => x"59",
          1069 => x"8a",
          1070 => x"b8",
          1071 => x"05",
          1072 => x"08",
          1073 => x"83",
          1074 => x"5a",
          1075 => x"2e",
          1076 => x"52",
          1077 => x"fa",
          1078 => x"53",
          1079 => x"84",
          1080 => x"38",
          1081 => x"bf",
          1082 => x"fe",
          1083 => x"e9",
          1084 => x"2e",
          1085 => x"11",
          1086 => x"3f",
          1087 => x"64",
          1088 => x"d6",
          1089 => x"c4",
          1090 => x"d0",
          1091 => x"78",
          1092 => x"26",
          1093 => x"46",
          1094 => x"11",
          1095 => x"3f",
          1096 => x"fe",
          1097 => x"ff",
          1098 => x"b8",
          1099 => x"78",
          1100 => x"51",
          1101 => x"53",
          1102 => x"3f",
          1103 => x"2e",
          1104 => x"ca",
          1105 => x"cf",
          1106 => x"ff",
          1107 => x"b8",
          1108 => x"b8",
          1109 => x"05",
          1110 => x"08",
          1111 => x"fe",
          1112 => x"e9",
          1113 => x"2e",
          1114 => x"ce",
          1115 => x"7c",
          1116 => x"7a",
          1117 => x"95",
          1118 => x"53",
          1119 => x"8f",
          1120 => x"81",
          1121 => x"ff",
          1122 => x"e8",
          1123 => x"2e",
          1124 => x"11",
          1125 => x"3f",
          1126 => x"8e",
          1127 => x"ff",
          1128 => x"b8",
          1129 => x"83",
          1130 => x"5a",
          1131 => x"5c",
          1132 => x"34",
          1133 => x"3d",
          1134 => x"51",
          1135 => x"80",
          1136 => x"fc",
          1137 => x"fd",
          1138 => x"68",
          1139 => x"51",
          1140 => x"53",
          1141 => x"3f",
          1142 => x"2e",
          1143 => x"97",
          1144 => x"68",
          1145 => x"34",
          1146 => x"fc",
          1147 => x"ad",
          1148 => x"f5",
          1149 => x"05",
          1150 => x"b8",
          1151 => x"05",
          1152 => x"08",
          1153 => x"3d",
          1154 => x"51",
          1155 => x"80",
          1156 => x"fc",
          1157 => x"dd",
          1158 => x"f5",
          1159 => x"53",
          1160 => x"84",
          1161 => x"e4",
          1162 => x"b7",
          1163 => x"27",
          1164 => x"84",
          1165 => x"38",
          1166 => x"39",
          1167 => x"96",
          1168 => x"ff",
          1169 => x"81",
          1170 => x"51",
          1171 => x"80",
          1172 => x"08",
          1173 => x"b8",
          1174 => x"05",
          1175 => x"08",
          1176 => x"79",
          1177 => x"a0",
          1178 => x"53",
          1179 => x"84",
          1180 => x"e8",
          1181 => x"38",
          1182 => x"fe",
          1183 => x"e5",
          1184 => x"2e",
          1185 => x"88",
          1186 => x"32",
          1187 => x"7e",
          1188 => x"88",
          1189 => x"46",
          1190 => x"80",
          1191 => x"68",
          1192 => x"51",
          1193 => x"64",
          1194 => x"b8",
          1195 => x"05",
          1196 => x"08",
          1197 => x"71",
          1198 => x"3d",
          1199 => x"51",
          1200 => x"c6",
          1201 => x"80",
          1202 => x"40",
          1203 => x"11",
          1204 => x"3f",
          1205 => x"96",
          1206 => x"22",
          1207 => x"45",
          1208 => x"80",
          1209 => x"e4",
          1210 => x"b8",
          1211 => x"05",
          1212 => x"08",
          1213 => x"02",
          1214 => x"81",
          1215 => x"fe",
          1216 => x"e1",
          1217 => x"2e",
          1218 => x"5d",
          1219 => x"e1",
          1220 => x"f3",
          1221 => x"54",
          1222 => x"51",
          1223 => x"52",
          1224 => x"39",
          1225 => x"f0",
          1226 => x"53",
          1227 => x"84",
          1228 => x"64",
          1229 => x"70",
          1230 => x"e7",
          1231 => x"80",
          1232 => x"08",
          1233 => x"33",
          1234 => x"f1",
          1235 => x"d8",
          1236 => x"f7",
          1237 => x"ca",
          1238 => x"f1",
          1239 => x"38",
          1240 => x"39",
          1241 => x"f9",
          1242 => x"78",
          1243 => x"08",
          1244 => x"33",
          1245 => x"f1",
          1246 => x"f1",
          1247 => x"38",
          1248 => x"39",
          1249 => x"2e",
          1250 => x"fb",
          1251 => x"7c",
          1252 => x"08",
          1253 => x"08",
          1254 => x"83",
          1255 => x"b5",
          1256 => x"b9",
          1257 => x"08",
          1258 => x"51",
          1259 => x"90",
          1260 => x"80",
          1261 => x"84",
          1262 => x"c0",
          1263 => x"84",
          1264 => x"84",
          1265 => x"57",
          1266 => x"da",
          1267 => x"07",
          1268 => x"c0",
          1269 => x"87",
          1270 => x"5c",
          1271 => x"05",
          1272 => x"c4",
          1273 => x"70",
          1274 => x"b6",
          1275 => x"3f",
          1276 => x"d2",
          1277 => x"9f",
          1278 => x"55",
          1279 => x"83",
          1280 => x"83",
          1281 => x"97",
          1282 => x"3d",
          1283 => x"75",
          1284 => x"38",
          1285 => x"52",
          1286 => x"38",
          1287 => x"06",
          1288 => x"38",
          1289 => x"2e",
          1290 => x"2e",
          1291 => x"81",
          1292 => x"2e",
          1293 => x"8b",
          1294 => x"12",
          1295 => x"06",
          1296 => x"06",
          1297 => x"70",
          1298 => x"52",
          1299 => x"72",
          1300 => x"0c",
          1301 => x"87",
          1302 => x"38",
          1303 => x"12",
          1304 => x"06",
          1305 => x"38",
          1306 => x"81",
          1307 => x"81",
          1308 => x"3d",
          1309 => x"80",
          1310 => x"0d",
          1311 => x"51",
          1312 => x"80",
          1313 => x"0c",
          1314 => x"76",
          1315 => x"81",
          1316 => x"83",
          1317 => x"73",
          1318 => x"33",
          1319 => x"fe",
          1320 => x"73",
          1321 => x"33",
          1322 => x"e6",
          1323 => x"74",
          1324 => x"13",
          1325 => x"26",
          1326 => x"98",
          1327 => x"bc",
          1328 => x"b8",
          1329 => x"b4",
          1330 => x"b0",
          1331 => x"ac",
          1332 => x"a8",
          1333 => x"73",
          1334 => x"87",
          1335 => x"84",
          1336 => x"f3",
          1337 => x"9c",
          1338 => x"bc",
          1339 => x"98",
          1340 => x"87",
          1341 => x"1c",
          1342 => x"7b",
          1343 => x"08",
          1344 => x"98",
          1345 => x"87",
          1346 => x"1c",
          1347 => x"79",
          1348 => x"83",
          1349 => x"ff",
          1350 => x"1b",
          1351 => x"1b",
          1352 => x"83",
          1353 => x"51",
          1354 => x"04",
          1355 => x"53",
          1356 => x"80",
          1357 => x"98",
          1358 => x"ff",
          1359 => x"83",
          1360 => x"0c",
          1361 => x"e8",
          1362 => x"2b",
          1363 => x"2e",
          1364 => x"80",
          1365 => x"98",
          1366 => x"ff",
          1367 => x"0d",
          1368 => x"54",
          1369 => x"b8",
          1370 => x"51",
          1371 => x"72",
          1372 => x"25",
          1373 => x"85",
          1374 => x"9b",
          1375 => x"81",
          1376 => x"2e",
          1377 => x"08",
          1378 => x"54",
          1379 => x"91",
          1380 => x"e3",
          1381 => x"72",
          1382 => x"81",
          1383 => x"ff",
          1384 => x"70",
          1385 => x"90",
          1386 => x"e4",
          1387 => x"2a",
          1388 => x"38",
          1389 => x"80",
          1390 => x"06",
          1391 => x"c0",
          1392 => x"81",
          1393 => x"d8",
          1394 => x"33",
          1395 => x"52",
          1396 => x"0d",
          1397 => x"75",
          1398 => x"2e",
          1399 => x"9c",
          1400 => x"55",
          1401 => x"c0",
          1402 => x"81",
          1403 => x"8c",
          1404 => x"51",
          1405 => x"81",
          1406 => x"71",
          1407 => x"38",
          1408 => x"94",
          1409 => x"87",
          1410 => x"81",
          1411 => x"9b",
          1412 => x"3d",
          1413 => x"06",
          1414 => x"32",
          1415 => x"38",
          1416 => x"80",
          1417 => x"84",
          1418 => x"53",
          1419 => x"ff",
          1420 => x"70",
          1421 => x"80",
          1422 => x"a4",
          1423 => x"9e",
          1424 => x"c0",
          1425 => x"87",
          1426 => x"0c",
          1427 => x"b0",
          1428 => x"f1",
          1429 => x"83",
          1430 => x"08",
          1431 => x"b4",
          1432 => x"9e",
          1433 => x"c0",
          1434 => x"87",
          1435 => x"0c",
          1436 => x"d0",
          1437 => x"71",
          1438 => x"84",
          1439 => x"9e",
          1440 => x"c0",
          1441 => x"81",
          1442 => x"87",
          1443 => x"0a",
          1444 => x"38",
          1445 => x"87",
          1446 => x"0a",
          1447 => x"83",
          1448 => x"34",
          1449 => x"70",
          1450 => x"70",
          1451 => x"83",
          1452 => x"9e",
          1453 => x"51",
          1454 => x"81",
          1455 => x"0b",
          1456 => x"80",
          1457 => x"2e",
          1458 => x"e9",
          1459 => x"08",
          1460 => x"52",
          1461 => x"71",
          1462 => x"c0",
          1463 => x"06",
          1464 => x"38",
          1465 => x"80",
          1466 => x"82",
          1467 => x"80",
          1468 => x"f1",
          1469 => x"90",
          1470 => x"52",
          1471 => x"52",
          1472 => x"87",
          1473 => x"80",
          1474 => x"83",
          1475 => x"34",
          1476 => x"70",
          1477 => x"80",
          1478 => x"f1",
          1479 => x"98",
          1480 => x"71",
          1481 => x"c0",
          1482 => x"51",
          1483 => x"81",
          1484 => x"c0",
          1485 => x"84",
          1486 => x"34",
          1487 => x"70",
          1488 => x"2e",
          1489 => x"f3",
          1490 => x"06",
          1491 => x"3d",
          1492 => x"fb",
          1493 => x"b6",
          1494 => x"73",
          1495 => x"c3",
          1496 => x"74",
          1497 => x"54",
          1498 => x"33",
          1499 => x"e9",
          1500 => x"f1",
          1501 => x"83",
          1502 => x"38",
          1503 => x"90",
          1504 => x"83",
          1505 => x"75",
          1506 => x"54",
          1507 => x"33",
          1508 => x"ed",
          1509 => x"f1",
          1510 => x"83",
          1511 => x"f1",
          1512 => x"ff",
          1513 => x"52",
          1514 => x"3f",
          1515 => x"a8",
          1516 => x"d0",
          1517 => x"22",
          1518 => x"97",
          1519 => x"84",
          1520 => x"84",
          1521 => x"76",
          1522 => x"08",
          1523 => x"ef",
          1524 => x"80",
          1525 => x"74",
          1526 => x"87",
          1527 => x"56",
          1528 => x"e4",
          1529 => x"c0",
          1530 => x"b8",
          1531 => x"ff",
          1532 => x"3f",
          1533 => x"08",
          1534 => x"c9",
          1535 => x"84",
          1536 => x"84",
          1537 => x"51",
          1538 => x"33",
          1539 => x"ff",
          1540 => x"d2",
          1541 => x"3f",
          1542 => x"d8",
          1543 => x"cc",
          1544 => x"b3",
          1545 => x"83",
          1546 => x"83",
          1547 => x"f1",
          1548 => x"ff",
          1549 => x"56",
          1550 => x"b4",
          1551 => x"c0",
          1552 => x"b8",
          1553 => x"ff",
          1554 => x"55",
          1555 => x"cc",
          1556 => x"d2",
          1557 => x"80",
          1558 => x"83",
          1559 => x"83",
          1560 => x"fc",
          1561 => x"51",
          1562 => x"33",
          1563 => x"d7",
          1564 => x"92",
          1565 => x"80",
          1566 => x"f1",
          1567 => x"ff",
          1568 => x"56",
          1569 => x"39",
          1570 => x"e0",
          1571 => x"f1",
          1572 => x"38",
          1573 => x"83",
          1574 => x"83",
          1575 => x"fb",
          1576 => x"08",
          1577 => x"83",
          1578 => x"83",
          1579 => x"fb",
          1580 => x"08",
          1581 => x"83",
          1582 => x"83",
          1583 => x"fa",
          1584 => x"08",
          1585 => x"83",
          1586 => x"83",
          1587 => x"fa",
          1588 => x"08",
          1589 => x"83",
          1590 => x"83",
          1591 => x"fa",
          1592 => x"08",
          1593 => x"83",
          1594 => x"83",
          1595 => x"f9",
          1596 => x"51",
          1597 => x"51",
          1598 => x"33",
          1599 => x"c4",
          1600 => x"33",
          1601 => x"10",
          1602 => x"08",
          1603 => x"ef",
          1604 => x"c8",
          1605 => x"0d",
          1606 => x"d7",
          1607 => x"d8",
          1608 => x"0d",
          1609 => x"bf",
          1610 => x"e8",
          1611 => x"0d",
          1612 => x"0b",
          1613 => x"f1",
          1614 => x"04",
          1615 => x"3d",
          1616 => x"80",
          1617 => x"88",
          1618 => x"ed",
          1619 => x"f2",
          1620 => x"76",
          1621 => x"e4",
          1622 => x"c0",
          1623 => x"17",
          1624 => x"08",
          1625 => x"ff",
          1626 => x"34",
          1627 => x"9f",
          1628 => x"85",
          1629 => x"d0",
          1630 => x"87",
          1631 => x"38",
          1632 => x"b8",
          1633 => x"e1",
          1634 => x"76",
          1635 => x"52",
          1636 => x"c0",
          1637 => x"b8",
          1638 => x"e1",
          1639 => x"0b",
          1640 => x"04",
          1641 => x"3d",
          1642 => x"57",
          1643 => x"38",
          1644 => x"10",
          1645 => x"08",
          1646 => x"b8",
          1647 => x"51",
          1648 => x"90",
          1649 => x"2e",
          1650 => x"38",
          1651 => x"54",
          1652 => x"73",
          1653 => x"04",
          1654 => x"11",
          1655 => x"3f",
          1656 => x"38",
          1657 => x"fd",
          1658 => x"ff",
          1659 => x"81",
          1660 => x"82",
          1661 => x"39",
          1662 => x"27",
          1663 => x"70",
          1664 => x"81",
          1665 => x"eb",
          1666 => x"fe",
          1667 => x"53",
          1668 => x"84",
          1669 => x"d0",
          1670 => x"f8",
          1671 => x"84",
          1672 => x"77",
          1673 => x"e4",
          1674 => x"08",
          1675 => x"ff",
          1676 => x"34",
          1677 => x"e1",
          1678 => x"74",
          1679 => x"38",
          1680 => x"3d",
          1681 => x"08",
          1682 => x"41",
          1683 => x"f2",
          1684 => x"5d",
          1685 => x"33",
          1686 => x"38",
          1687 => x"70",
          1688 => x"38",
          1689 => x"3d",
          1690 => x"80",
          1691 => x"70",
          1692 => x"ec",
          1693 => x"a0",
          1694 => x"84",
          1695 => x"97",
          1696 => x"10",
          1697 => x"70",
          1698 => x"5b",
          1699 => x"2e",
          1700 => x"87",
          1701 => x"ff",
          1702 => x"80",
          1703 => x"16",
          1704 => x"83",
          1705 => x"61",
          1706 => x"08",
          1707 => x"2e",
          1708 => x"38",
          1709 => x"76",
          1710 => x"70",
          1711 => x"9c",
          1712 => x"71",
          1713 => x"dd",
          1714 => x"58",
          1715 => x"90",
          1716 => x"ac",
          1717 => x"75",
          1718 => x"05",
          1719 => x"59",
          1720 => x"38",
          1721 => x"55",
          1722 => x"42",
          1723 => x"dd",
          1724 => x"55",
          1725 => x"80",
          1726 => x"81",
          1727 => x"fe",
          1728 => x"80",
          1729 => x"d0",
          1730 => x"79",
          1731 => x"74",
          1732 => x"10",
          1733 => x"04",
          1734 => x"80",
          1735 => x"84",
          1736 => x"a8",
          1737 => x"38",
          1738 => x"ff",
          1739 => x"ff",
          1740 => x"fc",
          1741 => x"81",
          1742 => x"57",
          1743 => x"84",
          1744 => x"77",
          1745 => x"33",
          1746 => x"bc",
          1747 => x"7c",
          1748 => x"08",
          1749 => x"84",
          1750 => x"d0",
          1751 => x"56",
          1752 => x"c8",
          1753 => x"3f",
          1754 => x"ff",
          1755 => x"52",
          1756 => x"d0",
          1757 => x"d0",
          1758 => x"74",
          1759 => x"3f",
          1760 => x"39",
          1761 => x"56",
          1762 => x"83",
          1763 => x"55",
          1764 => x"75",
          1765 => x"ff",
          1766 => x"84",
          1767 => x"81",
          1768 => x"7b",
          1769 => x"a4",
          1770 => x"74",
          1771 => x"c8",
          1772 => x"3f",
          1773 => x"ff",
          1774 => x"52",
          1775 => x"d0",
          1776 => x"d0",
          1777 => x"c7",
          1778 => x"ff",
          1779 => x"55",
          1780 => x"d4",
          1781 => x"84",
          1782 => x"52",
          1783 => x"a8",
          1784 => x"a4",
          1785 => x"fa",
          1786 => x"81",
          1787 => x"7b",
          1788 => x"8d",
          1789 => x"ff",
          1790 => x"55",
          1791 => x"d4",
          1792 => x"a4",
          1793 => x"c4",
          1794 => x"a4",
          1795 => x"7c",
          1796 => x"76",
          1797 => x"08",
          1798 => x"84",
          1799 => x"98",
          1800 => x"57",
          1801 => x"84",
          1802 => x"b2",
          1803 => x"81",
          1804 => x"d0",
          1805 => x"24",
          1806 => x"52",
          1807 => x"81",
          1808 => x"70",
          1809 => x"56",
          1810 => x"f8",
          1811 => x"33",
          1812 => x"77",
          1813 => x"81",
          1814 => x"70",
          1815 => x"57",
          1816 => x"7b",
          1817 => x"84",
          1818 => x"ff",
          1819 => x"29",
          1820 => x"84",
          1821 => x"76",
          1822 => x"84",
          1823 => x"f7",
          1824 => x"88",
          1825 => x"a8",
          1826 => x"a8",
          1827 => x"39",
          1828 => x"80",
          1829 => x"8a",
          1830 => x"a4",
          1831 => x"b8",
          1832 => x"89",
          1833 => x"76",
          1834 => x"d4",
          1835 => x"05",
          1836 => x"a0",
          1837 => x"83",
          1838 => x"57",
          1839 => x"e4",
          1840 => x"70",
          1841 => x"08",
          1842 => x"83",
          1843 => x"8c",
          1844 => x"80",
          1845 => x"d0",
          1846 => x"34",
          1847 => x"0d",
          1848 => x"80",
          1849 => x"52",
          1850 => x"d4",
          1851 => x"95",
          1852 => x"51",
          1853 => x"33",
          1854 => x"34",
          1855 => x"38",
          1856 => x"3f",
          1857 => x"0b",
          1858 => x"83",
          1859 => x"84",
          1860 => x"b6",
          1861 => x"51",
          1862 => x"08",
          1863 => x"84",
          1864 => x"ae",
          1865 => x"05",
          1866 => x"81",
          1867 => x"d1",
          1868 => x"0b",
          1869 => x"d0",
          1870 => x"b4",
          1871 => x"70",
          1872 => x"2e",
          1873 => x"ff",
          1874 => x"ff",
          1875 => x"84",
          1876 => x"ad",
          1877 => x"98",
          1878 => x"33",
          1879 => x"80",
          1880 => x"a0",
          1881 => x"a8",
          1882 => x"84",
          1883 => x"74",
          1884 => x"c8",
          1885 => x"3f",
          1886 => x"0a",
          1887 => x"33",
          1888 => x"cc",
          1889 => x"51",
          1890 => x"0a",
          1891 => x"2c",
          1892 => x"78",
          1893 => x"39",
          1894 => x"34",
          1895 => x"51",
          1896 => x"0a",
          1897 => x"2c",
          1898 => x"75",
          1899 => x"57",
          1900 => x"c8",
          1901 => x"85",
          1902 => x"80",
          1903 => x"a4",
          1904 => x"ff",
          1905 => x"a8",
          1906 => x"76",
          1907 => x"a4",
          1908 => x"74",
          1909 => x"76",
          1910 => x"7a",
          1911 => x"0a",
          1912 => x"2c",
          1913 => x"75",
          1914 => x"74",
          1915 => x"06",
          1916 => x"34",
          1917 => x"25",
          1918 => x"d0",
          1919 => x"33",
          1920 => x"0a",
          1921 => x"06",
          1922 => x"81",
          1923 => x"2c",
          1924 => x"75",
          1925 => x"c8",
          1926 => x"3f",
          1927 => x"0a",
          1928 => x"33",
          1929 => x"84",
          1930 => x"51",
          1931 => x"0a",
          1932 => x"2c",
          1933 => x"74",
          1934 => x"39",
          1935 => x"2e",
          1936 => x"a7",
          1937 => x"a4",
          1938 => x"06",
          1939 => x"ff",
          1940 => x"84",
          1941 => x"2e",
          1942 => x"52",
          1943 => x"d4",
          1944 => x"ad",
          1945 => x"51",
          1946 => x"33",
          1947 => x"34",
          1948 => x"a8",
          1949 => x"e4",
          1950 => x"e4",
          1951 => x"cc",
          1952 => x"39",
          1953 => x"70",
          1954 => x"75",
          1955 => x"05",
          1956 => x"52",
          1957 => x"84",
          1958 => x"98",
          1959 => x"5a",
          1960 => x"fd",
          1961 => x"2e",
          1962 => x"93",
          1963 => x"ff",
          1964 => x"25",
          1965 => x"34",
          1966 => x"2e",
          1967 => x"f6",
          1968 => x"d9",
          1969 => x"0c",
          1970 => x"bc",
          1971 => x"80",
          1972 => x"56",
          1973 => x"ba",
          1974 => x"84",
          1975 => x"84",
          1976 => x"05",
          1977 => x"a1",
          1978 => x"84",
          1979 => x"80",
          1980 => x"08",
          1981 => x"84",
          1982 => x"a6",
          1983 => x"88",
          1984 => x"a8",
          1985 => x"a8",
          1986 => x"39",
          1987 => x"a8",
          1988 => x"7b",
          1989 => x"04",
          1990 => x"b8",
          1991 => x"b8",
          1992 => x"53",
          1993 => x"3f",
          1994 => x"d0",
          1995 => x"52",
          1996 => x"38",
          1997 => x"ff",
          1998 => x"52",
          1999 => x"d4",
          2000 => x"ed",
          2001 => x"57",
          2002 => x"ff",
          2003 => x"a9",
          2004 => x"d0",
          2005 => x"ff",
          2006 => x"51",
          2007 => x"81",
          2008 => x"d0",
          2009 => x"80",
          2010 => x"08",
          2011 => x"84",
          2012 => x"a5",
          2013 => x"88",
          2014 => x"a8",
          2015 => x"a8",
          2016 => x"39",
          2017 => x"f2",
          2018 => x"06",
          2019 => x"54",
          2020 => x"84",
          2021 => x"d4",
          2022 => x"05",
          2023 => x"2e",
          2024 => x"74",
          2025 => x"d4",
          2026 => x"5a",
          2027 => x"77",
          2028 => x"b4",
          2029 => x"7b",
          2030 => x"83",
          2031 => x"ba",
          2032 => x"81",
          2033 => x"a8",
          2034 => x"7b",
          2035 => x"04",
          2036 => x"08",
          2037 => x"e4",
          2038 => x"08",
          2039 => x"08",
          2040 => x"b7",
          2041 => x"84",
          2042 => x"06",
          2043 => x"51",
          2044 => x"08",
          2045 => x"25",
          2046 => x"ff",
          2047 => x"34",
          2048 => x"33",
          2049 => x"70",
          2050 => x"f2",
          2051 => x"83",
          2052 => x"58",
          2053 => x"e4",
          2054 => x"70",
          2055 => x"08",
          2056 => x"1d",
          2057 => x"7d",
          2058 => x"2e",
          2059 => x"e8",
          2060 => x"79",
          2061 => x"83",
          2062 => x"ff",
          2063 => x"c8",
          2064 => x"ff",
          2065 => x"3f",
          2066 => x"87",
          2067 => x"1b",
          2068 => x"cf",
          2069 => x"83",
          2070 => x"f1",
          2071 => x"74",
          2072 => x"39",
          2073 => x"39",
          2074 => x"39",
          2075 => x"3f",
          2076 => x"f2",
          2077 => x"02",
          2078 => x"53",
          2079 => x"81",
          2080 => x"83",
          2081 => x"38",
          2082 => x"b0",
          2083 => x"a0",
          2084 => x"83",
          2085 => x"34",
          2086 => x"90",
          2087 => x"07",
          2088 => x"7f",
          2089 => x"94",
          2090 => x"0c",
          2091 => x"76",
          2092 => x"a2",
          2093 => x"b6",
          2094 => x"a0",
          2095 => x"70",
          2096 => x"72",
          2097 => x"a7",
          2098 => x"70",
          2099 => x"71",
          2100 => x"58",
          2101 => x"84",
          2102 => x"84",
          2103 => x"83",
          2104 => x"06",
          2105 => x"5e",
          2106 => x"38",
          2107 => x"81",
          2108 => x"81",
          2109 => x"62",
          2110 => x"5d",
          2111 => x"26",
          2112 => x"76",
          2113 => x"5f",
          2114 => x"fe",
          2115 => x"77",
          2116 => x"81",
          2117 => x"74",
          2118 => x"86",
          2119 => x"80",
          2120 => x"ff",
          2121 => x"ff",
          2122 => x"29",
          2123 => x"57",
          2124 => x"81",
          2125 => x"71",
          2126 => x"2e",
          2127 => x"94",
          2128 => x"83",
          2129 => x"90",
          2130 => x"07",
          2131 => x"79",
          2132 => x"72",
          2133 => x"70",
          2134 => x"83",
          2135 => x"86",
          2136 => x"56",
          2137 => x"14",
          2138 => x"06",
          2139 => x"06",
          2140 => x"ff",
          2141 => x"5a",
          2142 => x"79",
          2143 => x"15",
          2144 => x"81",
          2145 => x"71",
          2146 => x"81",
          2147 => x"5b",
          2148 => x"38",
          2149 => x"16",
          2150 => x"e2",
          2151 => x"da",
          2152 => x"7b",
          2153 => x"0d",
          2154 => x"73",
          2155 => x"81",
          2156 => x"80",
          2157 => x"86",
          2158 => x"80",
          2159 => x"8a",
          2160 => x"75",
          2161 => x"3f",
          2162 => x"54",
          2163 => x"73",
          2164 => x"75",
          2165 => x"80",
          2166 => x"86",
          2167 => x"81",
          2168 => x"f3",
          2169 => x"07",
          2170 => x"84",
          2171 => x"e4",
          2172 => x"d8",
          2173 => x"3d",
          2174 => x"05",
          2175 => x"5b",
          2176 => x"82",
          2177 => x"f8",
          2178 => x"71",
          2179 => x"83",
          2180 => x"71",
          2181 => x"06",
          2182 => x"53",
          2183 => x"f8",
          2184 => x"f8",
          2185 => x"05",
          2186 => x"06",
          2187 => x"8c",
          2188 => x"94",
          2189 => x"ff",
          2190 => x"55",
          2191 => x"84",
          2192 => x"58",
          2193 => x"38",
          2194 => x"e0",
          2195 => x"72",
          2196 => x"81",
          2197 => x"b6",
          2198 => x"9f",
          2199 => x"84",
          2200 => x"e0",
          2201 => x"05",
          2202 => x"74",
          2203 => x"ff",
          2204 => x"75",
          2205 => x"ff",
          2206 => x"81",
          2207 => x"84",
          2208 => x"55",
          2209 => x"58",
          2210 => x"06",
          2211 => x"19",
          2212 => x"b9",
          2213 => x"e0",
          2214 => x"33",
          2215 => x"70",
          2216 => x"05",
          2217 => x"33",
          2218 => x"19",
          2219 => x"ce",
          2220 => x"0c",
          2221 => x"94",
          2222 => x"ff",
          2223 => x"55",
          2224 => x"77",
          2225 => x"ff",
          2226 => x"56",
          2227 => x"fe",
          2228 => x"84",
          2229 => x"72",
          2230 => x"73",
          2231 => x"33",
          2232 => x"55",
          2233 => x"34",
          2234 => x"ff",
          2235 => x"38",
          2236 => x"75",
          2237 => x"53",
          2238 => x"0b",
          2239 => x"89",
          2240 => x"84",
          2241 => x"b6",
          2242 => x"3d",
          2243 => x"33",
          2244 => x"70",
          2245 => x"70",
          2246 => x"71",
          2247 => x"95",
          2248 => x"86",
          2249 => x"95",
          2250 => x"ff",
          2251 => x"38",
          2252 => x"34",
          2253 => x"3d",
          2254 => x"73",
          2255 => x"06",
          2256 => x"94",
          2257 => x"72",
          2258 => x"55",
          2259 => x"70",
          2260 => x"0b",
          2261 => x"04",
          2262 => x"70",
          2263 => x"56",
          2264 => x"80",
          2265 => x"0d",
          2266 => x"84",
          2267 => x"51",
          2268 => x"72",
          2269 => x"b8",
          2270 => x"0b",
          2271 => x"33",
          2272 => x"52",
          2273 => x"12",
          2274 => x"d0",
          2275 => x"33",
          2276 => x"10",
          2277 => x"08",
          2278 => x"f0",
          2279 => x"70",
          2280 => x"51",
          2281 => x"9c",
          2282 => x"34",
          2283 => x"3d",
          2284 => x"9f",
          2285 => x"90",
          2286 => x"83",
          2287 => x"80",
          2288 => x"34",
          2289 => x"fe",
          2290 => x"90",
          2291 => x"f8",
          2292 => x"0c",
          2293 => x"33",
          2294 => x"83",
          2295 => x"f8",
          2296 => x"f8",
          2297 => x"90",
          2298 => x"70",
          2299 => x"83",
          2300 => x"07",
          2301 => x"81",
          2302 => x"06",
          2303 => x"34",
          2304 => x"81",
          2305 => x"34",
          2306 => x"81",
          2307 => x"83",
          2308 => x"f8",
          2309 => x"51",
          2310 => x"39",
          2311 => x"80",
          2312 => x"34",
          2313 => x"81",
          2314 => x"83",
          2315 => x"f8",
          2316 => x"51",
          2317 => x"39",
          2318 => x"51",
          2319 => x"39",
          2320 => x"82",
          2321 => x"fd",
          2322 => x"05",
          2323 => x"33",
          2324 => x"33",
          2325 => x"33",
          2326 => x"82",
          2327 => x"a5",
          2328 => x"7d",
          2329 => x"b6",
          2330 => x"7b",
          2331 => x"95",
          2332 => x"2e",
          2333 => x"84",
          2334 => x"dc",
          2335 => x"a8",
          2336 => x"83",
          2337 => x"d8",
          2338 => x"84",
          2339 => x"53",
          2340 => x"81",
          2341 => x"80",
          2342 => x"f8",
          2343 => x"7c",
          2344 => x"04",
          2345 => x"0b",
          2346 => x"f8",
          2347 => x"34",
          2348 => x"b7",
          2349 => x"57",
          2350 => x"7b",
          2351 => x"f4",
          2352 => x"84",
          2353 => x"27",
          2354 => x"05",
          2355 => x"51",
          2356 => x"81",
          2357 => x"5b",
          2358 => x"d2",
          2359 => x"84",
          2360 => x"dc",
          2361 => x"83",
          2362 => x"34",
          2363 => x"b6",
          2364 => x"34",
          2365 => x"0b",
          2366 => x"f8",
          2367 => x"92",
          2368 => x"83",
          2369 => x"80",
          2370 => x"97",
          2371 => x"fd",
          2372 => x"52",
          2373 => x"3f",
          2374 => x"5a",
          2375 => x"84",
          2376 => x"33",
          2377 => x"33",
          2378 => x"80",
          2379 => x"59",
          2380 => x"ff",
          2381 => x"59",
          2382 => x"81",
          2383 => x"38",
          2384 => x"81",
          2385 => x"82",
          2386 => x"f8",
          2387 => x"72",
          2388 => x"e0",
          2389 => x"34",
          2390 => x"33",
          2391 => x"12",
          2392 => x"96",
          2393 => x"71",
          2394 => x"33",
          2395 => x"b6",
          2396 => x"f8",
          2397 => x"72",
          2398 => x"83",
          2399 => x"34",
          2400 => x"55",
          2401 => x"b6",
          2402 => x"ff",
          2403 => x"84",
          2404 => x"8c",
          2405 => x"80",
          2406 => x"b8",
          2407 => x"8d",
          2408 => x"f7",
          2409 => x"fe",
          2410 => x"96",
          2411 => x"ff",
          2412 => x"53",
          2413 => x"75",
          2414 => x"38",
          2415 => x"ba",
          2416 => x"54",
          2417 => x"76",
          2418 => x"13",
          2419 => x"73",
          2420 => x"83",
          2421 => x"52",
          2422 => x"84",
          2423 => x"75",
          2424 => x"ca",
          2425 => x"ff",
          2426 => x"38",
          2427 => x"76",
          2428 => x"f8",
          2429 => x"ff",
          2430 => x"53",
          2431 => x"39",
          2432 => x"52",
          2433 => x"39",
          2434 => x"fe",
          2435 => x"f3",
          2436 => x"59",
          2437 => x"82",
          2438 => x"84",
          2439 => x"38",
          2440 => x"89",
          2441 => x"33",
          2442 => x"33",
          2443 => x"84",
          2444 => x"80",
          2445 => x"f8",
          2446 => x"71",
          2447 => x"83",
          2448 => x"33",
          2449 => x"83",
          2450 => x"80",
          2451 => x"81",
          2452 => x"f8",
          2453 => x"40",
          2454 => x"84",
          2455 => x"81",
          2456 => x"81",
          2457 => x"79",
          2458 => x"83",
          2459 => x"e4",
          2460 => x"2e",
          2461 => x"fd",
          2462 => x"78",
          2463 => x"0b",
          2464 => x"33",
          2465 => x"33",
          2466 => x"84",
          2467 => x"80",
          2468 => x"f8",
          2469 => x"71",
          2470 => x"83",
          2471 => x"33",
          2472 => x"f8",
          2473 => x"34",
          2474 => x"06",
          2475 => x"33",
          2476 => x"58",
          2477 => x"97",
          2478 => x"81",
          2479 => x"ca",
          2480 => x"0b",
          2481 => x"04",
          2482 => x"9b",
          2483 => x"09",
          2484 => x"83",
          2485 => x"e4",
          2486 => x"2e",
          2487 => x"89",
          2488 => x"33",
          2489 => x"e4",
          2490 => x"77",
          2491 => x"b7",
          2492 => x"e4",
          2493 => x"2e",
          2494 => x"e0",
          2495 => x"94",
          2496 => x"29",
          2497 => x"19",
          2498 => x"84",
          2499 => x"83",
          2500 => x"41",
          2501 => x"1f",
          2502 => x"29",
          2503 => x"86",
          2504 => x"d8",
          2505 => x"92",
          2506 => x"29",
          2507 => x"f8",
          2508 => x"34",
          2509 => x"52",
          2510 => x"83",
          2511 => x"b6",
          2512 => x"81",
          2513 => x"71",
          2514 => x"83",
          2515 => x"7e",
          2516 => x"83",
          2517 => x"5c",
          2518 => x"81",
          2519 => x"fc",
          2520 => x"95",
          2521 => x"b7",
          2522 => x"34",
          2523 => x"0b",
          2524 => x"b7",
          2525 => x"0c",
          2526 => x"33",
          2527 => x"33",
          2528 => x"33",
          2529 => x"b7",
          2530 => x"0c",
          2531 => x"2e",
          2532 => x"f8",
          2533 => x"81",
          2534 => x"81",
          2535 => x"a7",
          2536 => x"5c",
          2537 => x"ff",
          2538 => x"5c",
          2539 => x"2e",
          2540 => x"ff",
          2541 => x"57",
          2542 => x"ff",
          2543 => x"ff",
          2544 => x"5b",
          2545 => x"80",
          2546 => x"f8",
          2547 => x"71",
          2548 => x"0b",
          2549 => x"94",
          2550 => x"56",
          2551 => x"80",
          2552 => x"81",
          2553 => x"f8",
          2554 => x"5d",
          2555 => x"7f",
          2556 => x"70",
          2557 => x"26",
          2558 => x"5a",
          2559 => x"77",
          2560 => x"33",
          2561 => x"56",
          2562 => x"d8",
          2563 => x"78",
          2564 => x"e4",
          2565 => x"bf",
          2566 => x"38",
          2567 => x"58",
          2568 => x"95",
          2569 => x"3f",
          2570 => x"3d",
          2571 => x"b6",
          2572 => x"f8",
          2573 => x"75",
          2574 => x"83",
          2575 => x"29",
          2576 => x"f6",
          2577 => x"5b",
          2578 => x"80",
          2579 => x"ff",
          2580 => x"29",
          2581 => x"33",
          2582 => x"b6",
          2583 => x"f8",
          2584 => x"41",
          2585 => x"1c",
          2586 => x"29",
          2587 => x"86",
          2588 => x"d8",
          2589 => x"92",
          2590 => x"29",
          2591 => x"f8",
          2592 => x"60",
          2593 => x"58",
          2594 => x"b6",
          2595 => x"ff",
          2596 => x"81",
          2597 => x"7b",
          2598 => x"94",
          2599 => x"95",
          2600 => x"ff",
          2601 => x"29",
          2602 => x"84",
          2603 => x"1b",
          2604 => x"95",
          2605 => x"29",
          2606 => x"83",
          2607 => x"33",
          2608 => x"f8",
          2609 => x"34",
          2610 => x"06",
          2611 => x"33",
          2612 => x"40",
          2613 => x"b6",
          2614 => x"ff",
          2615 => x"d6",
          2616 => x"df",
          2617 => x"80",
          2618 => x"0d",
          2619 => x"84",
          2620 => x"f8",
          2621 => x"ff",
          2622 => x"84",
          2623 => x"e4",
          2624 => x"96",
          2625 => x"33",
          2626 => x"b6",
          2627 => x"5b",
          2628 => x"b7",
          2629 => x"d8",
          2630 => x"b8",
          2631 => x"84",
          2632 => x"75",
          2633 => x"fe",
          2634 => x"61",
          2635 => x"39",
          2636 => x"b6",
          2637 => x"94",
          2638 => x"95",
          2639 => x"84",
          2640 => x"83",
          2641 => x"41",
          2642 => x"7f",
          2643 => x"b6",
          2644 => x"f8",
          2645 => x"43",
          2646 => x"34",
          2647 => x"1b",
          2648 => x"86",
          2649 => x"d8",
          2650 => x"92",
          2651 => x"29",
          2652 => x"f8",
          2653 => x"81",
          2654 => x"60",
          2655 => x"d9",
          2656 => x"1a",
          2657 => x"0b",
          2658 => x"33",
          2659 => x"84",
          2660 => x"38",
          2661 => x"80",
          2662 => x"0d",
          2663 => x"94",
          2664 => x"95",
          2665 => x"83",
          2666 => x"f8",
          2667 => x"f8",
          2668 => x"f8",
          2669 => x"9e",
          2670 => x"80",
          2671 => x"22",
          2672 => x"ff",
          2673 => x"05",
          2674 => x"54",
          2675 => x"3d",
          2676 => x"76",
          2677 => x"e4",
          2678 => x"33",
          2679 => x"fe",
          2680 => x"51",
          2681 => x"80",
          2682 => x"79",
          2683 => x"fe",
          2684 => x"05",
          2685 => x"26",
          2686 => x"c7",
          2687 => x"b7",
          2688 => x"a4",
          2689 => x"b9",
          2690 => x"9f",
          2691 => x"5c",
          2692 => x"39",
          2693 => x"2e",
          2694 => x"ff",
          2695 => x"d8",
          2696 => x"fd",
          2697 => x"fd",
          2698 => x"34",
          2699 => x"06",
          2700 => x"38",
          2701 => x"34",
          2702 => x"95",
          2703 => x"d7",
          2704 => x"25",
          2705 => x"83",
          2706 => x"b7",
          2707 => x"e0",
          2708 => x"b9",
          2709 => x"9f",
          2710 => x"5a",
          2711 => x"39",
          2712 => x"2e",
          2713 => x"41",
          2714 => x"b6",
          2715 => x"95",
          2716 => x"29",
          2717 => x"f8",
          2718 => x"60",
          2719 => x"83",
          2720 => x"06",
          2721 => x"80",
          2722 => x"f6",
          2723 => x"e5",
          2724 => x"38",
          2725 => x"2e",
          2726 => x"0b",
          2727 => x"84",
          2728 => x"90",
          2729 => x"f8",
          2730 => x"d8",
          2731 => x"7d",
          2732 => x"f8",
          2733 => x"e5",
          2734 => x"38",
          2735 => x"33",
          2736 => x"ff",
          2737 => x"83",
          2738 => x"34",
          2739 => x"fe",
          2740 => x"e5",
          2741 => x"c7",
          2742 => x"70",
          2743 => x"fe",
          2744 => x"ff",
          2745 => x"58",
          2746 => x"33",
          2747 => x"84",
          2748 => x"83",
          2749 => x"ff",
          2750 => x"39",
          2751 => x"27",
          2752 => x"ff",
          2753 => x"b9",
          2754 => x"84",
          2755 => x"ff",
          2756 => x"5c",
          2757 => x"79",
          2758 => x"06",
          2759 => x"83",
          2760 => x"34",
          2761 => x"40",
          2762 => x"56",
          2763 => x"39",
          2764 => x"2e",
          2765 => x"84",
          2766 => x"26",
          2767 => x"84",
          2768 => x"83",
          2769 => x"86",
          2770 => x"22",
          2771 => x"83",
          2772 => x"46",
          2773 => x"2e",
          2774 => x"06",
          2775 => x"24",
          2776 => x"56",
          2777 => x"16",
          2778 => x"81",
          2779 => x"80",
          2780 => x"d7",
          2781 => x"38",
          2782 => x"34",
          2783 => x"22",
          2784 => x"90",
          2785 => x"81",
          2786 => x"5b",
          2787 => x"86",
          2788 => x"7f",
          2789 => x"42",
          2790 => x"d6",
          2791 => x"e0",
          2792 => x"33",
          2793 => x"70",
          2794 => x"05",
          2795 => x"33",
          2796 => x"1d",
          2797 => x"f7",
          2798 => x"84",
          2799 => x"05",
          2800 => x"33",
          2801 => x"18",
          2802 => x"33",
          2803 => x"58",
          2804 => x"e6",
          2805 => x"80",
          2806 => x"b8",
          2807 => x"ce",
          2808 => x"ff",
          2809 => x"40",
          2810 => x"b8",
          2811 => x"81",
          2812 => x"33",
          2813 => x"94",
          2814 => x"2e",
          2815 => x"40",
          2816 => x"81",
          2817 => x"fe",
          2818 => x"07",
          2819 => x"10",
          2820 => x"a7",
          2821 => x"86",
          2822 => x"58",
          2823 => x"83",
          2824 => x"f8",
          2825 => x"2b",
          2826 => x"79",
          2827 => x"27",
          2828 => x"59",
          2829 => x"0c",
          2830 => x"d8",
          2831 => x"7e",
          2832 => x"83",
          2833 => x"05",
          2834 => x"8c",
          2835 => x"29",
          2836 => x"57",
          2837 => x"83",
          2838 => x"59",
          2839 => x"79",
          2840 => x"17",
          2841 => x"a0",
          2842 => x"70",
          2843 => x"75",
          2844 => x"ff",
          2845 => x"fe",
          2846 => x"80",
          2847 => x"06",
          2848 => x"7b",
          2849 => x"38",
          2850 => x"81",
          2851 => x"f5",
          2852 => x"5e",
          2853 => x"83",
          2854 => x"83",
          2855 => x"42",
          2856 => x"f8",
          2857 => x"f8",
          2858 => x"06",
          2859 => x"90",
          2860 => x"75",
          2861 => x"f8",
          2862 => x"56",
          2863 => x"83",
          2864 => x"07",
          2865 => x"39",
          2866 => x"90",
          2867 => x"ff",
          2868 => x"90",
          2869 => x"59",
          2870 => x"33",
          2871 => x"90",
          2872 => x"33",
          2873 => x"83",
          2874 => x"f8",
          2875 => x"07",
          2876 => x"ea",
          2877 => x"06",
          2878 => x"90",
          2879 => x"33",
          2880 => x"83",
          2881 => x"f8",
          2882 => x"56",
          2883 => x"39",
          2884 => x"84",
          2885 => x"fe",
          2886 => x"fa",
          2887 => x"90",
          2888 => x"33",
          2889 => x"90",
          2890 => x"33",
          2891 => x"90",
          2892 => x"33",
          2893 => x"90",
          2894 => x"33",
          2895 => x"75",
          2896 => x"83",
          2897 => x"07",
          2898 => x"ba",
          2899 => x"80",
          2900 => x"ff",
          2901 => x"94",
          2902 => x"95",
          2903 => x"83",
          2904 => x"e0",
          2905 => x"b7",
          2906 => x"0c",
          2907 => x"95",
          2908 => x"ff",
          2909 => x"39",
          2910 => x"11",
          2911 => x"3f",
          2912 => x"b8",
          2913 => x"0b",
          2914 => x"b8",
          2915 => x"83",
          2916 => x"b7",
          2917 => x"84",
          2918 => x"06",
          2919 => x"b8",
          2920 => x"e4",
          2921 => x"95",
          2922 => x"3f",
          2923 => x"06",
          2924 => x"80",
          2925 => x"81",
          2926 => x"8a",
          2927 => x"39",
          2928 => x"09",
          2929 => x"57",
          2930 => x"d9",
          2931 => x"60",
          2932 => x"95",
          2933 => x"33",
          2934 => x"72",
          2935 => x"83",
          2936 => x"d7",
          2937 => x"78",
          2938 => x"bb",
          2939 => x"ff",
          2940 => x"a6",
          2941 => x"d8",
          2942 => x"95",
          2943 => x"a0",
          2944 => x"5f",
          2945 => x"ff",
          2946 => x"44",
          2947 => x"f5",
          2948 => x"11",
          2949 => x"38",
          2950 => x"27",
          2951 => x"83",
          2952 => x"ff",
          2953 => x"df",
          2954 => x"76",
          2955 => x"75",
          2956 => x"06",
          2957 => x"5a",
          2958 => x"31",
          2959 => x"71",
          2960 => x"a7",
          2961 => x"7c",
          2962 => x"71",
          2963 => x"79",
          2964 => x"b6",
          2965 => x"84",
          2966 => x"05",
          2967 => x"33",
          2968 => x"18",
          2969 => x"33",
          2970 => x"58",
          2971 => x"e0",
          2972 => x"33",
          2973 => x"70",
          2974 => x"05",
          2975 => x"33",
          2976 => x"1d",
          2977 => x"ff",
          2978 => x"96",
          2979 => x"33",
          2980 => x"b6",
          2981 => x"b6",
          2982 => x"e9",
          2983 => x"d7",
          2984 => x"5c",
          2985 => x"76",
          2986 => x"81",
          2987 => x"7a",
          2988 => x"f8",
          2989 => x"81",
          2990 => x"80",
          2991 => x"75",
          2992 => x"83",
          2993 => x"d8",
          2994 => x"7f",
          2995 => x"c5",
          2996 => x"f4",
          2997 => x"81",
          2998 => x"44",
          2999 => x"81",
          3000 => x"ff",
          3001 => x"fd",
          3002 => x"f8",
          3003 => x"31",
          3004 => x"90",
          3005 => x"26",
          3006 => x"05",
          3007 => x"70",
          3008 => x"f4",
          3009 => x"58",
          3010 => x"81",
          3011 => x"38",
          3012 => x"75",
          3013 => x"80",
          3014 => x"39",
          3015 => x"39",
          3016 => x"8e",
          3017 => x"f1",
          3018 => x"5a",
          3019 => x"80",
          3020 => x"39",
          3021 => x"84",
          3022 => x"2e",
          3023 => x"80",
          3024 => x"0d",
          3025 => x"3f",
          3026 => x"3d",
          3027 => x"05",
          3028 => x"33",
          3029 => x"11",
          3030 => x"2e",
          3031 => x"83",
          3032 => x"b8",
          3033 => x"f6",
          3034 => x"2e",
          3035 => x"71",
          3036 => x"5d",
          3037 => x"ff",
          3038 => x"81",
          3039 => x"32",
          3040 => x"5c",
          3041 => x"38",
          3042 => x"33",
          3043 => x"12",
          3044 => x"92",
          3045 => x"05",
          3046 => x"e9",
          3047 => x"2e",
          3048 => x"86",
          3049 => x"c0",
          3050 => x"08",
          3051 => x"ee",
          3052 => x"94",
          3053 => x"06",
          3054 => x"38",
          3055 => x"70",
          3056 => x"33",
          3057 => x"c1",
          3058 => x"38",
          3059 => x"81",
          3060 => x"85",
          3061 => x"34",
          3062 => x"8e",
          3063 => x"06",
          3064 => x"38",
          3065 => x"70",
          3066 => x"f6",
          3067 => x"86",
          3068 => x"54",
          3069 => x"81",
          3070 => x"81",
          3071 => x"38",
          3072 => x"0b",
          3073 => x"08",
          3074 => x"c0",
          3075 => x"42",
          3076 => x"16",
          3077 => x"38",
          3078 => x"80",
          3079 => x"16",
          3080 => x"38",
          3081 => x"81",
          3082 => x"73",
          3083 => x"ac",
          3084 => x"da",
          3085 => x"81",
          3086 => x"ac",
          3087 => x"80",
          3088 => x"05",
          3089 => x"73",
          3090 => x"87",
          3091 => x"0c",
          3092 => x"57",
          3093 => x"76",
          3094 => x"c0",
          3095 => x"26",
          3096 => x"c8",
          3097 => x"f6",
          3098 => x"38",
          3099 => x"08",
          3100 => x"38",
          3101 => x"54",
          3102 => x"73",
          3103 => x"9c",
          3104 => x"ff",
          3105 => x"83",
          3106 => x"e0",
          3107 => x"fc",
          3108 => x"72",
          3109 => x"2e",
          3110 => x"81",
          3111 => x"fe",
          3112 => x"59",
          3113 => x"2e",
          3114 => x"81",
          3115 => x"80",
          3116 => x"87",
          3117 => x"72",
          3118 => x"9c",
          3119 => x"76",
          3120 => x"71",
          3121 => x"80",
          3122 => x"10",
          3123 => x"78",
          3124 => x"5b",
          3125 => x"08",
          3126 => x"39",
          3127 => x"38",
          3128 => x"39",
          3129 => x"2e",
          3130 => x"da",
          3131 => x"e8",
          3132 => x"80",
          3133 => x"8a",
          3134 => x"f9",
          3135 => x"38",
          3136 => x"f6",
          3137 => x"7c",
          3138 => x"81",
          3139 => x"e2",
          3140 => x"80",
          3141 => x"33",
          3142 => x"ff",
          3143 => x"78",
          3144 => x"04",
          3145 => x"f6",
          3146 => x"83",
          3147 => x"7a",
          3148 => x"39",
          3149 => x"ff",
          3150 => x"0b",
          3151 => x"39",
          3152 => x"ff",
          3153 => x"16",
          3154 => x"38",
          3155 => x"2e",
          3156 => x"f6",
          3157 => x"98",
          3158 => x"fb",
          3159 => x"83",
          3160 => x"59",
          3161 => x"98",
          3162 => x"f6",
          3163 => x"72",
          3164 => x"34",
          3165 => x"f6",
          3166 => x"83",
          3167 => x"5d",
          3168 => x"9c",
          3169 => x"fc",
          3170 => x"fc",
          3171 => x"06",
          3172 => x"76",
          3173 => x"80",
          3174 => x"75",
          3175 => x"db",
          3176 => x"0b",
          3177 => x"83",
          3178 => x"34",
          3179 => x"83",
          3180 => x"38",
          3181 => x"ff",
          3182 => x"ff",
          3183 => x"79",
          3184 => x"f8",
          3185 => x"15",
          3186 => x"80",
          3187 => x"b6",
          3188 => x"ff",
          3189 => x"80",
          3190 => x"59",
          3191 => x"ff",
          3192 => x"39",
          3193 => x"08",
          3194 => x"f6",
          3195 => x"83",
          3196 => x"80",
          3197 => x"82",
          3198 => x"0b",
          3199 => x"a3",
          3200 => x"f0",
          3201 => x"0b",
          3202 => x"0b",
          3203 => x"80",
          3204 => x"83",
          3205 => x"05",
          3206 => x"87",
          3207 => x"2e",
          3208 => x"98",
          3209 => x"87",
          3210 => x"87",
          3211 => x"70",
          3212 => x"71",
          3213 => x"98",
          3214 => x"87",
          3215 => x"98",
          3216 => x"38",
          3217 => x"08",
          3218 => x"71",
          3219 => x"98",
          3220 => x"38",
          3221 => x"81",
          3222 => x"98",
          3223 => x"fe",
          3224 => x"76",
          3225 => x"04",
          3226 => x"3d",
          3227 => x"84",
          3228 => x"0b",
          3229 => x"87",
          3230 => x"2a",
          3231 => x"15",
          3232 => x"15",
          3233 => x"15",
          3234 => x"f0",
          3235 => x"f2",
          3236 => x"85",
          3237 => x"fe",
          3238 => x"f0",
          3239 => x"08",
          3240 => x"90",
          3241 => x"52",
          3242 => x"72",
          3243 => x"c0",
          3244 => x"27",
          3245 => x"38",
          3246 => x"55",
          3247 => x"55",
          3248 => x"c0",
          3249 => x"53",
          3250 => x"c0",
          3251 => x"f6",
          3252 => x"9c",
          3253 => x"38",
          3254 => x"c0",
          3255 => x"83",
          3256 => x"70",
          3257 => x"2e",
          3258 => x"52",
          3259 => x"81",
          3260 => x"c6",
          3261 => x"52",
          3262 => x"81",
          3263 => x"53",
          3264 => x"84",
          3265 => x"81",
          3266 => x"0d",
          3267 => x"0d",
          3268 => x"56",
          3269 => x"77",
          3270 => x"70",
          3271 => x"57",
          3272 => x"51",
          3273 => x"52",
          3274 => x"34",
          3275 => x"11",
          3276 => x"70",
          3277 => x"05",
          3278 => x"34",
          3279 => x"f0",
          3280 => x"f2",
          3281 => x"85",
          3282 => x"fe",
          3283 => x"f0",
          3284 => x"08",
          3285 => x"90",
          3286 => x"52",
          3287 => x"72",
          3288 => x"c0",
          3289 => x"27",
          3290 => x"38",
          3291 => x"55",
          3292 => x"55",
          3293 => x"c0",
          3294 => x"53",
          3295 => x"c0",
          3296 => x"f6",
          3297 => x"9c",
          3298 => x"38",
          3299 => x"c0",
          3300 => x"83",
          3301 => x"70",
          3302 => x"2e",
          3303 => x"71",
          3304 => x"ff",
          3305 => x"81",
          3306 => x"3d",
          3307 => x"3d",
          3308 => x"d0",
          3309 => x"08",
          3310 => x"80",
          3311 => x"c0",
          3312 => x"56",
          3313 => x"98",
          3314 => x"08",
          3315 => x"15",
          3316 => x"52",
          3317 => x"fe",
          3318 => x"08",
          3319 => x"c8",
          3320 => x"c0",
          3321 => x"ce",
          3322 => x"08",
          3323 => x"70",
          3324 => x"87",
          3325 => x"73",
          3326 => x"db",
          3327 => x"72",
          3328 => x"53",
          3329 => x"52",
          3330 => x"ff",
          3331 => x"39",
          3332 => x"fe",
          3333 => x"f9",
          3334 => x"71",
          3335 => x"06",
          3336 => x"81",
          3337 => x"2b",
          3338 => x"33",
          3339 => x"5c",
          3340 => x"52",
          3341 => x"af",
          3342 => x"12",
          3343 => x"07",
          3344 => x"71",
          3345 => x"53",
          3346 => x"24",
          3347 => x"14",
          3348 => x"07",
          3349 => x"56",
          3350 => x"ff",
          3351 => x"b8",
          3352 => x"85",
          3353 => x"88",
          3354 => x"84",
          3355 => x"b8",
          3356 => x"13",
          3357 => x"b8",
          3358 => x"73",
          3359 => x"16",
          3360 => x"2b",
          3361 => x"2a",
          3362 => x"75",
          3363 => x"86",
          3364 => x"2b",
          3365 => x"16",
          3366 => x"07",
          3367 => x"53",
          3368 => x"85",
          3369 => x"16",
          3370 => x"8b",
          3371 => x"5a",
          3372 => x"13",
          3373 => x"2a",
          3374 => x"34",
          3375 => x"08",
          3376 => x"88",
          3377 => x"88",
          3378 => x"34",
          3379 => x"08",
          3380 => x"71",
          3381 => x"05",
          3382 => x"2b",
          3383 => x"06",
          3384 => x"53",
          3385 => x"82",
          3386 => x"b8",
          3387 => x"12",
          3388 => x"07",
          3389 => x"71",
          3390 => x"70",
          3391 => x"57",
          3392 => x"14",
          3393 => x"82",
          3394 => x"2b",
          3395 => x"33",
          3396 => x"90",
          3397 => x"57",
          3398 => x"38",
          3399 => x"2b",
          3400 => x"2a",
          3401 => x"81",
          3402 => x"17",
          3403 => x"2b",
          3404 => x"14",
          3405 => x"07",
          3406 => x"58",
          3407 => x"75",
          3408 => x"f9",
          3409 => x"58",
          3410 => x"80",
          3411 => x"3f",
          3412 => x"0b",
          3413 => x"84",
          3414 => x"76",
          3415 => x"c6",
          3416 => x"75",
          3417 => x"b8",
          3418 => x"81",
          3419 => x"08",
          3420 => x"87",
          3421 => x"b8",
          3422 => x"07",
          3423 => x"2a",
          3424 => x"34",
          3425 => x"22",
          3426 => x"08",
          3427 => x"15",
          3428 => x"ee",
          3429 => x"53",
          3430 => x"fb",
          3431 => x"ff",
          3432 => x"ff",
          3433 => x"33",
          3434 => x"70",
          3435 => x"ff",
          3436 => x"75",
          3437 => x"12",
          3438 => x"ff",
          3439 => x"ff",
          3440 => x"5c",
          3441 => x"70",
          3442 => x"58",
          3443 => x"88",
          3444 => x"73",
          3445 => x"74",
          3446 => x"11",
          3447 => x"2b",
          3448 => x"56",
          3449 => x"83",
          3450 => x"26",
          3451 => x"2e",
          3452 => x"88",
          3453 => x"11",
          3454 => x"2a",
          3455 => x"34",
          3456 => x"08",
          3457 => x"82",
          3458 => x"b8",
          3459 => x"12",
          3460 => x"2b",
          3461 => x"83",
          3462 => x"58",
          3463 => x"12",
          3464 => x"83",
          3465 => x"54",
          3466 => x"84",
          3467 => x"33",
          3468 => x"83",
          3469 => x"53",
          3470 => x"15",
          3471 => x"55",
          3472 => x"33",
          3473 => x"54",
          3474 => x"71",
          3475 => x"70",
          3476 => x"71",
          3477 => x"05",
          3478 => x"15",
          3479 => x"d4",
          3480 => x"11",
          3481 => x"07",
          3482 => x"70",
          3483 => x"84",
          3484 => x"70",
          3485 => x"04",
          3486 => x"8b",
          3487 => x"84",
          3488 => x"2b",
          3489 => x"53",
          3490 => x"85",
          3491 => x"19",
          3492 => x"8b",
          3493 => x"86",
          3494 => x"2b",
          3495 => x"52",
          3496 => x"34",
          3497 => x"08",
          3498 => x"88",
          3499 => x"88",
          3500 => x"34",
          3501 => x"08",
          3502 => x"f9",
          3503 => x"58",
          3504 => x"54",
          3505 => x"0c",
          3506 => x"91",
          3507 => x"e4",
          3508 => x"f4",
          3509 => x"0b",
          3510 => x"53",
          3511 => x"cd",
          3512 => x"76",
          3513 => x"84",
          3514 => x"34",
          3515 => x"d4",
          3516 => x"0b",
          3517 => x"84",
          3518 => x"80",
          3519 => x"88",
          3520 => x"17",
          3521 => x"d0",
          3522 => x"d4",
          3523 => x"82",
          3524 => x"77",
          3525 => x"fe",
          3526 => x"41",
          3527 => x"59",
          3528 => x"38",
          3529 => x"80",
          3530 => x"60",
          3531 => x"2a",
          3532 => x"55",
          3533 => x"78",
          3534 => x"06",
          3535 => x"81",
          3536 => x"75",
          3537 => x"10",
          3538 => x"61",
          3539 => x"88",
          3540 => x"2c",
          3541 => x"43",
          3542 => x"42",
          3543 => x"15",
          3544 => x"07",
          3545 => x"81",
          3546 => x"2b",
          3547 => x"80",
          3548 => x"27",
          3549 => x"62",
          3550 => x"85",
          3551 => x"25",
          3552 => x"79",
          3553 => x"33",
          3554 => x"83",
          3555 => x"12",
          3556 => x"07",
          3557 => x"58",
          3558 => x"1e",
          3559 => x"8b",
          3560 => x"86",
          3561 => x"2b",
          3562 => x"14",
          3563 => x"07",
          3564 => x"5b",
          3565 => x"84",
          3566 => x"b8",
          3567 => x"85",
          3568 => x"2b",
          3569 => x"15",
          3570 => x"2a",
          3571 => x"57",
          3572 => x"34",
          3573 => x"81",
          3574 => x"ff",
          3575 => x"5e",
          3576 => x"34",
          3577 => x"11",
          3578 => x"71",
          3579 => x"81",
          3580 => x"88",
          3581 => x"55",
          3582 => x"34",
          3583 => x"33",
          3584 => x"83",
          3585 => x"83",
          3586 => x"88",
          3587 => x"55",
          3588 => x"1a",
          3589 => x"82",
          3590 => x"2b",
          3591 => x"2b",
          3592 => x"05",
          3593 => x"d4",
          3594 => x"1c",
          3595 => x"5f",
          3596 => x"54",
          3597 => x"0d",
          3598 => x"d4",
          3599 => x"23",
          3600 => x"ff",
          3601 => x"b8",
          3602 => x"0b",
          3603 => x"5d",
          3604 => x"1e",
          3605 => x"86",
          3606 => x"84",
          3607 => x"ff",
          3608 => x"ff",
          3609 => x"5b",
          3610 => x"18",
          3611 => x"10",
          3612 => x"05",
          3613 => x"0b",
          3614 => x"57",
          3615 => x"82",
          3616 => x"fe",
          3617 => x"84",
          3618 => x"95",
          3619 => x"d4",
          3620 => x"44",
          3621 => x"71",
          3622 => x"70",
          3623 => x"63",
          3624 => x"84",
          3625 => x"57",
          3626 => x"19",
          3627 => x"70",
          3628 => x"07",
          3629 => x"74",
          3630 => x"88",
          3631 => x"5d",
          3632 => x"ff",
          3633 => x"84",
          3634 => x"34",
          3635 => x"d4",
          3636 => x"3f",
          3637 => x"31",
          3638 => x"fa",
          3639 => x"76",
          3640 => x"17",
          3641 => x"07",
          3642 => x"81",
          3643 => x"2b",
          3644 => x"45",
          3645 => x"ff",
          3646 => x"38",
          3647 => x"83",
          3648 => x"fc",
          3649 => x"f4",
          3650 => x"0b",
          3651 => x"53",
          3652 => x"c4",
          3653 => x"7e",
          3654 => x"84",
          3655 => x"34",
          3656 => x"d4",
          3657 => x"0b",
          3658 => x"84",
          3659 => x"80",
          3660 => x"88",
          3661 => x"88",
          3662 => x"84",
          3663 => x"84",
          3664 => x"43",
          3665 => x"83",
          3666 => x"24",
          3667 => x"06",
          3668 => x"fc",
          3669 => x"38",
          3670 => x"73",
          3671 => x"04",
          3672 => x"33",
          3673 => x"7a",
          3674 => x"71",
          3675 => x"05",
          3676 => x"88",
          3677 => x"45",
          3678 => x"56",
          3679 => x"85",
          3680 => x"17",
          3681 => x"8b",
          3682 => x"86",
          3683 => x"2b",
          3684 => x"48",
          3685 => x"05",
          3686 => x"b8",
          3687 => x"33",
          3688 => x"06",
          3689 => x"7b",
          3690 => x"b8",
          3691 => x"83",
          3692 => x"2b",
          3693 => x"33",
          3694 => x"5e",
          3695 => x"76",
          3696 => x"b8",
          3697 => x"12",
          3698 => x"07",
          3699 => x"33",
          3700 => x"40",
          3701 => x"78",
          3702 => x"84",
          3703 => x"33",
          3704 => x"66",
          3705 => x"52",
          3706 => x"fe",
          3707 => x"1e",
          3708 => x"5c",
          3709 => x"0b",
          3710 => x"84",
          3711 => x"7f",
          3712 => x"fe",
          3713 => x"76",
          3714 => x"b8",
          3715 => x"81",
          3716 => x"08",
          3717 => x"87",
          3718 => x"b8",
          3719 => x"07",
          3720 => x"2a",
          3721 => x"34",
          3722 => x"22",
          3723 => x"08",
          3724 => x"1c",
          3725 => x"51",
          3726 => x"39",
          3727 => x"8b",
          3728 => x"84",
          3729 => x"2b",
          3730 => x"43",
          3731 => x"63",
          3732 => x"08",
          3733 => x"33",
          3734 => x"74",
          3735 => x"71",
          3736 => x"5f",
          3737 => x"64",
          3738 => x"34",
          3739 => x"81",
          3740 => x"ff",
          3741 => x"58",
          3742 => x"34",
          3743 => x"33",
          3744 => x"83",
          3745 => x"12",
          3746 => x"2b",
          3747 => x"88",
          3748 => x"5d",
          3749 => x"83",
          3750 => x"1f",
          3751 => x"2b",
          3752 => x"33",
          3753 => x"81",
          3754 => x"5d",
          3755 => x"60",
          3756 => x"83",
          3757 => x"86",
          3758 => x"2b",
          3759 => x"18",
          3760 => x"07",
          3761 => x"41",
          3762 => x"1e",
          3763 => x"84",
          3764 => x"2b",
          3765 => x"14",
          3766 => x"07",
          3767 => x"5a",
          3768 => x"34",
          3769 => x"d4",
          3770 => x"71",
          3771 => x"70",
          3772 => x"75",
          3773 => x"d4",
          3774 => x"33",
          3775 => x"74",
          3776 => x"88",
          3777 => x"f8",
          3778 => x"54",
          3779 => x"7f",
          3780 => x"84",
          3781 => x"81",
          3782 => x"2b",
          3783 => x"33",
          3784 => x"06",
          3785 => x"5b",
          3786 => x"81",
          3787 => x"1f",
          3788 => x"8b",
          3789 => x"86",
          3790 => x"2b",
          3791 => x"14",
          3792 => x"07",
          3793 => x"5c",
          3794 => x"77",
          3795 => x"84",
          3796 => x"33",
          3797 => x"83",
          3798 => x"87",
          3799 => x"88",
          3800 => x"41",
          3801 => x"16",
          3802 => x"33",
          3803 => x"81",
          3804 => x"5c",
          3805 => x"1a",
          3806 => x"82",
          3807 => x"2b",
          3808 => x"33",
          3809 => x"70",
          3810 => x"5a",
          3811 => x"1a",
          3812 => x"70",
          3813 => x"71",
          3814 => x"33",
          3815 => x"70",
          3816 => x"5a",
          3817 => x"83",
          3818 => x"1f",
          3819 => x"88",
          3820 => x"83",
          3821 => x"84",
          3822 => x"b8",
          3823 => x"05",
          3824 => x"44",
          3825 => x"87",
          3826 => x"2b",
          3827 => x"1d",
          3828 => x"2a",
          3829 => x"61",
          3830 => x"34",
          3831 => x"11",
          3832 => x"71",
          3833 => x"33",
          3834 => x"70",
          3835 => x"59",
          3836 => x"7a",
          3837 => x"08",
          3838 => x"88",
          3839 => x"88",
          3840 => x"34",
          3841 => x"08",
          3842 => x"71",
          3843 => x"05",
          3844 => x"2b",
          3845 => x"06",
          3846 => x"5c",
          3847 => x"82",
          3848 => x"b8",
          3849 => x"12",
          3850 => x"07",
          3851 => x"71",
          3852 => x"70",
          3853 => x"59",
          3854 => x"1e",
          3855 => x"f3",
          3856 => x"a1",
          3857 => x"b8",
          3858 => x"53",
          3859 => x"fe",
          3860 => x"3f",
          3861 => x"38",
          3862 => x"7a",
          3863 => x"76",
          3864 => x"8a",
          3865 => x"3d",
          3866 => x"84",
          3867 => x"08",
          3868 => x"52",
          3869 => x"96",
          3870 => x"3d",
          3871 => x"b8",
          3872 => x"d0",
          3873 => x"84",
          3874 => x"84",
          3875 => x"81",
          3876 => x"08",
          3877 => x"85",
          3878 => x"76",
          3879 => x"34",
          3880 => x"22",
          3881 => x"83",
          3882 => x"51",
          3883 => x"89",
          3884 => x"10",
          3885 => x"f8",
          3886 => x"81",
          3887 => x"80",
          3888 => x"ff",
          3889 => x"81",
          3890 => x"b8",
          3891 => x"e4",
          3892 => x"0d",
          3893 => x"71",
          3894 => x"bb",
          3895 => x"06",
          3896 => x"e0",
          3897 => x"53",
          3898 => x"0d",
          3899 => x"02",
          3900 => x"57",
          3901 => x"38",
          3902 => x"81",
          3903 => x"73",
          3904 => x"0c",
          3905 => x"ca",
          3906 => x"06",
          3907 => x"c0",
          3908 => x"79",
          3909 => x"80",
          3910 => x"81",
          3911 => x"0c",
          3912 => x"81",
          3913 => x"56",
          3914 => x"39",
          3915 => x"8c",
          3916 => x"59",
          3917 => x"84",
          3918 => x"06",
          3919 => x"58",
          3920 => x"78",
          3921 => x"3f",
          3922 => x"55",
          3923 => x"98",
          3924 => x"78",
          3925 => x"06",
          3926 => x"54",
          3927 => x"8b",
          3928 => x"19",
          3929 => x"79",
          3930 => x"fc",
          3931 => x"05",
          3932 => x"53",
          3933 => x"87",
          3934 => x"72",
          3935 => x"38",
          3936 => x"81",
          3937 => x"71",
          3938 => x"38",
          3939 => x"86",
          3940 => x"0c",
          3941 => x"0d",
          3942 => x"84",
          3943 => x"71",
          3944 => x"53",
          3945 => x"81",
          3946 => x"2e",
          3947 => x"55",
          3948 => x"08",
          3949 => x"87",
          3950 => x"82",
          3951 => x"38",
          3952 => x"38",
          3953 => x"58",
          3954 => x"56",
          3955 => x"a8",
          3956 => x"81",
          3957 => x"18",
          3958 => x"e4",
          3959 => x"78",
          3960 => x"04",
          3961 => x"18",
          3962 => x"fc",
          3963 => x"08",
          3964 => x"84",
          3965 => x"18",
          3966 => x"1a",
          3967 => x"56",
          3968 => x"82",
          3969 => x"81",
          3970 => x"1b",
          3971 => x"fc",
          3972 => x"75",
          3973 => x"38",
          3974 => x"09",
          3975 => x"5a",
          3976 => x"70",
          3977 => x"76",
          3978 => x"19",
          3979 => x"34",
          3980 => x"b9",
          3981 => x"34",
          3982 => x"f2",
          3983 => x"0b",
          3984 => x"84",
          3985 => x"9f",
          3986 => x"84",
          3987 => x"7a",
          3988 => x"56",
          3989 => x"2a",
          3990 => x"18",
          3991 => x"7a",
          3992 => x"34",
          3993 => x"19",
          3994 => x"a7",
          3995 => x"70",
          3996 => x"53",
          3997 => x"e8",
          3998 => x"80",
          3999 => x"3f",
          4000 => x"b7",
          4001 => x"60",
          4002 => x"76",
          4003 => x"26",
          4004 => x"e4",
          4005 => x"33",
          4006 => x"38",
          4007 => x"81",
          4008 => x"81",
          4009 => x"08",
          4010 => x"08",
          4011 => x"5c",
          4012 => x"de",
          4013 => x"52",
          4014 => x"84",
          4015 => x"ff",
          4016 => x"7a",
          4017 => x"17",
          4018 => x"2a",
          4019 => x"59",
          4020 => x"80",
          4021 => x"5d",
          4022 => x"b5",
          4023 => x"52",
          4024 => x"84",
          4025 => x"ff",
          4026 => x"79",
          4027 => x"17",
          4028 => x"07",
          4029 => x"5d",
          4030 => x"76",
          4031 => x"8f",
          4032 => x"18",
          4033 => x"2e",
          4034 => x"71",
          4035 => x"81",
          4036 => x"53",
          4037 => x"f7",
          4038 => x"2e",
          4039 => x"b4",
          4040 => x"10",
          4041 => x"81",
          4042 => x"07",
          4043 => x"3d",
          4044 => x"06",
          4045 => x"18",
          4046 => x"2e",
          4047 => x"71",
          4048 => x"81",
          4049 => x"53",
          4050 => x"f6",
          4051 => x"2e",
          4052 => x"b4",
          4053 => x"82",
          4054 => x"05",
          4055 => x"90",
          4056 => x"33",
          4057 => x"71",
          4058 => x"84",
          4059 => x"5a",
          4060 => x"b4",
          4061 => x"81",
          4062 => x"81",
          4063 => x"09",
          4064 => x"e4",
          4065 => x"a8",
          4066 => x"5b",
          4067 => x"84",
          4068 => x"2e",
          4069 => x"54",
          4070 => x"53",
          4071 => x"98",
          4072 => x"54",
          4073 => x"53",
          4074 => x"3f",
          4075 => x"81",
          4076 => x"08",
          4077 => x"18",
          4078 => x"27",
          4079 => x"82",
          4080 => x"08",
          4081 => x"17",
          4082 => x"18",
          4083 => x"5a",
          4084 => x"81",
          4085 => x"08",
          4086 => x"18",
          4087 => x"5e",
          4088 => x"38",
          4089 => x"09",
          4090 => x"b4",
          4091 => x"7b",
          4092 => x"3f",
          4093 => x"b4",
          4094 => x"81",
          4095 => x"81",
          4096 => x"09",
          4097 => x"e4",
          4098 => x"a8",
          4099 => x"5b",
          4100 => x"91",
          4101 => x"2e",
          4102 => x"54",
          4103 => x"53",
          4104 => x"90",
          4105 => x"54",
          4106 => x"53",
          4107 => x"f8",
          4108 => x"f9",
          4109 => x"0d",
          4110 => x"58",
          4111 => x"1a",
          4112 => x"74",
          4113 => x"81",
          4114 => x"38",
          4115 => x"0d",
          4116 => x"05",
          4117 => x"5c",
          4118 => x"19",
          4119 => x"09",
          4120 => x"77",
          4121 => x"51",
          4122 => x"80",
          4123 => x"77",
          4124 => x"b0",
          4125 => x"05",
          4126 => x"76",
          4127 => x"79",
          4128 => x"34",
          4129 => x"0d",
          4130 => x"fe",
          4131 => x"08",
          4132 => x"58",
          4133 => x"83",
          4134 => x"2e",
          4135 => x"54",
          4136 => x"33",
          4137 => x"08",
          4138 => x"5a",
          4139 => x"fe",
          4140 => x"06",
          4141 => x"70",
          4142 => x"0a",
          4143 => x"7d",
          4144 => x"1d",
          4145 => x"1d",
          4146 => x"1d",
          4147 => x"e8",
          4148 => x"2a",
          4149 => x"59",
          4150 => x"80",
          4151 => x"5d",
          4152 => x"d4",
          4153 => x"52",
          4154 => x"84",
          4155 => x"ff",
          4156 => x"7b",
          4157 => x"ff",
          4158 => x"81",
          4159 => x"80",
          4160 => x"f0",
          4161 => x"56",
          4162 => x"1a",
          4163 => x"05",
          4164 => x"5f",
          4165 => x"54",
          4166 => x"1a",
          4167 => x"58",
          4168 => x"81",
          4169 => x"08",
          4170 => x"a8",
          4171 => x"b8",
          4172 => x"7a",
          4173 => x"74",
          4174 => x"75",
          4175 => x"ee",
          4176 => x"2e",
          4177 => x"b4",
          4178 => x"83",
          4179 => x"2a",
          4180 => x"2a",
          4181 => x"06",
          4182 => x"0b",
          4183 => x"54",
          4184 => x"1a",
          4185 => x"5a",
          4186 => x"81",
          4187 => x"08",
          4188 => x"a8",
          4189 => x"b8",
          4190 => x"77",
          4191 => x"55",
          4192 => x"bd",
          4193 => x"52",
          4194 => x"7b",
          4195 => x"53",
          4196 => x"52",
          4197 => x"b8",
          4198 => x"fd",
          4199 => x"1a",
          4200 => x"08",
          4201 => x"08",
          4202 => x"fc",
          4203 => x"82",
          4204 => x"81",
          4205 => x"19",
          4206 => x"fc",
          4207 => x"19",
          4208 => x"ed",
          4209 => x"08",
          4210 => x"38",
          4211 => x"b4",
          4212 => x"a0",
          4213 => x"5f",
          4214 => x"38",
          4215 => x"09",
          4216 => x"7c",
          4217 => x"51",
          4218 => x"39",
          4219 => x"81",
          4220 => x"58",
          4221 => x"fe",
          4222 => x"06",
          4223 => x"76",
          4224 => x"f9",
          4225 => x"7b",
          4226 => x"05",
          4227 => x"2b",
          4228 => x"07",
          4229 => x"34",
          4230 => x"34",
          4231 => x"34",
          4232 => x"34",
          4233 => x"7e",
          4234 => x"8a",
          4235 => x"2e",
          4236 => x"27",
          4237 => x"56",
          4238 => x"76",
          4239 => x"81",
          4240 => x"89",
          4241 => x"b2",
          4242 => x"3f",
          4243 => x"d0",
          4244 => x"81",
          4245 => x"09",
          4246 => x"70",
          4247 => x"82",
          4248 => x"06",
          4249 => x"b8",
          4250 => x"57",
          4251 => x"58",
          4252 => x"a4",
          4253 => x"08",
          4254 => x"55",
          4255 => x"38",
          4256 => x"26",
          4257 => x"81",
          4258 => x"83",
          4259 => x"ef",
          4260 => x"08",
          4261 => x"e4",
          4262 => x"80",
          4263 => x"08",
          4264 => x"85",
          4265 => x"9a",
          4266 => x"27",
          4267 => x"27",
          4268 => x"fe",
          4269 => x"38",
          4270 => x"f5",
          4271 => x"e4",
          4272 => x"07",
          4273 => x"c4",
          4274 => x"1a",
          4275 => x"1a",
          4276 => x"38",
          4277 => x"33",
          4278 => x"75",
          4279 => x"3d",
          4280 => x"0c",
          4281 => x"08",
          4282 => x"ff",
          4283 => x"51",
          4284 => x"55",
          4285 => x"84",
          4286 => x"ff",
          4287 => x"81",
          4288 => x"7a",
          4289 => x"f0",
          4290 => x"9f",
          4291 => x"90",
          4292 => x"80",
          4293 => x"26",
          4294 => x"82",
          4295 => x"79",
          4296 => x"19",
          4297 => x"08",
          4298 => x"38",
          4299 => x"73",
          4300 => x"19",
          4301 => x"0c",
          4302 => x"b8",
          4303 => x"17",
          4304 => x"38",
          4305 => x"59",
          4306 => x"08",
          4307 => x"80",
          4308 => x"17",
          4309 => x"05",
          4310 => x"91",
          4311 => x"3f",
          4312 => x"e4",
          4313 => x"84",
          4314 => x"9c",
          4315 => x"73",
          4316 => x"54",
          4317 => x"39",
          4318 => x"3d",
          4319 => x"08",
          4320 => x"57",
          4321 => x"80",
          4322 => x"55",
          4323 => x"79",
          4324 => x"81",
          4325 => x"a9",
          4326 => x"57",
          4327 => x"77",
          4328 => x"78",
          4329 => x"56",
          4330 => x"0d",
          4331 => x"22",
          4332 => x"7b",
          4333 => x"9c",
          4334 => x"56",
          4335 => x"d0",
          4336 => x"ff",
          4337 => x"b8",
          4338 => x"80",
          4339 => x"52",
          4340 => x"e4",
          4341 => x"08",
          4342 => x"84",
          4343 => x"38",
          4344 => x"2e",
          4345 => x"83",
          4346 => x"38",
          4347 => x"59",
          4348 => x"38",
          4349 => x"1b",
          4350 => x"0c",
          4351 => x"55",
          4352 => x"ff",
          4353 => x"8a",
          4354 => x"80",
          4355 => x"52",
          4356 => x"84",
          4357 => x"16",
          4358 => x"84",
          4359 => x"0d",
          4360 => x"b8",
          4361 => x"56",
          4362 => x"80",
          4363 => x"1a",
          4364 => x"31",
          4365 => x"e8",
          4366 => x"2e",
          4367 => x"54",
          4368 => x"53",
          4369 => x"c8",
          4370 => x"55",
          4371 => x"76",
          4372 => x"94",
          4373 => x"fe",
          4374 => x"27",
          4375 => x"71",
          4376 => x"0c",
          4377 => x"b8",
          4378 => x"3d",
          4379 => x"08",
          4380 => x"08",
          4381 => x"d2",
          4382 => x"58",
          4383 => x"38",
          4384 => x"78",
          4385 => x"81",
          4386 => x"19",
          4387 => x"e4",
          4388 => x"81",
          4389 => x"76",
          4390 => x"33",
          4391 => x"38",
          4392 => x"ff",
          4393 => x"76",
          4394 => x"32",
          4395 => x"25",
          4396 => x"93",
          4397 => x"61",
          4398 => x"2e",
          4399 => x"52",
          4400 => x"e4",
          4401 => x"b2",
          4402 => x"dc",
          4403 => x"3d",
          4404 => x"53",
          4405 => x"a8",
          4406 => x"78",
          4407 => x"84",
          4408 => x"19",
          4409 => x"e4",
          4410 => x"27",
          4411 => x"60",
          4412 => x"38",
          4413 => x"08",
          4414 => x"51",
          4415 => x"39",
          4416 => x"e7",
          4417 => x"7a",
          4418 => x"77",
          4419 => x"7f",
          4420 => x"7d",
          4421 => x"5d",
          4422 => x"2e",
          4423 => x"39",
          4424 => x"7a",
          4425 => x"04",
          4426 => x"33",
          4427 => x"cb",
          4428 => x"9a",
          4429 => x"56",
          4430 => x"70",
          4431 => x"51",
          4432 => x"e4",
          4433 => x"71",
          4434 => x"56",
          4435 => x"81",
          4436 => x"61",
          4437 => x"81",
          4438 => x"27",
          4439 => x"81",
          4440 => x"38",
          4441 => x"79",
          4442 => x"ff",
          4443 => x"fd",
          4444 => x"ca",
          4445 => x"7c",
          4446 => x"81",
          4447 => x"70",
          4448 => x"70",
          4449 => x"59",
          4450 => x"81",
          4451 => x"84",
          4452 => x"ef",
          4453 => x"80",
          4454 => x"b8",
          4455 => x"82",
          4456 => x"ff",
          4457 => x"98",
          4458 => x"08",
          4459 => x"33",
          4460 => x"81",
          4461 => x"53",
          4462 => x"dc",
          4463 => x"2e",
          4464 => x"b4",
          4465 => x"38",
          4466 => x"76",
          4467 => x"33",
          4468 => x"58",
          4469 => x"2e",
          4470 => x"06",
          4471 => x"74",
          4472 => x"e5",
          4473 => x"58",
          4474 => x"80",
          4475 => x"33",
          4476 => x"ff",
          4477 => x"74",
          4478 => x"33",
          4479 => x"0b",
          4480 => x"05",
          4481 => x"33",
          4482 => x"42",
          4483 => x"75",
          4484 => x"ff",
          4485 => x"51",
          4486 => x"5a",
          4487 => x"8f",
          4488 => x"3d",
          4489 => x"53",
          4490 => x"80",
          4491 => x"78",
          4492 => x"84",
          4493 => x"1b",
          4494 => x"e4",
          4495 => x"27",
          4496 => x"79",
          4497 => x"38",
          4498 => x"08",
          4499 => x"51",
          4500 => x"39",
          4501 => x"33",
          4502 => x"60",
          4503 => x"06",
          4504 => x"19",
          4505 => x"1f",
          4506 => x"5f",
          4507 => x"55",
          4508 => x"92",
          4509 => x"b8",
          4510 => x"fe",
          4511 => x"38",
          4512 => x"0c",
          4513 => x"7e",
          4514 => x"8c",
          4515 => x"33",
          4516 => x"76",
          4517 => x"06",
          4518 => x"77",
          4519 => x"79",
          4520 => x"88",
          4521 => x"2e",
          4522 => x"ff",
          4523 => x"3f",
          4524 => x"05",
          4525 => x"56",
          4526 => x"e4",
          4527 => x"38",
          4528 => x"27",
          4529 => x"2a",
          4530 => x"92",
          4531 => x"10",
          4532 => x"fe",
          4533 => x"06",
          4534 => x"84",
          4535 => x"76",
          4536 => x"81",
          4537 => x"0d",
          4538 => x"81",
          4539 => x"56",
          4540 => x"08",
          4541 => x"2e",
          4542 => x"70",
          4543 => x"95",
          4544 => x"7b",
          4545 => x"57",
          4546 => x"ff",
          4547 => x"db",
          4548 => x"76",
          4549 => x"0b",
          4550 => x"40",
          4551 => x"8b",
          4552 => x"81",
          4553 => x"58",
          4554 => x"85",
          4555 => x"22",
          4556 => x"74",
          4557 => x"81",
          4558 => x"70",
          4559 => x"81",
          4560 => x"2e",
          4561 => x"57",
          4562 => x"38",
          4563 => x"02",
          4564 => x"76",
          4565 => x"27",
          4566 => x"34",
          4567 => x"59",
          4568 => x"59",
          4569 => x"56",
          4570 => x"55",
          4571 => x"56",
          4572 => x"1a",
          4573 => x"09",
          4574 => x"a0",
          4575 => x"3d",
          4576 => x"33",
          4577 => x"76",
          4578 => x"8f",
          4579 => x"81",
          4580 => x"91",
          4581 => x"82",
          4582 => x"84",
          4583 => x"06",
          4584 => x"33",
          4585 => x"05",
          4586 => x"81",
          4587 => x"80",
          4588 => x"51",
          4589 => x"08",
          4590 => x"8c",
          4591 => x"b8",
          4592 => x"e4",
          4593 => x"08",
          4594 => x"2e",
          4595 => x"7f",
          4596 => x"38",
          4597 => x"81",
          4598 => x"b8",
          4599 => x"56",
          4600 => x"56",
          4601 => x"33",
          4602 => x"c9",
          4603 => x"07",
          4604 => x"38",
          4605 => x"89",
          4606 => x"3f",
          4607 => x"e4",
          4608 => x"58",
          4609 => x"58",
          4610 => x"7f",
          4611 => x"b4",
          4612 => x"1c",
          4613 => x"38",
          4614 => x"81",
          4615 => x"b8",
          4616 => x"57",
          4617 => x"58",
          4618 => x"1f",
          4619 => x"05",
          4620 => x"38",
          4621 => x"58",
          4622 => x"77",
          4623 => x"55",
          4624 => x"1f",
          4625 => x"1b",
          4626 => x"56",
          4627 => x"0d",
          4628 => x"72",
          4629 => x"38",
          4630 => x"c2",
          4631 => x"b8",
          4632 => x"fe",
          4633 => x"53",
          4634 => x"80",
          4635 => x"09",
          4636 => x"e4",
          4637 => x"a8",
          4638 => x"08",
          4639 => x"60",
          4640 => x"e4",
          4641 => x"2b",
          4642 => x"7d",
          4643 => x"08",
          4644 => x"38",
          4645 => x"8b",
          4646 => x"29",
          4647 => x"57",
          4648 => x"19",
          4649 => x"81",
          4650 => x"1e",
          4651 => x"77",
          4652 => x"7a",
          4653 => x"38",
          4654 => x"81",
          4655 => x"b8",
          4656 => x"57",
          4657 => x"58",
          4658 => x"9c",
          4659 => x"5c",
          4660 => x"8b",
          4661 => x"9a",
          4662 => x"8d",
          4663 => x"59",
          4664 => x"78",
          4665 => x"58",
          4666 => x"05",
          4667 => x"34",
          4668 => x"76",
          4669 => x"18",
          4670 => x"83",
          4671 => x"10",
          4672 => x"2e",
          4673 => x"0b",
          4674 => x"e9",
          4675 => x"84",
          4676 => x"ff",
          4677 => x"eb",
          4678 => x"b8",
          4679 => x"59",
          4680 => x"e4",
          4681 => x"08",
          4682 => x"1d",
          4683 => x"41",
          4684 => x"38",
          4685 => x"09",
          4686 => x"b4",
          4687 => x"78",
          4688 => x"3f",
          4689 => x"1f",
          4690 => x"81",
          4691 => x"38",
          4692 => x"76",
          4693 => x"39",
          4694 => x"39",
          4695 => x"52",
          4696 => x"84",
          4697 => x"06",
          4698 => x"1d",
          4699 => x"31",
          4700 => x"38",
          4701 => x"aa",
          4702 => x"f8",
          4703 => x"80",
          4704 => x"75",
          4705 => x"59",
          4706 => x"fa",
          4707 => x"a0",
          4708 => x"1c",
          4709 => x"39",
          4710 => x"08",
          4711 => x"51",
          4712 => x"3d",
          4713 => x"5c",
          4714 => x"08",
          4715 => x"08",
          4716 => x"71",
          4717 => x"58",
          4718 => x"38",
          4719 => x"1b",
          4720 => x"80",
          4721 => x"06",
          4722 => x"83",
          4723 => x"22",
          4724 => x"7a",
          4725 => x"06",
          4726 => x"57",
          4727 => x"89",
          4728 => x"16",
          4729 => x"74",
          4730 => x"81",
          4731 => x"70",
          4732 => x"77",
          4733 => x"8b",
          4734 => x"34",
          4735 => x"05",
          4736 => x"27",
          4737 => x"55",
          4738 => x"33",
          4739 => x"38",
          4740 => x"7c",
          4741 => x"17",
          4742 => x"55",
          4743 => x"34",
          4744 => x"88",
          4745 => x"83",
          4746 => x"2b",
          4747 => x"70",
          4748 => x"07",
          4749 => x"17",
          4750 => x"5b",
          4751 => x"1e",
          4752 => x"71",
          4753 => x"1e",
          4754 => x"55",
          4755 => x"81",
          4756 => x"b5",
          4757 => x"81",
          4758 => x"83",
          4759 => x"27",
          4760 => x"38",
          4761 => x"74",
          4762 => x"80",
          4763 => x"19",
          4764 => x"79",
          4765 => x"30",
          4766 => x"72",
          4767 => x"80",
          4768 => x"05",
          4769 => x"5b",
          4770 => x"5a",
          4771 => x"38",
          4772 => x"89",
          4773 => x"78",
          4774 => x"8c",
          4775 => x"b4",
          4776 => x"06",
          4777 => x"14",
          4778 => x"73",
          4779 => x"16",
          4780 => x"33",
          4781 => x"b7",
          4782 => x"53",
          4783 => x"25",
          4784 => x"58",
          4785 => x"70",
          4786 => x"70",
          4787 => x"83",
          4788 => x"81",
          4789 => x"38",
          4790 => x"33",
          4791 => x"9f",
          4792 => x"8c",
          4793 => x"70",
          4794 => x"81",
          4795 => x"2e",
          4796 => x"27",
          4797 => x"76",
          4798 => x"ff",
          4799 => x"73",
          4800 => x"5b",
          4801 => x"dc",
          4802 => x"26",
          4803 => x"e4",
          4804 => x"54",
          4805 => x"73",
          4806 => x"33",
          4807 => x"73",
          4808 => x"7a",
          4809 => x"80",
          4810 => x"7d",
          4811 => x"05",
          4812 => x"2e",
          4813 => x"73",
          4814 => x"25",
          4815 => x"80",
          4816 => x"54",
          4817 => x"2e",
          4818 => x"30",
          4819 => x"57",
          4820 => x"73",
          4821 => x"55",
          4822 => x"39",
          4823 => x"e7",
          4824 => x"ff",
          4825 => x"54",
          4826 => x"0d",
          4827 => x"ff",
          4828 => x"e3",
          4829 => x"1d",
          4830 => x"3f",
          4831 => x"0c",
          4832 => x"dc",
          4833 => x"07",
          4834 => x"a1",
          4835 => x"33",
          4836 => x"38",
          4837 => x"80",
          4838 => x"e1",
          4839 => x"82",
          4840 => x"38",
          4841 => x"17",
          4842 => x"17",
          4843 => x"a0",
          4844 => x"42",
          4845 => x"84",
          4846 => x"76",
          4847 => x"80",
          4848 => x"38",
          4849 => x"06",
          4850 => x"2e",
          4851 => x"06",
          4852 => x"76",
          4853 => x"05",
          4854 => x"9d",
          4855 => x"ff",
          4856 => x"fe",
          4857 => x"2e",
          4858 => x"a0",
          4859 => x"05",
          4860 => x"38",
          4861 => x"70",
          4862 => x"74",
          4863 => x"2e",
          4864 => x"30",
          4865 => x"77",
          4866 => x"38",
          4867 => x"81",
          4868 => x"72",
          4869 => x"51",
          4870 => x"38",
          4871 => x"77",
          4872 => x"75",
          4873 => x"5b",
          4874 => x"77",
          4875 => x"22",
          4876 => x"95",
          4877 => x"e5",
          4878 => x"82",
          4879 => x"8c",
          4880 => x"55",
          4881 => x"81",
          4882 => x"7d",
          4883 => x"38",
          4884 => x"81",
          4885 => x"79",
          4886 => x"7b",
          4887 => x"08",
          4888 => x"e4",
          4889 => x"b8",
          4890 => x"fb",
          4891 => x"5a",
          4892 => x"82",
          4893 => x"38",
          4894 => x"8c",
          4895 => x"39",
          4896 => x"22",
          4897 => x"f0",
          4898 => x"79",
          4899 => x"18",
          4900 => x"06",
          4901 => x"ae",
          4902 => x"76",
          4903 => x"0b",
          4904 => x"73",
          4905 => x"70",
          4906 => x"8a",
          4907 => x"58",
          4908 => x"bf",
          4909 => x"33",
          4910 => x"d6",
          4911 => x"77",
          4912 => x"84",
          4913 => x"2e",
          4914 => x"ff",
          4915 => x"80",
          4916 => x"62",
          4917 => x"2e",
          4918 => x"7b",
          4919 => x"77",
          4920 => x"38",
          4921 => x"fb",
          4922 => x"56",
          4923 => x"81",
          4924 => x"77",
          4925 => x"38",
          4926 => x"85",
          4927 => x"09",
          4928 => x"ff",
          4929 => x"84",
          4930 => x"74",
          4931 => x"75",
          4932 => x"78",
          4933 => x"07",
          4934 => x"a4",
          4935 => x"52",
          4936 => x"b8",
          4937 => x"87",
          4938 => x"2e",
          4939 => x"e4",
          4940 => x"ff",
          4941 => x"81",
          4942 => x"e4",
          4943 => x"54",
          4944 => x"73",
          4945 => x"33",
          4946 => x"73",
          4947 => x"78",
          4948 => x"73",
          4949 => x"70",
          4950 => x"15",
          4951 => x"81",
          4952 => x"70",
          4953 => x"53",
          4954 => x"34",
          4955 => x"fc",
          4956 => x"e4",
          4957 => x"53",
          4958 => x"df",
          4959 => x"5b",
          4960 => x"5b",
          4961 => x"cc",
          4962 => x"2b",
          4963 => x"57",
          4964 => x"75",
          4965 => x"81",
          4966 => x"74",
          4967 => x"39",
          4968 => x"5a",
          4969 => x"fa",
          4970 => x"2a",
          4971 => x"85",
          4972 => x"0d",
          4973 => x"88",
          4974 => x"5e",
          4975 => x"59",
          4976 => x"38",
          4977 => x"9f",
          4978 => x"d0",
          4979 => x"85",
          4980 => x"80",
          4981 => x"10",
          4982 => x"5a",
          4983 => x"38",
          4984 => x"77",
          4985 => x"38",
          4986 => x"3f",
          4987 => x"70",
          4988 => x"86",
          4989 => x"5d",
          4990 => x"34",
          4991 => x"bb",
          4992 => x"ff",
          4993 => x"58",
          4994 => x"8d",
          4995 => x"8a",
          4996 => x"7a",
          4997 => x"0c",
          4998 => x"53",
          4999 => x"52",
          5000 => x"e4",
          5001 => x"81",
          5002 => x"78",
          5003 => x"b6",
          5004 => x"56",
          5005 => x"85",
          5006 => x"84",
          5007 => x"bf",
          5008 => x"cd",
          5009 => x"c5",
          5010 => x"18",
          5011 => x"7c",
          5012 => x"ad",
          5013 => x"18",
          5014 => x"75",
          5015 => x"33",
          5016 => x"88",
          5017 => x"07",
          5018 => x"5a",
          5019 => x"18",
          5020 => x"34",
          5021 => x"81",
          5022 => x"7c",
          5023 => x"ff",
          5024 => x"33",
          5025 => x"77",
          5026 => x"ff",
          5027 => x"38",
          5028 => x"33",
          5029 => x"88",
          5030 => x"5a",
          5031 => x"cc",
          5032 => x"88",
          5033 => x"80",
          5034 => x"33",
          5035 => x"81",
          5036 => x"75",
          5037 => x"42",
          5038 => x"c6",
          5039 => x"58",
          5040 => x"38",
          5041 => x"79",
          5042 => x"74",
          5043 => x"84",
          5044 => x"08",
          5045 => x"e4",
          5046 => x"83",
          5047 => x"26",
          5048 => x"26",
          5049 => x"70",
          5050 => x"7b",
          5051 => x"b0",
          5052 => x"8a",
          5053 => x"58",
          5054 => x"16",
          5055 => x"82",
          5056 => x"81",
          5057 => x"83",
          5058 => x"78",
          5059 => x"0b",
          5060 => x"0c",
          5061 => x"83",
          5062 => x"84",
          5063 => x"84",
          5064 => x"84",
          5065 => x"0b",
          5066 => x"b8",
          5067 => x"0b",
          5068 => x"04",
          5069 => x"06",
          5070 => x"38",
          5071 => x"05",
          5072 => x"38",
          5073 => x"40",
          5074 => x"70",
          5075 => x"05",
          5076 => x"56",
          5077 => x"70",
          5078 => x"17",
          5079 => x"17",
          5080 => x"30",
          5081 => x"2e",
          5082 => x"be",
          5083 => x"72",
          5084 => x"55",
          5085 => x"1c",
          5086 => x"ff",
          5087 => x"78",
          5088 => x"2a",
          5089 => x"c5",
          5090 => x"78",
          5091 => x"09",
          5092 => x"81",
          5093 => x"7b",
          5094 => x"38",
          5095 => x"93",
          5096 => x"fa",
          5097 => x"2e",
          5098 => x"80",
          5099 => x"2b",
          5100 => x"07",
          5101 => x"07",
          5102 => x"7a",
          5103 => x"90",
          5104 => x"be",
          5105 => x"30",
          5106 => x"3d",
          5107 => x"b6",
          5108 => x"78",
          5109 => x"80",
          5110 => x"ff",
          5111 => x"56",
          5112 => x"7a",
          5113 => x"51",
          5114 => x"08",
          5115 => x"56",
          5116 => x"bf",
          5117 => x"88",
          5118 => x"82",
          5119 => x"38",
          5120 => x"75",
          5121 => x"81",
          5122 => x"7a",
          5123 => x"75",
          5124 => x"77",
          5125 => x"b8",
          5126 => x"2e",
          5127 => x"81",
          5128 => x"2e",
          5129 => x"5a",
          5130 => x"f8",
          5131 => x"83",
          5132 => x"81",
          5133 => x"40",
          5134 => x"52",
          5135 => x"38",
          5136 => x"81",
          5137 => x"58",
          5138 => x"70",
          5139 => x"ff",
          5140 => x"2e",
          5141 => x"38",
          5142 => x"7c",
          5143 => x"0c",
          5144 => x"80",
          5145 => x"8a",
          5146 => x"ff",
          5147 => x"0c",
          5148 => x"ee",
          5149 => x"78",
          5150 => x"81",
          5151 => x"1b",
          5152 => x"83",
          5153 => x"85",
          5154 => x"5c",
          5155 => x"33",
          5156 => x"71",
          5157 => x"77",
          5158 => x"2e",
          5159 => x"83",
          5160 => x"c6",
          5161 => x"18",
          5162 => x"75",
          5163 => x"38",
          5164 => x"08",
          5165 => x"5b",
          5166 => x"9b",
          5167 => x"52",
          5168 => x"3f",
          5169 => x"38",
          5170 => x"0c",
          5171 => x"34",
          5172 => x"33",
          5173 => x"82",
          5174 => x"fc",
          5175 => x"12",
          5176 => x"07",
          5177 => x"2b",
          5178 => x"45",
          5179 => x"a4",
          5180 => x"38",
          5181 => x"12",
          5182 => x"07",
          5183 => x"2b",
          5184 => x"5b",
          5185 => x"e4",
          5186 => x"38",
          5187 => x"12",
          5188 => x"07",
          5189 => x"2b",
          5190 => x"5d",
          5191 => x"12",
          5192 => x"07",
          5193 => x"2b",
          5194 => x"0c",
          5195 => x"45",
          5196 => x"d0",
          5197 => x"d0",
          5198 => x"d0",
          5199 => x"98",
          5200 => x"24",
          5201 => x"56",
          5202 => x"08",
          5203 => x"33",
          5204 => x"b8",
          5205 => x"81",
          5206 => x"18",
          5207 => x"31",
          5208 => x"38",
          5209 => x"81",
          5210 => x"fd",
          5211 => x"f3",
          5212 => x"83",
          5213 => x"39",
          5214 => x"33",
          5215 => x"58",
          5216 => x"42",
          5217 => x"83",
          5218 => x"2b",
          5219 => x"70",
          5220 => x"07",
          5221 => x"5a",
          5222 => x"39",
          5223 => x"38",
          5224 => x"2e",
          5225 => x"5a",
          5226 => x"79",
          5227 => x"54",
          5228 => x"53",
          5229 => x"ad",
          5230 => x"0d",
          5231 => x"43",
          5232 => x"5a",
          5233 => x"78",
          5234 => x"26",
          5235 => x"38",
          5236 => x"d9",
          5237 => x"74",
          5238 => x"84",
          5239 => x"73",
          5240 => x"62",
          5241 => x"74",
          5242 => x"54",
          5243 => x"93",
          5244 => x"81",
          5245 => x"84",
          5246 => x"8b",
          5247 => x"0d",
          5248 => x"ff",
          5249 => x"91",
          5250 => x"d0",
          5251 => x"f7",
          5252 => x"5e",
          5253 => x"79",
          5254 => x"81",
          5255 => x"57",
          5256 => x"15",
          5257 => x"9f",
          5258 => x"e0",
          5259 => x"74",
          5260 => x"76",
          5261 => x"ff",
          5262 => x"70",
          5263 => x"57",
          5264 => x"1b",
          5265 => x"ff",
          5266 => x"7a",
          5267 => x"0c",
          5268 => x"6c",
          5269 => x"56",
          5270 => x"38",
          5271 => x"cc",
          5272 => x"58",
          5273 => x"57",
          5274 => x"38",
          5275 => x"b8",
          5276 => x"40",
          5277 => x"e1",
          5278 => x"84",
          5279 => x"38",
          5280 => x"81",
          5281 => x"38",
          5282 => x"88",
          5283 => x"83",
          5284 => x"81",
          5285 => x"12",
          5286 => x"33",
          5287 => x"2e",
          5288 => x"34",
          5289 => x"90",
          5290 => x"34",
          5291 => x"7e",
          5292 => x"34",
          5293 => x"5d",
          5294 => x"5b",
          5295 => x"9d",
          5296 => x"80",
          5297 => x"0b",
          5298 => x"e2",
          5299 => x"08",
          5300 => x"89",
          5301 => x"8a",
          5302 => x"a3",
          5303 => x"98",
          5304 => x"b8",
          5305 => x"7c",
          5306 => x"02",
          5307 => x"81",
          5308 => x"77",
          5309 => x"2e",
          5310 => x"81",
          5311 => x"56",
          5312 => x"c0",
          5313 => x"1b",
          5314 => x"11",
          5315 => x"07",
          5316 => x"7b",
          5317 => x"1a",
          5318 => x"12",
          5319 => x"07",
          5320 => x"2b",
          5321 => x"05",
          5322 => x"59",
          5323 => x"1a",
          5324 => x"91",
          5325 => x"77",
          5326 => x"2e",
          5327 => x"f1",
          5328 => x"22",
          5329 => x"76",
          5330 => x"5b",
          5331 => x"70",
          5332 => x"84",
          5333 => x"ac",
          5334 => x"84",
          5335 => x"82",
          5336 => x"80",
          5337 => x"39",
          5338 => x"5e",
          5339 => x"06",
          5340 => x"88",
          5341 => x"87",
          5342 => x"84",
          5343 => x"79",
          5344 => x"08",
          5345 => x"c8",
          5346 => x"31",
          5347 => x"33",
          5348 => x"90",
          5349 => x"fd",
          5350 => x"81",
          5351 => x"ab",
          5352 => x"84",
          5353 => x"38",
          5354 => x"d9",
          5355 => x"83",
          5356 => x"51",
          5357 => x"08",
          5358 => x"11",
          5359 => x"75",
          5360 => x"18",
          5361 => x"74",
          5362 => x"26",
          5363 => x"0b",
          5364 => x"34",
          5365 => x"17",
          5366 => x"07",
          5367 => x"8e",
          5368 => x"a1",
          5369 => x"91",
          5370 => x"17",
          5371 => x"9a",
          5372 => x"7d",
          5373 => x"06",
          5374 => x"7f",
          5375 => x"16",
          5376 => x"33",
          5377 => x"b5",
          5378 => x"52",
          5379 => x"3f",
          5380 => x"38",
          5381 => x"0c",
          5382 => x"0c",
          5383 => x"80",
          5384 => x"b4",
          5385 => x"81",
          5386 => x"3f",
          5387 => x"81",
          5388 => x"08",
          5389 => x"17",
          5390 => x"55",
          5391 => x"38",
          5392 => x"09",
          5393 => x"b4",
          5394 => x"79",
          5395 => x"b8",
          5396 => x"94",
          5397 => x"77",
          5398 => x"75",
          5399 => x"f8",
          5400 => x"08",
          5401 => x"27",
          5402 => x"71",
          5403 => x"74",
          5404 => x"2a",
          5405 => x"ed",
          5406 => x"f7",
          5407 => x"f7",
          5408 => x"80",
          5409 => x"57",
          5410 => x"62",
          5411 => x"80",
          5412 => x"9f",
          5413 => x"97",
          5414 => x"8f",
          5415 => x"59",
          5416 => x"80",
          5417 => x"8c",
          5418 => x"84",
          5419 => x"87",
          5420 => x"94",
          5421 => x"56",
          5422 => x"7b",
          5423 => x"75",
          5424 => x"38",
          5425 => x"2a",
          5426 => x"d3",
          5427 => x"27",
          5428 => x"f0",
          5429 => x"98",
          5430 => x"fe",
          5431 => x"e7",
          5432 => x"b0",
          5433 => x"2e",
          5434 => x"2a",
          5435 => x"38",
          5436 => x"38",
          5437 => x"53",
          5438 => x"9f",
          5439 => x"98",
          5440 => x"75",
          5441 => x"77",
          5442 => x"84",
          5443 => x"58",
          5444 => x"33",
          5445 => x"15",
          5446 => x"58",
          5447 => x"0c",
          5448 => x"59",
          5449 => x"af",
          5450 => x"0c",
          5451 => x"e4",
          5452 => x"fe",
          5453 => x"83",
          5454 => x"5b",
          5455 => x"76",
          5456 => x"38",
          5457 => x"41",
          5458 => x"80",
          5459 => x"19",
          5460 => x"b1",
          5461 => x"85",
          5462 => x"1a",
          5463 => x"1b",
          5464 => x"5a",
          5465 => x"2e",
          5466 => x"56",
          5467 => x"ff",
          5468 => x"38",
          5469 => x"70",
          5470 => x"75",
          5471 => x"b4",
          5472 => x"81",
          5473 => x"3f",
          5474 => x"2e",
          5475 => x"b8",
          5476 => x"08",
          5477 => x"08",
          5478 => x"fe",
          5479 => x"82",
          5480 => x"81",
          5481 => x"05",
          5482 => x"ff",
          5483 => x"39",
          5484 => x"56",
          5485 => x"79",
          5486 => x"e4",
          5487 => x"33",
          5488 => x"e4",
          5489 => x"38",
          5490 => x"39",
          5491 => x"84",
          5492 => x"82",
          5493 => x"b8",
          5494 => x"3d",
          5495 => x"5c",
          5496 => x"80",
          5497 => x"80",
          5498 => x"80",
          5499 => x"1b",
          5500 => x"fd",
          5501 => x"76",
          5502 => x"74",
          5503 => x"81",
          5504 => x"76",
          5505 => x"08",
          5506 => x"84",
          5507 => x"82",
          5508 => x"7e",
          5509 => x"ff",
          5510 => x"78",
          5511 => x"1a",
          5512 => x"38",
          5513 => x"ff",
          5514 => x"0c",
          5515 => x"1b",
          5516 => x"1b",
          5517 => x"08",
          5518 => x"58",
          5519 => x"8a",
          5520 => x"08",
          5521 => x"de",
          5522 => x"5c",
          5523 => x"19",
          5524 => x"79",
          5525 => x"52",
          5526 => x"3f",
          5527 => x"60",
          5528 => x"74",
          5529 => x"b8",
          5530 => x"56",
          5531 => x"70",
          5532 => x"75",
          5533 => x"34",
          5534 => x"7e",
          5535 => x"1c",
          5536 => x"8c",
          5537 => x"75",
          5538 => x"8c",
          5539 => x"1a",
          5540 => x"7a",
          5541 => x"b8",
          5542 => x"84",
          5543 => x"83",
          5544 => x"60",
          5545 => x"08",
          5546 => x"80",
          5547 => x"83",
          5548 => x"08",
          5549 => x"17",
          5550 => x"2e",
          5551 => x"54",
          5552 => x"33",
          5553 => x"e4",
          5554 => x"81",
          5555 => x"bf",
          5556 => x"06",
          5557 => x"56",
          5558 => x"70",
          5559 => x"05",
          5560 => x"38",
          5561 => x"fe",
          5562 => x"53",
          5563 => x"52",
          5564 => x"84",
          5565 => x"06",
          5566 => x"83",
          5567 => x"08",
          5568 => x"74",
          5569 => x"82",
          5570 => x"81",
          5571 => x"16",
          5572 => x"52",
          5573 => x"3f",
          5574 => x"08",
          5575 => x"38",
          5576 => x"38",
          5577 => x"08",
          5578 => x"58",
          5579 => x"79",
          5580 => x"e4",
          5581 => x"d8",
          5582 => x"39",
          5583 => x"3f",
          5584 => x"e4",
          5585 => x"54",
          5586 => x"53",
          5587 => x"b8",
          5588 => x"38",
          5589 => x"b4",
          5590 => x"77",
          5591 => x"82",
          5592 => x"81",
          5593 => x"16",
          5594 => x"52",
          5595 => x"3f",
          5596 => x"33",
          5597 => x"e4",
          5598 => x"38",
          5599 => x"39",
          5600 => x"16",
          5601 => x"ff",
          5602 => x"80",
          5603 => x"17",
          5604 => x"31",
          5605 => x"98",
          5606 => x"2e",
          5607 => x"54",
          5608 => x"53",
          5609 => x"96",
          5610 => x"94",
          5611 => x"81",
          5612 => x"b8",
          5613 => x"0b",
          5614 => x"e4",
          5615 => x"0d",
          5616 => x"9f",
          5617 => x"97",
          5618 => x"8f",
          5619 => x"58",
          5620 => x"80",
          5621 => x"d8",
          5622 => x"81",
          5623 => x"c8",
          5624 => x"b4",
          5625 => x"17",
          5626 => x"54",
          5627 => x"33",
          5628 => x"e4",
          5629 => x"81",
          5630 => x"90",
          5631 => x"a0",
          5632 => x"77",
          5633 => x"ff",
          5634 => x"34",
          5635 => x"34",
          5636 => x"56",
          5637 => x"8c",
          5638 => x"88",
          5639 => x"90",
          5640 => x"98",
          5641 => x"7a",
          5642 => x"0b",
          5643 => x"18",
          5644 => x"0b",
          5645 => x"83",
          5646 => x"3f",
          5647 => x"81",
          5648 => x"34",
          5649 => x"0d",
          5650 => x"b8",
          5651 => x"5b",
          5652 => x"b8",
          5653 => x"e4",
          5654 => x"a8",
          5655 => x"57",
          5656 => x"8e",
          5657 => x"2e",
          5658 => x"54",
          5659 => x"53",
          5660 => x"92",
          5661 => x"78",
          5662 => x"74",
          5663 => x"8c",
          5664 => x"88",
          5665 => x"90",
          5666 => x"98",
          5667 => x"7a",
          5668 => x"0b",
          5669 => x"18",
          5670 => x"0b",
          5671 => x"83",
          5672 => x"3f",
          5673 => x"81",
          5674 => x"34",
          5675 => x"ff",
          5676 => x"81",
          5677 => x"78",
          5678 => x"3d",
          5679 => x"3f",
          5680 => x"e4",
          5681 => x"2e",
          5682 => x"2e",
          5683 => x"2e",
          5684 => x"22",
          5685 => x"80",
          5686 => x"38",
          5687 => x"0c",
          5688 => x"51",
          5689 => x"08",
          5690 => x"75",
          5691 => x"0d",
          5692 => x"80",
          5693 => x"57",
          5694 => x"ba",
          5695 => x"ba",
          5696 => x"51",
          5697 => x"d0",
          5698 => x"0c",
          5699 => x"b8",
          5700 => x"33",
          5701 => x"53",
          5702 => x"19",
          5703 => x"54",
          5704 => x"0b",
          5705 => x"79",
          5706 => x"33",
          5707 => x"9f",
          5708 => x"89",
          5709 => x"53",
          5710 => x"26",
          5711 => x"06",
          5712 => x"55",
          5713 => x"85",
          5714 => x"32",
          5715 => x"76",
          5716 => x"92",
          5717 => x"83",
          5718 => x"fe",
          5719 => x"77",
          5720 => x"3d",
          5721 => x"52",
          5722 => x"b8",
          5723 => x"80",
          5724 => x"0c",
          5725 => x"52",
          5726 => x"3f",
          5727 => x"e4",
          5728 => x"05",
          5729 => x"77",
          5730 => x"33",
          5731 => x"75",
          5732 => x"11",
          5733 => x"07",
          5734 => x"79",
          5735 => x"0c",
          5736 => x"0d",
          5737 => x"09",
          5738 => x"84",
          5739 => x"95",
          5740 => x"2b",
          5741 => x"1b",
          5742 => x"98",
          5743 => x"0c",
          5744 => x"0d",
          5745 => x"08",
          5746 => x"80",
          5747 => x"e5",
          5748 => x"e4",
          5749 => x"c8",
          5750 => x"61",
          5751 => x"58",
          5752 => x"80",
          5753 => x"98",
          5754 => x"ff",
          5755 => x"59",
          5756 => x"60",
          5757 => x"16",
          5758 => x"e4",
          5759 => x"83",
          5760 => x"16",
          5761 => x"c9",
          5762 => x"85",
          5763 => x"17",
          5764 => x"3d",
          5765 => x"71",
          5766 => x"40",
          5767 => x"da",
          5768 => x"52",
          5769 => x"b8",
          5770 => x"82",
          5771 => x"a8",
          5772 => x"84",
          5773 => x"3d",
          5774 => x"71",
          5775 => x"58",
          5776 => x"fd",
          5777 => x"b8",
          5778 => x"e2",
          5779 => x"b8",
          5780 => x"78",
          5781 => x"c8",
          5782 => x"52",
          5783 => x"7f",
          5784 => x"2e",
          5785 => x"81",
          5786 => x"f5",
          5787 => x"81",
          5788 => x"7e",
          5789 => x"e6",
          5790 => x"59",
          5791 => x"76",
          5792 => x"08",
          5793 => x"da",
          5794 => x"77",
          5795 => x"84",
          5796 => x"e4",
          5797 => x"59",
          5798 => x"38",
          5799 => x"5f",
          5800 => x"7a",
          5801 => x"7a",
          5802 => x"33",
          5803 => x"17",
          5804 => x"7c",
          5805 => x"2e",
          5806 => x"59",
          5807 => x"0c",
          5808 => x"33",
          5809 => x"90",
          5810 => x"fd",
          5811 => x"33",
          5812 => x"79",
          5813 => x"80",
          5814 => x"84",
          5815 => x"08",
          5816 => x"39",
          5817 => x"16",
          5818 => x"ff",
          5819 => x"e4",
          5820 => x"08",
          5821 => x"17",
          5822 => x"55",
          5823 => x"38",
          5824 => x"09",
          5825 => x"b4",
          5826 => x"7d",
          5827 => x"b8",
          5828 => x"18",
          5829 => x"af",
          5830 => x"33",
          5831 => x"70",
          5832 => x"5a",
          5833 => x"e8",
          5834 => x"08",
          5835 => x"7c",
          5836 => x"27",
          5837 => x"18",
          5838 => x"70",
          5839 => x"d4",
          5840 => x"7c",
          5841 => x"e4",
          5842 => x"7d",
          5843 => x"9f",
          5844 => x"97",
          5845 => x"8f",
          5846 => x"59",
          5847 => x"80",
          5848 => x"c2",
          5849 => x"ba",
          5850 => x"26",
          5851 => x"80",
          5852 => x"79",
          5853 => x"5a",
          5854 => x"75",
          5855 => x"3f",
          5856 => x"54",
          5857 => x"3f",
          5858 => x"d5",
          5859 => x"17",
          5860 => x"56",
          5861 => x"38",
          5862 => x"76",
          5863 => x"0c",
          5864 => x"06",
          5865 => x"fe",
          5866 => x"f3",
          5867 => x"b8",
          5868 => x"73",
          5869 => x"82",
          5870 => x"08",
          5871 => x"0c",
          5872 => x"34",
          5873 => x"8b",
          5874 => x"81",
          5875 => x"bb",
          5876 => x"80",
          5877 => x"fe",
          5878 => x"15",
          5879 => x"73",
          5880 => x"c0",
          5881 => x"83",
          5882 => x"38",
          5883 => x"77",
          5884 => x"e4",
          5885 => x"94",
          5886 => x"80",
          5887 => x"0c",
          5888 => x"a8",
          5889 => x"15",
          5890 => x"ff",
          5891 => x"79",
          5892 => x"5a",
          5893 => x"38",
          5894 => x"18",
          5895 => x"5a",
          5896 => x"8c",
          5897 => x"52",
          5898 => x"b8",
          5899 => x"14",
          5900 => x"b8",
          5901 => x"cf",
          5902 => x"c9",
          5903 => x"cb",
          5904 => x"b8",
          5905 => x"b8",
          5906 => x"84",
          5907 => x"98",
          5908 => x"91",
          5909 => x"0c",
          5910 => x"7c",
          5911 => x"38",
          5912 => x"8d",
          5913 => x"84",
          5914 => x"08",
          5915 => x"74",
          5916 => x"3d",
          5917 => x"75",
          5918 => x"e4",
          5919 => x"d1",
          5920 => x"59",
          5921 => x"16",
          5922 => x"54",
          5923 => x"16",
          5924 => x"71",
          5925 => x"5d",
          5926 => x"38",
          5927 => x"18",
          5928 => x"51",
          5929 => x"08",
          5930 => x"80",
          5931 => x"fe",
          5932 => x"fe",
          5933 => x"33",
          5934 => x"7a",
          5935 => x"bc",
          5936 => x"54",
          5937 => x"53",
          5938 => x"52",
          5939 => x"22",
          5940 => x"2e",
          5941 => x"84",
          5942 => x"e4",
          5943 => x"33",
          5944 => x"e4",
          5945 => x"71",
          5946 => x"3d",
          5947 => x"74",
          5948 => x"73",
          5949 => x"72",
          5950 => x"84",
          5951 => x"81",
          5952 => x"53",
          5953 => x"80",
          5954 => x"9d",
          5955 => x"84",
          5956 => x"84",
          5957 => x"74",
          5958 => x"74",
          5959 => x"e4",
          5960 => x"07",
          5961 => x"55",
          5962 => x"8a",
          5963 => x"52",
          5964 => x"74",
          5965 => x"e4",
          5966 => x"07",
          5967 => x"55",
          5968 => x"51",
          5969 => x"08",
          5970 => x"04",
          5971 => x"3f",
          5972 => x"72",
          5973 => x"56",
          5974 => x"57",
          5975 => x"3d",
          5976 => x"e4",
          5977 => x"2e",
          5978 => x"95",
          5979 => x"ff",
          5980 => x"55",
          5981 => x"80",
          5982 => x"58",
          5983 => x"2e",
          5984 => x"b0",
          5985 => x"95",
          5986 => x"e4",
          5987 => x"0d",
          5988 => x"3d",
          5989 => x"b9",
          5990 => x"b8",
          5991 => x"74",
          5992 => x"13",
          5993 => x"26",
          5994 => x"b8",
          5995 => x"b8",
          5996 => x"81",
          5997 => x"08",
          5998 => x"77",
          5999 => x"5c",
          6000 => x"82",
          6001 => x"5d",
          6002 => x"53",
          6003 => x"fe",
          6004 => x"80",
          6005 => x"79",
          6006 => x"7d",
          6007 => x"82",
          6008 => x"05",
          6009 => x"90",
          6010 => x"33",
          6011 => x"71",
          6012 => x"70",
          6013 => x"84",
          6014 => x"43",
          6015 => x"40",
          6016 => x"7f",
          6017 => x"33",
          6018 => x"79",
          6019 => x"04",
          6020 => x"17",
          6021 => x"fe",
          6022 => x"e4",
          6023 => x"08",
          6024 => x"18",
          6025 => x"55",
          6026 => x"38",
          6027 => x"09",
          6028 => x"b4",
          6029 => x"7c",
          6030 => x"e0",
          6031 => x"77",
          6032 => x"77",
          6033 => x"e4",
          6034 => x"b8",
          6035 => x"84",
          6036 => x"e4",
          6037 => x"18",
          6038 => x"08",
          6039 => x"7a",
          6040 => x"07",
          6041 => x"39",
          6042 => x"71",
          6043 => x"70",
          6044 => x"06",
          6045 => x"5f",
          6046 => x"39",
          6047 => x"58",
          6048 => x"0c",
          6049 => x"84",
          6050 => x"58",
          6051 => x"57",
          6052 => x"76",
          6053 => x"74",
          6054 => x"86",
          6055 => x"78",
          6056 => x"73",
          6057 => x"33",
          6058 => x"33",
          6059 => x"87",
          6060 => x"94",
          6061 => x"27",
          6062 => x"17",
          6063 => x"27",
          6064 => x"b3",
          6065 => x"0c",
          6066 => x"80",
          6067 => x"75",
          6068 => x"34",
          6069 => x"8b",
          6070 => x"27",
          6071 => x"fe",
          6072 => x"59",
          6073 => x"e9",
          6074 => x"82",
          6075 => x"2e",
          6076 => x"75",
          6077 => x"e4",
          6078 => x"fe",
          6079 => x"74",
          6080 => x"94",
          6081 => x"54",
          6082 => x"79",
          6083 => x"15",
          6084 => x"b8",
          6085 => x"95",
          6086 => x"8f",
          6087 => x"54",
          6088 => x"fe",
          6089 => x"51",
          6090 => x"08",
          6091 => x"e4",
          6092 => x"81",
          6093 => x"08",
          6094 => x"84",
          6095 => x"08",
          6096 => x"e4",
          6097 => x"e4",
          6098 => x"38",
          6099 => x"74",
          6100 => x"84",
          6101 => x"08",
          6102 => x"fe",
          6103 => x"59",
          6104 => x"cb",
          6105 => x"80",
          6106 => x"2e",
          6107 => x"75",
          6108 => x"e4",
          6109 => x"fe",
          6110 => x"74",
          6111 => x"17",
          6112 => x"73",
          6113 => x"26",
          6114 => x"90",
          6115 => x"56",
          6116 => x"33",
          6117 => x"e7",
          6118 => x"54",
          6119 => x"90",
          6120 => x"81",
          6121 => x"f0",
          6122 => x"39",
          6123 => x"0d",
          6124 => x"52",
          6125 => x"84",
          6126 => x"08",
          6127 => x"e4",
          6128 => x"a8",
          6129 => x"59",
          6130 => x"08",
          6131 => x"02",
          6132 => x"81",
          6133 => x"38",
          6134 => x"c4",
          6135 => x"81",
          6136 => x"b4",
          6137 => x"33",
          6138 => x"73",
          6139 => x"83",
          6140 => x"81",
          6141 => x"38",
          6142 => x"ff",
          6143 => x"b8",
          6144 => x"55",
          6145 => x"08",
          6146 => x"38",
          6147 => x"ff",
          6148 => x"56",
          6149 => x"0b",
          6150 => x"04",
          6151 => x"98",
          6152 => x"5d",
          6153 => x"e4",
          6154 => x"e4",
          6155 => x"a8",
          6156 => x"2e",
          6157 => x"ff",
          6158 => x"56",
          6159 => x"38",
          6160 => x"56",
          6161 => x"80",
          6162 => x"55",
          6163 => x"08",
          6164 => x"75",
          6165 => x"db",
          6166 => x"e4",
          6167 => x"5d",
          6168 => x"17",
          6169 => x"17",
          6170 => x"09",
          6171 => x"75",
          6172 => x"51",
          6173 => x"08",
          6174 => x"58",
          6175 => x"ab",
          6176 => x"34",
          6177 => x"08",
          6178 => x"78",
          6179 => x"e4",
          6180 => x"2e",
          6181 => x"81",
          6182 => x"c8",
          6183 => x"7c",
          6184 => x"90",
          6185 => x"7a",
          6186 => x"84",
          6187 => x"17",
          6188 => x"e4",
          6189 => x"27",
          6190 => x"74",
          6191 => x"38",
          6192 => x"08",
          6193 => x"51",
          6194 => x"c5",
          6195 => x"e1",
          6196 => x"e4",
          6197 => x"b8",
          6198 => x"84",
          6199 => x"38",
          6200 => x"cb",
          6201 => x"fe",
          6202 => x"b3",
          6203 => x"19",
          6204 => x"ff",
          6205 => x"84",
          6206 => x"18",
          6207 => x"a1",
          6208 => x"56",
          6209 => x"56",
          6210 => x"39",
          6211 => x"ff",
          6212 => x"b2",
          6213 => x"84",
          6214 => x"75",
          6215 => x"04",
          6216 => x"52",
          6217 => x"e4",
          6218 => x"38",
          6219 => x"3d",
          6220 => x"2e",
          6221 => x"f3",
          6222 => x"56",
          6223 => x"7d",
          6224 => x"5d",
          6225 => x"08",
          6226 => x"83",
          6227 => x"81",
          6228 => x"08",
          6229 => x"c9",
          6230 => x"12",
          6231 => x"38",
          6232 => x"5a",
          6233 => x"38",
          6234 => x"19",
          6235 => x"0c",
          6236 => x"55",
          6237 => x"ff",
          6238 => x"8a",
          6239 => x"f9",
          6240 => x"52",
          6241 => x"3f",
          6242 => x"81",
          6243 => x"84",
          6244 => x"b8",
          6245 => x"58",
          6246 => x"b8",
          6247 => x"08",
          6248 => x"18",
          6249 => x"27",
          6250 => x"7a",
          6251 => x"38",
          6252 => x"08",
          6253 => x"51",
          6254 => x"81",
          6255 => x"7c",
          6256 => x"08",
          6257 => x"51",
          6258 => x"08",
          6259 => x"fd",
          6260 => x"2e",
          6261 => x"ff",
          6262 => x"52",
          6263 => x"b8",
          6264 => x"08",
          6265 => x"59",
          6266 => x"94",
          6267 => x"5c",
          6268 => x"7a",
          6269 => x"e4",
          6270 => x"22",
          6271 => x"81",
          6272 => x"fe",
          6273 => x"56",
          6274 => x"ff",
          6275 => x"ae",
          6276 => x"0b",
          6277 => x"80",
          6278 => x"34",
          6279 => x"cc",
          6280 => x"83",
          6281 => x"d2",
          6282 => x"80",
          6283 => x"83",
          6284 => x"0b",
          6285 => x"56",
          6286 => x"70",
          6287 => x"75",
          6288 => x"d9",
          6289 => x"ff",
          6290 => x"17",
          6291 => x"f3",
          6292 => x"2e",
          6293 => x"83",
          6294 => x"3f",
          6295 => x"e4",
          6296 => x"b8",
          6297 => x"e4",
          6298 => x"17",
          6299 => x"7d",
          6300 => x"77",
          6301 => x"7c",
          6302 => x"38",
          6303 => x"7d",
          6304 => x"51",
          6305 => x"08",
          6306 => x"3d",
          6307 => x"80",
          6308 => x"76",
          6309 => x"7b",
          6310 => x"34",
          6311 => x"17",
          6312 => x"1a",
          6313 => x"39",
          6314 => x"34",
          6315 => x"34",
          6316 => x"7d",
          6317 => x"51",
          6318 => x"08",
          6319 => x"b3",
          6320 => x"5f",
          6321 => x"81",
          6322 => x"56",
          6323 => x"ed",
          6324 => x"82",
          6325 => x"b2",
          6326 => x"b8",
          6327 => x"80",
          6328 => x"0c",
          6329 => x"0c",
          6330 => x"52",
          6331 => x"e4",
          6332 => x"38",
          6333 => x"06",
          6334 => x"0b",
          6335 => x"55",
          6336 => x"70",
          6337 => x"74",
          6338 => x"7a",
          6339 => x"57",
          6340 => x"ff",
          6341 => x"08",
          6342 => x"84",
          6343 => x"08",
          6344 => x"2e",
          6345 => x"e4",
          6346 => x"d0",
          6347 => x"58",
          6348 => x"78",
          6349 => x"78",
          6350 => x"08",
          6351 => x"5e",
          6352 => x"5c",
          6353 => x"ff",
          6354 => x"26",
          6355 => x"06",
          6356 => x"99",
          6357 => x"ff",
          6358 => x"2a",
          6359 => x"06",
          6360 => x"7a",
          6361 => x"2a",
          6362 => x"2e",
          6363 => x"5c",
          6364 => x"08",
          6365 => x"83",
          6366 => x"82",
          6367 => x"b2",
          6368 => x"b8",
          6369 => x"fd",
          6370 => x"3d",
          6371 => x"38",
          6372 => x"b8",
          6373 => x"fd",
          6374 => x"19",
          6375 => x"56",
          6376 => x"75",
          6377 => x"5a",
          6378 => x"33",
          6379 => x"84",
          6380 => x"38",
          6381 => x"34",
          6382 => x"8b",
          6383 => x"57",
          6384 => x"a7",
          6385 => x"7f",
          6386 => x"88",
          6387 => x"57",
          6388 => x"16",
          6389 => x"75",
          6390 => x"22",
          6391 => x"57",
          6392 => x"75",
          6393 => x"2e",
          6394 => x"83",
          6395 => x"17",
          6396 => x"f1",
          6397 => x"85",
          6398 => x"18",
          6399 => x"56",
          6400 => x"33",
          6401 => x"bb",
          6402 => x"5d",
          6403 => x"88",
          6404 => x"76",
          6405 => x"06",
          6406 => x"80",
          6407 => x"75",
          6408 => x"0b",
          6409 => x"08",
          6410 => x"ff",
          6411 => x"fe",
          6412 => x"55",
          6413 => x"b8",
          6414 => x"5a",
          6415 => x"83",
          6416 => x"2e",
          6417 => x"54",
          6418 => x"33",
          6419 => x"e4",
          6420 => x"81",
          6421 => x"77",
          6422 => x"7a",
          6423 => x"19",
          6424 => x"78",
          6425 => x"e4",
          6426 => x"2e",
          6427 => x"2e",
          6428 => x"db",
          6429 => x"84",
          6430 => x"b1",
          6431 => x"e4",
          6432 => x"33",
          6433 => x"90",
          6434 => x"fd",
          6435 => x"2e",
          6436 => x"80",
          6437 => x"e4",
          6438 => x"b4",
          6439 => x"33",
          6440 => x"84",
          6441 => x"06",
          6442 => x"83",
          6443 => x"08",
          6444 => x"74",
          6445 => x"82",
          6446 => x"81",
          6447 => x"16",
          6448 => x"52",
          6449 => x"3f",
          6450 => x"b4",
          6451 => x"81",
          6452 => x"3f",
          6453 => x"c9",
          6454 => x"34",
          6455 => x"84",
          6456 => x"18",
          6457 => x"33",
          6458 => x"fc",
          6459 => x"a0",
          6460 => x"17",
          6461 => x"5c",
          6462 => x"80",
          6463 => x"e3",
          6464 => x"3d",
          6465 => x"a2",
          6466 => x"84",
          6467 => x"75",
          6468 => x"04",
          6469 => x"05",
          6470 => x"e4",
          6471 => x"38",
          6472 => x"06",
          6473 => x"a7",
          6474 => x"71",
          6475 => x"57",
          6476 => x"81",
          6477 => x"e2",
          6478 => x"b8",
          6479 => x"3d",
          6480 => x"cc",
          6481 => x"d9",
          6482 => x"b8",
          6483 => x"84",
          6484 => x"78",
          6485 => x"51",
          6486 => x"08",
          6487 => x"02",
          6488 => x"56",
          6489 => x"18",
          6490 => x"07",
          6491 => x"76",
          6492 => x"76",
          6493 => x"76",
          6494 => x"78",
          6495 => x"51",
          6496 => x"08",
          6497 => x"04",
          6498 => x"80",
          6499 => x"3d",
          6500 => x"e4",
          6501 => x"84",
          6502 => x"56",
          6503 => x"70",
          6504 => x"38",
          6505 => x"56",
          6506 => x"81",
          6507 => x"2e",
          6508 => x"58",
          6509 => x"2e",
          6510 => x"5a",
          6511 => x"81",
          6512 => x"16",
          6513 => x"c9",
          6514 => x"85",
          6515 => x"17",
          6516 => x"70",
          6517 => x"83",
          6518 => x"84",
          6519 => x"b8",
          6520 => x"71",
          6521 => x"14",
          6522 => x"33",
          6523 => x"57",
          6524 => x"9a",
          6525 => x"80",
          6526 => x"f4",
          6527 => x"84",
          6528 => x"38",
          6529 => x"b8",
          6530 => x"b0",
          6531 => x"b8",
          6532 => x"5b",
          6533 => x"b8",
          6534 => x"fe",
          6535 => x"17",
          6536 => x"31",
          6537 => x"a0",
          6538 => x"16",
          6539 => x"06",
          6540 => x"08",
          6541 => x"81",
          6542 => x"79",
          6543 => x"52",
          6544 => x"3f",
          6545 => x"8d",
          6546 => x"51",
          6547 => x"08",
          6548 => x"38",
          6549 => x"08",
          6550 => x"19",
          6551 => x"75",
          6552 => x"ec",
          6553 => x"76",
          6554 => x"ff",
          6555 => x"58",
          6556 => x"39",
          6557 => x"0d",
          6558 => x"52",
          6559 => x"84",
          6560 => x"08",
          6561 => x"7d",
          6562 => x"58",
          6563 => x"74",
          6564 => x"ff",
          6565 => x"27",
          6566 => x"5c",
          6567 => x"57",
          6568 => x"0c",
          6569 => x"38",
          6570 => x"52",
          6571 => x"3f",
          6572 => x"06",
          6573 => x"83",
          6574 => x"70",
          6575 => x"80",
          6576 => x"77",
          6577 => x"70",
          6578 => x"80",
          6579 => x"81",
          6580 => x"59",
          6581 => x"27",
          6582 => x"96",
          6583 => x"76",
          6584 => x"05",
          6585 => x"70",
          6586 => x"3d",
          6587 => x"5b",
          6588 => x"d1",
          6589 => x"76",
          6590 => x"2e",
          6591 => x"16",
          6592 => x"09",
          6593 => x"79",
          6594 => x"52",
          6595 => x"e4",
          6596 => x"b8",
          6597 => x"56",
          6598 => x"0d",
          6599 => x"e7",
          6600 => x"ff",
          6601 => x"56",
          6602 => x"0d",
          6603 => x"c3",
          6604 => x"ee",
          6605 => x"b8",
          6606 => x"2e",
          6607 => x"57",
          6608 => x"76",
          6609 => x"55",
          6610 => x"83",
          6611 => x"3f",
          6612 => x"ff",
          6613 => x"38",
          6614 => x"e4",
          6615 => x"ee",
          6616 => x"e6",
          6617 => x"58",
          6618 => x"08",
          6619 => x"09",
          6620 => x"e4",
          6621 => x"08",
          6622 => x"2e",
          6623 => x"79",
          6624 => x"81",
          6625 => x"18",
          6626 => x"b8",
          6627 => x"57",
          6628 => x"57",
          6629 => x"70",
          6630 => x"2e",
          6631 => x"25",
          6632 => x"81",
          6633 => x"2e",
          6634 => x"ef",
          6635 => x"84",
          6636 => x"38",
          6637 => x"38",
          6638 => x"6c",
          6639 => x"58",
          6640 => x"6b",
          6641 => x"6c",
          6642 => x"05",
          6643 => x"34",
          6644 => x"eb",
          6645 => x"76",
          6646 => x"55",
          6647 => x"5a",
          6648 => x"83",
          6649 => x"3f",
          6650 => x"39",
          6651 => x"b4",
          6652 => x"33",
          6653 => x"e4",
          6654 => x"c3",
          6655 => x"34",
          6656 => x"5c",
          6657 => x"82",
          6658 => x"38",
          6659 => x"39",
          6660 => x"ed",
          6661 => x"84",
          6662 => x"38",
          6663 => x"78",
          6664 => x"39",
          6665 => x"08",
          6666 => x"51",
          6667 => x"f2",
          6668 => x"80",
          6669 => x"56",
          6670 => x"55",
          6671 => x"54",
          6672 => x"22",
          6673 => x"2e",
          6674 => x"75",
          6675 => x"75",
          6676 => x"a2",
          6677 => x"90",
          6678 => x"56",
          6679 => x"7e",
          6680 => x"55",
          6681 => x"dc",
          6682 => x"70",
          6683 => x"08",
          6684 => x"5f",
          6685 => x"9c",
          6686 => x"58",
          6687 => x"52",
          6688 => x"15",
          6689 => x"26",
          6690 => x"08",
          6691 => x"e4",
          6692 => x"b8",
          6693 => x"59",
          6694 => x"2e",
          6695 => x"75",
          6696 => x"3d",
          6697 => x"0c",
          6698 => x"51",
          6699 => x"08",
          6700 => x"73",
          6701 => x"7b",
          6702 => x"56",
          6703 => x"18",
          6704 => x"73",
          6705 => x"dd",
          6706 => x"b8",
          6707 => x"19",
          6708 => x"38",
          6709 => x"80",
          6710 => x"0c",
          6711 => x"80",
          6712 => x"9c",
          6713 => x"58",
          6714 => x"76",
          6715 => x"33",
          6716 => x"75",
          6717 => x"97",
          6718 => x"39",
          6719 => x"fe",
          6720 => x"39",
          6721 => x"a3",
          6722 => x"05",
          6723 => x"ff",
          6724 => x"40",
          6725 => x"70",
          6726 => x"56",
          6727 => x"74",
          6728 => x"38",
          6729 => x"24",
          6730 => x"d0",
          6731 => x"80",
          6732 => x"16",
          6733 => x"d9",
          6734 => x"79",
          6735 => x"e4",
          6736 => x"5d",
          6737 => x"75",
          6738 => x"7f",
          6739 => x"53",
          6740 => x"3f",
          6741 => x"6d",
          6742 => x"74",
          6743 => x"ff",
          6744 => x"38",
          6745 => x"7f",
          6746 => x"0a",
          6747 => x"06",
          6748 => x"2a",
          6749 => x"2b",
          6750 => x"2e",
          6751 => x"25",
          6752 => x"83",
          6753 => x"38",
          6754 => x"51",
          6755 => x"b8",
          6756 => x"ff",
          6757 => x"71",
          6758 => x"77",
          6759 => x"82",
          6760 => x"83",
          6761 => x"2e",
          6762 => x"11",
          6763 => x"71",
          6764 => x"72",
          6765 => x"83",
          6766 => x"33",
          6767 => x"81",
          6768 => x"75",
          6769 => x"42",
          6770 => x"4e",
          6771 => x"78",
          6772 => x"82",
          6773 => x"26",
          6774 => x"81",
          6775 => x"f9",
          6776 => x"2e",
          6777 => x"83",
          6778 => x"46",
          6779 => x"c2",
          6780 => x"57",
          6781 => x"58",
          6782 => x"26",
          6783 => x"10",
          6784 => x"74",
          6785 => x"ee",
          6786 => x"94",
          6787 => x"05",
          6788 => x"26",
          6789 => x"08",
          6790 => x"11",
          6791 => x"83",
          6792 => x"a0",
          6793 => x"66",
          6794 => x"31",
          6795 => x"89",
          6796 => x"29",
          6797 => x"79",
          6798 => x"7d",
          6799 => x"56",
          6800 => x"08",
          6801 => x"62",
          6802 => x"38",
          6803 => x"08",
          6804 => x"38",
          6805 => x"89",
          6806 => x"8b",
          6807 => x"3d",
          6808 => x"4e",
          6809 => x"e4",
          6810 => x"0c",
          6811 => x"ff",
          6812 => x"91",
          6813 => x"d0",
          6814 => x"b2",
          6815 => x"5c",
          6816 => x"81",
          6817 => x"58",
          6818 => x"62",
          6819 => x"81",
          6820 => x"45",
          6821 => x"70",
          6822 => x"70",
          6823 => x"09",
          6824 => x"38",
          6825 => x"07",
          6826 => x"7a",
          6827 => x"84",
          6828 => x"98",
          6829 => x"3d",
          6830 => x"fe",
          6831 => x"e4",
          6832 => x"77",
          6833 => x"75",
          6834 => x"57",
          6835 => x"7f",
          6836 => x"fa",
          6837 => x"38",
          6838 => x"95",
          6839 => x"67",
          6840 => x"70",
          6841 => x"84",
          6842 => x"38",
          6843 => x"80",
          6844 => x"76",
          6845 => x"84",
          6846 => x"81",
          6847 => x"27",
          6848 => x"57",
          6849 => x"57",
          6850 => x"34",
          6851 => x"61",
          6852 => x"70",
          6853 => x"05",
          6854 => x"38",
          6855 => x"82",
          6856 => x"05",
          6857 => x"6a",
          6858 => x"5c",
          6859 => x"90",
          6860 => x"5a",
          6861 => x"9e",
          6862 => x"05",
          6863 => x"26",
          6864 => x"06",
          6865 => x"88",
          6866 => x"f8",
          6867 => x"05",
          6868 => x"61",
          6869 => x"34",
          6870 => x"2a",
          6871 => x"90",
          6872 => x"7e",
          6873 => x"b8",
          6874 => x"83",
          6875 => x"05",
          6876 => x"61",
          6877 => x"05",
          6878 => x"74",
          6879 => x"4b",
          6880 => x"61",
          6881 => x"34",
          6882 => x"59",
          6883 => x"33",
          6884 => x"15",
          6885 => x"05",
          6886 => x"ff",
          6887 => x"54",
          6888 => x"c6",
          6889 => x"08",
          6890 => x"83",
          6891 => x"55",
          6892 => x"ff",
          6893 => x"41",
          6894 => x"87",
          6895 => x"83",
          6896 => x"88",
          6897 => x"81",
          6898 => x"78",
          6899 => x"98",
          6900 => x"65",
          6901 => x"59",
          6902 => x"51",
          6903 => x"08",
          6904 => x"55",
          6905 => x"ff",
          6906 => x"77",
          6907 => x"7f",
          6908 => x"89",
          6909 => x"38",
          6910 => x"83",
          6911 => x"60",
          6912 => x"84",
          6913 => x"1b",
          6914 => x"38",
          6915 => x"86",
          6916 => x"38",
          6917 => x"81",
          6918 => x"2a",
          6919 => x"84",
          6920 => x"81",
          6921 => x"f4",
          6922 => x"6b",
          6923 => x"67",
          6924 => x"67",
          6925 => x"34",
          6926 => x"80",
          6927 => x"f8",
          6928 => x"84",
          6929 => x"57",
          6930 => x"e4",
          6931 => x"83",
          6932 => x"05",
          6933 => x"84",
          6934 => x"34",
          6935 => x"88",
          6936 => x"34",
          6937 => x"cc",
          6938 => x"61",
          6939 => x"53",
          6940 => x"3f",
          6941 => x"c9",
          6942 => x"fe",
          6943 => x"e4",
          6944 => x"08",
          6945 => x"84",
          6946 => x"e4",
          6947 => x"f6",
          6948 => x"2a",
          6949 => x"56",
          6950 => x"77",
          6951 => x"77",
          6952 => x"58",
          6953 => x"27",
          6954 => x"f6",
          6955 => x"10",
          6956 => x"5c",
          6957 => x"08",
          6958 => x"ff",
          6959 => x"8e",
          6960 => x"08",
          6961 => x"7a",
          6962 => x"7a",
          6963 => x"39",
          6964 => x"f8",
          6965 => x"75",
          6966 => x"49",
          6967 => x"2a",
          6968 => x"98",
          6969 => x"f9",
          6970 => x"34",
          6971 => x"61",
          6972 => x"80",
          6973 => x"34",
          6974 => x"05",
          6975 => x"a6",
          6976 => x"61",
          6977 => x"34",
          6978 => x"ae",
          6979 => x"81",
          6980 => x"05",
          6981 => x"61",
          6982 => x"c0",
          6983 => x"34",
          6984 => x"c0",
          6985 => x"58",
          6986 => x"ff",
          6987 => x"38",
          6988 => x"70",
          6989 => x"74",
          6990 => x"80",
          6991 => x"d9",
          6992 => x"f4",
          6993 => x"42",
          6994 => x"54",
          6995 => x"79",
          6996 => x"39",
          6997 => x"3d",
          6998 => x"61",
          6999 => x"05",
          7000 => x"4c",
          7001 => x"05",
          7002 => x"61",
          7003 => x"34",
          7004 => x"89",
          7005 => x"8f",
          7006 => x"76",
          7007 => x"51",
          7008 => x"56",
          7009 => x"34",
          7010 => x"5c",
          7011 => x"34",
          7012 => x"05",
          7013 => x"05",
          7014 => x"f2",
          7015 => x"61",
          7016 => x"83",
          7017 => x"e7",
          7018 => x"61",
          7019 => x"59",
          7020 => x"90",
          7021 => x"34",
          7022 => x"eb",
          7023 => x"34",
          7024 => x"61",
          7025 => x"ef",
          7026 => x"aa",
          7027 => x"60",
          7028 => x"81",
          7029 => x"51",
          7030 => x"55",
          7031 => x"61",
          7032 => x"5a",
          7033 => x"8d",
          7034 => x"81",
          7035 => x"b4",
          7036 => x"9e",
          7037 => x"2e",
          7038 => x"58",
          7039 => x"86",
          7040 => x"76",
          7041 => x"55",
          7042 => x"0d",
          7043 => x"05",
          7044 => x"2e",
          7045 => x"80",
          7046 => x"77",
          7047 => x"34",
          7048 => x"38",
          7049 => x"18",
          7050 => x"fc",
          7051 => x"76",
          7052 => x"7a",
          7053 => x"2a",
          7054 => x"88",
          7055 => x"8d",
          7056 => x"a3",
          7057 => x"05",
          7058 => x"77",
          7059 => x"58",
          7060 => x"a1",
          7061 => x"80",
          7062 => x"80",
          7063 => x"56",
          7064 => x"74",
          7065 => x"0c",
          7066 => x"80",
          7067 => x"ac",
          7068 => x"76",
          7069 => x"b8",
          7070 => x"ba",
          7071 => x"9f",
          7072 => x"11",
          7073 => x"08",
          7074 => x"32",
          7075 => x"70",
          7076 => x"39",
          7077 => x"ff",
          7078 => x"9f",
          7079 => x"02",
          7080 => x"80",
          7081 => x"72",
          7082 => x"b8",
          7083 => x"ff",
          7084 => x"2e",
          7085 => x"2e",
          7086 => x"72",
          7087 => x"83",
          7088 => x"ff",
          7089 => x"a8",
          7090 => x"81",
          7091 => x"b8",
          7092 => x"fe",
          7093 => x"84",
          7094 => x"53",
          7095 => x"53",
          7096 => x"0d",
          7097 => x"06",
          7098 => x"38",
          7099 => x"22",
          7100 => x"0d",
          7101 => x"83",
          7102 => x"83",
          7103 => x"56",
          7104 => x"74",
          7105 => x"30",
          7106 => x"54",
          7107 => x"70",
          7108 => x"2a",
          7109 => x"52",
          7110 => x"cf",
          7111 => x"05",
          7112 => x"25",
          7113 => x"70",
          7114 => x"84",
          7115 => x"83",
          7116 => x"88",
          7117 => x"c9",
          7118 => x"a0",
          7119 => x"51",
          7120 => x"70",
          7121 => x"39",
          7122 => x"57",
          7123 => x"ff",
          7124 => x"16",
          7125 => x"d0",
          7126 => x"06",
          7127 => x"83",
          7128 => x"39",
          7129 => x"31",
          7130 => x"55",
          7131 => x"75",
          7132 => x"39",
          7133 => x"ff",
          7134 => x"ff",
          7135 => x"00",
          7136 => x"00",
          7137 => x"00",
          7138 => x"00",
          7139 => x"00",
          7140 => x"00",
          7141 => x"00",
          7142 => x"00",
          7143 => x"00",
          7144 => x"00",
          7145 => x"00",
          7146 => x"00",
          7147 => x"00",
          7148 => x"00",
          7149 => x"00",
          7150 => x"00",
          7151 => x"00",
          7152 => x"00",
          7153 => x"00",
          7154 => x"00",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"64",
          7372 => x"64",
          7373 => x"66",
          7374 => x"66",
          7375 => x"66",
          7376 => x"6d",
          7377 => x"6d",
          7378 => x"6d",
          7379 => x"6d",
          7380 => x"6d",
          7381 => x"6d",
          7382 => x"68",
          7383 => x"68",
          7384 => x"00",
          7385 => x"72",
          7386 => x"72",
          7387 => x"69",
          7388 => x"74",
          7389 => x"63",
          7390 => x"74",
          7391 => x"6d",
          7392 => x"6b",
          7393 => x"65",
          7394 => x"6f",
          7395 => x"72",
          7396 => x"6d",
          7397 => x"6e",
          7398 => x"2e",
          7399 => x"6d",
          7400 => x"6e",
          7401 => x"00",
          7402 => x"66",
          7403 => x"20",
          7404 => x"00",
          7405 => x"20",
          7406 => x"65",
          7407 => x"6f",
          7408 => x"72",
          7409 => x"61",
          7410 => x"2e",
          7411 => x"61",
          7412 => x"65",
          7413 => x"6f",
          7414 => x"65",
          7415 => x"73",
          7416 => x"6e",
          7417 => x"73",
          7418 => x"20",
          7419 => x"62",
          7420 => x"44",
          7421 => x"6d",
          7422 => x"69",
          7423 => x"00",
          7424 => x"73",
          7425 => x"70",
          7426 => x"64",
          7427 => x"20",
          7428 => x"69",
          7429 => x"00",
          7430 => x"20",
          7431 => x"20",
          7432 => x"00",
          7433 => x"73",
          7434 => x"64",
          7435 => x"6c",
          7436 => x"6e",
          7437 => x"4e",
          7438 => x"66",
          7439 => x"4e",
          7440 => x"66",
          7441 => x"44",
          7442 => x"20",
          7443 => x"49",
          7444 => x"20",
          7445 => x"44",
          7446 => x"6f",
          7447 => x"65",
          7448 => x"0a",
          7449 => x"65",
          7450 => x"20",
          7451 => x"65",
          7452 => x"00",
          7453 => x"00",
          7454 => x"58",
          7455 => x"25",
          7456 => x"20",
          7457 => x"20",
          7458 => x"00",
          7459 => x"20",
          7460 => x"7a",
          7461 => x"73",
          7462 => x"33",
          7463 => x"76",
          7464 => x"20",
          7465 => x"76",
          7466 => x"25",
          7467 => x"0a",
          7468 => x"49",
          7469 => x"74",
          7470 => x"72",
          7471 => x"31",
          7472 => x"65",
          7473 => x"55",
          7474 => x"20",
          7475 => x"70",
          7476 => x"30",
          7477 => x"65",
          7478 => x"55",
          7479 => x"20",
          7480 => x"70",
          7481 => x"4c",
          7482 => x"65",
          7483 => x"49",
          7484 => x"20",
          7485 => x"70",
          7486 => x"69",
          7487 => x"74",
          7488 => x"72",
          7489 => x"75",
          7490 => x"69",
          7491 => x"69",
          7492 => x"45",
          7493 => x"20",
          7494 => x"2e",
          7495 => x"65",
          7496 => x"00",
          7497 => x"7a",
          7498 => x"46",
          7499 => x"6f",
          7500 => x"6c",
          7501 => x"63",
          7502 => x"70",
          7503 => x"6e",
          7504 => x"61",
          7505 => x"2a",
          7506 => x"25",
          7507 => x"42",
          7508 => x"61",
          7509 => x"5a",
          7510 => x"25",
          7511 => x"73",
          7512 => x"43",
          7513 => x"6f",
          7514 => x"2e",
          7515 => x"61",
          7516 => x"70",
          7517 => x"6f",
          7518 => x"43",
          7519 => x"63",
          7520 => x"30",
          7521 => x"0a",
          7522 => x"20",
          7523 => x"64",
          7524 => x"25",
          7525 => x"45",
          7526 => x"67",
          7527 => x"20",
          7528 => x"2e",
          7529 => x"58",
          7530 => x"00",
          7531 => x"58",
          7532 => x"43",
          7533 => x"67",
          7534 => x"25",
          7535 => x"38",
          7536 => x"6c",
          7537 => x"0a",
          7538 => x"69",
          7539 => x"25",
          7540 => x"32",
          7541 => x"72",
          7542 => x"00",
          7543 => x"20",
          7544 => x"0a",
          7545 => x"65",
          7546 => x"25",
          7547 => x"4d",
          7548 => x"78",
          7549 => x"2c",
          7550 => x"20",
          7551 => x"20",
          7552 => x"2e",
          7553 => x"25",
          7554 => x"20",
          7555 => x"64",
          7556 => x"53",
          7557 => x"69",
          7558 => x"6e",
          7559 => x"76",
          7560 => x"70",
          7561 => x"64",
          7562 => x"65",
          7563 => x"20",
          7564 => x"52",
          7565 => x"63",
          7566 => x"72",
          7567 => x"30",
          7568 => x"20",
          7569 => x"4d",
          7570 => x"74",
          7571 => x"72",
          7572 => x"30",
          7573 => x"20",
          7574 => x"6b",
          7575 => x"41",
          7576 => x"20",
          7577 => x"30",
          7578 => x"4d",
          7579 => x"20",
          7580 => x"49",
          7581 => x"20",
          7582 => x"20",
          7583 => x"30",
          7584 => x"20",
          7585 => x"65",
          7586 => x"20",
          7587 => x"20",
          7588 => x"64",
          7589 => x"7a",
          7590 => x"57",
          7591 => x"20",
          7592 => x"6c",
          7593 => x"71",
          7594 => x"34",
          7595 => x"20",
          7596 => x"4d",
          7597 => x"46",
          7598 => x"20",
          7599 => x"64",
          7600 => x"7a",
          7601 => x"53",
          7602 => x"50",
          7603 => x"49",
          7604 => x"20",
          7605 => x"32",
          7606 => x"57",
          7607 => x"20",
          7608 => x"20",
          7609 => x"20",
          7610 => x"68",
          7611 => x"25",
          7612 => x"20",
          7613 => x"52",
          7614 => x"69",
          7615 => x"25",
          7616 => x"20",
          7617 => x"41",
          7618 => x"65",
          7619 => x"25",
          7620 => x"20",
          7621 => x"20",
          7622 => x"30",
          7623 => x"29",
          7624 => x"42",
          7625 => x"20",
          7626 => x"25",
          7627 => x"20",
          7628 => x"20",
          7629 => x"30",
          7630 => x"29",
          7631 => x"53",
          7632 => x"20",
          7633 => x"25",
          7634 => x"20",
          7635 => x"44",
          7636 => x"30",
          7637 => x"29",
          7638 => x"6f",
          7639 => x"6f",
          7640 => x"55",
          7641 => x"45",
          7642 => x"53",
          7643 => x"4d",
          7644 => x"46",
          7645 => x"45",
          7646 => x"01",
          7647 => x"00",
          7648 => x"00",
          7649 => x"01",
          7650 => x"00",
          7651 => x"00",
          7652 => x"01",
          7653 => x"00",
          7654 => x"00",
          7655 => x"01",
          7656 => x"00",
          7657 => x"00",
          7658 => x"01",
          7659 => x"00",
          7660 => x"00",
          7661 => x"01",
          7662 => x"00",
          7663 => x"00",
          7664 => x"04",
          7665 => x"00",
          7666 => x"00",
          7667 => x"03",
          7668 => x"00",
          7669 => x"00",
          7670 => x"04",
          7671 => x"00",
          7672 => x"00",
          7673 => x"03",
          7674 => x"00",
          7675 => x"00",
          7676 => x"03",
          7677 => x"00",
          7678 => x"00",
          7679 => x"1b",
          7680 => x"1b",
          7681 => x"1b",
          7682 => x"1b",
          7683 => x"1b",
          7684 => x"10",
          7685 => x"0d",
          7686 => x"08",
          7687 => x"05",
          7688 => x"03",
          7689 => x"01",
          7690 => x"6f",
          7691 => x"63",
          7692 => x"69",
          7693 => x"69",
          7694 => x"61",
          7695 => x"68",
          7696 => x"68",
          7697 => x"21",
          7698 => x"75",
          7699 => x"46",
          7700 => x"6f",
          7701 => x"74",
          7702 => x"6f",
          7703 => x"20",
          7704 => x"00",
          7705 => x"00",
          7706 => x"00",
          7707 => x"1b",
          7708 => x"1b",
          7709 => x"7e",
          7710 => x"7e",
          7711 => x"7e",
          7712 => x"7e",
          7713 => x"7e",
          7714 => x"7e",
          7715 => x"7e",
          7716 => x"7e",
          7717 => x"7e",
          7718 => x"7e",
          7719 => x"00",
          7720 => x"00",
          7721 => x"1b",
          7722 => x"1b",
          7723 => x"58",
          7724 => x"25",
          7725 => x"2c",
          7726 => x"00",
          7727 => x"2d",
          7728 => x"63",
          7729 => x"25",
          7730 => x"4b",
          7731 => x"25",
          7732 => x"25",
          7733 => x"52",
          7734 => x"72",
          7735 => x"72",
          7736 => x"30",
          7737 => x"00",
          7738 => x"30",
          7739 => x"00",
          7740 => x"30",
          7741 => x"4e",
          7742 => x"64",
          7743 => x"00",
          7744 => x"22",
          7745 => x"00",
          7746 => x"5b",
          7747 => x"46",
          7748 => x"eb",
          7749 => x"35",
          7750 => x"41",
          7751 => x"41",
          7752 => x"4e",
          7753 => x"20",
          7754 => x"20",
          7755 => x"00",
          7756 => x"00",
          7757 => x"09",
          7758 => x"1e",
          7759 => x"8e",
          7760 => x"49",
          7761 => x"99",
          7762 => x"9c",
          7763 => x"a5",
          7764 => x"ac",
          7765 => x"b4",
          7766 => x"bc",
          7767 => x"c4",
          7768 => x"cc",
          7769 => x"d4",
          7770 => x"dc",
          7771 => x"e4",
          7772 => x"ec",
          7773 => x"f4",
          7774 => x"fc",
          7775 => x"3d",
          7776 => x"3c",
          7777 => x"00",
          7778 => x"01",
          7779 => x"00",
          7780 => x"00",
          7781 => x"00",
          7782 => x"00",
          7783 => x"00",
          7784 => x"00",
          7785 => x"00",
          7786 => x"00",
          7787 => x"00",
          7788 => x"00",
          7789 => x"00",
          7790 => x"00",
          7791 => x"00",
          7792 => x"00",
          7793 => x"25",
          7794 => x"25",
          7795 => x"25",
          7796 => x"25",
          7797 => x"25",
          7798 => x"25",
          7799 => x"25",
          7800 => x"25",
          7801 => x"25",
          7802 => x"25",
          7803 => x"25",
          7804 => x"25",
          7805 => x"03",
          7806 => x"03",
          7807 => x"03",
          7808 => x"22",
          7809 => x"22",
          7810 => x"23",
          7811 => x"00",
          7812 => x"20",
          7813 => x"00",
          7814 => x"00",
          7815 => x"01",
          7816 => x"01",
          7817 => x"01",
          7818 => x"00",
          7819 => x"01",
          7820 => x"01",
          7821 => x"01",
          7822 => x"01",
          7823 => x"01",
          7824 => x"01",
          7825 => x"01",
          7826 => x"01",
          7827 => x"01",
          7828 => x"01",
          7829 => x"01",
          7830 => x"01",
          7831 => x"01",
          7832 => x"01",
          7833 => x"01",
          7834 => x"01",
          7835 => x"01",
          7836 => x"01",
          7837 => x"01",
          7838 => x"01",
          7839 => x"01",
          7840 => x"01",
          7841 => x"02",
          7842 => x"2c",
          7843 => x"2c",
          7844 => x"02",
          7845 => x"00",
          7846 => x"01",
          7847 => x"02",
          7848 => x"02",
          7849 => x"02",
          7850 => x"02",
          7851 => x"02",
          7852 => x"02",
          7853 => x"01",
          7854 => x"02",
          7855 => x"02",
          7856 => x"02",
          7857 => x"02",
          7858 => x"02",
          7859 => x"01",
          7860 => x"02",
          7861 => x"01",
          7862 => x"03",
          7863 => x"03",
          7864 => x"03",
          7865 => x"03",
          7866 => x"03",
          7867 => x"03",
          7868 => x"00",
          7869 => x"03",
          7870 => x"03",
          7871 => x"03",
          7872 => x"01",
          7873 => x"01",
          7874 => x"04",
          7875 => x"00",
          7876 => x"2c",
          7877 => x"01",
          7878 => x"06",
          7879 => x"06",
          7880 => x"00",
          7881 => x"1f",
          7882 => x"1f",
          7883 => x"1f",
          7884 => x"1f",
          7885 => x"1f",
          7886 => x"1f",
          7887 => x"1f",
          7888 => x"1f",
          7889 => x"1f",
          7890 => x"1f",
          7891 => x"06",
          7892 => x"1f",
          7893 => x"00",
          7894 => x"21",
          7895 => x"05",
          7896 => x"01",
          7897 => x"01",
          7898 => x"08",
          7899 => x"00",
          7900 => x"01",
          7901 => x"00",
          7902 => x"01",
          7903 => x"00",
          7904 => x"01",
          7905 => x"00",
          7906 => x"01",
          7907 => x"00",
          7908 => x"01",
          7909 => x"00",
          7910 => x"01",
          7911 => x"00",
          7912 => x"01",
          7913 => x"00",
          7914 => x"01",
          7915 => x"00",
          7916 => x"01",
          7917 => x"00",
          7918 => x"01",
          7919 => x"00",
          7920 => x"01",
          7921 => x"00",
          7922 => x"01",
          7923 => x"00",
          7924 => x"01",
          7925 => x"00",
          7926 => x"01",
          7927 => x"00",
          7928 => x"01",
          7929 => x"00",
          7930 => x"01",
          7931 => x"00",
          7932 => x"01",
          7933 => x"00",
          7934 => x"01",
          7935 => x"00",
          7936 => x"01",
          7937 => x"00",
          7938 => x"01",
          7939 => x"00",
          7940 => x"01",
          7941 => x"00",
          7942 => x"01",
          7943 => x"00",
          7944 => x"01",
          7945 => x"00",
          7946 => x"01",
          7947 => x"00",
          7948 => x"01",
          7949 => x"00",
          7950 => x"01",
          7951 => x"00",
          7952 => x"01",
          7953 => x"00",
          7954 => x"01",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"00",
          7959 => x"00",
          7960 => x"01",
          7961 => x"00",
          7962 => x"00",
          7963 => x"05",
          7964 => x"05",
          7965 => x"01",
          7966 => x"01",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"00",
          7983 => x"f0",
          7984 => x"5d",
          7985 => x"75",
          7986 => x"6d",
          7987 => x"65",
          7988 => x"35",
          7989 => x"30",
          7990 => x"f1",
          7991 => x"f0",
          7992 => x"84",
          7993 => x"f0",
          7994 => x"5d",
          7995 => x"55",
          7996 => x"4d",
          7997 => x"45",
          7998 => x"35",
          7999 => x"30",
          8000 => x"f1",
          8001 => x"f0",
          8002 => x"84",
          8003 => x"f0",
          8004 => x"7d",
          8005 => x"55",
          8006 => x"4d",
          8007 => x"45",
          8008 => x"25",
          8009 => x"20",
          8010 => x"f9",
          8011 => x"f0",
          8012 => x"89",
          8013 => x"f0",
          8014 => x"1d",
          8015 => x"15",
          8016 => x"0d",
          8017 => x"05",
          8018 => x"f0",
          8019 => x"f0",
          8020 => x"f0",
          8021 => x"f0",
          8022 => x"84",
          8023 => x"f0",
          8024 => x"b7",
          8025 => x"39",
          8026 => x"1d",
          8027 => x"74",
          8028 => x"7a",
          8029 => x"9d",
          8030 => x"c3",
          8031 => x"f0",
          8032 => x"84",
          8033 => x"00",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"00",
          8045 => x"00",
          8046 => x"f8",
          8047 => x"f3",
          8048 => x"f4",
          8049 => x"f1",
          8050 => x"f2",
          8051 => x"80",
          8052 => x"81",
          8053 => x"82",
          8054 => x"83",
          8055 => x"84",
          8056 => x"85",
          8057 => x"86",
          8058 => x"87",
          8059 => x"88",
          8060 => x"89",
          8061 => x"f6",
          8062 => x"7f",
          8063 => x"f9",
          8064 => x"e0",
          8065 => x"e1",
          8066 => x"71",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"50",
          9068 => x"cc",
          9069 => x"f8",
          9070 => x"e1",
          9071 => x"e3",
          9072 => x"00",
          9073 => x"68",
          9074 => x"20",
          9075 => x"28",
          9076 => x"55",
          9077 => x"08",
          9078 => x"10",
          9079 => x"18",
          9080 => x"c7",
          9081 => x"88",
          9082 => x"90",
          9083 => x"98",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"01",
        others => X"00"
    );

    shared variable RAM4 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"80",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"09",
             9 => x"83",
            10 => x"00",
            11 => x"00",
            12 => x"73",
            13 => x"83",
            14 => x"ff",
            15 => x"00",
            16 => x"73",
            17 => x"06",
            18 => x"00",
            19 => x"00",
            20 => x"53",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"72",
            26 => x"06",
            27 => x"00",
            28 => x"53",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"00",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"04",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"0b",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"2a",
            49 => x"05",
            50 => x"00",
            51 => x"00",
            52 => x"83",
            53 => x"2b",
            54 => x"51",
            55 => x"00",
            56 => x"70",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"70",
            61 => x"06",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"51",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"06",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"09",
            77 => x"2a",
            78 => x"00",
            79 => x"00",
            80 => x"bd",
            81 => x"08",
            82 => x"00",
            83 => x"00",
            84 => x"75",
            85 => x"50",
            86 => x"88",
            87 => x"00",
            88 => x"75",
            89 => x"50",
            90 => x"88",
            91 => x"00",
            92 => x"0a",
            93 => x"06",
            94 => x"06",
            95 => x"00",
            96 => x"0a",
            97 => x"71",
            98 => x"05",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"52",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"51",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"8c",
           134 => x"04",
           135 => x"0b",
           136 => x"8c",
           137 => x"04",
           138 => x"0b",
           139 => x"8d",
           140 => x"04",
           141 => x"0b",
           142 => x"8d",
           143 => x"04",
           144 => x"0b",
           145 => x"8e",
           146 => x"04",
           147 => x"0b",
           148 => x"8e",
           149 => x"04",
           150 => x"0b",
           151 => x"8f",
           152 => x"04",
           153 => x"0b",
           154 => x"8f",
           155 => x"04",
           156 => x"0b",
           157 => x"90",
           158 => x"04",
           159 => x"0b",
           160 => x"90",
           161 => x"04",
           162 => x"0b",
           163 => x"91",
           164 => x"04",
           165 => x"0b",
           166 => x"91",
           167 => x"04",
           168 => x"0b",
           169 => x"92",
           170 => x"04",
           171 => x"0b",
           172 => x"92",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"f0",
           193 => x"f0",
           194 => x"b8",
           195 => x"f0",
           196 => x"b8",
           197 => x"f0",
           198 => x"b8",
           199 => x"f0",
           200 => x"b8",
           201 => x"f0",
           202 => x"b8",
           203 => x"f0",
           204 => x"b8",
           205 => x"f0",
           206 => x"b8",
           207 => x"f0",
           208 => x"b8",
           209 => x"f0",
           210 => x"b8",
           211 => x"f0",
           212 => x"b8",
           213 => x"f0",
           214 => x"b8",
           215 => x"f0",
           216 => x"b8",
           217 => x"b8",
           218 => x"84",
           219 => x"84",
           220 => x"04",
           221 => x"2d",
           222 => x"90",
           223 => x"c0",
           224 => x"80",
           225 => x"c9",
           226 => x"c0",
           227 => x"82",
           228 => x"80",
           229 => x"0c",
           230 => x"08",
           231 => x"f0",
           232 => x"f0",
           233 => x"b8",
           234 => x"b8",
           235 => x"84",
           236 => x"84",
           237 => x"04",
           238 => x"2d",
           239 => x"90",
           240 => x"ad",
           241 => x"80",
           242 => x"f2",
           243 => x"c0",
           244 => x"82",
           245 => x"80",
           246 => x"0c",
           247 => x"08",
           248 => x"f0",
           249 => x"f0",
           250 => x"b8",
           251 => x"b8",
           252 => x"84",
           253 => x"84",
           254 => x"04",
           255 => x"2d",
           256 => x"90",
           257 => x"f7",
           258 => x"80",
           259 => x"e5",
           260 => x"c0",
           261 => x"82",
           262 => x"80",
           263 => x"0c",
           264 => x"08",
           265 => x"f0",
           266 => x"f0",
           267 => x"b8",
           268 => x"b8",
           269 => x"84",
           270 => x"84",
           271 => x"04",
           272 => x"2d",
           273 => x"90",
           274 => x"ee",
           275 => x"80",
           276 => x"a4",
           277 => x"c0",
           278 => x"83",
           279 => x"80",
           280 => x"0c",
           281 => x"08",
           282 => x"f0",
           283 => x"f0",
           284 => x"b8",
           285 => x"b8",
           286 => x"84",
           287 => x"84",
           288 => x"04",
           289 => x"2d",
           290 => x"90",
           291 => x"df",
           292 => x"80",
           293 => x"d7",
           294 => x"c0",
           295 => x"b1",
           296 => x"c0",
           297 => x"81",
           298 => x"80",
           299 => x"0c",
           300 => x"08",
           301 => x"f0",
           302 => x"f0",
           303 => x"b8",
           304 => x"b8",
           305 => x"3c",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"ff",
           311 => x"83",
           312 => x"fc",
           313 => x"80",
           314 => x"06",
           315 => x"0a",
           316 => x"51",
           317 => x"d0",
           318 => x"05",
           319 => x"04",
           320 => x"00",
           321 => x"84",
           322 => x"84",
           323 => x"86",
           324 => x"7a",
           325 => x"06",
           326 => x"57",
           327 => x"06",
           328 => x"8a",
           329 => x"2a",
           330 => x"25",
           331 => x"75",
           332 => x"08",
           333 => x"ae",
           334 => x"81",
           335 => x"32",
           336 => x"51",
           337 => x"38",
           338 => x"b8",
           339 => x"0b",
           340 => x"04",
           341 => x"84",
           342 => x"0a",
           343 => x"52",
           344 => x"73",
           345 => x"0d",
           346 => x"05",
           347 => x"85",
           348 => x"63",
           349 => x"1f",
           350 => x"81",
           351 => x"54",
           352 => x"d2",
           353 => x"80",
           354 => x"54",
           355 => x"d0",
           356 => x"38",
           357 => x"25",
           358 => x"80",
           359 => x"81",
           360 => x"2e",
           361 => x"7b",
           362 => x"1d",
           363 => x"91",
           364 => x"78",
           365 => x"98",
           366 => x"80",
           367 => x"2c",
           368 => x"24",
           369 => x"72",
           370 => x"58",
           371 => x"76",
           372 => x"81",
           373 => x"33",
           374 => x"9e",
           375 => x"3f",
           376 => x"ff",
           377 => x"06",
           378 => x"74",
           379 => x"17",
           380 => x"72",
           381 => x"73",
           382 => x"80",
           383 => x"76",
           384 => x"58",
           385 => x"39",
           386 => x"5a",
           387 => x"83",
           388 => x"84",
           389 => x"93",
           390 => x"ff",
           391 => x"05",
           392 => x"84",
           393 => x"7e",
           394 => x"75",
           395 => x"08",
           396 => x"7d",
           397 => x"b2",
           398 => x"38",
           399 => x"80",
           400 => x"86",
           401 => x"80",
           402 => x"29",
           403 => x"2e",
           404 => x"fc",
           405 => x"58",
           406 => x"55",
           407 => x"2c",
           408 => x"73",
           409 => x"f7",
           410 => x"41",
           411 => x"80",
           412 => x"90",
           413 => x"06",
           414 => x"96",
           415 => x"73",
           416 => x"06",
           417 => x"2a",
           418 => x"7e",
           419 => x"7a",
           420 => x"2e",
           421 => x"29",
           422 => x"5a",
           423 => x"7c",
           424 => x"78",
           425 => x"05",
           426 => x"80",
           427 => x"72",
           428 => x"80",
           429 => x"98",
           430 => x"9d",
           431 => x"3f",
           432 => x"ff",
           433 => x"55",
           434 => x"2a",
           435 => x"2e",
           436 => x"84",
           437 => x"ca",
           438 => x"38",
           439 => x"7c",
           440 => x"87",
           441 => x"09",
           442 => x"5b",
           443 => x"78",
           444 => x"05",
           445 => x"75",
           446 => x"51",
           447 => x"07",
           448 => x"5b",
           449 => x"7a",
           450 => x"90",
           451 => x"83",
           452 => x"5a",
           453 => x"77",
           454 => x"70",
           455 => x"80",
           456 => x"2c",
           457 => x"7a",
           458 => x"7a",
           459 => x"80",
           460 => x"2c",
           461 => x"b3",
           462 => x"3f",
           463 => x"ff",
           464 => x"2e",
           465 => x"81",
           466 => x"e2",
           467 => x"06",
           468 => x"fe",
           469 => x"05",
           470 => x"39",
           471 => x"07",
           472 => x"80",
           473 => x"80",
           474 => x"5d",
           475 => x"fb",
           476 => x"70",
           477 => x"82",
           478 => x"5b",
           479 => x"7a",
           480 => x"f8",
           481 => x"07",
           482 => x"f7",
           483 => x"84",
           484 => x"58",
           485 => x"51",
           486 => x"83",
           487 => x"2b",
           488 => x"87",
           489 => x"58",
           490 => x"39",
           491 => x"81",
           492 => x"cf",
           493 => x"b8",
           494 => x"71",
           495 => x"7a",
           496 => x"76",
           497 => x"78",
           498 => x"05",
           499 => x"74",
           500 => x"51",
           501 => x"b0",
           502 => x"09",
           503 => x"76",
           504 => x"81",
           505 => x"38",
           506 => x"71",
           507 => x"83",
           508 => x"fa",
           509 => x"ad",
           510 => x"54",
           511 => x"ad",
           512 => x"82",
           513 => x"80",
           514 => x"78",
           515 => x"5a",
           516 => x"51",
           517 => x"a0",
           518 => x"78",
           519 => x"b8",
           520 => x"71",
           521 => x"39",
           522 => x"ff",
           523 => x"39",
           524 => x"53",
           525 => x"84",
           526 => x"55",
           527 => x"11",
           528 => x"81",
           529 => x"56",
           530 => x"d5",
           531 => x"53",
           532 => x"c8",
           533 => x"53",
           534 => x"2e",
           535 => x"05",
           536 => x"38",
           537 => x"84",
           538 => x"08",
           539 => x"74",
           540 => x"83",
           541 => x"b8",
           542 => x"3d",
           543 => x"85",
           544 => x"70",
           545 => x"56",
           546 => x"38",
           547 => x"72",
           548 => x"76",
           549 => x"3d",
           550 => x"33",
           551 => x"52",
           552 => x"2d",
           553 => x"38",
           554 => x"54",
           555 => x"3d",
           556 => x"51",
           557 => x"3d",
           558 => x"81",
           559 => x"56",
           560 => x"82",
           561 => x"ac",
           562 => x"16",
           563 => x"76",
           564 => x"0c",
           565 => x"16",
           566 => x"0c",
           567 => x"81",
           568 => x"73",
           569 => x"e3",
           570 => x"16",
           571 => x"0d",
           572 => x"06",
           573 => x"56",
           574 => x"86",
           575 => x"72",
           576 => x"2e",
           577 => x"53",
           578 => x"81",
           579 => x"05",
           580 => x"54",
           581 => x"0d",
           582 => x"85",
           583 => x"8c",
           584 => x"e4",
           585 => x"94",
           586 => x"e4",
           587 => x"25",
           588 => x"90",
           589 => x"ff",
           590 => x"72",
           591 => x"b8",
           592 => x"a0",
           593 => x"54",
           594 => x"71",
           595 => x"53",
           596 => x"52",
           597 => x"70",
           598 => x"f0",
           599 => x"3d",
           600 => x"71",
           601 => x"2e",
           602 => x"70",
           603 => x"05",
           604 => x"34",
           605 => x"84",
           606 => x"70",
           607 => x"70",
           608 => x"13",
           609 => x"11",
           610 => x"13",
           611 => x"34",
           612 => x"39",
           613 => x"71",
           614 => x"f7",
           615 => x"b8",
           616 => x"fd",
           617 => x"54",
           618 => x"70",
           619 => x"f0",
           620 => x"3d",
           621 => x"71",
           622 => x"2e",
           623 => x"33",
           624 => x"11",
           625 => x"e4",
           626 => x"0d",
           627 => x"80",
           628 => x"81",
           629 => x"2e",
           630 => x"54",
           631 => x"53",
           632 => x"b8",
           633 => x"80",
           634 => x"51",
           635 => x"33",
           636 => x"38",
           637 => x"86",
           638 => x"0c",
           639 => x"77",
           640 => x"3f",
           641 => x"08",
           642 => x"3f",
           643 => x"e4",
           644 => x"e4",
           645 => x"53",
           646 => x"fe",
           647 => x"73",
           648 => x"04",
           649 => x"54",
           650 => x"38",
           651 => x"70",
           652 => x"71",
           653 => x"ff",
           654 => x"84",
           655 => x"fd",
           656 => x"53",
           657 => x"72",
           658 => x"11",
           659 => x"e4",
           660 => x"0d",
           661 => x"80",
           662 => x"3f",
           663 => x"53",
           664 => x"80",
           665 => x"31",
           666 => x"cb",
           667 => x"c3",
           668 => x"72",
           669 => x"55",
           670 => x"72",
           671 => x"77",
           672 => x"2c",
           673 => x"71",
           674 => x"55",
           675 => x"10",
           676 => x"0c",
           677 => x"76",
           678 => x"70",
           679 => x"90",
           680 => x"fe",
           681 => x"83",
           682 => x"70",
           683 => x"25",
           684 => x"2a",
           685 => x"06",
           686 => x"71",
           687 => x"81",
           688 => x"74",
           689 => x"e4",
           690 => x"56",
           691 => x"56",
           692 => x"86",
           693 => x"77",
           694 => x"94",
           695 => x"74",
           696 => x"85",
           697 => x"7a",
           698 => x"8b",
           699 => x"b8",
           700 => x"80",
           701 => x"3f",
           702 => x"73",
           703 => x"80",
           704 => x"12",
           705 => x"71",
           706 => x"74",
           707 => x"9f",
           708 => x"72",
           709 => x"06",
           710 => x"1c",
           711 => x"53",
           712 => x"0c",
           713 => x"78",
           714 => x"2c",
           715 => x"73",
           716 => x"75",
           717 => x"fc",
           718 => x"32",
           719 => x"3d",
           720 => x"5b",
           721 => x"70",
           722 => x"09",
           723 => x"78",
           724 => x"2e",
           725 => x"38",
           726 => x"14",
           727 => x"db",
           728 => x"27",
           729 => x"89",
           730 => x"55",
           731 => x"51",
           732 => x"13",
           733 => x"73",
           734 => x"81",
           735 => x"16",
           736 => x"56",
           737 => x"80",
           738 => x"7a",
           739 => x"0c",
           740 => x"70",
           741 => x"73",
           742 => x"38",
           743 => x"55",
           744 => x"90",
           745 => x"81",
           746 => x"14",
           747 => x"27",
           748 => x"0c",
           749 => x"15",
           750 => x"80",
           751 => x"b8",
           752 => x"3d",
           753 => x"7b",
           754 => x"59",
           755 => x"38",
           756 => x"55",
           757 => x"ad",
           758 => x"81",
           759 => x"77",
           760 => x"80",
           761 => x"80",
           762 => x"70",
           763 => x"70",
           764 => x"27",
           765 => x"06",
           766 => x"38",
           767 => x"76",
           768 => x"70",
           769 => x"ff",
           770 => x"75",
           771 => x"75",
           772 => x"04",
           773 => x"33",
           774 => x"81",
           775 => x"78",
           776 => x"e2",
           777 => x"f8",
           778 => x"27",
           779 => x"88",
           780 => x"75",
           781 => x"04",
           782 => x"70",
           783 => x"39",
           784 => x"3d",
           785 => x"b8",
           786 => x"e4",
           787 => x"71",
           788 => x"83",
           789 => x"83",
           790 => x"3d",
           791 => x"b3",
           792 => x"b4",
           793 => x"04",
           794 => x"83",
           795 => x"ef",
           796 => x"ce",
           797 => x"0d",
           798 => x"3f",
           799 => x"51",
           800 => x"83",
           801 => x"3d",
           802 => x"db",
           803 => x"fc",
           804 => x"04",
           805 => x"83",
           806 => x"ee",
           807 => x"d0",
           808 => x"0d",
           809 => x"3f",
           810 => x"51",
           811 => x"83",
           812 => x"3d",
           813 => x"83",
           814 => x"98",
           815 => x"04",
           816 => x"83",
           817 => x"ed",
           818 => x"3d",
           819 => x"05",
           820 => x"70",
           821 => x"59",
           822 => x"38",
           823 => x"ff",
           824 => x"e2",
           825 => x"70",
           826 => x"b8",
           827 => x"80",
           828 => x"af",
           829 => x"80",
           830 => x"06",
           831 => x"aa",
           832 => x"74",
           833 => x"52",
           834 => x"3f",
           835 => x"e4",
           836 => x"df",
           837 => x"96",
           838 => x"87",
           839 => x"08",
           840 => x"80",
           841 => x"bd",
           842 => x"b8",
           843 => x"74",
           844 => x"75",
           845 => x"52",
           846 => x"e4",
           847 => x"84",
           848 => x"53",
           849 => x"f8",
           850 => x"7c",
           851 => x"59",
           852 => x"51",
           853 => x"8b",
           854 => x"81",
           855 => x"0c",
           856 => x"d4",
           857 => x"b8",
           858 => x"2d",
           859 => x"0c",
           860 => x"7f",
           861 => x"05",
           862 => x"5c",
           863 => x"83",
           864 => x"51",
           865 => x"dd",
           866 => x"b2",
           867 => x"7c",
           868 => x"53",
           869 => x"33",
           870 => x"3f",
           871 => x"54",
           872 => x"26",
           873 => x"b8",
           874 => x"c0",
           875 => x"80",
           876 => x"55",
           877 => x"81",
           878 => x"06",
           879 => x"80",
           880 => x"d4",
           881 => x"3f",
           882 => x"38",
           883 => x"78",
           884 => x"9d",
           885 => x"2b",
           886 => x"2e",
           887 => x"c3",
           888 => x"fe",
           889 => x"0c",
           890 => x"51",
           891 => x"c8",
           892 => x"3f",
           893 => x"da",
           894 => x"3f",
           895 => x"54",
           896 => x"27",
           897 => x"7a",
           898 => x"d2",
           899 => x"84",
           900 => x"ea",
           901 => x"fe",
           902 => x"d0",
           903 => x"53",
           904 => x"79",
           905 => x"72",
           906 => x"83",
           907 => x"14",
           908 => x"51",
           909 => x"38",
           910 => x"52",
           911 => x"56",
           912 => x"84",
           913 => x"88",
           914 => x"a0",
           915 => x"06",
           916 => x"39",
           917 => x"e4",
           918 => x"a0",
           919 => x"30",
           920 => x"51",
           921 => x"80",
           922 => x"f9",
           923 => x"70",
           924 => x"72",
           925 => x"73",
           926 => x"57",
           927 => x"38",
           928 => x"e4",
           929 => x"0d",
           930 => x"c7",
           931 => x"d2",
           932 => x"9c",
           933 => x"06",
           934 => x"82",
           935 => x"82",
           936 => x"06",
           937 => x"84",
           938 => x"81",
           939 => x"06",
           940 => x"86",
           941 => x"80",
           942 => x"06",
           943 => x"2a",
           944 => x"df",
           945 => x"9b",
           946 => x"8a",
           947 => x"c7",
           948 => x"9b",
           949 => x"f2",
           950 => x"88",
           951 => x"c6",
           952 => x"3f",
           953 => x"80",
           954 => x"70",
           955 => x"ff",
           956 => x"a2",
           957 => x"3f",
           958 => x"2a",
           959 => x"2e",
           960 => x"51",
           961 => x"9b",
           962 => x"72",
           963 => x"71",
           964 => x"39",
           965 => x"d8",
           966 => x"d2",
           967 => x"51",
           968 => x"ff",
           969 => x"83",
           970 => x"51",
           971 => x"81",
           972 => x"e6",
           973 => x"9a",
           974 => x"3f",
           975 => x"2a",
           976 => x"2e",
           977 => x"3d",
           978 => x"84",
           979 => x"51",
           980 => x"08",
           981 => x"78",
           982 => x"d0",
           983 => x"83",
           984 => x"48",
           985 => x"eb",
           986 => x"33",
           987 => x"80",
           988 => x"83",
           989 => x"7d",
           990 => x"5a",
           991 => x"79",
           992 => x"06",
           993 => x"5a",
           994 => x"7b",
           995 => x"83",
           996 => x"e7",
           997 => x"b8",
           998 => x"52",
           999 => x"08",
          1000 => x"81",
          1001 => x"81",
          1002 => x"c4",
          1003 => x"2e",
          1004 => x"51",
          1005 => x"5e",
          1006 => x"c9",
          1007 => x"3d",
          1008 => x"84",
          1009 => x"5c",
          1010 => x"b8",
          1011 => x"b8",
          1012 => x"81",
          1013 => x"2e",
          1014 => x"e2",
          1015 => x"7b",
          1016 => x"7c",
          1017 => x"58",
          1018 => x"55",
          1019 => x"80",
          1020 => x"84",
          1021 => x"09",
          1022 => x"51",
          1023 => x"26",
          1024 => x"59",
          1025 => x"70",
          1026 => x"95",
          1027 => x"07",
          1028 => x"2e",
          1029 => x"d0",
          1030 => x"3f",
          1031 => x"7e",
          1032 => x"ed",
          1033 => x"59",
          1034 => x"d4",
          1035 => x"88",
          1036 => x"c5",
          1037 => x"d8",
          1038 => x"52",
          1039 => x"b8",
          1040 => x"b8",
          1041 => x"0b",
          1042 => x"06",
          1043 => x"06",
          1044 => x"f4",
          1045 => x"0b",
          1046 => x"c4",
          1047 => x"c3",
          1048 => x"b7",
          1049 => x"85",
          1050 => x"fd",
          1051 => x"c4",
          1052 => x"83",
          1053 => x"3f",
          1054 => x"51",
          1055 => x"08",
          1056 => x"38",
          1057 => x"fb",
          1058 => x"db",
          1059 => x"fe",
          1060 => x"55",
          1061 => x"d5",
          1062 => x"fd",
          1063 => x"ff",
          1064 => x"81",
          1065 => x"ef",
          1066 => x"39",
          1067 => x"80",
          1068 => x"de",
          1069 => x"39",
          1070 => x"80",
          1071 => x"e4",
          1072 => x"52",
          1073 => x"68",
          1074 => x"80",
          1075 => x"08",
          1076 => x"3f",
          1077 => x"11",
          1078 => x"3f",
          1079 => x"ff",
          1080 => x"d0",
          1081 => x"3d",
          1082 => x"51",
          1083 => x"80",
          1084 => x"f0",
          1085 => x"92",
          1086 => x"38",
          1087 => x"83",
          1088 => x"d4",
          1089 => x"51",
          1090 => x"59",
          1091 => x"9f",
          1092 => x"70",
          1093 => x"f4",
          1094 => x"ca",
          1095 => x"f8",
          1096 => x"53",
          1097 => x"84",
          1098 => x"59",
          1099 => x"d4",
          1100 => x"08",
          1101 => x"b3",
          1102 => x"ae",
          1103 => x"87",
          1104 => x"59",
          1105 => x"53",
          1106 => x"84",
          1107 => x"38",
          1108 => x"80",
          1109 => x"e4",
          1110 => x"3d",
          1111 => x"51",
          1112 => x"80",
          1113 => x"51",
          1114 => x"78",
          1115 => x"33",
          1116 => x"2e",
          1117 => x"33",
          1118 => x"ce",
          1119 => x"19",
          1120 => x"3d",
          1121 => x"51",
          1122 => x"80",
          1123 => x"fc",
          1124 => x"de",
          1125 => x"f7",
          1126 => x"53",
          1127 => x"84",
          1128 => x"38",
          1129 => x"68",
          1130 => x"65",
          1131 => x"7c",
          1132 => x"b8",
          1133 => x"05",
          1134 => x"08",
          1135 => x"fe",
          1136 => x"e7",
          1137 => x"38",
          1138 => x"98",
          1139 => x"08",
          1140 => x"fb",
          1141 => x"ae",
          1142 => x"84",
          1143 => x"39",
          1144 => x"79",
          1145 => x"fe",
          1146 => x"e7",
          1147 => x"2e",
          1148 => x"db",
          1149 => x"49",
          1150 => x"80",
          1151 => x"e4",
          1152 => x"b8",
          1153 => x"05",
          1154 => x"08",
          1155 => x"fe",
          1156 => x"e6",
          1157 => x"2e",
          1158 => x"11",
          1159 => x"3f",
          1160 => x"b8",
          1161 => x"cb",
          1162 => x"7a",
          1163 => x"70",
          1164 => x"f5",
          1165 => x"cf",
          1166 => x"87",
          1167 => x"3d",
          1168 => x"3f",
          1169 => x"78",
          1170 => x"08",
          1171 => x"e4",
          1172 => x"39",
          1173 => x"80",
          1174 => x"e4",
          1175 => x"5a",
          1176 => x"f1",
          1177 => x"11",
          1178 => x"3f",
          1179 => x"f1",
          1180 => x"8a",
          1181 => x"3d",
          1182 => x"51",
          1183 => x"80",
          1184 => x"7a",
          1185 => x"90",
          1186 => x"2a",
          1187 => x"2e",
          1188 => x"88",
          1189 => x"3f",
          1190 => x"52",
          1191 => x"c0",
          1192 => x"64",
          1193 => x"45",
          1194 => x"80",
          1195 => x"e4",
          1196 => x"64",
          1197 => x"b8",
          1198 => x"05",
          1199 => x"08",
          1200 => x"02",
          1201 => x"05",
          1202 => x"f0",
          1203 => x"e2",
          1204 => x"f2",
          1205 => x"05",
          1206 => x"7d",
          1207 => x"ff",
          1208 => x"b8",
          1209 => x"39",
          1210 => x"80",
          1211 => x"e4",
          1212 => x"5c",
          1213 => x"68",
          1214 => x"3d",
          1215 => x"51",
          1216 => x"80",
          1217 => x"0c",
          1218 => x"f7",
          1219 => x"06",
          1220 => x"ac",
          1221 => x"7c",
          1222 => x"7b",
          1223 => x"8c",
          1224 => x"3f",
          1225 => x"11",
          1226 => x"3f",
          1227 => x"38",
          1228 => x"79",
          1229 => x"f7",
          1230 => x"7b",
          1231 => x"ac",
          1232 => x"e9",
          1233 => x"83",
          1234 => x"83",
          1235 => x"59",
          1236 => x"d3",
          1237 => x"83",
          1238 => x"a5",
          1239 => x"8b",
          1240 => x"3f",
          1241 => x"59",
          1242 => x"b4",
          1243 => x"eb",
          1244 => x"83",
          1245 => x"83",
          1246 => x"9b",
          1247 => x"ee",
          1248 => x"80",
          1249 => x"49",
          1250 => x"5d",
          1251 => x"c4",
          1252 => x"d0",
          1253 => x"39",
          1254 => x"fb",
          1255 => x"84",
          1256 => x"70",
          1257 => x"74",
          1258 => x"08",
          1259 => x"84",
          1260 => x"74",
          1261 => x"87",
          1262 => x"87",
          1263 => x"3f",
          1264 => x"08",
          1265 => x"51",
          1266 => x"08",
          1267 => x"87",
          1268 => x"0b",
          1269 => x"e1",
          1270 => x"84",
          1271 => x"d4",
          1272 => x"0c",
          1273 => x"56",
          1274 => x"87",
          1275 => x"83",
          1276 => x"c4",
          1277 => x"52",
          1278 => x"54",
          1279 => x"52",
          1280 => x"8d",
          1281 => x"fb",
          1282 => x"80",
          1283 => x"83",
          1284 => x"52",
          1285 => x"91",
          1286 => x"ff",
          1287 => x"f1",
          1288 => x"a2",
          1289 => x"81",
          1290 => x"70",
          1291 => x"a0",
          1292 => x"2e",
          1293 => x"81",
          1294 => x"ff",
          1295 => x"81",
          1296 => x"32",
          1297 => x"52",
          1298 => x"80",
          1299 => x"76",
          1300 => x"0c",
          1301 => x"c4",
          1302 => x"81",
          1303 => x"ff",
          1304 => x"e4",
          1305 => x"55",
          1306 => x"09",
          1307 => x"fc",
          1308 => x"38",
          1309 => x"3d",
          1310 => x"72",
          1311 => x"08",
          1312 => x"e4",
          1313 => x"0d",
          1314 => x"53",
          1315 => x"38",
          1316 => x"52",
          1317 => x"13",
          1318 => x"80",
          1319 => x"52",
          1320 => x"13",
          1321 => x"80",
          1322 => x"52",
          1323 => x"8a",
          1324 => x"e7",
          1325 => x"c0",
          1326 => x"98",
          1327 => x"98",
          1328 => x"98",
          1329 => x"98",
          1330 => x"98",
          1331 => x"98",
          1332 => x"0c",
          1333 => x"0b",
          1334 => x"71",
          1335 => x"04",
          1336 => x"98",
          1337 => x"98",
          1338 => x"c0",
          1339 => x"34",
          1340 => x"83",
          1341 => x"5c",
          1342 => x"ac",
          1343 => x"c0",
          1344 => x"34",
          1345 => x"88",
          1346 => x"5a",
          1347 => x"79",
          1348 => x"ff",
          1349 => x"85",
          1350 => x"83",
          1351 => x"7d",
          1352 => x"88",
          1353 => x"0d",
          1354 => x"33",
          1355 => x"51",
          1356 => x"08",
          1357 => x"71",
          1358 => x"72",
          1359 => x"e4",
          1360 => x"80",
          1361 => x"98",
          1362 => x"ff",
          1363 => x"51",
          1364 => x"08",
          1365 => x"71",
          1366 => x"3d",
          1367 => x"2b",
          1368 => x"84",
          1369 => x"2c",
          1370 => x"73",
          1371 => x"73",
          1372 => x"0c",
          1373 => x"02",
          1374 => x"70",
          1375 => x"80",
          1376 => x"94",
          1377 => x"53",
          1378 => x"71",
          1379 => x"70",
          1380 => x"53",
          1381 => x"2a",
          1382 => x"81",
          1383 => x"52",
          1384 => x"94",
          1385 => x"b8",
          1386 => x"91",
          1387 => x"97",
          1388 => x"72",
          1389 => x"81",
          1390 => x"87",
          1391 => x"70",
          1392 => x"38",
          1393 => x"05",
          1394 => x"52",
          1395 => x"3d",
          1396 => x"80",
          1397 => x"77",
          1398 => x"f1",
          1399 => x"57",
          1400 => x"87",
          1401 => x"70",
          1402 => x"2e",
          1403 => x"06",
          1404 => x"32",
          1405 => x"38",
          1406 => x"cf",
          1407 => x"c0",
          1408 => x"38",
          1409 => x"0c",
          1410 => x"ff",
          1411 => x"88",
          1412 => x"81",
          1413 => x"81",
          1414 => x"c1",
          1415 => x"71",
          1416 => x"94",
          1417 => x"06",
          1418 => x"39",
          1419 => x"08",
          1420 => x"70",
          1421 => x"9e",
          1422 => x"c0",
          1423 => x"87",
          1424 => x"0c",
          1425 => x"ac",
          1426 => x"f1",
          1427 => x"83",
          1428 => x"08",
          1429 => x"b0",
          1430 => x"9e",
          1431 => x"c0",
          1432 => x"87",
          1433 => x"0c",
          1434 => x"cc",
          1435 => x"f1",
          1436 => x"52",
          1437 => x"9e",
          1438 => x"c0",
          1439 => x"87",
          1440 => x"0c",
          1441 => x"0b",
          1442 => x"80",
          1443 => x"fb",
          1444 => x"0b",
          1445 => x"80",
          1446 => x"2e",
          1447 => x"e6",
          1448 => x"08",
          1449 => x"52",
          1450 => x"71",
          1451 => x"c0",
          1452 => x"06",
          1453 => x"38",
          1454 => x"80",
          1455 => x"a0",
          1456 => x"80",
          1457 => x"f1",
          1458 => x"90",
          1459 => x"52",
          1460 => x"52",
          1461 => x"87",
          1462 => x"80",
          1463 => x"83",
          1464 => x"34",
          1465 => x"70",
          1466 => x"70",
          1467 => x"83",
          1468 => x"9e",
          1469 => x"51",
          1470 => x"81",
          1471 => x"0b",
          1472 => x"c0",
          1473 => x"2e",
          1474 => x"ee",
          1475 => x"08",
          1476 => x"70",
          1477 => x"83",
          1478 => x"08",
          1479 => x"51",
          1480 => x"87",
          1481 => x"06",
          1482 => x"38",
          1483 => x"87",
          1484 => x"70",
          1485 => x"f2",
          1486 => x"08",
          1487 => x"80",
          1488 => x"f1",
          1489 => x"87",
          1490 => x"83",
          1491 => x"39",
          1492 => x"ff",
          1493 => x"54",
          1494 => x"51",
          1495 => x"55",
          1496 => x"33",
          1497 => x"e8",
          1498 => x"f1",
          1499 => x"83",
          1500 => x"38",
          1501 => x"b3",
          1502 => x"84",
          1503 => x"74",
          1504 => x"56",
          1505 => x"33",
          1506 => x"ec",
          1507 => x"f1",
          1508 => x"83",
          1509 => x"38",
          1510 => x"83",
          1511 => x"51",
          1512 => x"08",
          1513 => x"b8",
          1514 => x"d9",
          1515 => x"d9",
          1516 => x"d4",
          1517 => x"b5",
          1518 => x"bd",
          1519 => x"3f",
          1520 => x"29",
          1521 => x"e4",
          1522 => x"b4",
          1523 => x"74",
          1524 => x"55",
          1525 => x"3f",
          1526 => x"08",
          1527 => x"c9",
          1528 => x"84",
          1529 => x"84",
          1530 => x"51",
          1531 => x"fe",
          1532 => x"dc",
          1533 => x"51",
          1534 => x"bd",
          1535 => x"54",
          1536 => x"d8",
          1537 => x"e6",
          1538 => x"38",
          1539 => x"c0",
          1540 => x"cb",
          1541 => x"d8",
          1542 => x"f1",
          1543 => x"ff",
          1544 => x"52",
          1545 => x"3f",
          1546 => x"83",
          1547 => x"51",
          1548 => x"08",
          1549 => x"c8",
          1550 => x"84",
          1551 => x"84",
          1552 => x"51",
          1553 => x"33",
          1554 => x"fe",
          1555 => x"bf",
          1556 => x"73",
          1557 => x"39",
          1558 => x"3f",
          1559 => x"2e",
          1560 => x"a0",
          1561 => x"ec",
          1562 => x"38",
          1563 => x"bf",
          1564 => x"73",
          1565 => x"83",
          1566 => x"51",
          1567 => x"33",
          1568 => x"d2",
          1569 => x"db",
          1570 => x"f1",
          1571 => x"e3",
          1572 => x"52",
          1573 => x"3f",
          1574 => x"2e",
          1575 => x"b0",
          1576 => x"52",
          1577 => x"3f",
          1578 => x"2e",
          1579 => x"a8",
          1580 => x"52",
          1581 => x"3f",
          1582 => x"2e",
          1583 => x"a0",
          1584 => x"52",
          1585 => x"3f",
          1586 => x"2e",
          1587 => x"b8",
          1588 => x"52",
          1589 => x"3f",
          1590 => x"2e",
          1591 => x"c0",
          1592 => x"52",
          1593 => x"3f",
          1594 => x"2e",
          1595 => x"ac",
          1596 => x"b4",
          1597 => x"e6",
          1598 => x"38",
          1599 => x"05",
          1600 => x"71",
          1601 => x"71",
          1602 => x"af",
          1603 => x"dd",
          1604 => x"3d",
          1605 => x"af",
          1606 => x"dd",
          1607 => x"3d",
          1608 => x"af",
          1609 => x"dd",
          1610 => x"3d",
          1611 => x"80",
          1612 => x"83",
          1613 => x"0c",
          1614 => x"ad",
          1615 => x"58",
          1616 => x"82",
          1617 => x"80",
          1618 => x"83",
          1619 => x"52",
          1620 => x"b8",
          1621 => x"51",
          1622 => x"81",
          1623 => x"e4",
          1624 => x"08",
          1625 => x"74",
          1626 => x"07",
          1627 => x"2e",
          1628 => x"f2",
          1629 => x"82",
          1630 => x"8f",
          1631 => x"84",
          1632 => x"83",
          1633 => x"78",
          1634 => x"76",
          1635 => x"51",
          1636 => x"84",
          1637 => x"83",
          1638 => x"80",
          1639 => x"0d",
          1640 => x"ad",
          1641 => x"57",
          1642 => x"91",
          1643 => x"75",
          1644 => x"70",
          1645 => x"84",
          1646 => x"08",
          1647 => x"08",
          1648 => x"81",
          1649 => x"99",
          1650 => x"57",
          1651 => x"54",
          1652 => x"0d",
          1653 => x"84",
          1654 => x"ce",
          1655 => x"d1",
          1656 => x"51",
          1657 => x"81",
          1658 => x"38",
          1659 => x"54",
          1660 => x"b6",
          1661 => x"76",
          1662 => x"5b",
          1663 => x"09",
          1664 => x"26",
          1665 => x"56",
          1666 => x"08",
          1667 => x"82",
          1668 => x"80",
          1669 => x"80",
          1670 => x"3f",
          1671 => x"38",
          1672 => x"b8",
          1673 => x"e4",
          1674 => x"08",
          1675 => x"77",
          1676 => x"83",
          1677 => x"3f",
          1678 => x"b2",
          1679 => x"aa",
          1680 => x"3d",
          1681 => x"5a",
          1682 => x"83",
          1683 => x"56",
          1684 => x"cc",
          1685 => x"cb",
          1686 => x"81",
          1687 => x"a0",
          1688 => x"93",
          1689 => x"eb",
          1690 => x"2b",
          1691 => x"2e",
          1692 => x"d0",
          1693 => x"2c",
          1694 => x"70",
          1695 => x"10",
          1696 => x"15",
          1697 => x"52",
          1698 => x"79",
          1699 => x"81",
          1700 => x"81",
          1701 => x"55",
          1702 => x"10",
          1703 => x"0b",
          1704 => x"77",
          1705 => x"15",
          1706 => x"75",
          1707 => x"c2",
          1708 => x"57",
          1709 => x"1b",
          1710 => x"d0",
          1711 => x"2c",
          1712 => x"83",
          1713 => x"5d",
          1714 => x"81",
          1715 => x"fe",
          1716 => x"38",
          1717 => x"0a",
          1718 => x"06",
          1719 => x"c0",
          1720 => x"51",
          1721 => x"33",
          1722 => x"83",
          1723 => x"42",
          1724 => x"76",
          1725 => x"39",
          1726 => x"38",
          1727 => x"39",
          1728 => x"84",
          1729 => x"34",
          1730 => x"55",
          1731 => x"10",
          1732 => x"08",
          1733 => x"0c",
          1734 => x"0b",
          1735 => x"d0",
          1736 => x"85",
          1737 => x"51",
          1738 => x"33",
          1739 => x"34",
          1740 => x"70",
          1741 => x"5b",
          1742 => x"38",
          1743 => x"58",
          1744 => x"70",
          1745 => x"fc",
          1746 => x"38",
          1747 => x"70",
          1748 => x"75",
          1749 => x"84",
          1750 => x"56",
          1751 => x"d4",
          1752 => x"a6",
          1753 => x"51",
          1754 => x"08",
          1755 => x"84",
          1756 => x"84",
          1757 => x"55",
          1758 => x"90",
          1759 => x"cd",
          1760 => x"08",
          1761 => x"10",
          1762 => x"57",
          1763 => x"56",
          1764 => x"51",
          1765 => x"08",
          1766 => x"08",
          1767 => x"52",
          1768 => x"d0",
          1769 => x"56",
          1770 => x"d4",
          1771 => x"8e",
          1772 => x"51",
          1773 => x"08",
          1774 => x"84",
          1775 => x"84",
          1776 => x"55",
          1777 => x"81",
          1778 => x"57",
          1779 => x"84",
          1780 => x"76",
          1781 => x"33",
          1782 => x"d0",
          1783 => x"d0",
          1784 => x"27",
          1785 => x"52",
          1786 => x"34",
          1787 => x"b3",
          1788 => x"81",
          1789 => x"57",
          1790 => x"f9",
          1791 => x"d0",
          1792 => x"f9",
          1793 => x"d0",
          1794 => x"2c",
          1795 => x"60",
          1796 => x"c8",
          1797 => x"3f",
          1798 => x"70",
          1799 => x"57",
          1800 => x"38",
          1801 => x"ff",
          1802 => x"29",
          1803 => x"84",
          1804 => x"7b",
          1805 => x"08",
          1806 => x"74",
          1807 => x"05",
          1808 => x"5d",
          1809 => x"38",
          1810 => x"18",
          1811 => x"52",
          1812 => x"75",
          1813 => x"05",
          1814 => x"5b",
          1815 => x"38",
          1816 => x"34",
          1817 => x"51",
          1818 => x"0a",
          1819 => x"2c",
          1820 => x"78",
          1821 => x"39",
          1822 => x"2e",
          1823 => x"52",
          1824 => x"d0",
          1825 => x"d0",
          1826 => x"dd",
          1827 => x"5f",
          1828 => x"52",
          1829 => x"d0",
          1830 => x"84",
          1831 => x"77",
          1832 => x"57",
          1833 => x"f2",
          1834 => x"fc",
          1835 => x"8b",
          1836 => x"06",
          1837 => x"53",
          1838 => x"b8",
          1839 => x"33",
          1840 => x"70",
          1841 => x"38",
          1842 => x"2e",
          1843 => x"77",
          1844 => x"84",
          1845 => x"a4",
          1846 => x"3d",
          1847 => x"74",
          1848 => x"08",
          1849 => x"84",
          1850 => x"af",
          1851 => x"88",
          1852 => x"a8",
          1853 => x"a8",
          1854 => x"cc",
          1855 => x"88",
          1856 => x"80",
          1857 => x"39",
          1858 => x"34",
          1859 => x"2e",
          1860 => x"88",
          1861 => x"c8",
          1862 => x"3f",
          1863 => x"ff",
          1864 => x"ff",
          1865 => x"7c",
          1866 => x"83",
          1867 => x"80",
          1868 => x"84",
          1869 => x"0c",
          1870 => x"33",
          1871 => x"80",
          1872 => x"33",
          1873 => x"34",
          1874 => x"34",
          1875 => x"ff",
          1876 => x"70",
          1877 => x"a4",
          1878 => x"24",
          1879 => x"52",
          1880 => x"d0",
          1881 => x"2c",
          1882 => x"56",
          1883 => x"d4",
          1884 => x"86",
          1885 => x"80",
          1886 => x"a4",
          1887 => x"f3",
          1888 => x"88",
          1889 => x"80",
          1890 => x"98",
          1891 => x"55",
          1892 => x"a5",
          1893 => x"77",
          1894 => x"33",
          1895 => x"80",
          1896 => x"98",
          1897 => x"5b",
          1898 => x"16",
          1899 => x"d4",
          1900 => x"ac",
          1901 => x"81",
          1902 => x"d0",
          1903 => x"24",
          1904 => x"d0",
          1905 => x"58",
          1906 => x"d0",
          1907 => x"38",
          1908 => x"41",
          1909 => x"5b",
          1910 => x"80",
          1911 => x"98",
          1912 => x"58",
          1913 => x"55",
          1914 => x"ff",
          1915 => x"7a",
          1916 => x"60",
          1917 => x"84",
          1918 => x"a8",
          1919 => x"ff",
          1920 => x"ff",
          1921 => x"24",
          1922 => x"98",
          1923 => x"59",
          1924 => x"d4",
          1925 => x"be",
          1926 => x"80",
          1927 => x"a4",
          1928 => x"f1",
          1929 => x"88",
          1930 => x"80",
          1931 => x"98",
          1932 => x"41",
          1933 => x"dd",
          1934 => x"80",
          1935 => x"ad",
          1936 => x"d0",
          1937 => x"ff",
          1938 => x"51",
          1939 => x"33",
          1940 => x"80",
          1941 => x"08",
          1942 => x"84",
          1943 => x"a9",
          1944 => x"88",
          1945 => x"a8",
          1946 => x"a8",
          1947 => x"39",
          1948 => x"b8",
          1949 => x"b8",
          1950 => x"f2",
          1951 => x"c3",
          1952 => x"16",
          1953 => x"3f",
          1954 => x"0a",
          1955 => x"33",
          1956 => x"38",
          1957 => x"70",
          1958 => x"58",
          1959 => x"38",
          1960 => x"80",
          1961 => x"57",
          1962 => x"38",
          1963 => x"80",
          1964 => x"d4",
          1965 => x"80",
          1966 => x"e7",
          1967 => x"80",
          1968 => x"d0",
          1969 => x"ee",
          1970 => x"3f",
          1971 => x"58",
          1972 => x"ff",
          1973 => x"3f",
          1974 => x"34",
          1975 => x"81",
          1976 => x"ab",
          1977 => x"33",
          1978 => x"74",
          1979 => x"c8",
          1980 => x"3f",
          1981 => x"ff",
          1982 => x"52",
          1983 => x"d0",
          1984 => x"d0",
          1985 => x"c7",
          1986 => x"d0",
          1987 => x"34",
          1988 => x"0d",
          1989 => x"84",
          1990 => x"84",
          1991 => x"05",
          1992 => x"a2",
          1993 => x"84",
          1994 => x"58",
          1995 => x"93",
          1996 => x"51",
          1997 => x"08",
          1998 => x"84",
          1999 => x"a5",
          2000 => x"05",
          2001 => x"81",
          2002 => x"ff",
          2003 => x"84",
          2004 => x"81",
          2005 => x"7b",
          2006 => x"70",
          2007 => x"84",
          2008 => x"74",
          2009 => x"c8",
          2010 => x"3f",
          2011 => x"ff",
          2012 => x"52",
          2013 => x"d0",
          2014 => x"d0",
          2015 => x"c7",
          2016 => x"83",
          2017 => x"fc",
          2018 => x"70",
          2019 => x"3f",
          2020 => x"f2",
          2021 => x"fc",
          2022 => x"80",
          2023 => x"52",
          2024 => x"f2",
          2025 => x"06",
          2026 => x"38",
          2027 => x"39",
          2028 => x"53",
          2029 => x"3f",
          2030 => x"82",
          2031 => x"51",
          2032 => x"d0",
          2033 => x"34",
          2034 => x"0d",
          2035 => x"e4",
          2036 => x"b8",
          2037 => x"e4",
          2038 => x"d0",
          2039 => x"82",
          2040 => x"5a",
          2041 => x"81",
          2042 => x"08",
          2043 => x"e4",
          2044 => x"08",
          2045 => x"08",
          2046 => x"77",
          2047 => x"d4",
          2048 => x"05",
          2049 => x"80",
          2050 => x"06",
          2051 => x"53",
          2052 => x"b8",
          2053 => x"33",
          2054 => x"70",
          2055 => x"81",
          2056 => x"93",
          2057 => x"ff",
          2058 => x"77",
          2059 => x"53",
          2060 => x"3f",
          2061 => x"81",
          2062 => x"80",
          2063 => x"34",
          2064 => x"f8",
          2065 => x"2b",
          2066 => x"81",
          2067 => x"d9",
          2068 => x"0c",
          2069 => x"83",
          2070 => x"41",
          2071 => x"9e",
          2072 => x"f7",
          2073 => x"c0",
          2074 => x"9b",
          2075 => x"39",
          2076 => x"33",
          2077 => x"5b",
          2078 => x"72",
          2079 => x"25",
          2080 => x"a8",
          2081 => x"a7",
          2082 => x"9f",
          2083 => x"75",
          2084 => x"95",
          2085 => x"f8",
          2086 => x"2b",
          2087 => x"7a",
          2088 => x"27",
          2089 => x"56",
          2090 => x"0c",
          2091 => x"27",
          2092 => x"97",
          2093 => x"55",
          2094 => x"74",
          2095 => x"53",
          2096 => x"86",
          2097 => x"33",
          2098 => x"33",
          2099 => x"41",
          2100 => x"0b",
          2101 => x"06",
          2102 => x"06",
          2103 => x"ff",
          2104 => x"58",
          2105 => x"87",
          2106 => x"79",
          2107 => x"7c",
          2108 => x"06",
          2109 => x"14",
          2110 => x"74",
          2111 => x"74",
          2112 => x"59",
          2113 => x"2e",
          2114 => x"72",
          2115 => x"70",
          2116 => x"33",
          2117 => x"39",
          2118 => x"b0",
          2119 => x"81",
          2120 => x"81",
          2121 => x"74",
          2122 => x"5e",
          2123 => x"73",
          2124 => x"71",
          2125 => x"80",
          2126 => x"f8",
          2127 => x"34",
          2128 => x"71",
          2129 => x"71",
          2130 => x"76",
          2131 => x"39",
          2132 => x"33",
          2133 => x"11",
          2134 => x"11",
          2135 => x"5b",
          2136 => x"70",
          2137 => x"ff",
          2138 => x"ff",
          2139 => x"ff",
          2140 => x"5e",
          2141 => x"57",
          2142 => x"31",
          2143 => x"7d",
          2144 => x"71",
          2145 => x"62",
          2146 => x"5f",
          2147 => x"85",
          2148 => x"31",
          2149 => x"fd",
          2150 => x"fd",
          2151 => x"31",
          2152 => x"3d",
          2153 => x"8a",
          2154 => x"34",
          2155 => x"55",
          2156 => x"34",
          2157 => x"34",
          2158 => x"54",
          2159 => x"80",
          2160 => x"d8",
          2161 => x"54",
          2162 => x"f8",
          2163 => x"72",
          2164 => x"06",
          2165 => x"34",
          2166 => x"06",
          2167 => x"81",
          2168 => x"88",
          2169 => x"0b",
          2170 => x"b8",
          2171 => x"b6",
          2172 => x"f7",
          2173 => x"84",
          2174 => x"33",
          2175 => x"26",
          2176 => x"83",
          2177 => x"72",
          2178 => x"11",
          2179 => x"59",
          2180 => x"ff",
          2181 => x"58",
          2182 => x"83",
          2183 => x"83",
          2184 => x"76",
          2185 => x"ff",
          2186 => x"82",
          2187 => x"f8",
          2188 => x"83",
          2189 => x"5c",
          2190 => x"38",
          2191 => x"54",
          2192 => x"ac",
          2193 => x"55",
          2194 => x"34",
          2195 => x"70",
          2196 => x"84",
          2197 => x"9f",
          2198 => x"33",
          2199 => x"0b",
          2200 => x"81",
          2201 => x"9f",
          2202 => x"33",
          2203 => x"23",
          2204 => x"83",
          2205 => x"26",
          2206 => x"05",
          2207 => x"58",
          2208 => x"80",
          2209 => x"ff",
          2210 => x"29",
          2211 => x"27",
          2212 => x"e0",
          2213 => x"13",
          2214 => x"73",
          2215 => x"81",
          2216 => x"d8",
          2217 => x"29",
          2218 => x"26",
          2219 => x"e4",
          2220 => x"f8",
          2221 => x"83",
          2222 => x"5c",
          2223 => x"38",
          2224 => x"81",
          2225 => x"33",
          2226 => x"06",
          2227 => x"05",
          2228 => x"78",
          2229 => x"73",
          2230 => x"90",
          2231 => x"31",
          2232 => x"16",
          2233 => x"34",
          2234 => x"8a",
          2235 => x"75",
          2236 => x"13",
          2237 => x"80",
          2238 => x"fe",
          2239 => x"59",
          2240 => x"84",
          2241 => x"fc",
          2242 => x"05",
          2243 => x"38",
          2244 => x"51",
          2245 => x"51",
          2246 => x"f8",
          2247 => x"0c",
          2248 => x"f8",
          2249 => x"81",
          2250 => x"e2",
          2251 => x"94",
          2252 => x"86",
          2253 => x"70",
          2254 => x"72",
          2255 => x"f8",
          2256 => x"33",
          2257 => x"11",
          2258 => x"38",
          2259 => x"80",
          2260 => x"0d",
          2261 => x"31",
          2262 => x"54",
          2263 => x"34",
          2264 => x"3d",
          2265 => x"05",
          2266 => x"55",
          2267 => x"53",
          2268 => x"84",
          2269 => x"80",
          2270 => x"94",
          2271 => x"56",
          2272 => x"81",
          2273 => x"fe",
          2274 => x"05",
          2275 => x"70",
          2276 => x"70",
          2277 => x"80",
          2278 => x"06",
          2279 => x"53",
          2280 => x"06",
          2281 => x"90",
          2282 => x"83",
          2283 => x"81",
          2284 => x"f8",
          2285 => x"0c",
          2286 => x"33",
          2287 => x"90",
          2288 => x"81",
          2289 => x"f8",
          2290 => x"83",
          2291 => x"e4",
          2292 => x"90",
          2293 => x"70",
          2294 => x"83",
          2295 => x"83",
          2296 => x"f8",
          2297 => x"51",
          2298 => x"39",
          2299 => x"83",
          2300 => x"ff",
          2301 => x"f9",
          2302 => x"90",
          2303 => x"33",
          2304 => x"90",
          2305 => x"33",
          2306 => x"70",
          2307 => x"83",
          2308 => x"07",
          2309 => x"ba",
          2310 => x"06",
          2311 => x"90",
          2312 => x"33",
          2313 => x"70",
          2314 => x"83",
          2315 => x"07",
          2316 => x"82",
          2317 => x"06",
          2318 => x"f2",
          2319 => x"06",
          2320 => x"34",
          2321 => x"bf",
          2322 => x"05",
          2323 => x"93",
          2324 => x"da",
          2325 => x"78",
          2326 => x"24",
          2327 => x"38",
          2328 => x"84",
          2329 => x"34",
          2330 => x"f8",
          2331 => x"83",
          2332 => x"0b",
          2333 => x"b6",
          2334 => x"34",
          2335 => x"0b",
          2336 => x"b6",
          2337 => x"56",
          2338 => x"7c",
          2339 => x"ff",
          2340 => x"34",
          2341 => x"83",
          2342 => x"23",
          2343 => x"0d",
          2344 => x"81",
          2345 => x"83",
          2346 => x"95",
          2347 => x"84",
          2348 => x"33",
          2349 => x"55",
          2350 => x"e2",
          2351 => x"0b",
          2352 => x"79",
          2353 => x"b8",
          2354 => x"8c",
          2355 => x"70",
          2356 => x"52",
          2357 => x"83",
          2358 => x"7d",
          2359 => x"b6",
          2360 => x"7b",
          2361 => x"95",
          2362 => x"84",
          2363 => x"dc",
          2364 => x"a8",
          2365 => x"83",
          2366 => x"ff",
          2367 => x"52",
          2368 => x"3f",
          2369 => x"92",
          2370 => x"27",
          2371 => x"33",
          2372 => x"e0",
          2373 => x"5a",
          2374 => x"02",
          2375 => x"d8",
          2376 => x"94",
          2377 => x"a0",
          2378 => x"51",
          2379 => x"83",
          2380 => x"52",
          2381 => x"2e",
          2382 => x"f9",
          2383 => x"75",
          2384 => x"2e",
          2385 => x"83",
          2386 => x"72",
          2387 => x"b6",
          2388 => x"14",
          2389 => x"95",
          2390 => x"29",
          2391 => x"f8",
          2392 => x"73",
          2393 => x"90",
          2394 => x"84",
          2395 => x"83",
          2396 => x"72",
          2397 => x"57",
          2398 => x"14",
          2399 => x"59",
          2400 => x"84",
          2401 => x"38",
          2402 => x"34",
          2403 => x"2e",
          2404 => x"76",
          2405 => x"84",
          2406 => x"75",
          2407 => x"80",
          2408 => x"06",
          2409 => x"f1",
          2410 => x"34",
          2411 => x"33",
          2412 => x"34",
          2413 => x"89",
          2414 => x"fd",
          2415 => x"06",
          2416 => x"38",
          2417 => x"81",
          2418 => x"83",
          2419 => x"74",
          2420 => x"75",
          2421 => x"0b",
          2422 => x"04",
          2423 => x"fd",
          2424 => x"81",
          2425 => x"83",
          2426 => x"34",
          2427 => x"83",
          2428 => x"55",
          2429 => x"73",
          2430 => x"a0",
          2431 => x"81",
          2432 => x"90",
          2433 => x"3f",
          2434 => x"80",
          2435 => x"57",
          2436 => x"75",
          2437 => x"2e",
          2438 => x"d1",
          2439 => x"78",
          2440 => x"d8",
          2441 => x"95",
          2442 => x"5c",
          2443 => x"a0",
          2444 => x"83",
          2445 => x"72",
          2446 => x"78",
          2447 => x"94",
          2448 => x"5a",
          2449 => x"b0",
          2450 => x"70",
          2451 => x"83",
          2452 => x"42",
          2453 => x"33",
          2454 => x"70",
          2455 => x"26",
          2456 => x"5a",
          2457 => x"75",
          2458 => x"b8",
          2459 => x"b7",
          2460 => x"81",
          2461 => x"38",
          2462 => x"80",
          2463 => x"d8",
          2464 => x"95",
          2465 => x"40",
          2466 => x"a0",
          2467 => x"83",
          2468 => x"72",
          2469 => x"78",
          2470 => x"94",
          2471 => x"83",
          2472 => x"1b",
          2473 => x"ff",
          2474 => x"95",
          2475 => x"43",
          2476 => x"84",
          2477 => x"77",
          2478 => x"fe",
          2479 => x"80",
          2480 => x"0d",
          2481 => x"78",
          2482 => x"2e",
          2483 => x"0b",
          2484 => x"b8",
          2485 => x"9b",
          2486 => x"75",
          2487 => x"e4",
          2488 => x"b7",
          2489 => x"34",
          2490 => x"84",
          2491 => x"b8",
          2492 => x"9b",
          2493 => x"b7",
          2494 => x"f8",
          2495 => x"72",
          2496 => x"e0",
          2497 => x"34",
          2498 => x"33",
          2499 => x"12",
          2500 => x"96",
          2501 => x"71",
          2502 => x"33",
          2503 => x"b6",
          2504 => x"f8",
          2505 => x"72",
          2506 => x"83",
          2507 => x"05",
          2508 => x"81",
          2509 => x"0b",
          2510 => x"84",
          2511 => x"70",
          2512 => x"73",
          2513 => x"05",
          2514 => x"72",
          2515 => x"06",
          2516 => x"5a",
          2517 => x"78",
          2518 => x"76",
          2519 => x"f8",
          2520 => x"84",
          2521 => x"e5",
          2522 => x"80",
          2523 => x"84",
          2524 => x"e4",
          2525 => x"94",
          2526 => x"95",
          2527 => x"93",
          2528 => x"84",
          2529 => x"e4",
          2530 => x"ff",
          2531 => x"83",
          2532 => x"70",
          2533 => x"70",
          2534 => x"86",
          2535 => x"22",
          2536 => x"83",
          2537 => x"44",
          2538 => x"81",
          2539 => x"06",
          2540 => x"75",
          2541 => x"81",
          2542 => x"81",
          2543 => x"40",
          2544 => x"a0",
          2545 => x"83",
          2546 => x"72",
          2547 => x"a0",
          2548 => x"f8",
          2549 => x"5a",
          2550 => x"b0",
          2551 => x"70",
          2552 => x"83",
          2553 => x"43",
          2554 => x"33",
          2555 => x"1a",
          2556 => x"7b",
          2557 => x"33",
          2558 => x"58",
          2559 => x"95",
          2560 => x"05",
          2561 => x"95",
          2562 => x"38",
          2563 => x"b7",
          2564 => x"ff",
          2565 => x"c8",
          2566 => x"05",
          2567 => x"f8",
          2568 => x"9f",
          2569 => x"9c",
          2570 => x"84",
          2571 => x"83",
          2572 => x"72",
          2573 => x"05",
          2574 => x"7b",
          2575 => x"83",
          2576 => x"59",
          2577 => x"38",
          2578 => x"81",
          2579 => x"72",
          2580 => x"80",
          2581 => x"84",
          2582 => x"83",
          2583 => x"5e",
          2584 => x"96",
          2585 => x"71",
          2586 => x"33",
          2587 => x"b6",
          2588 => x"f8",
          2589 => x"72",
          2590 => x"83",
          2591 => x"34",
          2592 => x"5b",
          2593 => x"84",
          2594 => x"38",
          2595 => x"34",
          2596 => x"59",
          2597 => x"f8",
          2598 => x"f8",
          2599 => x"81",
          2600 => x"72",
          2601 => x"5b",
          2602 => x"80",
          2603 => x"f8",
          2604 => x"71",
          2605 => x"0b",
          2606 => x"94",
          2607 => x"83",
          2608 => x"1a",
          2609 => x"ff",
          2610 => x"95",
          2611 => x"5a",
          2612 => x"97",
          2613 => x"81",
          2614 => x"fe",
          2615 => x"fe",
          2616 => x"0c",
          2617 => x"3d",
          2618 => x"59",
          2619 => x"83",
          2620 => x"58",
          2621 => x"0b",
          2622 => x"b8",
          2623 => x"f8",
          2624 => x"1b",
          2625 => x"84",
          2626 => x"5b",
          2627 => x"84",
          2628 => x"53",
          2629 => x"84",
          2630 => x"38",
          2631 => x"5a",
          2632 => x"83",
          2633 => x"22",
          2634 => x"cf",
          2635 => x"84",
          2636 => x"f8",
          2637 => x"f8",
          2638 => x"39",
          2639 => x"33",
          2640 => x"05",
          2641 => x"33",
          2642 => x"84",
          2643 => x"83",
          2644 => x"5a",
          2645 => x"18",
          2646 => x"29",
          2647 => x"60",
          2648 => x"b6",
          2649 => x"f8",
          2650 => x"72",
          2651 => x"83",
          2652 => x"34",
          2653 => x"58",
          2654 => x"b6",
          2655 => x"ff",
          2656 => x"80",
          2657 => x"db",
          2658 => x"38",
          2659 => x"b4",
          2660 => x"3f",
          2661 => x"3d",
          2662 => x"f8",
          2663 => x"f8",
          2664 => x"76",
          2665 => x"83",
          2666 => x"83",
          2667 => x"83",
          2668 => x"ff",
          2669 => x"7a",
          2670 => x"b8",
          2671 => x"06",
          2672 => x"81",
          2673 => x"05",
          2674 => x"94",
          2675 => x"3f",
          2676 => x"b8",
          2677 => x"e8",
          2678 => x"24",
          2679 => x"c8",
          2680 => x"39",
          2681 => x"58",
          2682 => x"27",
          2683 => x"b8",
          2684 => x"b1",
          2685 => x"83",
          2686 => x"84",
          2687 => x"8f",
          2688 => x"b8",
          2689 => x"70",
          2690 => x"5e",
          2691 => x"e7",
          2692 => x"80",
          2693 => x"33",
          2694 => x"b6",
          2695 => x"27",
          2696 => x"34",
          2697 => x"95",
          2698 => x"ff",
          2699 => x"a7",
          2700 => x"94",
          2701 => x"f8",
          2702 => x"b6",
          2703 => x"76",
          2704 => x"75",
          2705 => x"84",
          2706 => x"8d",
          2707 => x"b8",
          2708 => x"70",
          2709 => x"42",
          2710 => x"cf",
          2711 => x"80",
          2712 => x"22",
          2713 => x"fc",
          2714 => x"f8",
          2715 => x"71",
          2716 => x"83",
          2717 => x"71",
          2718 => x"06",
          2719 => x"80",
          2720 => x"82",
          2721 => x"83",
          2722 => x"b7",
          2723 => x"e7",
          2724 => x"99",
          2725 => x"81",
          2726 => x"39",
          2727 => x"2e",
          2728 => x"83",
          2729 => x"b6",
          2730 => x"75",
          2731 => x"83",
          2732 => x"b7",
          2733 => x"c8",
          2734 => x"94",
          2735 => x"33",
          2736 => x"25",
          2737 => x"94",
          2738 => x"51",
          2739 => x"b7",
          2740 => x"8b",
          2741 => x"05",
          2742 => x"51",
          2743 => x"81",
          2744 => x"58",
          2745 => x"e5",
          2746 => x"38",
          2747 => x"26",
          2748 => x"81",
          2749 => x"97",
          2750 => x"77",
          2751 => x"33",
          2752 => x"b8",
          2753 => x"06",
          2754 => x"06",
          2755 => x"5c",
          2756 => x"5a",
          2757 => x"ff",
          2758 => x"27",
          2759 => x"94",
          2760 => x"57",
          2761 => x"7a",
          2762 => x"af",
          2763 => x"80",
          2764 => x"33",
          2765 => x"7f",
          2766 => x"33",
          2767 => x"06",
          2768 => x"11",
          2769 => x"92",
          2770 => x"70",
          2771 => x"33",
          2772 => x"81",
          2773 => x"ff",
          2774 => x"7c",
          2775 => x"33",
          2776 => x"ff",
          2777 => x"7c",
          2778 => x"57",
          2779 => x"b6",
          2780 => x"ee",
          2781 => x"94",
          2782 => x"92",
          2783 => x"26",
          2784 => x"7e",
          2785 => x"5e",
          2786 => x"5b",
          2787 => x"06",
          2788 => x"1d",
          2789 => x"f7",
          2790 => x"e0",
          2791 => x"1f",
          2792 => x"76",
          2793 => x"81",
          2794 => x"d8",
          2795 => x"29",
          2796 => x"27",
          2797 => x"5f",
          2798 => x"81",
          2799 => x"58",
          2800 => x"81",
          2801 => x"d7",
          2802 => x"5e",
          2803 => x"f6",
          2804 => x"75",
          2805 => x"84",
          2806 => x"f6",
          2807 => x"33",
          2808 => x"59",
          2809 => x"84",
          2810 => x"09",
          2811 => x"95",
          2812 => x"f8",
          2813 => x"ff",
          2814 => x"33",
          2815 => x"7e",
          2816 => x"f5",
          2817 => x"27",
          2818 => x"10",
          2819 => x"86",
          2820 => x"5a",
          2821 => x"06",
          2822 => x"79",
          2823 => x"83",
          2824 => x"90",
          2825 => x"07",
          2826 => x"7a",
          2827 => x"05",
          2828 => x"58",
          2829 => x"b6",
          2830 => x"5f",
          2831 => x"06",
          2832 => x"64",
          2833 => x"26",
          2834 => x"7b",
          2835 => x"1d",
          2836 => x"38",
          2837 => x"18",
          2838 => x"34",
          2839 => x"81",
          2840 => x"38",
          2841 => x"78",
          2842 => x"57",
          2843 => x"39",
          2844 => x"58",
          2845 => x"70",
          2846 => x"f0",
          2847 => x"57",
          2848 => x"be",
          2849 => x"34",
          2850 => x"56",
          2851 => x"33",
          2852 => x"34",
          2853 => x"33",
          2854 => x"33",
          2855 => x"83",
          2856 => x"83",
          2857 => x"ff",
          2858 => x"f8",
          2859 => x"56",
          2860 => x"83",
          2861 => x"07",
          2862 => x"39",
          2863 => x"81",
          2864 => x"c3",
          2865 => x"06",
          2866 => x"34",
          2867 => x"f8",
          2868 => x"06",
          2869 => x"90",
          2870 => x"f8",
          2871 => x"90",
          2872 => x"75",
          2873 => x"83",
          2874 => x"e0",
          2875 => x"fe",
          2876 => x"cf",
          2877 => x"f8",
          2878 => x"90",
          2879 => x"75",
          2880 => x"83",
          2881 => x"07",
          2882 => x"b3",
          2883 => x"06",
          2884 => x"34",
          2885 => x"81",
          2886 => x"f8",
          2887 => x"90",
          2888 => x"f8",
          2889 => x"90",
          2890 => x"f8",
          2891 => x"90",
          2892 => x"f8",
          2893 => x"90",
          2894 => x"56",
          2895 => x"39",
          2896 => x"b0",
          2897 => x"fd",
          2898 => x"34",
          2899 => x"ec",
          2900 => x"f8",
          2901 => x"f8",
          2902 => x"78",
          2903 => x"b7",
          2904 => x"84",
          2905 => x"e4",
          2906 => x"f8",
          2907 => x"81",
          2908 => x"cf",
          2909 => x"dc",
          2910 => x"8e",
          2911 => x"84",
          2912 => x"80",
          2913 => x"84",
          2914 => x"77",
          2915 => x"84",
          2916 => x"7a",
          2917 => x"fe",
          2918 => x"84",
          2919 => x"b7",
          2920 => x"f8",
          2921 => x"97",
          2922 => x"ff",
          2923 => x"39",
          2924 => x"52",
          2925 => x"39",
          2926 => x"8f",
          2927 => x"70",
          2928 => x"5f",
          2929 => x"51",
          2930 => x"75",
          2931 => x"f8",
          2932 => x"94",
          2933 => x"2c",
          2934 => x"39",
          2935 => x"b6",
          2936 => x"75",
          2937 => x"f3",
          2938 => x"81",
          2939 => x"ee",
          2940 => x"b6",
          2941 => x"f8",
          2942 => x"a7",
          2943 => x"5f",
          2944 => x"ff",
          2945 => x"5b",
          2946 => x"81",
          2947 => x"ff",
          2948 => x"89",
          2949 => x"76",
          2950 => x"75",
          2951 => x"06",
          2952 => x"83",
          2953 => x"76",
          2954 => x"56",
          2955 => x"ff",
          2956 => x"80",
          2957 => x"77",
          2958 => x"71",
          2959 => x"86",
          2960 => x"80",
          2961 => x"06",
          2962 => x"5d",
          2963 => x"97",
          2964 => x"5e",
          2965 => x"81",
          2966 => x"58",
          2967 => x"81",
          2968 => x"d7",
          2969 => x"5d",
          2970 => x"e0",
          2971 => x"1e",
          2972 => x"76",
          2973 => x"81",
          2974 => x"d8",
          2975 => x"29",
          2976 => x"26",
          2977 => x"f8",
          2978 => x"1c",
          2979 => x"84",
          2980 => x"84",
          2981 => x"fd",
          2982 => x"b6",
          2983 => x"11",
          2984 => x"38",
          2985 => x"77",
          2986 => x"80",
          2987 => x"83",
          2988 => x"70",
          2989 => x"56",
          2990 => x"56",
          2991 => x"39",
          2992 => x"b6",
          2993 => x"75",
          2994 => x"ef",
          2995 => x"06",
          2996 => x"70",
          2997 => x"7a",
          2998 => x"09",
          2999 => x"39",
          3000 => x"34",
          3001 => x"83",
          3002 => x"7b",
          3003 => x"f2",
          3004 => x"7a",
          3005 => x"81",
          3006 => x"77",
          3007 => x"26",
          3008 => x"05",
          3009 => x"70",
          3010 => x"d4",
          3011 => x"56",
          3012 => x"39",
          3013 => x"ad",
          3014 => x"84",
          3015 => x"f1",
          3016 => x"34",
          3017 => x"33",
          3018 => x"34",
          3019 => x"a7",
          3020 => x"33",
          3021 => x"80",
          3022 => x"3f",
          3023 => x"3d",
          3024 => x"ab",
          3025 => x"85",
          3026 => x"bf",
          3027 => x"e8",
          3028 => x"c8",
          3029 => x"80",
          3030 => x"75",
          3031 => x"84",
          3032 => x"83",
          3033 => x"80",
          3034 => x"30",
          3035 => x"56",
          3036 => x"0c",
          3037 => x"09",
          3038 => x"83",
          3039 => x"07",
          3040 => x"c4",
          3041 => x"95",
          3042 => x"29",
          3043 => x"f8",
          3044 => x"29",
          3045 => x"f6",
          3046 => x"81",
          3047 => x"73",
          3048 => x"87",
          3049 => x"88",
          3050 => x"86",
          3051 => x"f4",
          3052 => x"ff",
          3053 => x"cf",
          3054 => x"33",
          3055 => x"16",
          3056 => x"85",
          3057 => x"b4",
          3058 => x"75",
          3059 => x"2e",
          3060 => x"15",
          3061 => x"f6",
          3062 => x"ff",
          3063 => x"b3",
          3064 => x"2b",
          3065 => x"83",
          3066 => x"70",
          3067 => x"51",
          3068 => x"38",
          3069 => x"09",
          3070 => x"e4",
          3071 => x"80",
          3072 => x"c4",
          3073 => x"f6",
          3074 => x"5d",
          3075 => x"98",
          3076 => x"8d",
          3077 => x"73",
          3078 => x"a2",
          3079 => x"8b",
          3080 => x"73",
          3081 => x"54",
          3082 => x"f6",
          3083 => x"81",
          3084 => x"72",
          3085 => x"f6",
          3086 => x"84",
          3087 => x"e8",
          3088 => x"54",
          3089 => x"0b",
          3090 => x"b8",
          3091 => x"06",
          3092 => x"38",
          3093 => x"f6",
          3094 => x"9c",
          3095 => x"83",
          3096 => x"83",
          3097 => x"91",
          3098 => x"9c",
          3099 => x"dc",
          3100 => x"54",
          3101 => x"54",
          3102 => x"98",
          3103 => x"81",
          3104 => x"38",
          3105 => x"b6",
          3106 => x"54",
          3107 => x"53",
          3108 => x"81",
          3109 => x"34",
          3110 => x"58",
          3111 => x"83",
          3112 => x"77",
          3113 => x"7d",
          3114 => x"2e",
          3115 => x"59",
          3116 => x"54",
          3117 => x"2e",
          3118 => x"06",
          3119 => x"27",
          3120 => x"54",
          3121 => x"10",
          3122 => x"2b",
          3123 => x"33",
          3124 => x"9c",
          3125 => x"ea",
          3126 => x"a8",
          3127 => x"a0",
          3128 => x"ff",
          3129 => x"b6",
          3130 => x"83",
          3131 => x"70",
          3132 => x"7d",
          3133 => x"06",
          3134 => x"c6",
          3135 => x"83",
          3136 => x"78",
          3137 => x"70",
          3138 => x"27",
          3139 => x"72",
          3140 => x"dc",
          3141 => x"81",
          3142 => x"3f",
          3143 => x"0d",
          3144 => x"f9",
          3145 => x"38",
          3146 => x"5b",
          3147 => x"c9",
          3148 => x"34",
          3149 => x"ff",
          3150 => x"b1",
          3151 => x"81",
          3152 => x"ac",
          3153 => x"8a",
          3154 => x"81",
          3155 => x"83",
          3156 => x"c0",
          3157 => x"27",
          3158 => x"08",
          3159 => x"06",
          3160 => x"f6",
          3161 => x"83",
          3162 => x"53",
          3163 => x"be",
          3164 => x"83",
          3165 => x"70",
          3166 => x"33",
          3167 => x"fa",
          3168 => x"06",
          3169 => x"2e",
          3170 => x"81",
          3171 => x"ef",
          3172 => x"39",
          3173 => x"54",
          3174 => x"b6",
          3175 => x"80",
          3176 => x"76",
          3177 => x"da",
          3178 => x"53",
          3179 => x"83",
          3180 => x"f6",
          3181 => x"81",
          3182 => x"80",
          3183 => x"83",
          3184 => x"ff",
          3185 => x"38",
          3186 => x"84",
          3187 => x"56",
          3188 => x"38",
          3189 => x"ff",
          3190 => x"51",
          3191 => x"aa",
          3192 => x"14",
          3193 => x"de",
          3194 => x"34",
          3195 => x"39",
          3196 => x"3f",
          3197 => x"80",
          3198 => x"02",
          3199 => x"f2",
          3200 => x"85",
          3201 => x"fe",
          3202 => x"f0",
          3203 => x"08",
          3204 => x"90",
          3205 => x"52",
          3206 => x"72",
          3207 => x"c0",
          3208 => x"27",
          3209 => x"38",
          3210 => x"55",
          3211 => x"55",
          3212 => x"c0",
          3213 => x"53",
          3214 => x"c0",
          3215 => x"f6",
          3216 => x"9c",
          3217 => x"38",
          3218 => x"c0",
          3219 => x"83",
          3220 => x"70",
          3221 => x"2e",
          3222 => x"71",
          3223 => x"38",
          3224 => x"0d",
          3225 => x"88",
          3226 => x"02",
          3227 => x"80",
          3228 => x"2b",
          3229 => x"98",
          3230 => x"83",
          3231 => x"84",
          3232 => x"85",
          3233 => x"f2",
          3234 => x"83",
          3235 => x"34",
          3236 => x"56",
          3237 => x"86",
          3238 => x"9c",
          3239 => x"ce",
          3240 => x"08",
          3241 => x"70",
          3242 => x"87",
          3243 => x"73",
          3244 => x"db",
          3245 => x"ff",
          3246 => x"71",
          3247 => x"87",
          3248 => x"05",
          3249 => x"87",
          3250 => x"2e",
          3251 => x"98",
          3252 => x"87",
          3253 => x"87",
          3254 => x"26",
          3255 => x"16",
          3256 => x"80",
          3257 => x"06",
          3258 => x"70",
          3259 => x"80",
          3260 => x"52",
          3261 => x"70",
          3262 => x"05",
          3263 => x"76",
          3264 => x"04",
          3265 => x"3d",
          3266 => x"3d",
          3267 => x"33",
          3268 => x"08",
          3269 => x"06",
          3270 => x"55",
          3271 => x"2a",
          3272 => x"2a",
          3273 => x"15",
          3274 => x"c6",
          3275 => x"51",
          3276 => x"81",
          3277 => x"54",
          3278 => x"f2",
          3279 => x"83",
          3280 => x"34",
          3281 => x"56",
          3282 => x"86",
          3283 => x"9c",
          3284 => x"ce",
          3285 => x"08",
          3286 => x"70",
          3287 => x"87",
          3288 => x"73",
          3289 => x"db",
          3290 => x"ff",
          3291 => x"71",
          3292 => x"87",
          3293 => x"05",
          3294 => x"87",
          3295 => x"2e",
          3296 => x"98",
          3297 => x"87",
          3298 => x"87",
          3299 => x"26",
          3300 => x"16",
          3301 => x"80",
          3302 => x"52",
          3303 => x"81",
          3304 => x"38",
          3305 => x"88",
          3306 => x"fb",
          3307 => x"80",
          3308 => x"f0",
          3309 => x"34",
          3310 => x"87",
          3311 => x"08",
          3312 => x"c0",
          3313 => x"9c",
          3314 => x"81",
          3315 => x"52",
          3316 => x"81",
          3317 => x"a4",
          3318 => x"80",
          3319 => x"80",
          3320 => x"80",
          3321 => x"9c",
          3322 => x"51",
          3323 => x"33",
          3324 => x"73",
          3325 => x"2e",
          3326 => x"51",
          3327 => x"71",
          3328 => x"57",
          3329 => x"81",
          3330 => x"ff",
          3331 => x"51",
          3332 => x"04",
          3333 => x"7a",
          3334 => x"ff",
          3335 => x"33",
          3336 => x"83",
          3337 => x"12",
          3338 => x"07",
          3339 => x"59",
          3340 => x"81",
          3341 => x"83",
          3342 => x"2b",
          3343 => x"33",
          3344 => x"57",
          3345 => x"71",
          3346 => x"85",
          3347 => x"2b",
          3348 => x"54",
          3349 => x"81",
          3350 => x"84",
          3351 => x"33",
          3352 => x"70",
          3353 => x"77",
          3354 => x"84",
          3355 => x"86",
          3356 => x"84",
          3357 => x"34",
          3358 => x"08",
          3359 => x"88",
          3360 => x"88",
          3361 => x"34",
          3362 => x"04",
          3363 => x"8b",
          3364 => x"84",
          3365 => x"2b",
          3366 => x"51",
          3367 => x"72",
          3368 => x"70",
          3369 => x"71",
          3370 => x"5a",
          3371 => x"87",
          3372 => x"88",
          3373 => x"13",
          3374 => x"d4",
          3375 => x"71",
          3376 => x"70",
          3377 => x"72",
          3378 => x"d4",
          3379 => x"33",
          3380 => x"74",
          3381 => x"88",
          3382 => x"f8",
          3383 => x"52",
          3384 => x"77",
          3385 => x"84",
          3386 => x"81",
          3387 => x"2b",
          3388 => x"33",
          3389 => x"06",
          3390 => x"5a",
          3391 => x"81",
          3392 => x"17",
          3393 => x"8b",
          3394 => x"70",
          3395 => x"71",
          3396 => x"5a",
          3397 => x"e4",
          3398 => x"88",
          3399 => x"88",
          3400 => x"77",
          3401 => x"70",
          3402 => x"8b",
          3403 => x"82",
          3404 => x"2b",
          3405 => x"52",
          3406 => x"34",
          3407 => x"04",
          3408 => x"08",
          3409 => x"77",
          3410 => x"90",
          3411 => x"f4",
          3412 => x"0b",
          3413 => x"53",
          3414 => x"d3",
          3415 => x"76",
          3416 => x"84",
          3417 => x"34",
          3418 => x"d4",
          3419 => x"0b",
          3420 => x"84",
          3421 => x"80",
          3422 => x"88",
          3423 => x"17",
          3424 => x"d0",
          3425 => x"d4",
          3426 => x"82",
          3427 => x"fe",
          3428 => x"80",
          3429 => x"38",
          3430 => x"83",
          3431 => x"ff",
          3432 => x"11",
          3433 => x"07",
          3434 => x"ff",
          3435 => x"38",
          3436 => x"81",
          3437 => x"81",
          3438 => x"ff",
          3439 => x"5c",
          3440 => x"38",
          3441 => x"55",
          3442 => x"71",
          3443 => x"38",
          3444 => x"77",
          3445 => x"78",
          3446 => x"88",
          3447 => x"56",
          3448 => x"2e",
          3449 => x"73",
          3450 => x"80",
          3451 => x"82",
          3452 => x"78",
          3453 => x"88",
          3454 => x"74",
          3455 => x"d4",
          3456 => x"71",
          3457 => x"84",
          3458 => x"81",
          3459 => x"83",
          3460 => x"7e",
          3461 => x"5c",
          3462 => x"82",
          3463 => x"72",
          3464 => x"18",
          3465 => x"34",
          3466 => x"11",
          3467 => x"71",
          3468 => x"5c",
          3469 => x"85",
          3470 => x"16",
          3471 => x"12",
          3472 => x"2a",
          3473 => x"34",
          3474 => x"08",
          3475 => x"33",
          3476 => x"74",
          3477 => x"86",
          3478 => x"b8",
          3479 => x"84",
          3480 => x"2b",
          3481 => x"59",
          3482 => x"34",
          3483 => x"51",
          3484 => x"0d",
          3485 => x"71",
          3486 => x"05",
          3487 => x"88",
          3488 => x"59",
          3489 => x"76",
          3490 => x"70",
          3491 => x"71",
          3492 => x"05",
          3493 => x"88",
          3494 => x"5f",
          3495 => x"1a",
          3496 => x"d4",
          3497 => x"71",
          3498 => x"70",
          3499 => x"77",
          3500 => x"d4",
          3501 => x"39",
          3502 => x"08",
          3503 => x"77",
          3504 => x"e4",
          3505 => x"fb",
          3506 => x"b8",
          3507 => x"ff",
          3508 => x"80",
          3509 => x"80",
          3510 => x"fe",
          3511 => x"55",
          3512 => x"34",
          3513 => x"15",
          3514 => x"b8",
          3515 => x"81",
          3516 => x"08",
          3517 => x"80",
          3518 => x"70",
          3519 => x"88",
          3520 => x"b8",
          3521 => x"b8",
          3522 => x"76",
          3523 => x"34",
          3524 => x"38",
          3525 => x"67",
          3526 => x"08",
          3527 => x"aa",
          3528 => x"7f",
          3529 => x"84",
          3530 => x"83",
          3531 => x"06",
          3532 => x"7f",
          3533 => x"ff",
          3534 => x"33",
          3535 => x"70",
          3536 => x"70",
          3537 => x"2b",
          3538 => x"71",
          3539 => x"90",
          3540 => x"54",
          3541 => x"5f",
          3542 => x"82",
          3543 => x"2b",
          3544 => x"33",
          3545 => x"90",
          3546 => x"56",
          3547 => x"62",
          3548 => x"77",
          3549 => x"2e",
          3550 => x"62",
          3551 => x"61",
          3552 => x"70",
          3553 => x"71",
          3554 => x"81",
          3555 => x"2b",
          3556 => x"5b",
          3557 => x"76",
          3558 => x"71",
          3559 => x"11",
          3560 => x"8b",
          3561 => x"84",
          3562 => x"2b",
          3563 => x"52",
          3564 => x"77",
          3565 => x"84",
          3566 => x"33",
          3567 => x"83",
          3568 => x"87",
          3569 => x"88",
          3570 => x"41",
          3571 => x"16",
          3572 => x"33",
          3573 => x"81",
          3574 => x"5c",
          3575 => x"1a",
          3576 => x"82",
          3577 => x"2b",
          3578 => x"33",
          3579 => x"70",
          3580 => x"5a",
          3581 => x"1a",
          3582 => x"70",
          3583 => x"71",
          3584 => x"33",
          3585 => x"70",
          3586 => x"5a",
          3587 => x"83",
          3588 => x"1f",
          3589 => x"88",
          3590 => x"83",
          3591 => x"84",
          3592 => x"b8",
          3593 => x"05",
          3594 => x"44",
          3595 => x"7e",
          3596 => x"3d",
          3597 => x"b8",
          3598 => x"d0",
          3599 => x"84",
          3600 => x"84",
          3601 => x"81",
          3602 => x"08",
          3603 => x"85",
          3604 => x"60",
          3605 => x"34",
          3606 => x"22",
          3607 => x"83",
          3608 => x"5a",
          3609 => x"89",
          3610 => x"10",
          3611 => x"f8",
          3612 => x"81",
          3613 => x"08",
          3614 => x"2e",
          3615 => x"2e",
          3616 => x"3f",
          3617 => x"0c",
          3618 => x"b8",
          3619 => x"5e",
          3620 => x"33",
          3621 => x"06",
          3622 => x"40",
          3623 => x"61",
          3624 => x"2a",
          3625 => x"83",
          3626 => x"1f",
          3627 => x"2b",
          3628 => x"06",
          3629 => x"70",
          3630 => x"5b",
          3631 => x"81",
          3632 => x"34",
          3633 => x"7b",
          3634 => x"b8",
          3635 => x"88",
          3636 => x"75",
          3637 => x"54",
          3638 => x"06",
          3639 => x"82",
          3640 => x"2b",
          3641 => x"33",
          3642 => x"90",
          3643 => x"58",
          3644 => x"38",
          3645 => x"83",
          3646 => x"77",
          3647 => x"27",
          3648 => x"ff",
          3649 => x"80",
          3650 => x"80",
          3651 => x"fe",
          3652 => x"5a",
          3653 => x"34",
          3654 => x"1a",
          3655 => x"b8",
          3656 => x"81",
          3657 => x"08",
          3658 => x"80",
          3659 => x"70",
          3660 => x"64",
          3661 => x"34",
          3662 => x"10",
          3663 => x"42",
          3664 => x"61",
          3665 => x"7a",
          3666 => x"ff",
          3667 => x"38",
          3668 => x"bd",
          3669 => x"54",
          3670 => x"0d",
          3671 => x"12",
          3672 => x"07",
          3673 => x"33",
          3674 => x"7e",
          3675 => x"71",
          3676 => x"44",
          3677 => x"45",
          3678 => x"64",
          3679 => x"70",
          3680 => x"71",
          3681 => x"05",
          3682 => x"88",
          3683 => x"42",
          3684 => x"86",
          3685 => x"84",
          3686 => x"12",
          3687 => x"ff",
          3688 => x"5d",
          3689 => x"84",
          3690 => x"33",
          3691 => x"83",
          3692 => x"15",
          3693 => x"2a",
          3694 => x"54",
          3695 => x"84",
          3696 => x"81",
          3697 => x"2b",
          3698 => x"15",
          3699 => x"2a",
          3700 => x"55",
          3701 => x"34",
          3702 => x"11",
          3703 => x"07",
          3704 => x"42",
          3705 => x"51",
          3706 => x"08",
          3707 => x"06",
          3708 => x"f4",
          3709 => x"0b",
          3710 => x"53",
          3711 => x"c0",
          3712 => x"7f",
          3713 => x"84",
          3714 => x"34",
          3715 => x"d4",
          3716 => x"0b",
          3717 => x"84",
          3718 => x"80",
          3719 => x"88",
          3720 => x"1f",
          3721 => x"d0",
          3722 => x"d4",
          3723 => x"82",
          3724 => x"7e",
          3725 => x"c0",
          3726 => x"71",
          3727 => x"05",
          3728 => x"88",
          3729 => x"5e",
          3730 => x"34",
          3731 => x"d4",
          3732 => x"12",
          3733 => x"07",
          3734 => x"33",
          3735 => x"41",
          3736 => x"79",
          3737 => x"05",
          3738 => x"33",
          3739 => x"81",
          3740 => x"42",
          3741 => x"19",
          3742 => x"70",
          3743 => x"71",
          3744 => x"81",
          3745 => x"83",
          3746 => x"63",
          3747 => x"40",
          3748 => x"7b",
          3749 => x"70",
          3750 => x"8b",
          3751 => x"70",
          3752 => x"07",
          3753 => x"48",
          3754 => x"60",
          3755 => x"61",
          3756 => x"39",
          3757 => x"8b",
          3758 => x"84",
          3759 => x"2b",
          3760 => x"52",
          3761 => x"85",
          3762 => x"19",
          3763 => x"8b",
          3764 => x"86",
          3765 => x"2b",
          3766 => x"52",
          3767 => x"05",
          3768 => x"b8",
          3769 => x"33",
          3770 => x"06",
          3771 => x"77",
          3772 => x"b8",
          3773 => x"12",
          3774 => x"07",
          3775 => x"71",
          3776 => x"ff",
          3777 => x"56",
          3778 => x"55",
          3779 => x"34",
          3780 => x"33",
          3781 => x"83",
          3782 => x"12",
          3783 => x"ff",
          3784 => x"58",
          3785 => x"76",
          3786 => x"70",
          3787 => x"71",
          3788 => x"11",
          3789 => x"8b",
          3790 => x"84",
          3791 => x"2b",
          3792 => x"52",
          3793 => x"57",
          3794 => x"34",
          3795 => x"11",
          3796 => x"71",
          3797 => x"33",
          3798 => x"70",
          3799 => x"57",
          3800 => x"87",
          3801 => x"70",
          3802 => x"07",
          3803 => x"5a",
          3804 => x"81",
          3805 => x"1f",
          3806 => x"8b",
          3807 => x"73",
          3808 => x"07",
          3809 => x"5f",
          3810 => x"81",
          3811 => x"1f",
          3812 => x"2b",
          3813 => x"14",
          3814 => x"07",
          3815 => x"5f",
          3816 => x"75",
          3817 => x"70",
          3818 => x"71",
          3819 => x"70",
          3820 => x"05",
          3821 => x"84",
          3822 => x"65",
          3823 => x"5d",
          3824 => x"33",
          3825 => x"83",
          3826 => x"85",
          3827 => x"88",
          3828 => x"7a",
          3829 => x"05",
          3830 => x"84",
          3831 => x"2b",
          3832 => x"14",
          3833 => x"07",
          3834 => x"5c",
          3835 => x"34",
          3836 => x"d4",
          3837 => x"71",
          3838 => x"70",
          3839 => x"75",
          3840 => x"d4",
          3841 => x"33",
          3842 => x"74",
          3843 => x"88",
          3844 => x"f8",
          3845 => x"44",
          3846 => x"74",
          3847 => x"84",
          3848 => x"81",
          3849 => x"2b",
          3850 => x"33",
          3851 => x"06",
          3852 => x"46",
          3853 => x"81",
          3854 => x"5b",
          3855 => x"e5",
          3856 => x"84",
          3857 => x"62",
          3858 => x"51",
          3859 => x"88",
          3860 => x"b7",
          3861 => x"7a",
          3862 => x"58",
          3863 => x"77",
          3864 => x"89",
          3865 => x"3f",
          3866 => x"e4",
          3867 => x"80",
          3868 => x"b7",
          3869 => x"89",
          3870 => x"84",
          3871 => x"b8",
          3872 => x"52",
          3873 => x"3f",
          3874 => x"34",
          3875 => x"d4",
          3876 => x"0b",
          3877 => x"56",
          3878 => x"17",
          3879 => x"d0",
          3880 => x"70",
          3881 => x"58",
          3882 => x"73",
          3883 => x"70",
          3884 => x"05",
          3885 => x"34",
          3886 => x"77",
          3887 => x"39",
          3888 => x"51",
          3889 => x"84",
          3890 => x"b8",
          3891 => x"3d",
          3892 => x"53",
          3893 => x"d4",
          3894 => x"ff",
          3895 => x"b8",
          3896 => x"33",
          3897 => x"3d",
          3898 => x"60",
          3899 => x"5c",
          3900 => x"87",
          3901 => x"73",
          3902 => x"38",
          3903 => x"8c",
          3904 => x"d5",
          3905 => x"ff",
          3906 => x"87",
          3907 => x"38",
          3908 => x"80",
          3909 => x"38",
          3910 => x"e4",
          3911 => x"16",
          3912 => x"55",
          3913 => x"d5",
          3914 => x"02",
          3915 => x"57",
          3916 => x"38",
          3917 => x"81",
          3918 => x"73",
          3919 => x"0c",
          3920 => x"8e",
          3921 => x"06",
          3922 => x"c0",
          3923 => x"79",
          3924 => x"80",
          3925 => x"81",
          3926 => x"0c",
          3927 => x"81",
          3928 => x"56",
          3929 => x"39",
          3930 => x"9b",
          3931 => x"33",
          3932 => x"26",
          3933 => x"53",
          3934 => x"9b",
          3935 => x"0c",
          3936 => x"72",
          3937 => x"9a",
          3938 => x"0c",
          3939 => x"75",
          3940 => x"3d",
          3941 => x"0b",
          3942 => x"04",
          3943 => x"11",
          3944 => x"70",
          3945 => x"80",
          3946 => x"08",
          3947 => x"8c",
          3948 => x"0c",
          3949 => x"08",
          3950 => x"9b",
          3951 => x"ee",
          3952 => x"7c",
          3953 => x"5b",
          3954 => x"06",
          3955 => x"2e",
          3956 => x"81",
          3957 => x"b8",
          3958 => x"59",
          3959 => x"0d",
          3960 => x"b8",
          3961 => x"5a",
          3962 => x"e4",
          3963 => x"38",
          3964 => x"b4",
          3965 => x"a0",
          3966 => x"58",
          3967 => x"38",
          3968 => x"09",
          3969 => x"75",
          3970 => x"51",
          3971 => x"59",
          3972 => x"fb",
          3973 => x"2e",
          3974 => x"18",
          3975 => x"75",
          3976 => x"57",
          3977 => x"b6",
          3978 => x"19",
          3979 => x"0b",
          3980 => x"19",
          3981 => x"80",
          3982 => x"f2",
          3983 => x"0b",
          3984 => x"84",
          3985 => x"74",
          3986 => x"5b",
          3987 => x"2a",
          3988 => x"98",
          3989 => x"90",
          3990 => x"34",
          3991 => x"19",
          3992 => x"a6",
          3993 => x"84",
          3994 => x"05",
          3995 => x"7a",
          3996 => x"fa",
          3997 => x"53",
          3998 => x"d8",
          3999 => x"fd",
          4000 => x"0d",
          4001 => x"81",
          4002 => x"76",
          4003 => x"b8",
          4004 => x"77",
          4005 => x"cc",
          4006 => x"74",
          4007 => x"75",
          4008 => x"19",
          4009 => x"17",
          4010 => x"33",
          4011 => x"83",
          4012 => x"17",
          4013 => x"3f",
          4014 => x"38",
          4015 => x"0c",
          4016 => x"06",
          4017 => x"89",
          4018 => x"5d",
          4019 => x"38",
          4020 => x"56",
          4021 => x"84",
          4022 => x"17",
          4023 => x"3f",
          4024 => x"38",
          4025 => x"0c",
          4026 => x"06",
          4027 => x"7e",
          4028 => x"53",
          4029 => x"38",
          4030 => x"0c",
          4031 => x"a8",
          4032 => x"79",
          4033 => x"33",
          4034 => x"09",
          4035 => x"78",
          4036 => x"51",
          4037 => x"80",
          4038 => x"78",
          4039 => x"75",
          4040 => x"05",
          4041 => x"2b",
          4042 => x"8f",
          4043 => x"81",
          4044 => x"a8",
          4045 => x"79",
          4046 => x"33",
          4047 => x"09",
          4048 => x"78",
          4049 => x"51",
          4050 => x"80",
          4051 => x"78",
          4052 => x"75",
          4053 => x"b8",
          4054 => x"71",
          4055 => x"14",
          4056 => x"33",
          4057 => x"07",
          4058 => x"59",
          4059 => x"54",
          4060 => x"53",
          4061 => x"3f",
          4062 => x"2e",
          4063 => x"b8",
          4064 => x"08",
          4065 => x"08",
          4066 => x"fe",
          4067 => x"82",
          4068 => x"81",
          4069 => x"05",
          4070 => x"f6",
          4071 => x"81",
          4072 => x"70",
          4073 => x"81",
          4074 => x"09",
          4075 => x"e4",
          4076 => x"a8",
          4077 => x"08",
          4078 => x"7d",
          4079 => x"e4",
          4080 => x"b4",
          4081 => x"81",
          4082 => x"81",
          4083 => x"09",
          4084 => x"e4",
          4085 => x"a8",
          4086 => x"5b",
          4087 => x"c5",
          4088 => x"2e",
          4089 => x"54",
          4090 => x"53",
          4091 => x"f1",
          4092 => x"54",
          4093 => x"53",
          4094 => x"3f",
          4095 => x"2e",
          4096 => x"b8",
          4097 => x"08",
          4098 => x"08",
          4099 => x"fb",
          4100 => x"82",
          4101 => x"81",
          4102 => x"05",
          4103 => x"f4",
          4104 => x"81",
          4105 => x"05",
          4106 => x"f3",
          4107 => x"7a",
          4108 => x"3d",
          4109 => x"82",
          4110 => x"9c",
          4111 => x"55",
          4112 => x"24",
          4113 => x"8a",
          4114 => x"3d",
          4115 => x"08",
          4116 => x"58",
          4117 => x"83",
          4118 => x"2e",
          4119 => x"54",
          4120 => x"33",
          4121 => x"08",
          4122 => x"5a",
          4123 => x"ff",
          4124 => x"79",
          4125 => x"5e",
          4126 => x"5a",
          4127 => x"1a",
          4128 => x"3d",
          4129 => x"06",
          4130 => x"1a",
          4131 => x"08",
          4132 => x"38",
          4133 => x"7c",
          4134 => x"81",
          4135 => x"19",
          4136 => x"e4",
          4137 => x"81",
          4138 => x"79",
          4139 => x"fc",
          4140 => x"33",
          4141 => x"f0",
          4142 => x"7d",
          4143 => x"b9",
          4144 => x"ba",
          4145 => x"bb",
          4146 => x"fe",
          4147 => x"89",
          4148 => x"08",
          4149 => x"38",
          4150 => x"56",
          4151 => x"82",
          4152 => x"19",
          4153 => x"3f",
          4154 => x"38",
          4155 => x"0c",
          4156 => x"83",
          4157 => x"77",
          4158 => x"7c",
          4159 => x"9f",
          4160 => x"07",
          4161 => x"83",
          4162 => x"08",
          4163 => x"56",
          4164 => x"81",
          4165 => x"81",
          4166 => x"81",
          4167 => x"09",
          4168 => x"e4",
          4169 => x"70",
          4170 => x"84",
          4171 => x"74",
          4172 => x"55",
          4173 => x"54",
          4174 => x"51",
          4175 => x"80",
          4176 => x"75",
          4177 => x"7d",
          4178 => x"84",
          4179 => x"88",
          4180 => x"8f",
          4181 => x"81",
          4182 => x"81",
          4183 => x"81",
          4184 => x"81",
          4185 => x"09",
          4186 => x"e4",
          4187 => x"70",
          4188 => x"84",
          4189 => x"7e",
          4190 => x"33",
          4191 => x"fb",
          4192 => x"7c",
          4193 => x"3f",
          4194 => x"76",
          4195 => x"33",
          4196 => x"84",
          4197 => x"06",
          4198 => x"83",
          4199 => x"1b",
          4200 => x"e4",
          4201 => x"27",
          4202 => x"74",
          4203 => x"38",
          4204 => x"81",
          4205 => x"5c",
          4206 => x"b8",
          4207 => x"57",
          4208 => x"e4",
          4209 => x"c5",
          4210 => x"34",
          4211 => x"31",
          4212 => x"5d",
          4213 => x"87",
          4214 => x"2e",
          4215 => x"54",
          4216 => x"33",
          4217 => x"e7",
          4218 => x"52",
          4219 => x"7e",
          4220 => x"83",
          4221 => x"ff",
          4222 => x"34",
          4223 => x"34",
          4224 => x"39",
          4225 => x"7a",
          4226 => x"98",
          4227 => x"06",
          4228 => x"7d",
          4229 => x"1d",
          4230 => x"1d",
          4231 => x"1d",
          4232 => x"7c",
          4233 => x"81",
          4234 => x"80",
          4235 => x"08",
          4236 => x"70",
          4237 => x"38",
          4238 => x"56",
          4239 => x"26",
          4240 => x"82",
          4241 => x"f5",
          4242 => x"81",
          4243 => x"08",
          4244 => x"08",
          4245 => x"25",
          4246 => x"73",
          4247 => x"81",
          4248 => x"84",
          4249 => x"81",
          4250 => x"08",
          4251 => x"f0",
          4252 => x"e4",
          4253 => x"08",
          4254 => x"ce",
          4255 => x"08",
          4256 => x"39",
          4257 => x"26",
          4258 => x"51",
          4259 => x"e4",
          4260 => x"b8",
          4261 => x"07",
          4262 => x"e4",
          4263 => x"ff",
          4264 => x"2e",
          4265 => x"74",
          4266 => x"08",
          4267 => x"57",
          4268 => x"8e",
          4269 => x"f5",
          4270 => x"b8",
          4271 => x"08",
          4272 => x"80",
          4273 => x"90",
          4274 => x"94",
          4275 => x"86",
          4276 => x"19",
          4277 => x"34",
          4278 => x"8c",
          4279 => x"e4",
          4280 => x"e4",
          4281 => x"2e",
          4282 => x"78",
          4283 => x"08",
          4284 => x"08",
          4285 => x"04",
          4286 => x"38",
          4287 => x"0d",
          4288 => x"73",
          4289 => x"73",
          4290 => x"73",
          4291 => x"74",
          4292 => x"82",
          4293 => x"53",
          4294 => x"72",
          4295 => x"98",
          4296 => x"18",
          4297 => x"94",
          4298 => x"0c",
          4299 => x"9c",
          4300 => x"e4",
          4301 => x"84",
          4302 => x"ac",
          4303 => x"ac",
          4304 => x"57",
          4305 => x"17",
          4306 => x"56",
          4307 => x"8a",
          4308 => x"08",
          4309 => x"ff",
          4310 => x"cd",
          4311 => x"b8",
          4312 => x"0b",
          4313 => x"38",
          4314 => x"08",
          4315 => x"31",
          4316 => x"aa",
          4317 => x"8a",
          4318 => x"70",
          4319 => x"5a",
          4320 => x"38",
          4321 => x"08",
          4322 => x"38",
          4323 => x"38",
          4324 => x"75",
          4325 => x"22",
          4326 => x"38",
          4327 => x"0c",
          4328 => x"80",
          4329 => x"3d",
          4330 => x"19",
          4331 => x"5c",
          4332 => x"eb",
          4333 => x"82",
          4334 => x"27",
          4335 => x"08",
          4336 => x"84",
          4337 => x"60",
          4338 => x"08",
          4339 => x"b8",
          4340 => x"e4",
          4341 => x"56",
          4342 => x"91",
          4343 => x"ff",
          4344 => x"08",
          4345 => x"ea",
          4346 => x"05",
          4347 => x"8d",
          4348 => x"b0",
          4349 => x"1a",
          4350 => x"57",
          4351 => x"34",
          4352 => x"56",
          4353 => x"81",
          4354 => x"77",
          4355 => x"3f",
          4356 => x"81",
          4357 => x"0c",
          4358 => x"3d",
          4359 => x"53",
          4360 => x"52",
          4361 => x"08",
          4362 => x"83",
          4363 => x"08",
          4364 => x"fe",
          4365 => x"82",
          4366 => x"81",
          4367 => x"05",
          4368 => x"e3",
          4369 => x"22",
          4370 => x"74",
          4371 => x"7c",
          4372 => x"08",
          4373 => x"7d",
          4374 => x"76",
          4375 => x"19",
          4376 => x"84",
          4377 => x"ee",
          4378 => x"7c",
          4379 => x"1e",
          4380 => x"82",
          4381 => x"80",
          4382 => x"d1",
          4383 => x"74",
          4384 => x"38",
          4385 => x"81",
          4386 => x"b8",
          4387 => x"5a",
          4388 => x"5b",
          4389 => x"70",
          4390 => x"81",
          4391 => x"81",
          4392 => x"34",
          4393 => x"ae",
          4394 => x"80",
          4395 => x"74",
          4396 => x"56",
          4397 => x"60",
          4398 => x"80",
          4399 => x"b8",
          4400 => x"81",
          4401 => x"fe",
          4402 => x"94",
          4403 => x"08",
          4404 => x"e1",
          4405 => x"08",
          4406 => x"38",
          4407 => x"b4",
          4408 => x"b8",
          4409 => x"08",
          4410 => x"41",
          4411 => x"a8",
          4412 => x"1a",
          4413 => x"33",
          4414 => x"90",
          4415 => x"81",
          4416 => x"5b",
          4417 => x"33",
          4418 => x"08",
          4419 => x"76",
          4420 => x"74",
          4421 => x"60",
          4422 => x"c1",
          4423 => x"0c",
          4424 => x"0d",
          4425 => x"18",
          4426 => x"06",
          4427 => x"33",
          4428 => x"58",
          4429 => x"33",
          4430 => x"05",
          4431 => x"e4",
          4432 => x"33",
          4433 => x"44",
          4434 => x"79",
          4435 => x"10",
          4436 => x"23",
          4437 => x"77",
          4438 => x"2a",
          4439 => x"90",
          4440 => x"38",
          4441 => x"23",
          4442 => x"41",
          4443 => x"2e",
          4444 => x"39",
          4445 => x"74",
          4446 => x"78",
          4447 => x"05",
          4448 => x"56",
          4449 => x"fd",
          4450 => x"7a",
          4451 => x"04",
          4452 => x"5c",
          4453 => x"84",
          4454 => x"08",
          4455 => x"5d",
          4456 => x"5e",
          4457 => x"1b",
          4458 => x"1b",
          4459 => x"09",
          4460 => x"75",
          4461 => x"51",
          4462 => x"80",
          4463 => x"75",
          4464 => x"b2",
          4465 => x"59",
          4466 => x"19",
          4467 => x"57",
          4468 => x"e5",
          4469 => x"81",
          4470 => x"38",
          4471 => x"81",
          4472 => x"56",
          4473 => x"81",
          4474 => x"5a",
          4475 => x"06",
          4476 => x"38",
          4477 => x"1c",
          4478 => x"8b",
          4479 => x"81",
          4480 => x"5a",
          4481 => x"58",
          4482 => x"38",
          4483 => x"5d",
          4484 => x"7b",
          4485 => x"08",
          4486 => x"fe",
          4487 => x"93",
          4488 => x"08",
          4489 => x"dc",
          4490 => x"08",
          4491 => x"38",
          4492 => x"b4",
          4493 => x"b8",
          4494 => x"08",
          4495 => x"5a",
          4496 => x"dd",
          4497 => x"1c",
          4498 => x"33",
          4499 => x"c5",
          4500 => x"1c",
          4501 => x"55",
          4502 => x"81",
          4503 => x"8d",
          4504 => x"90",
          4505 => x"5e",
          4506 => x"ff",
          4507 => x"f4",
          4508 => x"84",
          4509 => x"38",
          4510 => x"c2",
          4511 => x"1d",
          4512 => x"57",
          4513 => x"38",
          4514 => x"1b",
          4515 => x"40",
          4516 => x"bf",
          4517 => x"81",
          4518 => x"33",
          4519 => x"71",
          4520 => x"80",
          4521 => x"26",
          4522 => x"8a",
          4523 => x"61",
          4524 => x"5b",
          4525 => x"b8",
          4526 => x"de",
          4527 => x"78",
          4528 => x"86",
          4529 => x"2e",
          4530 => x"79",
          4531 => x"7f",
          4532 => x"ff",
          4533 => x"0b",
          4534 => x"04",
          4535 => x"38",
          4536 => x"3d",
          4537 => x"33",
          4538 => x"86",
          4539 => x"1d",
          4540 => x"80",
          4541 => x"17",
          4542 => x"38",
          4543 => x"60",
          4544 => x"05",
          4545 => x"34",
          4546 => x"80",
          4547 => x"56",
          4548 => x"c0",
          4549 => x"3d",
          4550 => x"59",
          4551 => x"70",
          4552 => x"05",
          4553 => x"38",
          4554 => x"79",
          4555 => x"38",
          4556 => x"75",
          4557 => x"2a",
          4558 => x"2a",
          4559 => x"80",
          4560 => x"32",
          4561 => x"d7",
          4562 => x"87",
          4563 => x"58",
          4564 => x"75",
          4565 => x"76",
          4566 => x"2a",
          4567 => x"1f",
          4568 => x"58",
          4569 => x"33",
          4570 => x"16",
          4571 => x"75",
          4572 => x"2e",
          4573 => x"56",
          4574 => x"98",
          4575 => x"71",
          4576 => x"87",
          4577 => x"f8",
          4578 => x"38",
          4579 => x"fe",
          4580 => x"2e",
          4581 => x"56",
          4582 => x"81",
          4583 => x"05",
          4584 => x"84",
          4585 => x"75",
          4586 => x"7e",
          4587 => x"1d",
          4588 => x"e4",
          4589 => x"ed",
          4590 => x"84",
          4591 => x"b8",
          4592 => x"1e",
          4593 => x"76",
          4594 => x"40",
          4595 => x"a3",
          4596 => x"52",
          4597 => x"84",
          4598 => x"ff",
          4599 => x"76",
          4600 => x"70",
          4601 => x"81",
          4602 => x"78",
          4603 => x"c9",
          4604 => x"86",
          4605 => x"83",
          4606 => x"b8",
          4607 => x"87",
          4608 => x"75",
          4609 => x"40",
          4610 => x"57",
          4611 => x"83",
          4612 => x"82",
          4613 => x"52",
          4614 => x"84",
          4615 => x"ff",
          4616 => x"75",
          4617 => x"9c",
          4618 => x"81",
          4619 => x"f4",
          4620 => x"58",
          4621 => x"33",
          4622 => x"15",
          4623 => x"ab",
          4624 => x"8c",
          4625 => x"77",
          4626 => x"3d",
          4627 => x"25",
          4628 => x"b9",
          4629 => x"ec",
          4630 => x"84",
          4631 => x"38",
          4632 => x"08",
          4633 => x"d3",
          4634 => x"2e",
          4635 => x"b8",
          4636 => x"08",
          4637 => x"19",
          4638 => x"41",
          4639 => x"b8",
          4640 => x"85",
          4641 => x"58",
          4642 => x"e4",
          4643 => x"ef",
          4644 => x"58",
          4645 => x"80",
          4646 => x"33",
          4647 => x"ff",
          4648 => x"74",
          4649 => x"98",
          4650 => x"08",
          4651 => x"5b",
          4652 => x"c9",
          4653 => x"52",
          4654 => x"84",
          4655 => x"ff",
          4656 => x"75",
          4657 => x"08",
          4658 => x"5f",
          4659 => x"0b",
          4660 => x"75",
          4661 => x"7c",
          4662 => x"58",
          4663 => x"38",
          4664 => x"5b",
          4665 => x"7b",
          4666 => x"57",
          4667 => x"34",
          4668 => x"81",
          4669 => x"76",
          4670 => x"78",
          4671 => x"80",
          4672 => x"81",
          4673 => x"51",
          4674 => x"58",
          4675 => x"7f",
          4676 => x"fb",
          4677 => x"53",
          4678 => x"52",
          4679 => x"b8",
          4680 => x"e4",
          4681 => x"a8",
          4682 => x"57",
          4683 => x"c9",
          4684 => x"2e",
          4685 => x"54",
          4686 => x"53",
          4687 => x"d1",
          4688 => x"9c",
          4689 => x"74",
          4690 => x"ba",
          4691 => x"57",
          4692 => x"d7",
          4693 => x"d4",
          4694 => x"61",
          4695 => x"3f",
          4696 => x"81",
          4697 => x"83",
          4698 => x"08",
          4699 => x"8a",
          4700 => x"2e",
          4701 => x"fc",
          4702 => x"7f",
          4703 => x"39",
          4704 => x"70",
          4705 => x"38",
          4706 => x"08",
          4707 => x"81",
          4708 => x"c1",
          4709 => x"19",
          4710 => x"33",
          4711 => x"f3",
          4712 => x"5e",
          4713 => x"1c",
          4714 => x"1c",
          4715 => x"70",
          4716 => x"57",
          4717 => x"bc",
          4718 => x"81",
          4719 => x"38",
          4720 => x"ff",
          4721 => x"82",
          4722 => x"70",
          4723 => x"38",
          4724 => x"7a",
          4725 => x"05",
          4726 => x"70",
          4727 => x"08",
          4728 => x"53",
          4729 => x"2e",
          4730 => x"30",
          4731 => x"54",
          4732 => x"2e",
          4733 => x"59",
          4734 => x"81",
          4735 => x"76",
          4736 => x"05",
          4737 => x"1d",
          4738 => x"f3",
          4739 => x"57",
          4740 => x"82",
          4741 => x"33",
          4742 => x"1e",
          4743 => x"33",
          4744 => x"11",
          4745 => x"90",
          4746 => x"33",
          4747 => x"71",
          4748 => x"96",
          4749 => x"41",
          4750 => x"86",
          4751 => x"33",
          4752 => x"84",
          4753 => x"e5",
          4754 => x"11",
          4755 => x"83",
          4756 => x"51",
          4757 => x"08",
          4758 => x"75",
          4759 => x"b3",
          4760 => x"34",
          4761 => x"58",
          4762 => x"78",
          4763 => x"54",
          4764 => x"74",
          4765 => x"25",
          4766 => x"75",
          4767 => x"78",
          4768 => x"56",
          4769 => x"33",
          4770 => x"88",
          4771 => x"54",
          4772 => x"54",
          4773 => x"08",
          4774 => x"27",
          4775 => x"81",
          4776 => x"a0",
          4777 => x"53",
          4778 => x"81",
          4779 => x"13",
          4780 => x"ff",
          4781 => x"2a",
          4782 => x"80",
          4783 => x"5f",
          4784 => x"63",
          4785 => x"65",
          4786 => x"2e",
          4787 => x"2e",
          4788 => x"d9",
          4789 => x"73",
          4790 => x"55",
          4791 => x"42",
          4792 => x"70",
          4793 => x"73",
          4794 => x"ff",
          4795 => x"74",
          4796 => x"80",
          4797 => x"ff",
          4798 => x"9f",
          4799 => x"5b",
          4800 => x"80",
          4801 => x"ff",
          4802 => x"83",
          4803 => x"56",
          4804 => x"38",
          4805 => x"70",
          4806 => x"56",
          4807 => x"5b",
          4808 => x"26",
          4809 => x"74",
          4810 => x"81",
          4811 => x"80",
          4812 => x"81",
          4813 => x"80",
          4814 => x"72",
          4815 => x"46",
          4816 => x"af",
          4817 => x"70",
          4818 => x"54",
          4819 => x"0c",
          4820 => x"42",
          4821 => x"b4",
          4822 => x"8d",
          4823 => x"ff",
          4824 => x"86",
          4825 => x"3d",
          4826 => x"81",
          4827 => x"fe",
          4828 => x"ab",
          4829 => x"8d",
          4830 => x"e4",
          4831 => x"80",
          4832 => x"73",
          4833 => x"2e",
          4834 => x"70",
          4835 => x"dd",
          4836 => x"70",
          4837 => x"7d",
          4838 => x"27",
          4839 => x"f8",
          4840 => x"76",
          4841 => x"76",
          4842 => x"70",
          4843 => x"52",
          4844 => x"2e",
          4845 => x"57",
          4846 => x"56",
          4847 => x"c7",
          4848 => x"ff",
          4849 => x"a0",
          4850 => x"ff",
          4851 => x"38",
          4852 => x"fe",
          4853 => x"2e",
          4854 => x"54",
          4855 => x"38",
          4856 => x"ae",
          4857 => x"0b",
          4858 => x"81",
          4859 => x"f4",
          4860 => x"16",
          4861 => x"5d",
          4862 => x"a0",
          4863 => x"70",
          4864 => x"75",
          4865 => x"bb",
          4866 => x"38",
          4867 => x"70",
          4868 => x"51",
          4869 => x"e0",
          4870 => x"75",
          4871 => x"5a",
          4872 => x"88",
          4873 => x"06",
          4874 => x"70",
          4875 => x"ff",
          4876 => x"81",
          4877 => x"2e",
          4878 => x"77",
          4879 => x"06",
          4880 => x"79",
          4881 => x"38",
          4882 => x"85",
          4883 => x"2a",
          4884 => x"38",
          4885 => x"34",
          4886 => x"e4",
          4887 => x"b8",
          4888 => x"84",
          4889 => x"06",
          4890 => x"06",
          4891 => x"74",
          4892 => x"98",
          4893 => x"42",
          4894 => x"ce",
          4895 => x"70",
          4896 => x"2e",
          4897 => x"38",
          4898 => x"82",
          4899 => x"81",
          4900 => x"73",
          4901 => x"38",
          4902 => x"80",
          4903 => x"76",
          4904 => x"75",
          4905 => x"53",
          4906 => x"07",
          4907 => x"e3",
          4908 => x"1d",
          4909 => x"fe",
          4910 => x"58",
          4911 => x"70",
          4912 => x"80",
          4913 => x"83",
          4914 => x"33",
          4915 => x"07",
          4916 => x"83",
          4917 => x"0c",
          4918 => x"39",
          4919 => x"f0",
          4920 => x"38",
          4921 => x"17",
          4922 => x"2b",
          4923 => x"5e",
          4924 => x"95",
          4925 => x"39",
          4926 => x"2e",
          4927 => x"39",
          4928 => x"0b",
          4929 => x"04",
          4930 => x"ff",
          4931 => x"59",
          4932 => x"83",
          4933 => x"fc",
          4934 => x"b5",
          4935 => x"84",
          4936 => x"70",
          4937 => x"80",
          4938 => x"83",
          4939 => x"81",
          4940 => x"2e",
          4941 => x"83",
          4942 => x"56",
          4943 => x"38",
          4944 => x"70",
          4945 => x"59",
          4946 => x"59",
          4947 => x"54",
          4948 => x"07",
          4949 => x"9f",
          4950 => x"7d",
          4951 => x"17",
          4952 => x"5f",
          4953 => x"79",
          4954 => x"fa",
          4955 => x"83",
          4956 => x"5a",
          4957 => x"80",
          4958 => x"05",
          4959 => x"1b",
          4960 => x"80",
          4961 => x"90",
          4962 => x"5a",
          4963 => x"05",
          4964 => x"34",
          4965 => x"5b",
          4966 => x"9c",
          4967 => x"58",
          4968 => x"06",
          4969 => x"82",
          4970 => x"38",
          4971 => x"3d",
          4972 => x"02",
          4973 => x"42",
          4974 => x"70",
          4975 => x"d7",
          4976 => x"70",
          4977 => x"85",
          4978 => x"2e",
          4979 => x"56",
          4980 => x"10",
          4981 => x"58",
          4982 => x"96",
          4983 => x"06",
          4984 => x"9b",
          4985 => x"b0",
          4986 => x"06",
          4987 => x"2e",
          4988 => x"16",
          4989 => x"18",
          4990 => x"ff",
          4991 => x"81",
          4992 => x"83",
          4993 => x"2e",
          4994 => x"41",
          4995 => x"5b",
          4996 => x"18",
          4997 => x"7a",
          4998 => x"33",
          4999 => x"b8",
          5000 => x"55",
          5001 => x"56",
          5002 => x"84",
          5003 => x"56",
          5004 => x"2e",
          5005 => x"38",
          5006 => x"85",
          5007 => x"83",
          5008 => x"83",
          5009 => x"c3",
          5010 => x"59",
          5011 => x"83",
          5012 => x"ce",
          5013 => x"5a",
          5014 => x"11",
          5015 => x"71",
          5016 => x"72",
          5017 => x"56",
          5018 => x"a0",
          5019 => x"18",
          5020 => x"70",
          5021 => x"58",
          5022 => x"81",
          5023 => x"19",
          5024 => x"23",
          5025 => x"38",
          5026 => x"bb",
          5027 => x"18",
          5028 => x"74",
          5029 => x"5e",
          5030 => x"80",
          5031 => x"71",
          5032 => x"38",
          5033 => x"12",
          5034 => x"07",
          5035 => x"2b",
          5036 => x"58",
          5037 => x"80",
          5038 => x"5d",
          5039 => x"ce",
          5040 => x"5a",
          5041 => x"52",
          5042 => x"3f",
          5043 => x"e4",
          5044 => x"b8",
          5045 => x"26",
          5046 => x"f5",
          5047 => x"f5",
          5048 => x"16",
          5049 => x"0c",
          5050 => x"1d",
          5051 => x"2e",
          5052 => x"8d",
          5053 => x"7d",
          5054 => x"7c",
          5055 => x"70",
          5056 => x"5a",
          5057 => x"58",
          5058 => x"ff",
          5059 => x"18",
          5060 => x"7c",
          5061 => x"34",
          5062 => x"7c",
          5063 => x"23",
          5064 => x"80",
          5065 => x"84",
          5066 => x"8b",
          5067 => x"0d",
          5068 => x"ff",
          5069 => x"91",
          5070 => x"d0",
          5071 => x"fe",
          5072 => x"5f",
          5073 => x"7a",
          5074 => x"81",
          5075 => x"58",
          5076 => x"16",
          5077 => x"9f",
          5078 => x"e0",
          5079 => x"75",
          5080 => x"77",
          5081 => x"ff",
          5082 => x"70",
          5083 => x"58",
          5084 => x"81",
          5085 => x"25",
          5086 => x"39",
          5087 => x"82",
          5088 => x"fe",
          5089 => x"7a",
          5090 => x"2e",
          5091 => x"75",
          5092 => x"25",
          5093 => x"ad",
          5094 => x"38",
          5095 => x"83",
          5096 => x"80",
          5097 => x"84",
          5098 => x"88",
          5099 => x"72",
          5100 => x"71",
          5101 => x"77",
          5102 => x"19",
          5103 => x"ff",
          5104 => x"70",
          5105 => x"9b",
          5106 => x"84",
          5107 => x"42",
          5108 => x"2e",
          5109 => x"34",
          5110 => x"80",
          5111 => x"54",
          5112 => x"33",
          5113 => x"e4",
          5114 => x"81",
          5115 => x"75",
          5116 => x"71",
          5117 => x"7b",
          5118 => x"a8",
          5119 => x"58",
          5120 => x"75",
          5121 => x"25",
          5122 => x"38",
          5123 => x"58",
          5124 => x"84",
          5125 => x"78",
          5126 => x"58",
          5127 => x"80",
          5128 => x"1a",
          5129 => x"38",
          5130 => x"18",
          5131 => x"70",
          5132 => x"05",
          5133 => x"5b",
          5134 => x"c5",
          5135 => x"0b",
          5136 => x"5d",
          5137 => x"7e",
          5138 => x"31",
          5139 => x"80",
          5140 => x"e1",
          5141 => x"58",
          5142 => x"e4",
          5143 => x"75",
          5144 => x"81",
          5145 => x"58",
          5146 => x"e4",
          5147 => x"80",
          5148 => x"58",
          5149 => x"70",
          5150 => x"ff",
          5151 => x"2e",
          5152 => x"38",
          5153 => x"98",
          5154 => x"5a",
          5155 => x"71",
          5156 => x"40",
          5157 => x"80",
          5158 => x"5a",
          5159 => x"fd",
          5160 => x"e8",
          5161 => x"55",
          5162 => x"d5",
          5163 => x"17",
          5164 => x"33",
          5165 => x"82",
          5166 => x"17",
          5167 => x"d2",
          5168 => x"85",
          5169 => x"18",
          5170 => x"18",
          5171 => x"18",
          5172 => x"75",
          5173 => x"f8",
          5174 => x"82",
          5175 => x"2b",
          5176 => x"88",
          5177 => x"59",
          5178 => x"85",
          5179 => x"cd",
          5180 => x"82",
          5181 => x"2b",
          5182 => x"88",
          5183 => x"40",
          5184 => x"85",
          5185 => x"9d",
          5186 => x"82",
          5187 => x"2b",
          5188 => x"88",
          5189 => x"0c",
          5190 => x"82",
          5191 => x"2b",
          5192 => x"88",
          5193 => x"05",
          5194 => x"40",
          5195 => x"84",
          5196 => x"84",
          5197 => x"84",
          5198 => x"0b",
          5199 => x"83",
          5200 => x"0c",
          5201 => x"17",
          5202 => x"18",
          5203 => x"84",
          5204 => x"06",
          5205 => x"83",
          5206 => x"08",
          5207 => x"8b",
          5208 => x"2e",
          5209 => x"5a",
          5210 => x"2e",
          5211 => x"18",
          5212 => x"ab",
          5213 => x"18",
          5214 => x"8d",
          5215 => x"22",
          5216 => x"17",
          5217 => x"90",
          5218 => x"33",
          5219 => x"71",
          5220 => x"2b",
          5221 => x"d8",
          5222 => x"e8",
          5223 => x"80",
          5224 => x"57",
          5225 => x"5a",
          5226 => x"75",
          5227 => x"05",
          5228 => x"ff",
          5229 => x"3d",
          5230 => x"70",
          5231 => x"76",
          5232 => x"38",
          5233 => x"9f",
          5234 => x"e2",
          5235 => x"80",
          5236 => x"80",
          5237 => x"10",
          5238 => x"55",
          5239 => x"34",
          5240 => x"80",
          5241 => x"7c",
          5242 => x"53",
          5243 => x"ef",
          5244 => x"73",
          5245 => x"04",
          5246 => x"3d",
          5247 => x"81",
          5248 => x"26",
          5249 => x"06",
          5250 => x"80",
          5251 => x"d4",
          5252 => x"5a",
          5253 => x"70",
          5254 => x"59",
          5255 => x"e0",
          5256 => x"ff",
          5257 => x"38",
          5258 => x"54",
          5259 => x"74",
          5260 => x"76",
          5261 => x"30",
          5262 => x"5c",
          5263 => x"81",
          5264 => x"25",
          5265 => x"39",
          5266 => x"60",
          5267 => x"0d",
          5268 => x"33",
          5269 => x"a6",
          5270 => x"3d",
          5271 => x"52",
          5272 => x"08",
          5273 => x"8f",
          5274 => x"84",
          5275 => x"7e",
          5276 => x"5a",
          5277 => x"57",
          5278 => x"ba",
          5279 => x"2e",
          5280 => x"c1",
          5281 => x"77",
          5282 => x"77",
          5283 => x"2e",
          5284 => x"9a",
          5285 => x"70",
          5286 => x"83",
          5287 => x"17",
          5288 => x"0b",
          5289 => x"17",
          5290 => x"34",
          5291 => x"17",
          5292 => x"33",
          5293 => x"66",
          5294 => x"0b",
          5295 => x"34",
          5296 => x"81",
          5297 => x"80",
          5298 => x"7c",
          5299 => x"27",
          5300 => x"83",
          5301 => x"fe",
          5302 => x"70",
          5303 => x"fe",
          5304 => x"57",
          5305 => x"38",
          5306 => x"2a",
          5307 => x"38",
          5308 => x"80",
          5309 => x"79",
          5310 => x"06",
          5311 => x"80",
          5312 => x"a0",
          5313 => x"9b",
          5314 => x"2b",
          5315 => x"5a",
          5316 => x"88",
          5317 => x"82",
          5318 => x"2b",
          5319 => x"88",
          5320 => x"8c",
          5321 => x"41",
          5322 => x"84",
          5323 => x"0b",
          5324 => x"0c",
          5325 => x"80",
          5326 => x"84",
          5327 => x"1a",
          5328 => x"58",
          5329 => x"56",
          5330 => x"81",
          5331 => x"2e",
          5332 => x"ff",
          5333 => x"58",
          5334 => x"38",
          5335 => x"2e",
          5336 => x"c0",
          5337 => x"06",
          5338 => x"81",
          5339 => x"38",
          5340 => x"39",
          5341 => x"39",
          5342 => x"39",
          5343 => x"e4",
          5344 => x"fb",
          5345 => x"7b",
          5346 => x"16",
          5347 => x"71",
          5348 => x"5c",
          5349 => x"27",
          5350 => x"ff",
          5351 => x"5d",
          5352 => x"a7",
          5353 => x"fc",
          5354 => x"2e",
          5355 => x"76",
          5356 => x"e4",
          5357 => x"fe",
          5358 => x"75",
          5359 => x"94",
          5360 => x"55",
          5361 => x"7d",
          5362 => x"80",
          5363 => x"17",
          5364 => x"94",
          5365 => x"2b",
          5366 => x"0b",
          5367 => x"34",
          5368 => x"0b",
          5369 => x"8b",
          5370 => x"0b",
          5371 => x"34",
          5372 => x"81",
          5373 => x"80",
          5374 => x"b4",
          5375 => x"16",
          5376 => x"06",
          5377 => x"16",
          5378 => x"ba",
          5379 => x"85",
          5380 => x"17",
          5381 => x"18",
          5382 => x"38",
          5383 => x"54",
          5384 => x"53",
          5385 => x"81",
          5386 => x"09",
          5387 => x"e4",
          5388 => x"a8",
          5389 => x"5c",
          5390 => x"92",
          5391 => x"2e",
          5392 => x"54",
          5393 => x"53",
          5394 => x"a3",
          5395 => x"74",
          5396 => x"39",
          5397 => x"38",
          5398 => x"2e",
          5399 => x"12",
          5400 => x"7d",
          5401 => x"78",
          5402 => x"5c",
          5403 => x"89",
          5404 => x"f7",
          5405 => x"56",
          5406 => x"0c",
          5407 => x"57",
          5408 => x"7f",
          5409 => x"0d",
          5410 => x"5a",
          5411 => x"2e",
          5412 => x"2e",
          5413 => x"2e",
          5414 => x"22",
          5415 => x"38",
          5416 => x"82",
          5417 => x"82",
          5418 => x"57",
          5419 => x"38",
          5420 => x"31",
          5421 => x"38",
          5422 => x"59",
          5423 => x"e3",
          5424 => x"89",
          5425 => x"83",
          5426 => x"75",
          5427 => x"83",
          5428 => x"59",
          5429 => x"08",
          5430 => x"83",
          5431 => x"29",
          5432 => x"80",
          5433 => x"89",
          5434 => x"81",
          5435 => x"85",
          5436 => x"76",
          5437 => x"ff",
          5438 => x"83",
          5439 => x"59",
          5440 => x"08",
          5441 => x"38",
          5442 => x"1b",
          5443 => x"57",
          5444 => x"ff",
          5445 => x"2b",
          5446 => x"7f",
          5447 => x"70",
          5448 => x"fe",
          5449 => x"e4",
          5450 => x"b8",
          5451 => x"5c",
          5452 => x"75",
          5453 => x"59",
          5454 => x"58",
          5455 => x"b6",
          5456 => x"5d",
          5457 => x"06",
          5458 => x"b8",
          5459 => x"9e",
          5460 => x"2e",
          5461 => x"b4",
          5462 => x"94",
          5463 => x"7f",
          5464 => x"80",
          5465 => x"05",
          5466 => x"34",
          5467 => x"d1",
          5468 => x"77",
          5469 => x"56",
          5470 => x"54",
          5471 => x"53",
          5472 => x"c9",
          5473 => x"7f",
          5474 => x"84",
          5475 => x"19",
          5476 => x"e4",
          5477 => x"27",
          5478 => x"74",
          5479 => x"38",
          5480 => x"08",
          5481 => x"51",
          5482 => x"bb",
          5483 => x"08",
          5484 => x"52",
          5485 => x"b8",
          5486 => x"16",
          5487 => x"b8",
          5488 => x"b8",
          5489 => x"b2",
          5490 => x"0b",
          5491 => x"04",
          5492 => x"84",
          5493 => x"f0",
          5494 => x"40",
          5495 => x"79",
          5496 => x"75",
          5497 => x"74",
          5498 => x"84",
          5499 => x"85",
          5500 => x"55",
          5501 => x"55",
          5502 => x"70",
          5503 => x"56",
          5504 => x"1a",
          5505 => x"27",
          5506 => x"2e",
          5507 => x"5f",
          5508 => x"22",
          5509 => x"56",
          5510 => x"88",
          5511 => x"b1",
          5512 => x"74",
          5513 => x"1b",
          5514 => x"88",
          5515 => x"9c",
          5516 => x"1a",
          5517 => x"05",
          5518 => x"38",
          5519 => x"18",
          5520 => x"85",
          5521 => x"59",
          5522 => x"77",
          5523 => x"76",
          5524 => x"7c",
          5525 => x"a1",
          5526 => x"38",
          5527 => x"57",
          5528 => x"0b",
          5529 => x"58",
          5530 => x"77",
          5531 => x"56",
          5532 => x"1a",
          5533 => x"31",
          5534 => x"94",
          5535 => x"0c",
          5536 => x"5b",
          5537 => x"75",
          5538 => x"90",
          5539 => x"5b",
          5540 => x"84",
          5541 => x"74",
          5542 => x"04",
          5543 => x"38",
          5544 => x"1b",
          5545 => x"84",
          5546 => x"27",
          5547 => x"16",
          5548 => x"83",
          5549 => x"7f",
          5550 => x"81",
          5551 => x"16",
          5552 => x"b8",
          5553 => x"57",
          5554 => x"83",
          5555 => x"ff",
          5556 => x"59",
          5557 => x"76",
          5558 => x"81",
          5559 => x"ef",
          5560 => x"34",
          5561 => x"08",
          5562 => x"33",
          5563 => x"5c",
          5564 => x"81",
          5565 => x"08",
          5566 => x"17",
          5567 => x"55",
          5568 => x"38",
          5569 => x"09",
          5570 => x"b4",
          5571 => x"7f",
          5572 => x"a9",
          5573 => x"1a",
          5574 => x"93",
          5575 => x"b9",
          5576 => x"1b",
          5577 => x"0c",
          5578 => x"52",
          5579 => x"b8",
          5580 => x"fb",
          5581 => x"ab",
          5582 => x"cc",
          5583 => x"b8",
          5584 => x"81",
          5585 => x"70",
          5586 => x"97",
          5587 => x"b8",
          5588 => x"34",
          5589 => x"58",
          5590 => x"38",
          5591 => x"09",
          5592 => x"b4",
          5593 => x"76",
          5594 => x"f9",
          5595 => x"16",
          5596 => x"b8",
          5597 => x"f2",
          5598 => x"ec",
          5599 => x"b8",
          5600 => x"57",
          5601 => x"08",
          5602 => x"83",
          5603 => x"08",
          5604 => x"fe",
          5605 => x"82",
          5606 => x"81",
          5607 => x"05",
          5608 => x"ff",
          5609 => x"0c",
          5610 => x"39",
          5611 => x"84",
          5612 => x"82",
          5613 => x"b8",
          5614 => x"3d",
          5615 => x"2e",
          5616 => x"2e",
          5617 => x"2e",
          5618 => x"22",
          5619 => x"38",
          5620 => x"81",
          5621 => x"2a",
          5622 => x"81",
          5623 => x"57",
          5624 => x"83",
          5625 => x"81",
          5626 => x"17",
          5627 => x"b8",
          5628 => x"59",
          5629 => x"81",
          5630 => x"33",
          5631 => x"34",
          5632 => x"ff",
          5633 => x"18",
          5634 => x"18",
          5635 => x"5c",
          5636 => x"38",
          5637 => x"74",
          5638 => x"74",
          5639 => x"74",
          5640 => x"80",
          5641 => x"a1",
          5642 => x"99",
          5643 => x"80",
          5644 => x"0b",
          5645 => x"94",
          5646 => x"33",
          5647 => x"19",
          5648 => x"3d",
          5649 => x"53",
          5650 => x"52",
          5651 => x"84",
          5652 => x"b8",
          5653 => x"08",
          5654 => x"08",
          5655 => x"fe",
          5656 => x"82",
          5657 => x"81",
          5658 => x"05",
          5659 => x"ff",
          5660 => x"39",
          5661 => x"34",
          5662 => x"34",
          5663 => x"74",
          5664 => x"74",
          5665 => x"74",
          5666 => x"80",
          5667 => x"a1",
          5668 => x"99",
          5669 => x"80",
          5670 => x"0b",
          5671 => x"c4",
          5672 => x"33",
          5673 => x"19",
          5674 => x"51",
          5675 => x"08",
          5676 => x"74",
          5677 => x"f9",
          5678 => x"fe",
          5679 => x"b8",
          5680 => x"80",
          5681 => x"80",
          5682 => x"80",
          5683 => x"16",
          5684 => x"38",
          5685 => x"84",
          5686 => x"e4",
          5687 => x"33",
          5688 => x"e4",
          5689 => x"73",
          5690 => x"3d",
          5691 => x"75",
          5692 => x"05",
          5693 => x"71",
          5694 => x"71",
          5695 => x"33",
          5696 => x"84",
          5697 => x"e4",
          5698 => x"84",
          5699 => x"78",
          5700 => x"53",
          5701 => x"82",
          5702 => x"59",
          5703 => x"80",
          5704 => x"08",
          5705 => x"58",
          5706 => x"ff",
          5707 => x"26",
          5708 => x"06",
          5709 => x"99",
          5710 => x"ff",
          5711 => x"2a",
          5712 => x"06",
          5713 => x"76",
          5714 => x"2a",
          5715 => x"2e",
          5716 => x"58",
          5717 => x"51",
          5718 => x"38",
          5719 => x"ea",
          5720 => x"05",
          5721 => x"84",
          5722 => x"08",
          5723 => x"e4",
          5724 => x"68",
          5725 => x"94",
          5726 => x"b8",
          5727 => x"d7",
          5728 => x"80",
          5729 => x"05",
          5730 => x"59",
          5731 => x"9b",
          5732 => x"2b",
          5733 => x"58",
          5734 => x"19",
          5735 => x"3d",
          5736 => x"2e",
          5737 => x"0b",
          5738 => x"04",
          5739 => x"98",
          5740 => x"98",
          5741 => x"7e",
          5742 => x"e4",
          5743 => x"3d",
          5744 => x"3d",
          5745 => x"53",
          5746 => x"80",
          5747 => x"b8",
          5748 => x"83",
          5749 => x"7f",
          5750 => x"0c",
          5751 => x"79",
          5752 => x"3d",
          5753 => x"51",
          5754 => x"08",
          5755 => x"38",
          5756 => x"b4",
          5757 => x"b8",
          5758 => x"7d",
          5759 => x"b8",
          5760 => x"8b",
          5761 => x"2e",
          5762 => x"b4",
          5763 => x"df",
          5764 => x"33",
          5765 => x"5d",
          5766 => x"82",
          5767 => x"80",
          5768 => x"84",
          5769 => x"08",
          5770 => x"ff",
          5771 => x"59",
          5772 => x"df",
          5773 => x"33",
          5774 => x"42",
          5775 => x"81",
          5776 => x"84",
          5777 => x"a4",
          5778 => x"84",
          5779 => x"38",
          5780 => x"81",
          5781 => x"05",
          5782 => x"78",
          5783 => x"80",
          5784 => x"17",
          5785 => x"7c",
          5786 => x"26",
          5787 => x"38",
          5788 => x"80",
          5789 => x"19",
          5790 => x"34",
          5791 => x"3d",
          5792 => x"80",
          5793 => x"38",
          5794 => x"0b",
          5795 => x"83",
          5796 => x"43",
          5797 => x"8d",
          5798 => x"57",
          5799 => x"5b",
          5800 => x"76",
          5801 => x"7e",
          5802 => x"81",
          5803 => x"ba",
          5804 => x"ff",
          5805 => x"91",
          5806 => x"e4",
          5807 => x"16",
          5808 => x"71",
          5809 => x"5e",
          5810 => x"17",
          5811 => x"07",
          5812 => x"5d",
          5813 => x"3f",
          5814 => x"e4",
          5815 => x"b1",
          5816 => x"b8",
          5817 => x"5e",
          5818 => x"b8",
          5819 => x"e4",
          5820 => x"a8",
          5821 => x"5a",
          5822 => x"83",
          5823 => x"2e",
          5824 => x"54",
          5825 => x"53",
          5826 => x"88",
          5827 => x"ff",
          5828 => x"58",
          5829 => x"c0",
          5830 => x"05",
          5831 => x"5e",
          5832 => x"fd",
          5833 => x"3d",
          5834 => x"33",
          5835 => x"60",
          5836 => x"08",
          5837 => x"7c",
          5838 => x"26",
          5839 => x"80",
          5840 => x"80",
          5841 => x"7b",
          5842 => x"2e",
          5843 => x"2e",
          5844 => x"2e",
          5845 => x"22",
          5846 => x"38",
          5847 => x"81",
          5848 => x"81",
          5849 => x"76",
          5850 => x"54",
          5851 => x"38",
          5852 => x"52",
          5853 => x"38",
          5854 => x"ad",
          5855 => x"77",
          5856 => x"9d",
          5857 => x"81",
          5858 => x"94",
          5859 => x"08",
          5860 => x"98",
          5861 => x"76",
          5862 => x"17",
          5863 => x"81",
          5864 => x"81",
          5865 => x"99",
          5866 => x"84",
          5867 => x"38",
          5868 => x"27",
          5869 => x"14",
          5870 => x"16",
          5871 => x"16",
          5872 => x"0c",
          5873 => x"70",
          5874 => x"fe",
          5875 => x"57",
          5876 => x"06",
          5877 => x"94",
          5878 => x"38",
          5879 => x"80",
          5880 => x"73",
          5881 => x"8c",
          5882 => x"38",
          5883 => x"b8",
          5884 => x"0b",
          5885 => x"73",
          5886 => x"16",
          5887 => x"fe",
          5888 => x"94",
          5889 => x"83",
          5890 => x"38",
          5891 => x"05",
          5892 => x"f6",
          5893 => x"b0",
          5894 => x"5a",
          5895 => x"38",
          5896 => x"73",
          5897 => x"84",
          5898 => x"81",
          5899 => x"84",
          5900 => x"fc",
          5901 => x"fc",
          5902 => x"97",
          5903 => x"84",
          5904 => x"84",
          5905 => x"38",
          5906 => x"73",
          5907 => x"0b",
          5908 => x"e4",
          5909 => x"0d",
          5910 => x"a2",
          5911 => x"52",
          5912 => x"3f",
          5913 => x"e4",
          5914 => x"0c",
          5915 => x"8c",
          5916 => x"52",
          5917 => x"b8",
          5918 => x"80",
          5919 => x"2b",
          5920 => x"86",
          5921 => x"5b",
          5922 => x"9c",
          5923 => x"33",
          5924 => x"5d",
          5925 => x"b3",
          5926 => x"86",
          5927 => x"75",
          5928 => x"e4",
          5929 => x"74",
          5930 => x"0c",
          5931 => x"0c",
          5932 => x"18",
          5933 => x"07",
          5934 => x"ff",
          5935 => x"89",
          5936 => x"08",
          5937 => x"33",
          5938 => x"13",
          5939 => x"76",
          5940 => x"73",
          5941 => x"b8",
          5942 => x"13",
          5943 => x"b8",
          5944 => x"38",
          5945 => x"f8",
          5946 => x"56",
          5947 => x"54",
          5948 => x"53",
          5949 => x"22",
          5950 => x"2e",
          5951 => x"75",
          5952 => x"2e",
          5953 => x"ff",
          5954 => x"53",
          5955 => x"38",
          5956 => x"52",
          5957 => x"52",
          5958 => x"b8",
          5959 => x"72",
          5960 => x"06",
          5961 => x"0c",
          5962 => x"75",
          5963 => x"52",
          5964 => x"b8",
          5965 => x"72",
          5966 => x"06",
          5967 => x"74",
          5968 => x"e4",
          5969 => x"0d",
          5970 => x"e8",
          5971 => x"53",
          5972 => x"54",
          5973 => x"66",
          5974 => x"97",
          5975 => x"b8",
          5976 => x"80",
          5977 => x"0c",
          5978 => x"51",
          5979 => x"08",
          5980 => x"02",
          5981 => x"55",
          5982 => x"80",
          5983 => x"ff",
          5984 => x"0c",
          5985 => x"b8",
          5986 => x"3d",
          5987 => x"95",
          5988 => x"c0",
          5989 => x"84",
          5990 => x"0c",
          5991 => x"94",
          5992 => x"75",
          5993 => x"84",
          5994 => x"84",
          5995 => x"78",
          5996 => x"18",
          5997 => x"59",
          5998 => x"71",
          5999 => x"2e",
          6000 => x"5f",
          6001 => x"75",
          6002 => x"51",
          6003 => x"08",
          6004 => x"5e",
          6005 => x"57",
          6006 => x"7d",
          6007 => x"b8",
          6008 => x"71",
          6009 => x"14",
          6010 => x"33",
          6011 => x"07",
          6012 => x"60",
          6013 => x"05",
          6014 => x"58",
          6015 => x"7a",
          6016 => x"17",
          6017 => x"34",
          6018 => x"0d",
          6019 => x"b8",
          6020 => x"5d",
          6021 => x"b8",
          6022 => x"e4",
          6023 => x"a8",
          6024 => x"5f",
          6025 => x"bd",
          6026 => x"2e",
          6027 => x"54",
          6028 => x"53",
          6029 => x"fb",
          6030 => x"82",
          6031 => x"52",
          6032 => x"b8",
          6033 => x"84",
          6034 => x"38",
          6035 => x"b8",
          6036 => x"81",
          6037 => x"17",
          6038 => x"0c",
          6039 => x"81",
          6040 => x"c8",
          6041 => x"33",
          6042 => x"30",
          6043 => x"ff",
          6044 => x"5f",
          6045 => x"8f",
          6046 => x"60",
          6047 => x"18",
          6048 => x"77",
          6049 => x"60",
          6050 => x"7b",
          6051 => x"38",
          6052 => x"38",
          6053 => x"38",
          6054 => x"59",
          6055 => x"54",
          6056 => x"17",
          6057 => x"17",
          6058 => x"58",
          6059 => x"38",
          6060 => x"08",
          6061 => x"88",
          6062 => x"74",
          6063 => x"26",
          6064 => x"18",
          6065 => x"77",
          6066 => x"34",
          6067 => x"18",
          6068 => x"0c",
          6069 => x"78",
          6070 => x"51",
          6071 => x"08",
          6072 => x"80",
          6073 => x"2e",
          6074 => x"ff",
          6075 => x"52",
          6076 => x"b8",
          6077 => x"08",
          6078 => x"58",
          6079 => x"15",
          6080 => x"07",
          6081 => x"77",
          6082 => x"81",
          6083 => x"84",
          6084 => x"fe",
          6085 => x"fe",
          6086 => x"59",
          6087 => x"0c",
          6088 => x"76",
          6089 => x"e4",
          6090 => x"b8",
          6091 => x"75",
          6092 => x"e4",
          6093 => x"38",
          6094 => x"78",
          6095 => x"b8",
          6096 => x"b8",
          6097 => x"96",
          6098 => x"53",
          6099 => x"3f",
          6100 => x"e4",
          6101 => x"51",
          6102 => x"08",
          6103 => x"80",
          6104 => x"2e",
          6105 => x"ff",
          6106 => x"52",
          6107 => x"b8",
          6108 => x"08",
          6109 => x"58",
          6110 => x"94",
          6111 => x"54",
          6112 => x"79",
          6113 => x"56",
          6114 => x"81",
          6115 => x"18",
          6116 => x"56",
          6117 => x"59",
          6118 => x"08",
          6119 => x"39",
          6120 => x"fd",
          6121 => x"c0",
          6122 => x"3d",
          6123 => x"05",
          6124 => x"3f",
          6125 => x"e4",
          6126 => x"b8",
          6127 => x"4b",
          6128 => x"52",
          6129 => x"e4",
          6130 => x"38",
          6131 => x"2a",
          6132 => x"cd",
          6133 => x"24",
          6134 => x"70",
          6135 => x"ff",
          6136 => x"11",
          6137 => x"07",
          6138 => x"7c",
          6139 => x"2a",
          6140 => x"ed",
          6141 => x"2e",
          6142 => x"84",
          6143 => x"52",
          6144 => x"e4",
          6145 => x"e5",
          6146 => x"51",
          6147 => x"08",
          6148 => x"87",
          6149 => x"0d",
          6150 => x"71",
          6151 => x"07",
          6152 => x"b8",
          6153 => x"b8",
          6154 => x"6f",
          6155 => x"ff",
          6156 => x"51",
          6157 => x"08",
          6158 => x"be",
          6159 => x"25",
          6160 => x"74",
          6161 => x"58",
          6162 => x"17",
          6163 => x"56",
          6164 => x"f5",
          6165 => x"b8",
          6166 => x"17",
          6167 => x"b4",
          6168 => x"83",
          6169 => x"2e",
          6170 => x"54",
          6171 => x"33",
          6172 => x"e4",
          6173 => x"81",
          6174 => x"77",
          6175 => x"78",
          6176 => x"19",
          6177 => x"52",
          6178 => x"b8",
          6179 => x"80",
          6180 => x"09",
          6181 => x"fe",
          6182 => x"53",
          6183 => x"f2",
          6184 => x"08",
          6185 => x"38",
          6186 => x"b4",
          6187 => x"b8",
          6188 => x"08",
          6189 => x"55",
          6190 => x"de",
          6191 => x"18",
          6192 => x"33",
          6193 => x"fe",
          6194 => x"80",
          6195 => x"f6",
          6196 => x"84",
          6197 => x"38",
          6198 => x"e6",
          6199 => x"80",
          6200 => x"51",
          6201 => x"08",
          6202 => x"94",
          6203 => x"27",
          6204 => x"0c",
          6205 => x"84",
          6206 => x"ff",
          6207 => x"79",
          6208 => x"08",
          6209 => x"90",
          6210 => x"3d",
          6211 => x"ff",
          6212 => x"56",
          6213 => x"38",
          6214 => x"0d",
          6215 => x"70",
          6216 => x"b8",
          6217 => x"8b",
          6218 => x"9f",
          6219 => x"84",
          6220 => x"80",
          6221 => x"06",
          6222 => x"38",
          6223 => x"52",
          6224 => x"e4",
          6225 => x"08",
          6226 => x"08",
          6227 => x"e4",
          6228 => x"81",
          6229 => x"83",
          6230 => x"e2",
          6231 => x"05",
          6232 => x"8d",
          6233 => x"b0",
          6234 => x"18",
          6235 => x"57",
          6236 => x"34",
          6237 => x"58",
          6238 => x"81",
          6239 => x"78",
          6240 => x"c9",
          6241 => x"38",
          6242 => x"ff",
          6243 => x"53",
          6244 => x"52",
          6245 => x"84",
          6246 => x"e4",
          6247 => x"a8",
          6248 => x"08",
          6249 => x"5b",
          6250 => x"e1",
          6251 => x"18",
          6252 => x"33",
          6253 => x"39",
          6254 => x"81",
          6255 => x"18",
          6256 => x"7c",
          6257 => x"e4",
          6258 => x"2e",
          6259 => x"81",
          6260 => x"08",
          6261 => x"74",
          6262 => x"84",
          6263 => x"17",
          6264 => x"5c",
          6265 => x"18",
          6266 => x"07",
          6267 => x"78",
          6268 => x"b8",
          6269 => x"17",
          6270 => x"57",
          6271 => x"06",
          6272 => x"56",
          6273 => x"34",
          6274 => x"57",
          6275 => x"90",
          6276 => x"75",
          6277 => x"1a",
          6278 => x"80",
          6279 => x"7c",
          6280 => x"80",
          6281 => x"7a",
          6282 => x"74",
          6283 => x"a0",
          6284 => x"58",
          6285 => x"77",
          6286 => x"56",
          6287 => x"80",
          6288 => x"ff",
          6289 => x"f2",
          6290 => x"80",
          6291 => x"83",
          6292 => x"0b",
          6293 => x"96",
          6294 => x"b8",
          6295 => x"84",
          6296 => x"b8",
          6297 => x"98",
          6298 => x"34",
          6299 => x"34",
          6300 => x"34",
          6301 => x"d9",
          6302 => x"34",
          6303 => x"7d",
          6304 => x"e4",
          6305 => x"9f",
          6306 => x"74",
          6307 => x"57",
          6308 => x"39",
          6309 => x"17",
          6310 => x"cd",
          6311 => x"d8",
          6312 => x"a1",
          6313 => x"18",
          6314 => x"18",
          6315 => x"34",
          6316 => x"7d",
          6317 => x"e4",
          6318 => x"0d",
          6319 => x"5b",
          6320 => x"70",
          6321 => x"56",
          6322 => x"74",
          6323 => x"38",
          6324 => x"52",
          6325 => x"84",
          6326 => x"08",
          6327 => x"e4",
          6328 => x"3d",
          6329 => x"70",
          6330 => x"b8",
          6331 => x"dc",
          6332 => x"a0",
          6333 => x"a0",
          6334 => x"58",
          6335 => x"77",
          6336 => x"55",
          6337 => x"78",
          6338 => x"05",
          6339 => x"34",
          6340 => x"3d",
          6341 => x"3f",
          6342 => x"e4",
          6343 => x"08",
          6344 => x"b8",
          6345 => x"33",
          6346 => x"57",
          6347 => x"17",
          6348 => x"59",
          6349 => x"7f",
          6350 => x"5d",
          6351 => x"05",
          6352 => x"33",
          6353 => x"99",
          6354 => x"ff",
          6355 => x"77",
          6356 => x"81",
          6357 => x"9f",
          6358 => x"81",
          6359 => x"78",
          6360 => x"9f",
          6361 => x"80",
          6362 => x"5e",
          6363 => x"7c",
          6364 => x"7b",
          6365 => x"0c",
          6366 => x"52",
          6367 => x"84",
          6368 => x"08",
          6369 => x"aa",
          6370 => x"ac",
          6371 => x"84",
          6372 => x"08",
          6373 => x"8d",
          6374 => x"58",
          6375 => x"33",
          6376 => x"1a",
          6377 => x"05",
          6378 => x"70",
          6379 => x"89",
          6380 => x"19",
          6381 => x"34",
          6382 => x"06",
          6383 => x"38",
          6384 => x"38",
          6385 => x"71",
          6386 => x"5c",
          6387 => x"fe",
          6388 => x"56",
          6389 => x"17",
          6390 => x"05",
          6391 => x"38",
          6392 => x"76",
          6393 => x"7e",
          6394 => x"b8",
          6395 => x"e3",
          6396 => x"2e",
          6397 => x"b4",
          6398 => x"18",
          6399 => x"15",
          6400 => x"06",
          6401 => x"06",
          6402 => x"7b",
          6403 => x"34",
          6404 => x"81",
          6405 => x"7d",
          6406 => x"56",
          6407 => x"81",
          6408 => x"3d",
          6409 => x"74",
          6410 => x"51",
          6411 => x"08",
          6412 => x"38",
          6413 => x"80",
          6414 => x"38",
          6415 => x"7a",
          6416 => x"81",
          6417 => x"16",
          6418 => x"b8",
          6419 => x"57",
          6420 => x"55",
          6421 => x"e5",
          6422 => x"90",
          6423 => x"52",
          6424 => x"b8",
          6425 => x"80",
          6426 => x"84",
          6427 => x"f9",
          6428 => x"3f",
          6429 => x"0c",
          6430 => x"b8",
          6431 => x"18",
          6432 => x"71",
          6433 => x"5c",
          6434 => x"84",
          6435 => x"08",
          6436 => x"b8",
          6437 => x"54",
          6438 => x"16",
          6439 => x"58",
          6440 => x"81",
          6441 => x"08",
          6442 => x"17",
          6443 => x"55",
          6444 => x"38",
          6445 => x"09",
          6446 => x"b4",
          6447 => x"7b",
          6448 => x"c9",
          6449 => x"54",
          6450 => x"53",
          6451 => x"b1",
          6452 => x"fc",
          6453 => x"18",
          6454 => x"31",
          6455 => x"a0",
          6456 => x"17",
          6457 => x"06",
          6458 => x"08",
          6459 => x"81",
          6460 => x"79",
          6461 => x"02",
          6462 => x"80",
          6463 => x"96",
          6464 => x"ff",
          6465 => x"56",
          6466 => x"38",
          6467 => x"0d",
          6468 => x"d0",
          6469 => x"b8",
          6470 => x"e0",
          6471 => x"a0",
          6472 => x"74",
          6473 => x"33",
          6474 => x"56",
          6475 => x"55",
          6476 => x"fe",
          6477 => x"84",
          6478 => x"ec",
          6479 => x"3d",
          6480 => x"a1",
          6481 => x"84",
          6482 => x"74",
          6483 => x"04",
          6484 => x"05",
          6485 => x"e4",
          6486 => x"38",
          6487 => x"06",
          6488 => x"84",
          6489 => x"2b",
          6490 => x"34",
          6491 => x"34",
          6492 => x"34",
          6493 => x"34",
          6494 => x"78",
          6495 => x"e4",
          6496 => x"0d",
          6497 => x"5b",
          6498 => x"9b",
          6499 => x"b8",
          6500 => x"70",
          6501 => x"51",
          6502 => x"81",
          6503 => x"a4",
          6504 => x"25",
          6505 => x"38",
          6506 => x"80",
          6507 => x"08",
          6508 => x"77",
          6509 => x"7a",
          6510 => x"06",
          6511 => x"b8",
          6512 => x"dc",
          6513 => x"2e",
          6514 => x"b4",
          6515 => x"7c",
          6516 => x"74",
          6517 => x"74",
          6518 => x"18",
          6519 => x"33",
          6520 => x"81",
          6521 => x"75",
          6522 => x"5e",
          6523 => x"0c",
          6524 => x"40",
          6525 => x"fe",
          6526 => x"57",
          6527 => x"8d",
          6528 => x"fe",
          6529 => x"fe",
          6530 => x"53",
          6531 => x"52",
          6532 => x"84",
          6533 => x"06",
          6534 => x"83",
          6535 => x"08",
          6536 => x"74",
          6537 => x"82",
          6538 => x"81",
          6539 => x"16",
          6540 => x"52",
          6541 => x"3f",
          6542 => x"16",
          6543 => x"d2",
          6544 => x"fe",
          6545 => x"74",
          6546 => x"e4",
          6547 => x"e1",
          6548 => x"e4",
          6549 => x"81",
          6550 => x"33",
          6551 => x"27",
          6552 => x"80",
          6553 => x"38",
          6554 => x"57",
          6555 => x"e1",
          6556 => x"3d",
          6557 => x"05",
          6558 => x"3f",
          6559 => x"e4",
          6560 => x"8b",
          6561 => x"05",
          6562 => x"38",
          6563 => x"81",
          6564 => x"78",
          6565 => x"3d",
          6566 => x"18",
          6567 => x"7c",
          6568 => x"ff",
          6569 => x"b5",
          6570 => x"dc",
          6571 => x"ff",
          6572 => x"38",
          6573 => x"33",
          6574 => x"78",
          6575 => x"78",
          6576 => x"33",
          6577 => x"74",
          6578 => x"09",
          6579 => x"06",
          6580 => x"77",
          6581 => x"81",
          6582 => x"38",
          6583 => x"81",
          6584 => x"7b",
          6585 => x"a3",
          6586 => x"06",
          6587 => x"fe",
          6588 => x"56",
          6589 => x"80",
          6590 => x"79",
          6591 => x"2e",
          6592 => x"5a",
          6593 => x"80",
          6594 => x"ef",
          6595 => x"84",
          6596 => x"74",
          6597 => x"3d",
          6598 => x"9e",
          6599 => x"ff",
          6600 => x"86",
          6601 => x"3d",
          6602 => x"fe",
          6603 => x"f4",
          6604 => x"84",
          6605 => x"80",
          6606 => x"59",
          6607 => x"33",
          6608 => x"15",
          6609 => x"0b",
          6610 => x"ec",
          6611 => x"56",
          6612 => x"8a",
          6613 => x"b8",
          6614 => x"fe",
          6615 => x"fe",
          6616 => x"52",
          6617 => x"e4",
          6618 => x"2e",
          6619 => x"b8",
          6620 => x"16",
          6621 => x"77",
          6622 => x"74",
          6623 => x"38",
          6624 => x"81",
          6625 => x"84",
          6626 => x"ff",
          6627 => x"78",
          6628 => x"08",
          6629 => x"e5",
          6630 => x"80",
          6631 => x"2e",
          6632 => x"81",
          6633 => x"fe",
          6634 => x"57",
          6635 => x"86",
          6636 => x"bf",
          6637 => x"a0",
          6638 => x"05",
          6639 => x"38",
          6640 => x"8b",
          6641 => x"81",
          6642 => x"58",
          6643 => x"fd",
          6644 => x"33",
          6645 => x"15",
          6646 => x"6b",
          6647 => x"0b",
          6648 => x"bc",
          6649 => x"ce",
          6650 => x"54",
          6651 => x"18",
          6652 => x"b8",
          6653 => x"80",
          6654 => x"19",
          6655 => x"31",
          6656 => x"38",
          6657 => x"b1",
          6658 => x"e8",
          6659 => x"fe",
          6660 => x"57",
          6661 => x"b6",
          6662 => x"59",
          6663 => x"a1",
          6664 => x"19",
          6665 => x"33",
          6666 => x"39",
          6667 => x"05",
          6668 => x"89",
          6669 => x"08",
          6670 => x"33",
          6671 => x"15",
          6672 => x"78",
          6673 => x"5f",
          6674 => x"56",
          6675 => x"81",
          6676 => x"38",
          6677 => x"06",
          6678 => x"38",
          6679 => x"70",
          6680 => x"87",
          6681 => x"30",
          6682 => x"e4",
          6683 => x"53",
          6684 => x"38",
          6685 => x"82",
          6686 => x"74",
          6687 => x"81",
          6688 => x"75",
          6689 => x"e4",
          6690 => x"b8",
          6691 => x"84",
          6692 => x"19",
          6693 => x"78",
          6694 => x"56",
          6695 => x"90",
          6696 => x"e4",
          6697 => x"33",
          6698 => x"e4",
          6699 => x"38",
          6700 => x"39",
          6701 => x"7d",
          6702 => x"81",
          6703 => x"38",
          6704 => x"dd",
          6705 => x"84",
          6706 => x"81",
          6707 => x"d7",
          6708 => x"7b",
          6709 => x"18",
          6710 => x"33",
          6711 => x"34",
          6712 => x"08",
          6713 => x"38",
          6714 => x"15",
          6715 => x"34",
          6716 => x"ff",
          6717 => x"be",
          6718 => x"54",
          6719 => x"a1",
          6720 => x"0d",
          6721 => x"88",
          6722 => x"5f",
          6723 => x"5b",
          6724 => x"79",
          6725 => x"26",
          6726 => x"38",
          6727 => x"92",
          6728 => x"76",
          6729 => x"84",
          6730 => x"74",
          6731 => x"75",
          6732 => x"b8",
          6733 => x"52",
          6734 => x"b8",
          6735 => x"06",
          6736 => x"38",
          6737 => x"57",
          6738 => x"05",
          6739 => x"b0",
          6740 => x"38",
          6741 => x"38",
          6742 => x"38",
          6743 => x"ff",
          6744 => x"80",
          6745 => x"80",
          6746 => x"7f",
          6747 => x"89",
          6748 => x"89",
          6749 => x"80",
          6750 => x"80",
          6751 => x"74",
          6752 => x"df",
          6753 => x"79",
          6754 => x"84",
          6755 => x"83",
          6756 => x"33",
          6757 => x"57",
          6758 => x"06",
          6759 => x"05",
          6760 => x"80",
          6761 => x"83",
          6762 => x"2b",
          6763 => x"70",
          6764 => x"07",
          6765 => x"12",
          6766 => x"07",
          6767 => x"2b",
          6768 => x"0c",
          6769 => x"44",
          6770 => x"4b",
          6771 => x"27",
          6772 => x"80",
          6773 => x"70",
          6774 => x"83",
          6775 => x"82",
          6776 => x"66",
          6777 => x"4a",
          6778 => x"8a",
          6779 => x"2a",
          6780 => x"56",
          6781 => x"77",
          6782 => x"77",
          6783 => x"58",
          6784 => x"27",
          6785 => x"81",
          6786 => x"84",
          6787 => x"f5",
          6788 => x"e4",
          6789 => x"71",
          6790 => x"43",
          6791 => x"5c",
          6792 => x"05",
          6793 => x"72",
          6794 => x"2e",
          6795 => x"90",
          6796 => x"74",
          6797 => x"31",
          6798 => x"52",
          6799 => x"e4",
          6800 => x"38",
          6801 => x"dd",
          6802 => x"e4",
          6803 => x"f9",
          6804 => x"26",
          6805 => x"39",
          6806 => x"9f",
          6807 => x"81",
          6808 => x"b8",
          6809 => x"f0",
          6810 => x"81",
          6811 => x"26",
          6812 => x"06",
          6813 => x"81",
          6814 => x"5f",
          6815 => x"70",
          6816 => x"05",
          6817 => x"57",
          6818 => x"70",
          6819 => x"18",
          6820 => x"18",
          6821 => x"30",
          6822 => x"2e",
          6823 => x"be",
          6824 => x"72",
          6825 => x"4a",
          6826 => x"1c",
          6827 => x"ff",
          6828 => x"9f",
          6829 => x"51",
          6830 => x"b8",
          6831 => x"2a",
          6832 => x"56",
          6833 => x"8e",
          6834 => x"74",
          6835 => x"56",
          6836 => x"ba",
          6837 => x"f9",
          6838 => x"57",
          6839 => x"6e",
          6840 => x"39",
          6841 => x"9d",
          6842 => x"81",
          6843 => x"57",
          6844 => x"0d",
          6845 => x"62",
          6846 => x"60",
          6847 => x"8e",
          6848 => x"61",
          6849 => x"58",
          6850 => x"8b",
          6851 => x"76",
          6852 => x"81",
          6853 => x"ef",
          6854 => x"34",
          6855 => x"8d",
          6856 => x"4b",
          6857 => x"2a",
          6858 => x"61",
          6859 => x"30",
          6860 => x"78",
          6861 => x"92",
          6862 => x"ff",
          6863 => x"ff",
          6864 => x"74",
          6865 => x"34",
          6866 => x"98",
          6867 => x"ff",
          6868 => x"05",
          6869 => x"88",
          6870 => x"7e",
          6871 => x"34",
          6872 => x"84",
          6873 => x"62",
          6874 => x"a7",
          6875 => x"a1",
          6876 => x"aa",
          6877 => x"55",
          6878 => x"2a",
          6879 => x"80",
          6880 => x"05",
          6881 => x"ac",
          6882 => x"58",
          6883 => x"ff",
          6884 => x"fe",
          6885 => x"83",
          6886 => x"81",
          6887 => x"fe",
          6888 => x"e4",
          6889 => x"62",
          6890 => x"57",
          6891 => x"34",
          6892 => x"75",
          6893 => x"38",
          6894 => x"2e",
          6895 => x"76",
          6896 => x"70",
          6897 => x"59",
          6898 => x"76",
          6899 => x"57",
          6900 => x"76",
          6901 => x"79",
          6902 => x"e4",
          6903 => x"57",
          6904 => x"34",
          6905 => x"1b",
          6906 => x"38",
          6907 => x"ff",
          6908 => x"83",
          6909 => x"26",
          6910 => x"53",
          6911 => x"3f",
          6912 => x"74",
          6913 => x"db",
          6914 => x"38",
          6915 => x"8a",
          6916 => x"38",
          6917 => x"83",
          6918 => x"38",
          6919 => x"70",
          6920 => x"78",
          6921 => x"aa",
          6922 => x"78",
          6923 => x"81",
          6924 => x"05",
          6925 => x"43",
          6926 => x"fc",
          6927 => x"34",
          6928 => x"07",
          6929 => x"b8",
          6930 => x"61",
          6931 => x"c7",
          6932 => x"34",
          6933 => x"05",
          6934 => x"62",
          6935 => x"05",
          6936 => x"83",
          6937 => x"7e",
          6938 => x"78",
          6939 => x"f1",
          6940 => x"f7",
          6941 => x"51",
          6942 => x"b8",
          6943 => x"e4",
          6944 => x"0d",
          6945 => x"f9",
          6946 => x"5c",
          6947 => x"91",
          6948 => x"22",
          6949 => x"74",
          6950 => x"56",
          6951 => x"57",
          6952 => x"75",
          6953 => x"fc",
          6954 => x"10",
          6955 => x"5e",
          6956 => x"e4",
          6957 => x"fd",
          6958 => x"38",
          6959 => x"e4",
          6960 => x"38",
          6961 => x"5b",
          6962 => x"c8",
          6963 => x"2e",
          6964 => x"39",
          6965 => x"2a",
          6966 => x"90",
          6967 => x"75",
          6968 => x"34",
          6969 => x"05",
          6970 => x"a1",
          6971 => x"61",
          6972 => x"05",
          6973 => x"a5",
          6974 => x"61",
          6975 => x"75",
          6976 => x"05",
          6977 => x"61",
          6978 => x"34",
          6979 => x"b1",
          6980 => x"80",
          6981 => x"80",
          6982 => x"05",
          6983 => x"e4",
          6984 => x"05",
          6985 => x"34",
          6986 => x"cd",
          6987 => x"76",
          6988 => x"55",
          6989 => x"54",
          6990 => x"be",
          6991 => x"08",
          6992 => x"05",
          6993 => x"76",
          6994 => x"52",
          6995 => x"c3",
          6996 => x"9f",
          6997 => x"f8",
          6998 => x"81",
          6999 => x"05",
          7000 => x"84",
          7001 => x"ff",
          7002 => x"05",
          7003 => x"61",
          7004 => x"34",
          7005 => x"39",
          7006 => x"79",
          7007 => x"61",
          7008 => x"57",
          7009 => x"60",
          7010 => x"5e",
          7011 => x"81",
          7012 => x"81",
          7013 => x"80",
          7014 => x"f2",
          7015 => x"61",
          7016 => x"83",
          7017 => x"7a",
          7018 => x"2a",
          7019 => x"7a",
          7020 => x"05",
          7021 => x"83",
          7022 => x"05",
          7023 => x"76",
          7024 => x"83",
          7025 => x"ff",
          7026 => x"53",
          7027 => x"3f",
          7028 => x"79",
          7029 => x"57",
          7030 => x"7e",
          7031 => x"05",
          7032 => x"38",
          7033 => x"54",
          7034 => x"9a",
          7035 => x"06",
          7036 => x"8d",
          7037 => x"05",
          7038 => x"2e",
          7039 => x"80",
          7040 => x"76",
          7041 => x"3d",
          7042 => x"84",
          7043 => x"8a",
          7044 => x"56",
          7045 => x"08",
          7046 => x"75",
          7047 => x"8e",
          7048 => x"88",
          7049 => x"3d",
          7050 => x"52",
          7051 => x"74",
          7052 => x"9f",
          7053 => x"1c",
          7054 => x"39",
          7055 => x"ff",
          7056 => x"ff",
          7057 => x"cc",
          7058 => x"05",
          7059 => x"38",
          7060 => x"2e",
          7061 => x"24",
          7062 => x"05",
          7063 => x"55",
          7064 => x"18",
          7065 => x"55",
          7066 => x"ff",
          7067 => x"52",
          7068 => x"84",
          7069 => x"2e",
          7070 => x"0c",
          7071 => x"b0",
          7072 => x"76",
          7073 => x"7b",
          7074 => x"2a",
          7075 => x"a5",
          7076 => x"3f",
          7077 => x"0c",
          7078 => x"75",
          7079 => x"53",
          7080 => x"38",
          7081 => x"84",
          7082 => x"83",
          7083 => x"b5",
          7084 => x"80",
          7085 => x"51",
          7086 => x"70",
          7087 => x"80",
          7088 => x"e6",
          7089 => x"39",
          7090 => x"84",
          7091 => x"04",
          7092 => x"02",
          7093 => x"80",
          7094 => x"70",
          7095 => x"3d",
          7096 => x"81",
          7097 => x"e9",
          7098 => x"70",
          7099 => x"3d",
          7100 => x"70",
          7101 => x"70",
          7102 => x"56",
          7103 => x"38",
          7104 => x"71",
          7105 => x"07",
          7106 => x"71",
          7107 => x"88",
          7108 => x"14",
          7109 => x"71",
          7110 => x"82",
          7111 => x"80",
          7112 => x"52",
          7113 => x"70",
          7114 => x"04",
          7115 => x"71",
          7116 => x"83",
          7117 => x"c7",
          7118 => x"57",
          7119 => x"16",
          7120 => x"f1",
          7121 => x"06",
          7122 => x"83",
          7123 => x"d0",
          7124 => x"51",
          7125 => x"ff",
          7126 => x"70",
          7127 => x"b9",
          7128 => x"71",
          7129 => x"52",
          7130 => x"10",
          7131 => x"ef",
          7132 => x"ff",
          7133 => x"ff",
          7134 => x"8b",
          7135 => x"75",
          7136 => x"5f",
          7137 => x"49",
          7138 => x"33",
          7139 => x"1d",
          7140 => x"07",
          7141 => x"f1",
          7142 => x"db",
          7143 => x"c5",
          7144 => x"bf",
          7145 => x"59",
          7146 => x"59",
          7147 => x"59",
          7148 => x"59",
          7149 => x"59",
          7150 => x"59",
          7151 => x"59",
          7152 => x"59",
          7153 => x"59",
          7154 => x"59",
          7155 => x"59",
          7156 => x"59",
          7157 => x"59",
          7158 => x"59",
          7159 => x"59",
          7160 => x"59",
          7161 => x"59",
          7162 => x"59",
          7163 => x"59",
          7164 => x"59",
          7165 => x"59",
          7166 => x"59",
          7167 => x"59",
          7168 => x"59",
          7169 => x"59",
          7170 => x"59",
          7171 => x"59",
          7172 => x"59",
          7173 => x"59",
          7174 => x"07",
          7175 => x"59",
          7176 => x"a8",
          7177 => x"2c",
          7178 => x"59",
          7179 => x"59",
          7180 => x"59",
          7181 => x"59",
          7182 => x"59",
          7183 => x"59",
          7184 => x"59",
          7185 => x"59",
          7186 => x"59",
          7187 => x"59",
          7188 => x"59",
          7189 => x"59",
          7190 => x"59",
          7191 => x"59",
          7192 => x"59",
          7193 => x"59",
          7194 => x"59",
          7195 => x"59",
          7196 => x"59",
          7197 => x"59",
          7198 => x"59",
          7199 => x"59",
          7200 => x"59",
          7201 => x"59",
          7202 => x"59",
          7203 => x"59",
          7204 => x"ab",
          7205 => x"59",
          7206 => x"59",
          7207 => x"59",
          7208 => x"59",
          7209 => x"63",
          7210 => x"59",
          7211 => x"59",
          7212 => x"47",
          7213 => x"12",
          7214 => x"36",
          7215 => x"4e",
          7216 => x"86",
          7217 => x"f0",
          7218 => x"10",
          7219 => x"8a",
          7220 => x"ba",
          7221 => x"01",
          7222 => x"cd",
          7223 => x"fa",
          7224 => x"cd",
          7225 => x"01",
          7226 => x"63",
          7227 => x"6b",
          7228 => x"a9",
          7229 => x"2b",
          7230 => x"44",
          7231 => x"51",
          7232 => x"51",
          7233 => x"51",
          7234 => x"2a",
          7235 => x"51",
          7236 => x"51",
          7237 => x"51",
          7238 => x"51",
          7239 => x"51",
          7240 => x"51",
          7241 => x"51",
          7242 => x"51",
          7243 => x"51",
          7244 => x"51",
          7245 => x"51",
          7246 => x"57",
          7247 => x"31",
          7248 => x"1f",
          7249 => x"74",
          7250 => x"74",
          7251 => x"79",
          7252 => x"83",
          7253 => x"d8",
          7254 => x"b7",
          7255 => x"5b",
          7256 => x"66",
          7257 => x"8f",
          7258 => x"4b",
          7259 => x"f1",
          7260 => x"cb",
          7261 => x"78",
          7262 => x"78",
          7263 => x"78",
          7264 => x"94",
          7265 => x"59",
          7266 => x"78",
          7267 => x"78",
          7268 => x"78",
          7269 => x"78",
          7270 => x"78",
          7271 => x"78",
          7272 => x"78",
          7273 => x"78",
          7274 => x"78",
          7275 => x"16",
          7276 => x"78",
          7277 => x"b9",
          7278 => x"6a",
          7279 => x"78",
          7280 => x"78",
          7281 => x"78",
          7282 => x"9b",
          7283 => x"10",
          7284 => x"10",
          7285 => x"10",
          7286 => x"10",
          7287 => x"10",
          7288 => x"10",
          7289 => x"10",
          7290 => x"10",
          7291 => x"10",
          7292 => x"10",
          7293 => x"10",
          7294 => x"10",
          7295 => x"10",
          7296 => x"10",
          7297 => x"ad",
          7298 => x"e2",
          7299 => x"bd",
          7300 => x"6d",
          7301 => x"10",
          7302 => x"3d",
          7303 => x"19",
          7304 => x"78",
          7305 => x"56",
          7306 => x"10",
          7307 => x"6a",
          7308 => x"c6",
          7309 => x"c6",
          7310 => x"c6",
          7311 => x"c6",
          7312 => x"c6",
          7313 => x"c6",
          7314 => x"e8",
          7315 => x"c6",
          7316 => x"c6",
          7317 => x"c6",
          7318 => x"c6",
          7319 => x"3f",
          7320 => x"56",
          7321 => x"28",
          7322 => x"c1",
          7323 => x"aa",
          7324 => x"94",
          7325 => x"7d",
          7326 => x"01",
          7327 => x"fd",
          7328 => x"fd",
          7329 => x"fd",
          7330 => x"fd",
          7331 => x"fd",
          7332 => x"fd",
          7333 => x"0d",
          7334 => x"fd",
          7335 => x"fd",
          7336 => x"fd",
          7337 => x"fd",
          7338 => x"fd",
          7339 => x"fd",
          7340 => x"fd",
          7341 => x"fd",
          7342 => x"fd",
          7343 => x"fd",
          7344 => x"fd",
          7345 => x"fd",
          7346 => x"fd",
          7347 => x"fd",
          7348 => x"fd",
          7349 => x"fd",
          7350 => x"fd",
          7351 => x"fd",
          7352 => x"fd",
          7353 => x"fd",
          7354 => x"17",
          7355 => x"fd",
          7356 => x"fd",
          7357 => x"fd",
          7358 => x"fd",
          7359 => x"fd",
          7360 => x"e1",
          7361 => x"b8",
          7362 => x"fd",
          7363 => x"fd",
          7364 => x"ff",
          7365 => x"fd",
          7366 => x"0f",
          7367 => x"fd",
          7368 => x"fd",
          7369 => x"fd",
          7370 => x"17",
          7371 => x"00",
          7372 => x"00",
          7373 => x"00",
          7374 => x"00",
          7375 => x"00",
          7376 => x"00",
          7377 => x"00",
          7378 => x"00",
          7379 => x"00",
          7380 => x"00",
          7381 => x"00",
          7382 => x"00",
          7383 => x"6c",
          7384 => x"00",
          7385 => x"00",
          7386 => x"00",
          7387 => x"00",
          7388 => x"00",
          7389 => x"00",
          7390 => x"00",
          7391 => x"00",
          7392 => x"00",
          7393 => x"6e",
          7394 => x"6f",
          7395 => x"61",
          7396 => x"69",
          7397 => x"74",
          7398 => x"20",
          7399 => x"65",
          7400 => x"2e",
          7401 => x"75",
          7402 => x"74",
          7403 => x"2e",
          7404 => x"65",
          7405 => x"6b",
          7406 => x"65",
          7407 => x"65",
          7408 => x"63",
          7409 => x"64",
          7410 => x"6d",
          7411 => x"74",
          7412 => x"63",
          7413 => x"6c",
          7414 => x"79",
          7415 => x"75",
          7416 => x"69",
          7417 => x"6b",
          7418 => x"61",
          7419 => x"00",
          7420 => x"75",
          7421 => x"20",
          7422 => x"2e",
          7423 => x"69",
          7424 => x"20",
          7425 => x"65",
          7426 => x"65",
          7427 => x"20",
          7428 => x"2e",
          7429 => x"65",
          7430 => x"79",
          7431 => x"2e",
          7432 => x"65",
          7433 => x"65",
          7434 => x"61",
          7435 => x"65",
          7436 => x"00",
          7437 => x"20",
          7438 => x"00",
          7439 => x"20",
          7440 => x"00",
          7441 => x"74",
          7442 => x"00",
          7443 => x"6c",
          7444 => x"00",
          7445 => x"72",
          7446 => x"63",
          7447 => x"00",
          7448 => x"74",
          7449 => x"74",
          7450 => x"74",
          7451 => x"0a",
          7452 => x"64",
          7453 => x"6c",
          7454 => x"00",
          7455 => x"00",
          7456 => x"00",
          7457 => x"58",
          7458 => x"20",
          7459 => x"00",
          7460 => x"25",
          7461 => x"30",
          7462 => x"00",
          7463 => x"00",
          7464 => x"65",
          7465 => x"20",
          7466 => x"2a",
          7467 => x"20",
          7468 => x"70",
          7469 => x"65",
          7470 => x"54",
          7471 => x"74",
          7472 => x"00",
          7473 => x"58",
          7474 => x"75",
          7475 => x"54",
          7476 => x"74",
          7477 => x"00",
          7478 => x"58",
          7479 => x"75",
          7480 => x"54",
          7481 => x"74",
          7482 => x"00",
          7483 => x"44",
          7484 => x"75",
          7485 => x"20",
          7486 => x"70",
          7487 => x"65",
          7488 => x"72",
          7489 => x"74",
          7490 => x"74",
          7491 => x"00",
          7492 => x"67",
          7493 => x"2e",
          7494 => x"6f",
          7495 => x"74",
          7496 => x"5f",
          7497 => x"00",
          7498 => x"74",
          7499 => x"61",
          7500 => x"20",
          7501 => x"20",
          7502 => x"69",
          7503 => x"75",
          7504 => x"00",
          7505 => x"5c",
          7506 => x"00",
          7507 => x"6d",
          7508 => x"00",
          7509 => x"00",
          7510 => x"25",
          7511 => x"00",
          7512 => x"62",
          7513 => x"2e",
          7514 => x"74",
          7515 => x"61",
          7516 => x"69",
          7517 => x"00",
          7518 => x"20",
          7519 => x"25",
          7520 => x"2e",
          7521 => x"6c",
          7522 => x"65",
          7523 => x"28",
          7524 => x"00",
          7525 => x"6e",
          7526 => x"40",
          7527 => x"2e",
          7528 => x"6c",
          7529 => x"2d",
          7530 => x"6c",
          7531 => x"00",
          7532 => x"6e",
          7533 => x"00",
          7534 => x"30",
          7535 => x"38",
          7536 => x"29",
          7537 => x"79",
          7538 => x"00",
          7539 => x"30",
          7540 => x"61",
          7541 => x"2e",
          7542 => x"70",
          7543 => x"00",
          7544 => x"74",
          7545 => x"5c",
          7546 => x"00",
          7547 => x"65",
          7548 => x"64",
          7549 => x"74",
          7550 => x"73",
          7551 => x"64",
          7552 => x"00",
          7553 => x"64",
          7554 => x"25",
          7555 => x"00",
          7556 => x"66",
          7557 => x"6f",
          7558 => x"65",
          7559 => x"6d",
          7560 => x"65",
          7561 => x"72",
          7562 => x"00",
          7563 => x"20",
          7564 => x"65",
          7565 => x"64",
          7566 => x"25",
          7567 => x"00",
          7568 => x"20",
          7569 => x"53",
          7570 => x"64",
          7571 => x"25",
          7572 => x"00",
          7573 => x"63",
          7574 => x"20",
          7575 => x"20",
          7576 => x"25",
          7577 => x"00",
          7578 => x"00",
          7579 => x"20",
          7580 => x"20",
          7581 => x"20",
          7582 => x"25",
          7583 => x"00",
          7584 => x"74",
          7585 => x"6b",
          7586 => x"20",
          7587 => x"25",
          7588 => x"48",
          7589 => x"20",
          7590 => x"65",
          7591 => x"43",
          7592 => x"65",
          7593 => x"30",
          7594 => x"00",
          7595 => x"41",
          7596 => x"20",
          7597 => x"20",
          7598 => x"25",
          7599 => x"48",
          7600 => x"20",
          7601 => x"20",
          7602 => x"20",
          7603 => x"00",
          7604 => x"49",
          7605 => x"20",
          7606 => x"45",
          7607 => x"00",
          7608 => x"52",
          7609 => x"43",
          7610 => x"3d",
          7611 => x"00",
          7612 => x"45",
          7613 => x"54",
          7614 => x"3d",
          7615 => x"00",
          7616 => x"43",
          7617 => x"44",
          7618 => x"3d",
          7619 => x"00",
          7620 => x"20",
          7621 => x"25",
          7622 => x"58",
          7623 => x"20",
          7624 => x"20",
          7625 => x"3a",
          7626 => x"00",
          7627 => x"4e",
          7628 => x"25",
          7629 => x"58",
          7630 => x"20",
          7631 => x"20",
          7632 => x"3a",
          7633 => x"00",
          7634 => x"53",
          7635 => x"25",
          7636 => x"58",
          7637 => x"72",
          7638 => x"63",
          7639 => x"00",
          7640 => x"00",
          7641 => x"00",
          7642 => x"00",
          7643 => x"00",
          7644 => x"00",
          7645 => x"48",
          7646 => x"02",
          7647 => x"00",
          7648 => x"40",
          7649 => x"04",
          7650 => x"00",
          7651 => x"38",
          7652 => x"06",
          7653 => x"00",
          7654 => x"30",
          7655 => x"01",
          7656 => x"00",
          7657 => x"28",
          7658 => x"0b",
          7659 => x"00",
          7660 => x"20",
          7661 => x"0a",
          7662 => x"00",
          7663 => x"18",
          7664 => x"0c",
          7665 => x"00",
          7666 => x"10",
          7667 => x"0f",
          7668 => x"00",
          7669 => x"08",
          7670 => x"10",
          7671 => x"00",
          7672 => x"00",
          7673 => x"12",
          7674 => x"00",
          7675 => x"f8",
          7676 => x"14",
          7677 => x"00",
          7678 => x"00",
          7679 => x"00",
          7680 => x"7e",
          7681 => x"7e",
          7682 => x"7e",
          7683 => x"7e",
          7684 => x"00",
          7685 => x"00",
          7686 => x"00",
          7687 => x"00",
          7688 => x"00",
          7689 => x"6e",
          7690 => x"2f",
          7691 => x"68",
          7692 => x"66",
          7693 => x"73",
          7694 => x"00",
          7695 => x"00",
          7696 => x"00",
          7697 => x"6c",
          7698 => x"00",
          7699 => x"74",
          7700 => x"20",
          7701 => x"74",
          7702 => x"65",
          7703 => x"2e",
          7704 => x"0a",
          7705 => x"7e",
          7706 => x"00",
          7707 => x"00",
          7708 => x"30",
          7709 => x"31",
          7710 => x"32",
          7711 => x"33",
          7712 => x"34",
          7713 => x"35",
          7714 => x"37",
          7715 => x"38",
          7716 => x"39",
          7717 => x"30",
          7718 => x"7e",
          7719 => x"7e",
          7720 => x"00",
          7721 => x"00",
          7722 => x"00",
          7723 => x"2c",
          7724 => x"64",
          7725 => x"78",
          7726 => x"64",
          7727 => x"25",
          7728 => x"2c",
          7729 => x"00",
          7730 => x"00",
          7731 => x"00",
          7732 => x"64",
          7733 => x"6f",
          7734 => x"6f",
          7735 => x"25",
          7736 => x"78",
          7737 => x"25",
          7738 => x"78",
          7739 => x"25",
          7740 => x"00",
          7741 => x"20",
          7742 => x"2e",
          7743 => x"00",
          7744 => x"7f",
          7745 => x"3d",
          7746 => x"00",
          7747 => x"00",
          7748 => x"53",
          7749 => x"4e",
          7750 => x"46",
          7751 => x"00",
          7752 => x"20",
          7753 => x"32",
          7754 => x"fc",
          7755 => x"00",
          7756 => x"07",
          7757 => x"1c",
          7758 => x"41",
          7759 => x"49",
          7760 => x"4f",
          7761 => x"9b",
          7762 => x"55",
          7763 => x"ab",
          7764 => x"b3",
          7765 => x"bb",
          7766 => x"c3",
          7767 => x"cb",
          7768 => x"d3",
          7769 => x"db",
          7770 => x"e3",
          7771 => x"eb",
          7772 => x"f3",
          7773 => x"fb",
          7774 => x"3b",
          7775 => x"3a",
          7776 => x"00",
          7777 => x"40",
          7778 => x"00",
          7779 => x"08",
          7780 => x"00",
          7781 => x"e2",
          7782 => x"e7",
          7783 => x"ef",
          7784 => x"c5",
          7785 => x"f4",
          7786 => x"f9",
          7787 => x"a2",
          7788 => x"92",
          7789 => x"fa",
          7790 => x"ba",
          7791 => x"bd",
          7792 => x"bb",
          7793 => x"02",
          7794 => x"56",
          7795 => x"57",
          7796 => x"10",
          7797 => x"1c",
          7798 => x"5f",
          7799 => x"66",
          7800 => x"67",
          7801 => x"59",
          7802 => x"6b",
          7803 => x"88",
          7804 => x"80",
          7805 => x"c0",
          7806 => x"c4",
          7807 => x"b4",
          7808 => x"29",
          7809 => x"64",
          7810 => x"48",
          7811 => x"1a",
          7812 => x"a0",
          7813 => x"17",
          7814 => x"01",
          7815 => x"32",
          7816 => x"4a",
          7817 => x"80",
          7818 => x"82",
          7819 => x"86",
          7820 => x"8a",
          7821 => x"8e",
          7822 => x"91",
          7823 => x"96",
          7824 => x"3d",
          7825 => x"20",
          7826 => x"a2",
          7827 => x"a6",
          7828 => x"aa",
          7829 => x"ae",
          7830 => x"b2",
          7831 => x"b5",
          7832 => x"ba",
          7833 => x"be",
          7834 => x"c2",
          7835 => x"c4",
          7836 => x"ca",
          7837 => x"10",
          7838 => x"de",
          7839 => x"f1",
          7840 => x"28",
          7841 => x"09",
          7842 => x"3d",
          7843 => x"41",
          7844 => x"53",
          7845 => x"55",
          7846 => x"8f",
          7847 => x"5d",
          7848 => x"61",
          7849 => x"65",
          7850 => x"96",
          7851 => x"6d",
          7852 => x"71",
          7853 => x"9f",
          7854 => x"79",
          7855 => x"64",
          7856 => x"81",
          7857 => x"85",
          7858 => x"44",
          7859 => x"8d",
          7860 => x"91",
          7861 => x"fd",
          7862 => x"04",
          7863 => x"8a",
          7864 => x"02",
          7865 => x"08",
          7866 => x"8e",
          7867 => x"f2",
          7868 => x"f4",
          7869 => x"f7",
          7870 => x"30",
          7871 => x"60",
          7872 => x"c1",
          7873 => x"c0",
          7874 => x"26",
          7875 => x"01",
          7876 => x"a0",
          7877 => x"10",
          7878 => x"30",
          7879 => x"51",
          7880 => x"5b",
          7881 => x"5f",
          7882 => x"0e",
          7883 => x"c9",
          7884 => x"db",
          7885 => x"eb",
          7886 => x"08",
          7887 => x"08",
          7888 => x"b9",
          7889 => x"01",
          7890 => x"e0",
          7891 => x"ec",
          7892 => x"4e",
          7893 => x"10",
          7894 => x"d0",
          7895 => x"60",
          7896 => x"75",
          7897 => x"00",
          7898 => x"00",
          7899 => x"58",
          7900 => x"00",
          7901 => x"60",
          7902 => x"00",
          7903 => x"68",
          7904 => x"00",
          7905 => x"70",
          7906 => x"00",
          7907 => x"78",
          7908 => x"00",
          7909 => x"80",
          7910 => x"00",
          7911 => x"88",
          7912 => x"00",
          7913 => x"90",
          7914 => x"00",
          7915 => x"98",
          7916 => x"00",
          7917 => x"a0",
          7918 => x"00",
          7919 => x"a4",
          7920 => x"00",
          7921 => x"a8",
          7922 => x"00",
          7923 => x"ac",
          7924 => x"00",
          7925 => x"b0",
          7926 => x"00",
          7927 => x"b4",
          7928 => x"00",
          7929 => x"b8",
          7930 => x"00",
          7931 => x"bc",
          7932 => x"00",
          7933 => x"c4",
          7934 => x"00",
          7935 => x"c8",
          7936 => x"00",
          7937 => x"d0",
          7938 => x"00",
          7939 => x"d8",
          7940 => x"00",
          7941 => x"e0",
          7942 => x"00",
          7943 => x"e8",
          7944 => x"00",
          7945 => x"ec",
          7946 => x"00",
          7947 => x"f0",
          7948 => x"00",
          7949 => x"f8",
          7950 => x"00",
          7951 => x"00",
          7952 => x"00",
          7953 => x"08",
          7954 => x"00",
          7955 => x"00",
          7956 => x"ff",
          7957 => x"ff",
          7958 => x"ff",
          7959 => x"00",
          7960 => x"ff",
          7961 => x"00",
          7962 => x"00",
          7963 => x"00",
          7964 => x"00",
          7965 => x"01",
          7966 => x"00",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"fd",
          7983 => x"5b",
          7984 => x"74",
          7985 => x"6c",
          7986 => x"64",
          7987 => x"34",
          7988 => x"20",
          7989 => x"f4",
          7990 => x"f0",
          7991 => x"83",
          7992 => x"fd",
          7993 => x"5b",
          7994 => x"54",
          7995 => x"4c",
          7996 => x"44",
          7997 => x"34",
          7998 => x"20",
          7999 => x"f4",
          8000 => x"f0",
          8001 => x"83",
          8002 => x"fd",
          8003 => x"7b",
          8004 => x"54",
          8005 => x"4c",
          8006 => x"44",
          8007 => x"24",
          8008 => x"20",
          8009 => x"e1",
          8010 => x"f0",
          8011 => x"88",
          8012 => x"fa",
          8013 => x"1b",
          8014 => x"14",
          8015 => x"0c",
          8016 => x"04",
          8017 => x"f0",
          8018 => x"f0",
          8019 => x"f0",
          8020 => x"f0",
          8021 => x"83",
          8022 => x"c9",
          8023 => x"b3",
          8024 => x"31",
          8025 => x"56",
          8026 => x"48",
          8027 => x"3b",
          8028 => x"00",
          8029 => x"c1",
          8030 => x"f0",
          8031 => x"83",
          8032 => x"00",
          8033 => x"00",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"00",
          8045 => x"00",
          8046 => x"cc",
          8047 => x"d4",
          8048 => x"d8",
          8049 => x"dc",
          8050 => x"e0",
          8051 => x"e4",
          8052 => x"ec",
          8053 => x"f4",
          8054 => x"fc",
          8055 => x"04",
          8056 => x"0c",
          8057 => x"14",
          8058 => x"1c",
          8059 => x"24",
          8060 => x"2c",
          8061 => x"34",
          8062 => x"3c",
          8063 => x"44",
          8064 => x"48",
          8065 => x"50",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"19",
          9067 => x"00",
          9068 => x"f7",
          9069 => x"ff",
          9070 => x"e2",
          9071 => x"f4",
          9072 => x"67",
          9073 => x"2d",
          9074 => x"27",
          9075 => x"49",
          9076 => x"07",
          9077 => x"0f",
          9078 => x"17",
          9079 => x"3c",
          9080 => x"87",
          9081 => x"8f",
          9082 => x"97",
          9083 => x"c0",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"01",
          9100 => x"01",
        others => X"00"
    );

    shared variable RAM5 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"88",
             5 => x"88",
             6 => x"00",
             7 => x"00",
             8 => x"06",
             9 => x"2a",
            10 => x"00",
            11 => x"00",
            12 => x"ff",
            13 => x"05",
            14 => x"ff",
            15 => x"04",
            16 => x"73",
            17 => x"73",
            18 => x"04",
            19 => x"00",
            20 => x"07",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"81",
            25 => x"0a",
            26 => x"81",
            27 => x"00",
            28 => x"07",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"00",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"51",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"05",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"06",
            49 => x"ff",
            50 => x"00",
            51 => x"00",
            52 => x"73",
            53 => x"83",
            54 => x"0c",
            55 => x"00",
            56 => x"09",
            57 => x"06",
            58 => x"00",
            59 => x"00",
            60 => x"09",
            61 => x"81",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"53",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"09",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"06",
            77 => x"10",
            78 => x"00",
            79 => x"00",
            80 => x"83",
            81 => x"05",
            82 => x"04",
            83 => x"00",
            84 => x"75",
            85 => x"50",
            86 => x"0c",
            87 => x"00",
            88 => x"75",
            89 => x"50",
            90 => x"0c",
            91 => x"00",
            92 => x"06",
            93 => x"71",
            94 => x"05",
            95 => x"00",
            96 => x"06",
            97 => x"54",
            98 => x"ff",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"05",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"53",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"0b",
           134 => x"a6",
           135 => x"0b",
           136 => x"0b",
           137 => x"e6",
           138 => x"0b",
           139 => x"0b",
           140 => x"a6",
           141 => x"0b",
           142 => x"0b",
           143 => x"e8",
           144 => x"0b",
           145 => x"0b",
           146 => x"ac",
           147 => x"0b",
           148 => x"0b",
           149 => x"f0",
           150 => x"0b",
           151 => x"0b",
           152 => x"b4",
           153 => x"0b",
           154 => x"0b",
           155 => x"f8",
           156 => x"0b",
           157 => x"0b",
           158 => x"bc",
           159 => x"0b",
           160 => x"0b",
           161 => x"80",
           162 => x"0b",
           163 => x"0b",
           164 => x"c4",
           165 => x"0b",
           166 => x"0b",
           167 => x"88",
           168 => x"0b",
           169 => x"0b",
           170 => x"cb",
           171 => x"0b",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"b8",
           193 => x"b8",
           194 => x"84",
           195 => x"b8",
           196 => x"84",
           197 => x"b8",
           198 => x"84",
           199 => x"b8",
           200 => x"84",
           201 => x"b8",
           202 => x"84",
           203 => x"b8",
           204 => x"84",
           205 => x"b8",
           206 => x"84",
           207 => x"b8",
           208 => x"84",
           209 => x"b8",
           210 => x"84",
           211 => x"b8",
           212 => x"84",
           213 => x"b8",
           214 => x"84",
           215 => x"b8",
           216 => x"84",
           217 => x"84",
           218 => x"04",
           219 => x"2d",
           220 => x"90",
           221 => x"8d",
           222 => x"80",
           223 => x"d3",
           224 => x"c0",
           225 => x"82",
           226 => x"80",
           227 => x"0c",
           228 => x"08",
           229 => x"f0",
           230 => x"f0",
           231 => x"b8",
           232 => x"b8",
           233 => x"84",
           234 => x"84",
           235 => x"04",
           236 => x"2d",
           237 => x"90",
           238 => x"f6",
           239 => x"80",
           240 => x"f1",
           241 => x"c0",
           242 => x"82",
           243 => x"80",
           244 => x"0c",
           245 => x"08",
           246 => x"f0",
           247 => x"f0",
           248 => x"b8",
           249 => x"b8",
           250 => x"84",
           251 => x"84",
           252 => x"04",
           253 => x"2d",
           254 => x"90",
           255 => x"ec",
           256 => x"80",
           257 => x"94",
           258 => x"c0",
           259 => x"82",
           260 => x"80",
           261 => x"0c",
           262 => x"08",
           263 => x"f0",
           264 => x"f0",
           265 => x"b8",
           266 => x"b8",
           267 => x"84",
           268 => x"84",
           269 => x"04",
           270 => x"2d",
           271 => x"90",
           272 => x"d8",
           273 => x"80",
           274 => x"c6",
           275 => x"c0",
           276 => x"83",
           277 => x"80",
           278 => x"0c",
           279 => x"08",
           280 => x"f0",
           281 => x"f0",
           282 => x"b8",
           283 => x"b8",
           284 => x"84",
           285 => x"84",
           286 => x"04",
           287 => x"2d",
           288 => x"90",
           289 => x"8f",
           290 => x"80",
           291 => x"d1",
           292 => x"c0",
           293 => x"80",
           294 => x"80",
           295 => x"0c",
           296 => x"80",
           297 => x"0c",
           298 => x"08",
           299 => x"f0",
           300 => x"f0",
           301 => x"b8",
           302 => x"b8",
           303 => x"84",
           304 => x"84",
           305 => x"04",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"81",
           311 => x"05",
           312 => x"72",
           313 => x"72",
           314 => x"72",
           315 => x"10",
           316 => x"53",
           317 => x"d4",
           318 => x"84",
           319 => x"ec",
           320 => x"04",
           321 => x"70",
           322 => x"52",
           323 => x"3f",
           324 => x"78",
           325 => x"81",
           326 => x"55",
           327 => x"81",
           328 => x"74",
           329 => x"9f",
           330 => x"74",
           331 => x"38",
           332 => x"e4",
           333 => x"2e",
           334 => x"70",
           335 => x"8a",
           336 => x"2a",
           337 => x"cb",
           338 => x"84",
           339 => x"80",
           340 => x"0d",
           341 => x"02",
           342 => x"fe",
           343 => x"7e",
           344 => x"3f",
           345 => x"3d",
           346 => x"88",
           347 => x"3f",
           348 => x"61",
           349 => x"8c",
           350 => x"2a",
           351 => x"ff",
           352 => x"80",
           353 => x"2e",
           354 => x"06",
           355 => x"38",
           356 => x"a3",
           357 => x"80",
           358 => x"72",
           359 => x"70",
           360 => x"80",
           361 => x"5b",
           362 => x"8c",
           363 => x"0c",
           364 => x"54",
           365 => x"70",
           366 => x"81",
           367 => x"98",
           368 => x"79",
           369 => x"53",
           370 => x"58",
           371 => x"39",
           372 => x"38",
           373 => x"7c",
           374 => x"ff",
           375 => x"af",
           376 => x"38",
           377 => x"81",
           378 => x"70",
           379 => x"e0",
           380 => x"38",
           381 => x"54",
           382 => x"59",
           383 => x"52",
           384 => x"33",
           385 => x"c7",
           386 => x"88",
           387 => x"7d",
           388 => x"54",
           389 => x"51",
           390 => x"81",
           391 => x"df",
           392 => x"38",
           393 => x"74",
           394 => x"52",
           395 => x"e4",
           396 => x"38",
           397 => x"7b",
           398 => x"8f",
           399 => x"80",
           400 => x"7a",
           401 => x"73",
           402 => x"80",
           403 => x"90",
           404 => x"29",
           405 => x"2c",
           406 => x"54",
           407 => x"98",
           408 => x"78",
           409 => x"ff",
           410 => x"2a",
           411 => x"73",
           412 => x"31",
           413 => x"80",
           414 => x"85",
           415 => x"54",
           416 => x"81",
           417 => x"85",
           418 => x"38",
           419 => x"38",
           420 => x"80",
           421 => x"80",
           422 => x"2c",
           423 => x"38",
           424 => x"77",
           425 => x"80",
           426 => x"73",
           427 => x"53",
           428 => x"81",
           429 => x"70",
           430 => x"25",
           431 => x"ef",
           432 => x"81",
           433 => x"55",
           434 => x"87",
           435 => x"80",
           436 => x"2e",
           437 => x"81",
           438 => x"e2",
           439 => x"38",
           440 => x"5e",
           441 => x"2e",
           442 => x"06",
           443 => x"77",
           444 => x"80",
           445 => x"80",
           446 => x"a0",
           447 => x"90",
           448 => x"58",
           449 => x"39",
           450 => x"57",
           451 => x"7e",
           452 => x"55",
           453 => x"05",
           454 => x"33",
           455 => x"80",
           456 => x"90",
           457 => x"5f",
           458 => x"55",
           459 => x"80",
           460 => x"90",
           461 => x"fe",
           462 => x"f7",
           463 => x"ff",
           464 => x"ff",
           465 => x"70",
           466 => x"3f",
           467 => x"ff",
           468 => x"2e",
           469 => x"81",
           470 => x"e2",
           471 => x"0a",
           472 => x"80",
           473 => x"56",
           474 => x"06",
           475 => x"fe",
           476 => x"08",
           477 => x"24",
           478 => x"06",
           479 => x"39",
           480 => x"76",
           481 => x"88",
           482 => x"76",
           483 => x"60",
           484 => x"56",
           485 => x"75",
           486 => x"08",
           487 => x"90",
           488 => x"fe",
           489 => x"33",
           490 => x"ff",
           491 => x"77",
           492 => x"81",
           493 => x"84",
           494 => x"78",
           495 => x"39",
           496 => x"5b",
           497 => x"77",
           498 => x"80",
           499 => x"80",
           500 => x"a0",
           501 => x"52",
           502 => x"2e",
           503 => x"52",
           504 => x"2a",
           505 => x"8c",
           506 => x"78",
           507 => x"7d",
           508 => x"73",
           509 => x"52",
           510 => x"06",
           511 => x"ff",
           512 => x"51",
           513 => x"7a",
           514 => x"39",
           515 => x"2c",
           516 => x"ab",
           517 => x"52",
           518 => x"39",
           519 => x"84",
           520 => x"78",
           521 => x"f3",
           522 => x"83",
           523 => x"99",
           524 => x"08",
           525 => x"3f",
           526 => x"78",
           527 => x"85",
           528 => x"70",
           529 => x"ff",
           530 => x"80",
           531 => x"33",
           532 => x"d4",
           533 => x"08",
           534 => x"80",
           535 => x"81",
           536 => x"88",
           537 => x"39",
           538 => x"c8",
           539 => x"55",
           540 => x"2e",
           541 => x"84",
           542 => x"fa",
           543 => x"0b",
           544 => x"32",
           545 => x"ff",
           546 => x"92",
           547 => x"53",
           548 => x"38",
           549 => x"88",
           550 => x"55",
           551 => x"74",
           552 => x"72",
           553 => x"e3",
           554 => x"33",
           555 => x"ff",
           556 => x"73",
           557 => x"fa",
           558 => x"70",
           559 => x"56",
           560 => x"73",
           561 => x"2e",
           562 => x"88",
           563 => x"56",
           564 => x"75",
           565 => x"8c",
           566 => x"e4",
           567 => x"76",
           568 => x"54",
           569 => x"08",
           570 => x"8c",
           571 => x"3d",
           572 => x"ff",
           573 => x"55",
           574 => x"72",
           575 => x"38",
           576 => x"80",
           577 => x"33",
           578 => x"38",
           579 => x"81",
           580 => x"06",
           581 => x"3d",
           582 => x"72",
           583 => x"05",
           584 => x"b8",
           585 => x"51",
           586 => x"b8",
           587 => x"80",
           588 => x"70",
           589 => x"08",
           590 => x"53",
           591 => x"84",
           592 => x"74",
           593 => x"ff",
           594 => x"77",
           595 => x"05",
           596 => x"12",
           597 => x"51",
           598 => x"70",
           599 => x"85",
           600 => x"79",
           601 => x"80",
           602 => x"38",
           603 => x"81",
           604 => x"55",
           605 => x"73",
           606 => x"04",
           607 => x"38",
           608 => x"ff",
           609 => x"ff",
           610 => x"ff",
           611 => x"73",
           612 => x"c7",
           613 => x"53",
           614 => x"70",
           615 => x"84",
           616 => x"04",
           617 => x"54",
           618 => x"51",
           619 => x"70",
           620 => x"85",
           621 => x"78",
           622 => x"80",
           623 => x"53",
           624 => x"ff",
           625 => x"b8",
           626 => x"3d",
           627 => x"72",
           628 => x"70",
           629 => x"71",
           630 => x"14",
           631 => x"13",
           632 => x"84",
           633 => x"72",
           634 => x"ff",
           635 => x"15",
           636 => x"de",
           637 => x"0c",
           638 => x"e4",
           639 => x"0d",
           640 => x"c1",
           641 => x"e4",
           642 => x"d9",
           643 => x"b8",
           644 => x"b8",
           645 => x"74",
           646 => x"51",
           647 => x"54",
           648 => x"0d",
           649 => x"71",
           650 => x"9f",
           651 => x"51",
           652 => x"52",
           653 => x"38",
           654 => x"70",
           655 => x"04",
           656 => x"55",
           657 => x"38",
           658 => x"ff",
           659 => x"b8",
           660 => x"3d",
           661 => x"76",
           662 => x"f5",
           663 => x"12",
           664 => x"51",
           665 => x"08",
           666 => x"80",
           667 => x"80",
           668 => x"a0",
           669 => x"54",
           670 => x"38",
           671 => x"10",
           672 => x"9f",
           673 => x"75",
           674 => x"52",
           675 => x"73",
           676 => x"e4",
           677 => x"0d",
           678 => x"30",
           679 => x"2b",
           680 => x"83",
           681 => x"25",
           682 => x"2a",
           683 => x"80",
           684 => x"71",
           685 => x"8c",
           686 => x"82",
           687 => x"2a",
           688 => x"82",
           689 => x"b8",
           690 => x"54",
           691 => x"56",
           692 => x"52",
           693 => x"75",
           694 => x"81",
           695 => x"29",
           696 => x"53",
           697 => x"78",
           698 => x"2e",
           699 => x"84",
           700 => x"73",
           701 => x"bd",
           702 => x"52",
           703 => x"38",
           704 => x"81",
           705 => x"76",
           706 => x"56",
           707 => x"74",
           708 => x"78",
           709 => x"81",
           710 => x"ff",
           711 => x"55",
           712 => x"e4",
           713 => x"0d",
           714 => x"9f",
           715 => x"32",
           716 => x"72",
           717 => x"56",
           718 => x"75",
           719 => x"88",
           720 => x"7d",
           721 => x"08",
           722 => x"2e",
           723 => x"70",
           724 => x"a0",
           725 => x"f5",
           726 => x"d0",
           727 => x"80",
           728 => x"74",
           729 => x"27",
           730 => x"06",
           731 => x"06",
           732 => x"f9",
           733 => x"89",
           734 => x"27",
           735 => x"81",
           736 => x"56",
           737 => x"78",
           738 => x"75",
           739 => x"e4",
           740 => x"16",
           741 => x"59",
           742 => x"ff",
           743 => x"33",
           744 => x"38",
           745 => x"38",
           746 => x"d0",
           747 => x"73",
           748 => x"e4",
           749 => x"81",
           750 => x"55",
           751 => x"84",
           752 => x"f7",
           753 => x"70",
           754 => x"56",
           755 => x"8f",
           756 => x"33",
           757 => x"73",
           758 => x"2e",
           759 => x"56",
           760 => x"58",
           761 => x"38",
           762 => x"14",
           763 => x"14",
           764 => x"73",
           765 => x"ff",
           766 => x"89",
           767 => x"77",
           768 => x"0c",
           769 => x"26",
           770 => x"38",
           771 => x"56",
           772 => x"0d",
           773 => x"70",
           774 => x"09",
           775 => x"70",
           776 => x"80",
           777 => x"80",
           778 => x"74",
           779 => x"56",
           780 => x"38",
           781 => x"0d",
           782 => x"0c",
           783 => x"ca",
           784 => x"8b",
           785 => x"84",
           786 => x"b8",
           787 => x"52",
           788 => x"10",
           789 => x"04",
           790 => x"83",
           791 => x"ef",
           792 => x"ce",
           793 => x"0d",
           794 => x"3f",
           795 => x"51",
           796 => x"83",
           797 => x"3d",
           798 => x"fc",
           799 => x"a4",
           800 => x"04",
           801 => x"83",
           802 => x"ee",
           803 => x"cf",
           804 => x"0d",
           805 => x"3f",
           806 => x"51",
           807 => x"83",
           808 => x"3d",
           809 => x"a4",
           810 => x"e8",
           811 => x"04",
           812 => x"83",
           813 => x"ee",
           814 => x"d1",
           815 => x"0d",
           816 => x"3f",
           817 => x"51",
           818 => x"ec",
           819 => x"e3",
           820 => x"30",
           821 => x"57",
           822 => x"83",
           823 => x"81",
           824 => x"80",
           825 => x"3d",
           826 => x"84",
           827 => x"08",
           828 => x"82",
           829 => x"07",
           830 => x"72",
           831 => x"2e",
           832 => x"55",
           833 => x"74",
           834 => x"8e",
           835 => x"d1",
           836 => x"51",
           837 => x"0c",
           838 => x"08",
           839 => x"e4",
           840 => x"84",
           841 => x"9d",
           842 => x"84",
           843 => x"55",
           844 => x"19",
           845 => x"e8",
           846 => x"b8",
           847 => x"3f",
           848 => x"e4",
           849 => x"de",
           850 => x"0d",
           851 => x"58",
           852 => x"7a",
           853 => x"08",
           854 => x"76",
           855 => x"e4",
           856 => x"84",
           857 => x"84",
           858 => x"78",
           859 => x"e4",
           860 => x"0d",
           861 => x"cf",
           862 => x"5f",
           863 => x"2e",
           864 => x"ec",
           865 => x"51",
           866 => x"27",
           867 => x"38",
           868 => x"18",
           869 => x"72",
           870 => x"d1",
           871 => x"53",
           872 => x"74",
           873 => x"dd",
           874 => x"80",
           875 => x"53",
           876 => x"81",
           877 => x"38",
           878 => x"ff",
           879 => x"38",
           880 => x"84",
           881 => x"df",
           882 => x"c2",
           883 => x"3f",
           884 => x"51",
           885 => x"98",
           886 => x"a0",
           887 => x"82",
           888 => x"26",
           889 => x"e4",
           890 => x"88",
           891 => x"d4",
           892 => x"87",
           893 => x"fe",
           894 => x"91",
           895 => x"53",
           896 => x"79",
           897 => x"72",
           898 => x"83",
           899 => x"14",
           900 => x"51",
           901 => x"38",
           902 => x"db",
           903 => x"08",
           904 => x"73",
           905 => x"53",
           906 => x"52",
           907 => x"84",
           908 => x"a0",
           909 => x"dd",
           910 => x"08",
           911 => x"16",
           912 => x"3f",
           913 => x"53",
           914 => x"38",
           915 => x"81",
           916 => x"db",
           917 => x"b8",
           918 => x"70",
           919 => x"70",
           920 => x"06",
           921 => x"72",
           922 => x"9a",
           923 => x"2b",
           924 => x"30",
           925 => x"07",
           926 => x"59",
           927 => x"a9",
           928 => x"b8",
           929 => x"3d",
           930 => x"aa",
           931 => x"83",
           932 => x"51",
           933 => x"81",
           934 => x"72",
           935 => x"71",
           936 => x"81",
           937 => x"72",
           938 => x"71",
           939 => x"81",
           940 => x"72",
           941 => x"71",
           942 => x"81",
           943 => x"88",
           944 => x"a9",
           945 => x"51",
           946 => x"9c",
           947 => x"a9",
           948 => x"51",
           949 => x"9b",
           950 => x"72",
           951 => x"2e",
           952 => x"c3",
           953 => x"3f",
           954 => x"2a",
           955 => x"2e",
           956 => x"9b",
           957 => x"b3",
           958 => x"86",
           959 => x"80",
           960 => x"81",
           961 => x"51",
           962 => x"3f",
           963 => x"52",
           964 => x"bd",
           965 => x"d3",
           966 => x"9a",
           967 => x"06",
           968 => x"38",
           969 => x"3f",
           970 => x"80",
           971 => x"70",
           972 => x"fd",
           973 => x"9a",
           974 => x"ab",
           975 => x"82",
           976 => x"80",
           977 => x"ca",
           978 => x"61",
           979 => x"60",
           980 => x"e4",
           981 => x"59",
           982 => x"d4",
           983 => x"43",
           984 => x"7e",
           985 => x"51",
           986 => x"d8",
           987 => x"79",
           988 => x"2e",
           989 => x"5e",
           990 => x"70",
           991 => x"38",
           992 => x"81",
           993 => x"5d",
           994 => x"5c",
           995 => x"29",
           996 => x"5b",
           997 => x"84",
           998 => x"08",
           999 => x"e4",
          1000 => x"7d",
          1001 => x"70",
          1002 => x"27",
          1003 => x"80",
          1004 => x"7e",
          1005 => x"08",
          1006 => x"8d",
          1007 => x"b8",
          1008 => x"3f",
          1009 => x"5c",
          1010 => x"84",
          1011 => x"84",
          1012 => x"38",
          1013 => x"82",
          1014 => x"8c",
          1015 => x"38",
          1016 => x"52",
          1017 => x"a0",
          1018 => x"67",
          1019 => x"90",
          1020 => x"3f",
          1021 => x"08",
          1022 => x"25",
          1023 => x"83",
          1024 => x"06",
          1025 => x"1b",
          1026 => x"ff",
          1027 => x"32",
          1028 => x"ff",
          1029 => x"94",
          1030 => x"d1",
          1031 => x"52",
          1032 => x"83",
          1033 => x"5b",
          1034 => x"83",
          1035 => x"82",
          1036 => x"80",
          1037 => x"ed",
          1038 => x"f8",
          1039 => x"84",
          1040 => x"84",
          1041 => x"0b",
          1042 => x"ff",
          1043 => x"81",
          1044 => x"cf",
          1045 => x"0b",
          1046 => x"d4",
          1047 => x"a7",
          1048 => x"fc",
          1049 => x"0c",
          1050 => x"26",
          1051 => x"be",
          1052 => x"53",
          1053 => x"fb",
          1054 => x"90",
          1055 => x"e4",
          1056 => x"ae",
          1057 => x"41",
          1058 => x"de",
          1059 => x"3f",
          1060 => x"7b",
          1061 => x"83",
          1062 => x"3f",
          1063 => x"fa",
          1064 => x"39",
          1065 => x"fa",
          1066 => x"e8",
          1067 => x"3f",
          1068 => x"51",
          1069 => x"d0",
          1070 => x"ff",
          1071 => x"b8",
          1072 => x"68",
          1073 => x"3f",
          1074 => x"08",
          1075 => x"e4",
          1076 => x"e1",
          1077 => x"84",
          1078 => x"cf",
          1079 => x"f9",
          1080 => x"51",
          1081 => x"b8",
          1082 => x"05",
          1083 => x"08",
          1084 => x"fe",
          1085 => x"e9",
          1086 => x"d0",
          1087 => x"52",
          1088 => x"84",
          1089 => x"7e",
          1090 => x"33",
          1091 => x"78",
          1092 => x"05",
          1093 => x"fe",
          1094 => x"e8",
          1095 => x"2e",
          1096 => x"11",
          1097 => x"3f",
          1098 => x"64",
          1099 => x"d6",
          1100 => x"c4",
          1101 => x"cf",
          1102 => x"78",
          1103 => x"26",
          1104 => x"46",
          1105 => x"11",
          1106 => x"3f",
          1107 => x"a0",
          1108 => x"ff",
          1109 => x"b8",
          1110 => x"b8",
          1111 => x"05",
          1112 => x"08",
          1113 => x"e0",
          1114 => x"59",
          1115 => x"70",
          1116 => x"7d",
          1117 => x"78",
          1118 => x"51",
          1119 => x"81",
          1120 => x"b8",
          1121 => x"05",
          1122 => x"08",
          1123 => x"fe",
          1124 => x"e8",
          1125 => x"2e",
          1126 => x"11",
          1127 => x"3f",
          1128 => x"f8",
          1129 => x"3f",
          1130 => x"38",
          1131 => x"33",
          1132 => x"39",
          1133 => x"80",
          1134 => x"e4",
          1135 => x"3d",
          1136 => x"51",
          1137 => x"b1",
          1138 => x"d7",
          1139 => x"c4",
          1140 => x"cc",
          1141 => x"78",
          1142 => x"26",
          1143 => x"d1",
          1144 => x"33",
          1145 => x"3d",
          1146 => x"51",
          1147 => x"80",
          1148 => x"80",
          1149 => x"05",
          1150 => x"ff",
          1151 => x"b8",
          1152 => x"39",
          1153 => x"80",
          1154 => x"e4",
          1155 => x"3d",
          1156 => x"51",
          1157 => x"80",
          1158 => x"f8",
          1159 => x"c7",
          1160 => x"84",
          1161 => x"51",
          1162 => x"78",
          1163 => x"79",
          1164 => x"26",
          1165 => x"f4",
          1166 => x"51",
          1167 => x"b9",
          1168 => x"d8",
          1169 => x"52",
          1170 => x"e4",
          1171 => x"b8",
          1172 => x"98",
          1173 => x"ff",
          1174 => x"b8",
          1175 => x"33",
          1176 => x"83",
          1177 => x"fc",
          1178 => x"af",
          1179 => x"83",
          1180 => x"83",
          1181 => x"b8",
          1182 => x"05",
          1183 => x"08",
          1184 => x"5c",
          1185 => x"7a",
          1186 => x"9f",
          1187 => x"80",
          1188 => x"38",
          1189 => x"c4",
          1190 => x"66",
          1191 => x"d7",
          1192 => x"39",
          1193 => x"05",
          1194 => x"ff",
          1195 => x"b8",
          1196 => x"64",
          1197 => x"45",
          1198 => x"80",
          1199 => x"e4",
          1200 => x"5e",
          1201 => x"82",
          1202 => x"fe",
          1203 => x"e1",
          1204 => x"2e",
          1205 => x"ce",
          1206 => x"23",
          1207 => x"53",
          1208 => x"84",
          1209 => x"f0",
          1210 => x"ff",
          1211 => x"b8",
          1212 => x"68",
          1213 => x"34",
          1214 => x"b8",
          1215 => x"05",
          1216 => x"08",
          1217 => x"71",
          1218 => x"59",
          1219 => x"81",
          1220 => x"d5",
          1221 => x"52",
          1222 => x"39",
          1223 => x"f3",
          1224 => x"ac",
          1225 => x"f0",
          1226 => x"ab",
          1227 => x"b8",
          1228 => x"22",
          1229 => x"45",
          1230 => x"5c",
          1231 => x"f1",
          1232 => x"f1",
          1233 => x"38",
          1234 => x"39",
          1235 => x"64",
          1236 => x"51",
          1237 => x"39",
          1238 => x"2e",
          1239 => x"fc",
          1240 => x"ac",
          1241 => x"33",
          1242 => x"f1",
          1243 => x"f1",
          1244 => x"38",
          1245 => x"39",
          1246 => x"2e",
          1247 => x"fb",
          1248 => x"7c",
          1249 => x"08",
          1250 => x"33",
          1251 => x"f1",
          1252 => x"f1",
          1253 => x"9c",
          1254 => x"47",
          1255 => x"0b",
          1256 => x"8c",
          1257 => x"52",
          1258 => x"e4",
          1259 => x"87",
          1260 => x"3f",
          1261 => x"0c",
          1262 => x"57",
          1263 => x"a6",
          1264 => x"77",
          1265 => x"75",
          1266 => x"e4",
          1267 => x"0b",
          1268 => x"83",
          1269 => x"bc",
          1270 => x"02",
          1271 => x"84",
          1272 => x"13",
          1273 => x"0c",
          1274 => x"95",
          1275 => x"3f",
          1276 => x"51",
          1277 => x"22",
          1278 => x"ac",
          1279 => x"33",
          1280 => x"3f",
          1281 => x"04",
          1282 => x"56",
          1283 => x"81",
          1284 => x"06",
          1285 => x"06",
          1286 => x"81",
          1287 => x"2e",
          1288 => x"73",
          1289 => x"72",
          1290 => x"33",
          1291 => x"70",
          1292 => x"80",
          1293 => x"38",
          1294 => x"81",
          1295 => x"09",
          1296 => x"a2",
          1297 => x"07",
          1298 => x"38",
          1299 => x"71",
          1300 => x"e4",
          1301 => x"2e",
          1302 => x"38",
          1303 => x"81",
          1304 => x"2e",
          1305 => x"15",
          1306 => x"2e",
          1307 => x"39",
          1308 => x"8b",
          1309 => x"86",
          1310 => x"52",
          1311 => x"e4",
          1312 => x"b8",
          1313 => x"3d",
          1314 => x"52",
          1315 => x"98",
          1316 => x"82",
          1317 => x"84",
          1318 => x"26",
          1319 => x"84",
          1320 => x"86",
          1321 => x"26",
          1322 => x"86",
          1323 => x"38",
          1324 => x"87",
          1325 => x"87",
          1326 => x"c0",
          1327 => x"c0",
          1328 => x"c0",
          1329 => x"c0",
          1330 => x"c0",
          1331 => x"c0",
          1332 => x"a4",
          1333 => x"80",
          1334 => x"52",
          1335 => x"0d",
          1336 => x"c0",
          1337 => x"c0",
          1338 => x"87",
          1339 => x"1c",
          1340 => x"79",
          1341 => x"08",
          1342 => x"98",
          1343 => x"87",
          1344 => x"1c",
          1345 => x"7b",
          1346 => x"08",
          1347 => x"0c",
          1348 => x"83",
          1349 => x"57",
          1350 => x"55",
          1351 => x"53",
          1352 => x"d8",
          1353 => x"3d",
          1354 => x"05",
          1355 => x"72",
          1356 => x"e4",
          1357 => x"52",
          1358 => x"38",
          1359 => x"b8",
          1360 => x"51",
          1361 => x"08",
          1362 => x"71",
          1363 => x"72",
          1364 => x"e4",
          1365 => x"52",
          1366 => x"fd",
          1367 => x"88",
          1368 => x"3f",
          1369 => x"98",
          1370 => x"38",
          1371 => x"83",
          1372 => x"e4",
          1373 => x"0d",
          1374 => x"33",
          1375 => x"70",
          1376 => x"94",
          1377 => x"06",
          1378 => x"38",
          1379 => x"51",
          1380 => x"06",
          1381 => x"93",
          1382 => x"73",
          1383 => x"80",
          1384 => x"c0",
          1385 => x"84",
          1386 => x"71",
          1387 => x"70",
          1388 => x"53",
          1389 => x"2a",
          1390 => x"38",
          1391 => x"2a",
          1392 => x"cf",
          1393 => x"8f",
          1394 => x"51",
          1395 => x"83",
          1396 => x"55",
          1397 => x"70",
          1398 => x"83",
          1399 => x"54",
          1400 => x"38",
          1401 => x"2a",
          1402 => x"80",
          1403 => x"81",
          1404 => x"81",
          1405 => x"8a",
          1406 => x"71",
          1407 => x"87",
          1408 => x"86",
          1409 => x"72",
          1410 => x"73",
          1411 => x"0c",
          1412 => x"70",
          1413 => x"72",
          1414 => x"2e",
          1415 => x"52",
          1416 => x"c0",
          1417 => x"81",
          1418 => x"d7",
          1419 => x"80",
          1420 => x"52",
          1421 => x"c0",
          1422 => x"87",
          1423 => x"0c",
          1424 => x"a8",
          1425 => x"f1",
          1426 => x"83",
          1427 => x"08",
          1428 => x"ac",
          1429 => x"9e",
          1430 => x"c0",
          1431 => x"87",
          1432 => x"0c",
          1433 => x"c8",
          1434 => x"f1",
          1435 => x"83",
          1436 => x"08",
          1437 => x"c0",
          1438 => x"87",
          1439 => x"0c",
          1440 => x"e0",
          1441 => x"80",
          1442 => x"84",
          1443 => x"82",
          1444 => x"80",
          1445 => x"88",
          1446 => x"80",
          1447 => x"f1",
          1448 => x"90",
          1449 => x"52",
          1450 => x"52",
          1451 => x"87",
          1452 => x"80",
          1453 => x"83",
          1454 => x"34",
          1455 => x"70",
          1456 => x"70",
          1457 => x"83",
          1458 => x"9e",
          1459 => x"51",
          1460 => x"81",
          1461 => x"0b",
          1462 => x"80",
          1463 => x"2e",
          1464 => x"eb",
          1465 => x"08",
          1466 => x"52",
          1467 => x"71",
          1468 => x"c0",
          1469 => x"06",
          1470 => x"38",
          1471 => x"80",
          1472 => x"80",
          1473 => x"80",
          1474 => x"f1",
          1475 => x"90",
          1476 => x"52",
          1477 => x"71",
          1478 => x"90",
          1479 => x"53",
          1480 => x"0b",
          1481 => x"80",
          1482 => x"83",
          1483 => x"34",
          1484 => x"06",
          1485 => x"f1",
          1486 => x"90",
          1487 => x"70",
          1488 => x"83",
          1489 => x"08",
          1490 => x"34",
          1491 => x"82",
          1492 => x"51",
          1493 => x"33",
          1494 => x"b4",
          1495 => x"33",
          1496 => x"eb",
          1497 => x"f1",
          1498 => x"83",
          1499 => x"38",
          1500 => x"d6",
          1501 => x"84",
          1502 => x"73",
          1503 => x"55",
          1504 => x"33",
          1505 => x"e7",
          1506 => x"f1",
          1507 => x"83",
          1508 => x"38",
          1509 => x"ec",
          1510 => x"3f",
          1511 => x"d8",
          1512 => x"cc",
          1513 => x"b5",
          1514 => x"83",
          1515 => x"83",
          1516 => x"f1",
          1517 => x"ff",
          1518 => x"56",
          1519 => x"a6",
          1520 => x"c0",
          1521 => x"b8",
          1522 => x"ff",
          1523 => x"55",
          1524 => x"33",
          1525 => x"af",
          1526 => x"e0",
          1527 => x"51",
          1528 => x"bd",
          1529 => x"54",
          1530 => x"ac",
          1531 => x"c2",
          1532 => x"f1",
          1533 => x"75",
          1534 => x"08",
          1535 => x"54",
          1536 => x"da",
          1537 => x"f1",
          1538 => x"94",
          1539 => x"51",
          1540 => x"c0",
          1541 => x"83",
          1542 => x"83",
          1543 => x"51",
          1544 => x"08",
          1545 => x"b9",
          1546 => x"3f",
          1547 => x"d8",
          1548 => x"d8",
          1549 => x"51",
          1550 => x"bd",
          1551 => x"54",
          1552 => x"80",
          1553 => x"eb",
          1554 => x"38",
          1555 => x"ff",
          1556 => x"54",
          1557 => x"ec",
          1558 => x"bc",
          1559 => x"80",
          1560 => x"db",
          1561 => x"f1",
          1562 => x"c7",
          1563 => x"ff",
          1564 => x"54",
          1565 => x"39",
          1566 => x"c0",
          1567 => x"e5",
          1568 => x"38",
          1569 => x"83",
          1570 => x"83",
          1571 => x"fb",
          1572 => x"33",
          1573 => x"d9",
          1574 => x"80",
          1575 => x"f1",
          1576 => x"54",
          1577 => x"b9",
          1578 => x"80",
          1579 => x"f1",
          1580 => x"54",
          1581 => x"99",
          1582 => x"80",
          1583 => x"f1",
          1584 => x"54",
          1585 => x"f9",
          1586 => x"80",
          1587 => x"f1",
          1588 => x"54",
          1589 => x"d9",
          1590 => x"80",
          1591 => x"f1",
          1592 => x"54",
          1593 => x"b9",
          1594 => x"80",
          1595 => x"dd",
          1596 => x"d8",
          1597 => x"f1",
          1598 => x"cd",
          1599 => x"8e",
          1600 => x"38",
          1601 => x"52",
          1602 => x"ff",
          1603 => x"83",
          1604 => x"83",
          1605 => x"ff",
          1606 => x"83",
          1607 => x"83",
          1608 => x"ff",
          1609 => x"83",
          1610 => x"83",
          1611 => x"04",
          1612 => x"04",
          1613 => x"84",
          1614 => x"08",
          1615 => x"57",
          1616 => x"51",
          1617 => x"08",
          1618 => x"0b",
          1619 => x"f8",
          1620 => x"84",
          1621 => x"76",
          1622 => x"08",
          1623 => x"b8",
          1624 => x"e4",
          1625 => x"80",
          1626 => x"72",
          1627 => x"76",
          1628 => x"83",
          1629 => x"51",
          1630 => x"08",
          1631 => x"77",
          1632 => x"04",
          1633 => x"3f",
          1634 => x"38",
          1635 => x"79",
          1636 => x"56",
          1637 => x"52",
          1638 => x"3f",
          1639 => x"3d",
          1640 => x"08",
          1641 => x"33",
          1642 => x"81",
          1643 => x"56",
          1644 => x"05",
          1645 => x"3f",
          1646 => x"73",
          1647 => x"e4",
          1648 => x"73",
          1649 => x"2e",
          1650 => x"06",
          1651 => x"80",
          1652 => x"3d",
          1653 => x"ff",
          1654 => x"c7",
          1655 => x"2e",
          1656 => x"76",
          1657 => x"08",
          1658 => x"c9",
          1659 => x"57",
          1660 => x"ff",
          1661 => x"76",
          1662 => x"70",
          1663 => x"2e",
          1664 => x"75",
          1665 => x"59",
          1666 => x"e4",
          1667 => x"56",
          1668 => x"08",
          1669 => x"53",
          1670 => x"fd",
          1671 => x"ba",
          1672 => x"84",
          1673 => x"b8",
          1674 => x"e4",
          1675 => x"80",
          1676 => x"16",
          1677 => x"99",
          1678 => x"ff",
          1679 => x"0c",
          1680 => x"b5",
          1681 => x"08",
          1682 => x"34",
          1683 => x"08",
          1684 => x"f2",
          1685 => x"82",
          1686 => x"38",
          1687 => x"90",
          1688 => x"38",
          1689 => x"51",
          1690 => x"98",
          1691 => x"ff",
          1692 => x"84",
          1693 => x"98",
          1694 => x"2b",
          1695 => x"70",
          1696 => x"08",
          1697 => x"46",
          1698 => x"74",
          1699 => x"27",
          1700 => x"29",
          1701 => x"57",
          1702 => x"75",
          1703 => x"80",
          1704 => x"57",
          1705 => x"ec",
          1706 => x"78",
          1707 => x"2e",
          1708 => x"81",
          1709 => x"81",
          1710 => x"84",
          1711 => x"97",
          1712 => x"2b",
          1713 => x"5f",
          1714 => x"2e",
          1715 => x"34",
          1716 => x"ba",
          1717 => x"80",
          1718 => x"ff",
          1719 => x"80",
          1720 => x"2b",
          1721 => x"16",
          1722 => x"38",
          1723 => x"33",
          1724 => x"38",
          1725 => x"f2",
          1726 => x"ab",
          1727 => x"b2",
          1728 => x"76",
          1729 => x"9c",
          1730 => x"62",
          1731 => x"74",
          1732 => x"76",
          1733 => x"7f",
          1734 => x"80",
          1735 => x"84",
          1736 => x"fd",
          1737 => x"88",
          1738 => x"a8",
          1739 => x"a8",
          1740 => x"33",
          1741 => x"33",
          1742 => x"d6",
          1743 => x"15",
          1744 => x"16",
          1745 => x"3f",
          1746 => x"da",
          1747 => x"05",
          1748 => x"38",
          1749 => x"34",
          1750 => x"33",
          1751 => x"84",
          1752 => x"b5",
          1753 => x"a0",
          1754 => x"c8",
          1755 => x"3f",
          1756 => x"7a",
          1757 => x"06",
          1758 => x"a6",
          1759 => x"fb",
          1760 => x"c8",
          1761 => x"10",
          1762 => x"08",
          1763 => x"08",
          1764 => x"75",
          1765 => x"e4",
          1766 => x"e4",
          1767 => x"75",
          1768 => x"84",
          1769 => x"56",
          1770 => x"84",
          1771 => x"b4",
          1772 => x"a0",
          1773 => x"c8",
          1774 => x"3f",
          1775 => x"74",
          1776 => x"06",
          1777 => x"70",
          1778 => x"5b",
          1779 => x"38",
          1780 => x"57",
          1781 => x"70",
          1782 => x"84",
          1783 => x"84",
          1784 => x"78",
          1785 => x"08",
          1786 => x"a8",
          1787 => x"ff",
          1788 => x"70",
          1789 => x"5a",
          1790 => x"38",
          1791 => x"84",
          1792 => x"2e",
          1793 => x"84",
          1794 => x"98",
          1795 => x"5a",
          1796 => x"d4",
          1797 => x"bf",
          1798 => x"2b",
          1799 => x"5a",
          1800 => x"86",
          1801 => x"51",
          1802 => x"0a",
          1803 => x"2c",
          1804 => x"74",
          1805 => x"c8",
          1806 => x"3f",
          1807 => x"0a",
          1808 => x"33",
          1809 => x"b9",
          1810 => x"81",
          1811 => x"08",
          1812 => x"3f",
          1813 => x"0a",
          1814 => x"33",
          1815 => x"e6",
          1816 => x"78",
          1817 => x"33",
          1818 => x"80",
          1819 => x"98",
          1820 => x"55",
          1821 => x"b6",
          1822 => x"80",
          1823 => x"08",
          1824 => x"84",
          1825 => x"84",
          1826 => x"55",
          1827 => x"05",
          1828 => x"08",
          1829 => x"84",
          1830 => x"3f",
          1831 => x"58",
          1832 => x"33",
          1833 => x"83",
          1834 => x"f1",
          1835 => x"74",
          1836 => x"fc",
          1837 => x"70",
          1838 => x"84",
          1839 => x"d4",
          1840 => x"05",
          1841 => x"ad",
          1842 => x"80",
          1843 => x"58",
          1844 => x"0b",
          1845 => x"d0",
          1846 => x"b4",
          1847 => x"55",
          1848 => x"c8",
          1849 => x"3f",
          1850 => x"ff",
          1851 => x"52",
          1852 => x"d0",
          1853 => x"d0",
          1854 => x"74",
          1855 => x"a0",
          1856 => x"34",
          1857 => x"be",
          1858 => x"1d",
          1859 => x"80",
          1860 => x"52",
          1861 => x"d4",
          1862 => x"b7",
          1863 => x"51",
          1864 => x"33",
          1865 => x"34",
          1866 => x"38",
          1867 => x"3f",
          1868 => x"0b",
          1869 => x"e4",
          1870 => x"a8",
          1871 => x"7a",
          1872 => x"a4",
          1873 => x"a4",
          1874 => x"a8",
          1875 => x"51",
          1876 => x"33",
          1877 => x"d0",
          1878 => x"76",
          1879 => x"08",
          1880 => x"84",
          1881 => x"98",
          1882 => x"59",
          1883 => x"84",
          1884 => x"ad",
          1885 => x"81",
          1886 => x"d0",
          1887 => x"24",
          1888 => x"52",
          1889 => x"81",
          1890 => x"70",
          1891 => x"51",
          1892 => x"f3",
          1893 => x"33",
          1894 => x"76",
          1895 => x"81",
          1896 => x"70",
          1897 => x"57",
          1898 => x"7b",
          1899 => x"84",
          1900 => x"ff",
          1901 => x"29",
          1902 => x"84",
          1903 => x"76",
          1904 => x"84",
          1905 => x"58",
          1906 => x"84",
          1907 => x"ae",
          1908 => x"57",
          1909 => x"16",
          1910 => x"81",
          1911 => x"70",
          1912 => x"57",
          1913 => x"18",
          1914 => x"81",
          1915 => x"33",
          1916 => x"76",
          1917 => x"75",
          1918 => x"d0",
          1919 => x"81",
          1920 => x"81",
          1921 => x"76",
          1922 => x"70",
          1923 => x"57",
          1924 => x"84",
          1925 => x"aa",
          1926 => x"81",
          1927 => x"d0",
          1928 => x"25",
          1929 => x"52",
          1930 => x"81",
          1931 => x"70",
          1932 => x"57",
          1933 => x"f0",
          1934 => x"75",
          1935 => x"ff",
          1936 => x"84",
          1937 => x"81",
          1938 => x"7b",
          1939 => x"a4",
          1940 => x"74",
          1941 => x"c8",
          1942 => x"3f",
          1943 => x"ff",
          1944 => x"52",
          1945 => x"d0",
          1946 => x"d0",
          1947 => x"c7",
          1948 => x"84",
          1949 => x"84",
          1950 => x"83",
          1951 => x"80",
          1952 => x"7b",
          1953 => x"df",
          1954 => x"80",
          1955 => x"a4",
          1956 => x"da",
          1957 => x"2b",
          1958 => x"5d",
          1959 => x"8e",
          1960 => x"08",
          1961 => x"fc",
          1962 => x"bb",
          1963 => x"75",
          1964 => x"f2",
          1965 => x"74",
          1966 => x"81",
          1967 => x"51",
          1968 => x"f2",
          1969 => x"5f",
          1970 => x"e9",
          1971 => x"18",
          1972 => x"38",
          1973 => x"f9",
          1974 => x"a4",
          1975 => x"06",
          1976 => x"ff",
          1977 => x"a4",
          1978 => x"5d",
          1979 => x"d4",
          1980 => x"87",
          1981 => x"51",
          1982 => x"08",
          1983 => x"84",
          1984 => x"84",
          1985 => x"55",
          1986 => x"84",
          1987 => x"a4",
          1988 => x"3d",
          1989 => x"3f",
          1990 => x"34",
          1991 => x"81",
          1992 => x"aa",
          1993 => x"06",
          1994 => x"33",
          1995 => x"f1",
          1996 => x"88",
          1997 => x"c8",
          1998 => x"3f",
          1999 => x"ff",
          2000 => x"ff",
          2001 => x"76",
          2002 => x"51",
          2003 => x"08",
          2004 => x"08",
          2005 => x"52",
          2006 => x"1d",
          2007 => x"33",
          2008 => x"58",
          2009 => x"d4",
          2010 => x"97",
          2011 => x"51",
          2012 => x"08",
          2013 => x"84",
          2014 => x"84",
          2015 => x"55",
          2016 => x"3f",
          2017 => x"87",
          2018 => x"19",
          2019 => x"d1",
          2020 => x"83",
          2021 => x"f1",
          2022 => x"74",
          2023 => x"7b",
          2024 => x"83",
          2025 => x"ff",
          2026 => x"f2",
          2027 => x"b1",
          2028 => x"76",
          2029 => x"c0",
          2030 => x"51",
          2031 => x"08",
          2032 => x"84",
          2033 => x"a4",
          2034 => x"3d",
          2035 => x"b8",
          2036 => x"84",
          2037 => x"b8",
          2038 => x"f2",
          2039 => x"51",
          2040 => x"08",
          2041 => x"09",
          2042 => x"e4",
          2043 => x"b8",
          2044 => x"e4",
          2045 => x"e4",
          2046 => x"80",
          2047 => x"f2",
          2048 => x"fc",
          2049 => x"74",
          2050 => x"fc",
          2051 => x"70",
          2052 => x"84",
          2053 => x"d4",
          2054 => x"05",
          2055 => x"38",
          2056 => x"57",
          2057 => x"75",
          2058 => x"38",
          2059 => x"76",
          2060 => x"83",
          2061 => x"70",
          2062 => x"27",
          2063 => x"d4",
          2064 => x"d3",
          2065 => x"82",
          2066 => x"05",
          2067 => x"80",
          2068 => x"75",
          2069 => x"10",
          2070 => x"40",
          2071 => x"ff",
          2072 => x"fe",
          2073 => x"f1",
          2074 => x"9f",
          2075 => x"e4",
          2076 => x"05",
          2077 => x"33",
          2078 => x"38",
          2079 => x"73",
          2080 => x"82",
          2081 => x"86",
          2082 => x"56",
          2083 => x"38",
          2084 => x"f8",
          2085 => x"83",
          2086 => x"90",
          2087 => x"07",
          2088 => x"77",
          2089 => x"05",
          2090 => x"55",
          2091 => x"78",
          2092 => x"84",
          2093 => x"55",
          2094 => x"74",
          2095 => x"13",
          2096 => x"04",
          2097 => x"94",
          2098 => x"95",
          2099 => x"5b",
          2100 => x"80",
          2101 => x"ff",
          2102 => x"ff",
          2103 => x"ff",
          2104 => x"5d",
          2105 => x"26",
          2106 => x"56",
          2107 => x"06",
          2108 => x"ff",
          2109 => x"29",
          2110 => x"74",
          2111 => x"33",
          2112 => x"1b",
          2113 => x"80",
          2114 => x"53",
          2115 => x"73",
          2116 => x"90",
          2117 => x"e8",
          2118 => x"a7",
          2119 => x"70",
          2120 => x"70",
          2121 => x"70",
          2122 => x"56",
          2123 => x"38",
          2124 => x"06",
          2125 => x"79",
          2126 => x"83",
          2127 => x"95",
          2128 => x"2b",
          2129 => x"07",
          2130 => x"5b",
          2131 => x"be",
          2132 => x"94",
          2133 => x"10",
          2134 => x"29",
          2135 => x"57",
          2136 => x"80",
          2137 => x"81",
          2138 => x"81",
          2139 => x"83",
          2140 => x"05",
          2141 => x"5e",
          2142 => x"7a",
          2143 => x"53",
          2144 => x"06",
          2145 => x"06",
          2146 => x"58",
          2147 => x"26",
          2148 => x"73",
          2149 => x"79",
          2150 => x"7b",
          2151 => x"78",
          2152 => x"fb",
          2153 => x"ff",
          2154 => x"73",
          2155 => x"9c",
          2156 => x"75",
          2157 => x"76",
          2158 => x"94",
          2159 => x"ff",
          2160 => x"fa",
          2161 => x"08",
          2162 => x"81",
          2163 => x"55",
          2164 => x"ff",
          2165 => x"75",
          2166 => x"77",
          2167 => x"a0",
          2168 => x"06",
          2169 => x"d0",
          2170 => x"84",
          2171 => x"84",
          2172 => x"04",
          2173 => x"02",
          2174 => x"d7",
          2175 => x"79",
          2176 => x"33",
          2177 => x"33",
          2178 => x"80",
          2179 => x"57",
          2180 => x"ff",
          2181 => x"57",
          2182 => x"38",
          2183 => x"74",
          2184 => x"33",
          2185 => x"81",
          2186 => x"26",
          2187 => x"83",
          2188 => x"70",
          2189 => x"33",
          2190 => x"89",
          2191 => x"29",
          2192 => x"26",
          2193 => x"54",
          2194 => x"16",
          2195 => x"75",
          2196 => x"54",
          2197 => x"73",
          2198 => x"90",
          2199 => x"a0",
          2200 => x"70",
          2201 => x"9f",
          2202 => x"d6",
          2203 => x"92",
          2204 => x"77",
          2205 => x"73",
          2206 => x"81",
          2207 => x"29",
          2208 => x"a0",
          2209 => x"81",
          2210 => x"71",
          2211 => x"79",
          2212 => x"54",
          2213 => x"e0",
          2214 => x"34",
          2215 => x"70",
          2216 => x"b6",
          2217 => x"71",
          2218 => x"75",
          2219 => x"b8",
          2220 => x"83",
          2221 => x"70",
          2222 => x"33",
          2223 => x"f9",
          2224 => x"78",
          2225 => x"94",
          2226 => x"81",
          2227 => x"81",
          2228 => x"29",
          2229 => x"54",
          2230 => x"f8",
          2231 => x"76",
          2232 => x"e0",
          2233 => x"57",
          2234 => x"fe",
          2235 => x"34",
          2236 => x"ff",
          2237 => x"39",
          2238 => x"56",
          2239 => x"33",
          2240 => x"34",
          2241 => x"39",
          2242 => x"9f",
          2243 => x"9b",
          2244 => x"05",
          2245 => x"33",
          2246 => x"83",
          2247 => x"e4",
          2248 => x"83",
          2249 => x"70",
          2250 => x"2e",
          2251 => x"f8",
          2252 => x"0c",
          2253 => x"33",
          2254 => x"2c",
          2255 => x"83",
          2256 => x"94",
          2257 => x"ff",
          2258 => x"83",
          2259 => x"34",
          2260 => x"3d",
          2261 => x"73",
          2262 => x"06",
          2263 => x"95",
          2264 => x"86",
          2265 => x"72",
          2266 => x"55",
          2267 => x"70",
          2268 => x"0b",
          2269 => x"04",
          2270 => x"f8",
          2271 => x"05",
          2272 => x"38",
          2273 => x"34",
          2274 => x"8f",
          2275 => x"38",
          2276 => x"51",
          2277 => x"70",
          2278 => x"f0",
          2279 => x"52",
          2280 => x"81",
          2281 => x"f8",
          2282 => x"0c",
          2283 => x"33",
          2284 => x"83",
          2285 => x"e4",
          2286 => x"90",
          2287 => x"f8",
          2288 => x"33",
          2289 => x"83",
          2290 => x"0b",
          2291 => x"b8",
          2292 => x"f8",
          2293 => x"51",
          2294 => x"39",
          2295 => x"70",
          2296 => x"83",
          2297 => x"07",
          2298 => x"93",
          2299 => x"06",
          2300 => x"34",
          2301 => x"81",
          2302 => x"f8",
          2303 => x"90",
          2304 => x"f8",
          2305 => x"90",
          2306 => x"51",
          2307 => x"39",
          2308 => x"b0",
          2309 => x"fe",
          2310 => x"ef",
          2311 => x"f8",
          2312 => x"90",
          2313 => x"51",
          2314 => x"39",
          2315 => x"a0",
          2316 => x"fe",
          2317 => x"8f",
          2318 => x"fd",
          2319 => x"fa",
          2320 => x"90",
          2321 => x"02",
          2322 => x"c3",
          2323 => x"f8",
          2324 => x"b6",
          2325 => x"59",
          2326 => x"82",
          2327 => x"82",
          2328 => x"0b",
          2329 => x"94",
          2330 => x"83",
          2331 => x"78",
          2332 => x"80",
          2333 => x"84",
          2334 => x"94",
          2335 => x"82",
          2336 => x"84",
          2337 => x"33",
          2338 => x"54",
          2339 => x"51",
          2340 => x"da",
          2341 => x"7a",
          2342 => x"92",
          2343 => x"3d",
          2344 => x"34",
          2345 => x"0b",
          2346 => x"f8",
          2347 => x"23",
          2348 => x"e6",
          2349 => x"79",
          2350 => x"83",
          2351 => x"80",
          2352 => x"79",
          2353 => x"b8",
          2354 => x"e3",
          2355 => x"1a",
          2356 => x"33",
          2357 => x"38",
          2358 => x"3f",
          2359 => x"84",
          2360 => x"34",
          2361 => x"f8",
          2362 => x"0b",
          2363 => x"b6",
          2364 => x"34",
          2365 => x"0b",
          2366 => x"51",
          2367 => x"08",
          2368 => x"81",
          2369 => x"ff",
          2370 => x"08",
          2371 => x"19",
          2372 => x"ff",
          2373 => x"06",
          2374 => x"7a",
          2375 => x"b6",
          2376 => x"f8",
          2377 => x"a7",
          2378 => x"53",
          2379 => x"70",
          2380 => x"33",
          2381 => x"81",
          2382 => x"81",
          2383 => x"38",
          2384 => x"88",
          2385 => x"33",
          2386 => x"33",
          2387 => x"84",
          2388 => x"80",
          2389 => x"f8",
          2390 => x"71",
          2391 => x"83",
          2392 => x"33",
          2393 => x"f8",
          2394 => x"34",
          2395 => x"06",
          2396 => x"33",
          2397 => x"55",
          2398 => x"b6",
          2399 => x"06",
          2400 => x"38",
          2401 => x"ea",
          2402 => x"95",
          2403 => x"80",
          2404 => x"57",
          2405 => x"0b",
          2406 => x"04",
          2407 => x"24",
          2408 => x"81",
          2409 => x"51",
          2410 => x"95",
          2411 => x"15",
          2412 => x"74",
          2413 => x"fe",
          2414 => x"51",
          2415 => x"ff",
          2416 => x"91",
          2417 => x"3f",
          2418 => x"54",
          2419 => x"39",
          2420 => x"39",
          2421 => x"80",
          2422 => x"0d",
          2423 => x"06",
          2424 => x"70",
          2425 => x"73",
          2426 => x"95",
          2427 => x"3f",
          2428 => x"06",
          2429 => x"38",
          2430 => x"fe",
          2431 => x"34",
          2432 => x"fe",
          2433 => x"d8",
          2434 => x"02",
          2435 => x"08",
          2436 => x"38",
          2437 => x"8a",
          2438 => x"82",
          2439 => x"38",
          2440 => x"b6",
          2441 => x"f8",
          2442 => x"5e",
          2443 => x"a7",
          2444 => x"33",
          2445 => x"22",
          2446 => x"40",
          2447 => x"f8",
          2448 => x"40",
          2449 => x"a7",
          2450 => x"33",
          2451 => x"22",
          2452 => x"11",
          2453 => x"90",
          2454 => x"1d",
          2455 => x"61",
          2456 => x"33",
          2457 => x"56",
          2458 => x"84",
          2459 => x"78",
          2460 => x"25",
          2461 => x"b3",
          2462 => x"38",
          2463 => x"b6",
          2464 => x"f8",
          2465 => x"40",
          2466 => x"a7",
          2467 => x"33",
          2468 => x"22",
          2469 => x"56",
          2470 => x"f8",
          2471 => x"57",
          2472 => x"80",
          2473 => x"81",
          2474 => x"f8",
          2475 => x"42",
          2476 => x"60",
          2477 => x"58",
          2478 => x"27",
          2479 => x"34",
          2480 => x"3d",
          2481 => x"38",
          2482 => x"8d",
          2483 => x"80",
          2484 => x"84",
          2485 => x"78",
          2486 => x"56",
          2487 => x"b7",
          2488 => x"84",
          2489 => x"18",
          2490 => x"0b",
          2491 => x"84",
          2492 => x"78",
          2493 => x"84",
          2494 => x"83",
          2495 => x"72",
          2496 => x"b6",
          2497 => x"1d",
          2498 => x"95",
          2499 => x"29",
          2500 => x"f8",
          2501 => x"76",
          2502 => x"90",
          2503 => x"84",
          2504 => x"83",
          2505 => x"72",
          2506 => x"59",
          2507 => x"b6",
          2508 => x"39",
          2509 => x"80",
          2510 => x"39",
          2511 => x"33",
          2512 => x"33",
          2513 => x"80",
          2514 => x"5d",
          2515 => x"ff",
          2516 => x"59",
          2517 => x"38",
          2518 => x"57",
          2519 => x"83",
          2520 => x"0b",
          2521 => x"b7",
          2522 => x"34",
          2523 => x"0b",
          2524 => x"b8",
          2525 => x"f8",
          2526 => x"f8",
          2527 => x"f8",
          2528 => x"0b",
          2529 => x"b8",
          2530 => x"80",
          2531 => x"38",
          2532 => x"33",
          2533 => x"33",
          2534 => x"11",
          2535 => x"92",
          2536 => x"70",
          2537 => x"33",
          2538 => x"7d",
          2539 => x"ff",
          2540 => x"38",
          2541 => x"7b",
          2542 => x"78",
          2543 => x"5f",
          2544 => x"a7",
          2545 => x"33",
          2546 => x"22",
          2547 => x"40",
          2548 => x"83",
          2549 => x"05",
          2550 => x"a7",
          2551 => x"33",
          2552 => x"22",
          2553 => x"11",
          2554 => x"90",
          2555 => x"81",
          2556 => x"7c",
          2557 => x"d9",
          2558 => x"19",
          2559 => x"f8",
          2560 => x"ff",
          2561 => x"2e",
          2562 => x"d7",
          2563 => x"84",
          2564 => x"38",
          2565 => x"84",
          2566 => x"c0",
          2567 => x"83",
          2568 => x"e7",
          2569 => x"0c",
          2570 => x"33",
          2571 => x"06",
          2572 => x"06",
          2573 => x"80",
          2574 => x"72",
          2575 => x"06",
          2576 => x"5c",
          2577 => x"ef",
          2578 => x"7a",
          2579 => x"72",
          2580 => x"b7",
          2581 => x"34",
          2582 => x"33",
          2583 => x"12",
          2584 => x"f8",
          2585 => x"76",
          2586 => x"90",
          2587 => x"84",
          2588 => x"83",
          2589 => x"72",
          2590 => x"59",
          2591 => x"18",
          2592 => x"06",
          2593 => x"38",
          2594 => x"fb",
          2595 => x"95",
          2596 => x"5d",
          2597 => x"83",
          2598 => x"83",
          2599 => x"72",
          2600 => x"72",
          2601 => x"5b",
          2602 => x"a0",
          2603 => x"83",
          2604 => x"72",
          2605 => x"a0",
          2606 => x"f8",
          2607 => x"5e",
          2608 => x"80",
          2609 => x"81",
          2610 => x"f8",
          2611 => x"44",
          2612 => x"84",
          2613 => x"70",
          2614 => x"27",
          2615 => x"34",
          2616 => x"e0",
          2617 => x"9c",
          2618 => x"33",
          2619 => x"34",
          2620 => x"06",
          2621 => x"81",
          2622 => x"84",
          2623 => x"83",
          2624 => x"e0",
          2625 => x"33",
          2626 => x"33",
          2627 => x"39",
          2628 => x"11",
          2629 => x"3f",
          2630 => x"f0",
          2631 => x"57",
          2632 => x"10",
          2633 => x"05",
          2634 => x"fb",
          2635 => x"5c",
          2636 => x"83",
          2637 => x"83",
          2638 => x"e5",
          2639 => x"94",
          2640 => x"29",
          2641 => x"19",
          2642 => x"34",
          2643 => x"33",
          2644 => x"12",
          2645 => x"96",
          2646 => x"71",
          2647 => x"33",
          2648 => x"84",
          2649 => x"83",
          2650 => x"72",
          2651 => x"5a",
          2652 => x"1e",
          2653 => x"5c",
          2654 => x"84",
          2655 => x"38",
          2656 => x"34",
          2657 => x"b6",
          2658 => x"bd",
          2659 => x"f3",
          2660 => x"e4",
          2661 => x"9c",
          2662 => x"83",
          2663 => x"83",
          2664 => x"57",
          2665 => x"39",
          2666 => x"34",
          2667 => x"34",
          2668 => x"34",
          2669 => x"5b",
          2670 => x"b8",
          2671 => x"81",
          2672 => x"33",
          2673 => x"81",
          2674 => x"52",
          2675 => x"89",
          2676 => x"84",
          2677 => x"f6",
          2678 => x"a0",
          2679 => x"f6",
          2680 => x"c0",
          2681 => x"5b",
          2682 => x"7b",
          2683 => x"b8",
          2684 => x"75",
          2685 => x"10",
          2686 => x"04",
          2687 => x"2e",
          2688 => x"84",
          2689 => x"09",
          2690 => x"59",
          2691 => x"fd",
          2692 => x"75",
          2693 => x"b9",
          2694 => x"84",
          2695 => x"7b",
          2696 => x"95",
          2697 => x"f8",
          2698 => x"81",
          2699 => x"fd",
          2700 => x"f8",
          2701 => x"83",
          2702 => x"84",
          2703 => x"76",
          2704 => x"56",
          2705 => x"39",
          2706 => x"2e",
          2707 => x"84",
          2708 => x"09",
          2709 => x"59",
          2710 => x"fc",
          2711 => x"7a",
          2712 => x"b8",
          2713 => x"06",
          2714 => x"83",
          2715 => x"72",
          2716 => x"11",
          2717 => x"58",
          2718 => x"ff",
          2719 => x"fe",
          2720 => x"84",
          2721 => x"0b",
          2722 => x"84",
          2723 => x"fb",
          2724 => x"77",
          2725 => x"38",
          2726 => x"d0",
          2727 => x"80",
          2728 => x"33",
          2729 => x"84",
          2730 => x"56",
          2731 => x"76",
          2732 => x"84",
          2733 => x"8c",
          2734 => x"f8",
          2735 => x"d7",
          2736 => x"60",
          2737 => x"f8",
          2738 => x"ac",
          2739 => x"84",
          2740 => x"27",
          2741 => x"b8",
          2742 => x"8c",
          2743 => x"70",
          2744 => x"58",
          2745 => x"b7",
          2746 => x"8d",
          2747 => x"83",
          2748 => x"76",
          2749 => x"fa",
          2750 => x"81",
          2751 => x"bb",
          2752 => x"84",
          2753 => x"ff",
          2754 => x"ff",
          2755 => x"59",
          2756 => x"77",
          2757 => x"81",
          2758 => x"7f",
          2759 => x"f8",
          2760 => x"11",
          2761 => x"38",
          2762 => x"f9",
          2763 => x"7e",
          2764 => x"b9",
          2765 => x"7a",
          2766 => x"94",
          2767 => x"ff",
          2768 => x"29",
          2769 => x"f8",
          2770 => x"05",
          2771 => x"ea",
          2772 => x"60",
          2773 => x"ff",
          2774 => x"80",
          2775 => x"d7",
          2776 => x"38",
          2777 => x"23",
          2778 => x"41",
          2779 => x"84",
          2780 => x"8d",
          2781 => x"f8",
          2782 => x"f8",
          2783 => x"76",
          2784 => x"05",
          2785 => x"5c",
          2786 => x"80",
          2787 => x"ff",
          2788 => x"29",
          2789 => x"27",
          2790 => x"57",
          2791 => x"e0",
          2792 => x"34",
          2793 => x"70",
          2794 => x"b6",
          2795 => x"71",
          2796 => x"60",
          2797 => x"33",
          2798 => x"70",
          2799 => x"05",
          2800 => x"34",
          2801 => x"b6",
          2802 => x"40",
          2803 => x"38",
          2804 => x"56",
          2805 => x"52",
          2806 => x"3f",
          2807 => x"d8",
          2808 => x"5d",
          2809 => x"38",
          2810 => x"2e",
          2811 => x"f8",
          2812 => x"83",
          2813 => x"76",
          2814 => x"d7",
          2815 => x"38",
          2816 => x"26",
          2817 => x"7d",
          2818 => x"7a",
          2819 => x"05",
          2820 => x"5d",
          2821 => x"83",
          2822 => x"38",
          2823 => x"38",
          2824 => x"71",
          2825 => x"71",
          2826 => x"77",
          2827 => x"84",
          2828 => x"05",
          2829 => x"84",
          2830 => x"41",
          2831 => x"ff",
          2832 => x"29",
          2833 => x"77",
          2834 => x"70",
          2835 => x"76",
          2836 => x"e0",
          2837 => x"b6",
          2838 => x"19",
          2839 => x"34",
          2840 => x"c0",
          2841 => x"79",
          2842 => x"17",
          2843 => x"a8",
          2844 => x"5d",
          2845 => x"33",
          2846 => x"80",
          2847 => x"5d",
          2848 => x"06",
          2849 => x"90",
          2850 => x"59",
          2851 => x"17",
          2852 => x"7c",
          2853 => x"d8",
          2854 => x"d7",
          2855 => x"39",
          2856 => x"75",
          2857 => x"81",
          2858 => x"83",
          2859 => x"07",
          2860 => x"39",
          2861 => x"83",
          2862 => x"d4",
          2863 => x"06",
          2864 => x"34",
          2865 => x"9f",
          2866 => x"90",
          2867 => x"83",
          2868 => x"ff",
          2869 => x"f8",
          2870 => x"83",
          2871 => x"f8",
          2872 => x"56",
          2873 => x"39",
          2874 => x"80",
          2875 => x"34",
          2876 => x"81",
          2877 => x"83",
          2878 => x"f8",
          2879 => x"56",
          2880 => x"39",
          2881 => x"86",
          2882 => x"fe",
          2883 => x"fc",
          2884 => x"90",
          2885 => x"33",
          2886 => x"83",
          2887 => x"f8",
          2888 => x"83",
          2889 => x"f8",
          2890 => x"83",
          2891 => x"f8",
          2892 => x"83",
          2893 => x"f8",
          2894 => x"07",
          2895 => x"cc",
          2896 => x"06",
          2897 => x"34",
          2898 => x"95",
          2899 => x"3f",
          2900 => x"83",
          2901 => x"83",
          2902 => x"59",
          2903 => x"84",
          2904 => x"0b",
          2905 => x"b8",
          2906 => x"83",
          2907 => x"70",
          2908 => x"e7",
          2909 => x"3d",
          2910 => x"f9",
          2911 => x"38",
          2912 => x"0c",
          2913 => x"0b",
          2914 => x"04",
          2915 => x"39",
          2916 => x"5c",
          2917 => x"83",
          2918 => x"22",
          2919 => x"84",
          2920 => x"83",
          2921 => x"d1",
          2922 => x"81",
          2923 => x"d8",
          2924 => x"80",
          2925 => x"98",
          2926 => x"ef",
          2927 => x"05",
          2928 => x"58",
          2929 => x"81",
          2930 => x"40",
          2931 => x"83",
          2932 => x"f8",
          2933 => x"9f",
          2934 => x"e2",
          2935 => x"84",
          2936 => x"56",
          2937 => x"57",
          2938 => x"70",
          2939 => x"26",
          2940 => x"84",
          2941 => x"83",
          2942 => x"86",
          2943 => x"22",
          2944 => x"83",
          2945 => x"5d",
          2946 => x"2e",
          2947 => x"06",
          2948 => x"84",
          2949 => x"76",
          2950 => x"56",
          2951 => x"ff",
          2952 => x"24",
          2953 => x"56",
          2954 => x"16",
          2955 => x"81",
          2956 => x"57",
          2957 => x"75",
          2958 => x"06",
          2959 => x"58",
          2960 => x"b0",
          2961 => x"ff",
          2962 => x"42",
          2963 => x"84",
          2964 => x"33",
          2965 => x"70",
          2966 => x"05",
          2967 => x"34",
          2968 => x"b6",
          2969 => x"41",
          2970 => x"38",
          2971 => x"e0",
          2972 => x"34",
          2973 => x"70",
          2974 => x"b6",
          2975 => x"71",
          2976 => x"78",
          2977 => x"83",
          2978 => x"e0",
          2979 => x"33",
          2980 => x"22",
          2981 => x"5d",
          2982 => x"84",
          2983 => x"ff",
          2984 => x"83",
          2985 => x"23",
          2986 => x"5a",
          2987 => x"76",
          2988 => x"33",
          2989 => x"59",
          2990 => x"80",
          2991 => x"88",
          2992 => x"84",
          2993 => x"56",
          2994 => x"57",
          2995 => x"81",
          2996 => x"33",
          2997 => x"33",
          2998 => x"2e",
          2999 => x"a1",
          3000 => x"94",
          3001 => x"75",
          3002 => x"7c",
          3003 => x"34",
          3004 => x"77",
          3005 => x"70",
          3006 => x"33",
          3007 => x"7a",
          3008 => x"81",
          3009 => x"77",
          3010 => x"27",
          3011 => x"31",
          3012 => x"a8",
          3013 => x"fc",
          3014 => x"fc",
          3015 => x"23",
          3016 => x"94",
          3017 => x"18",
          3018 => x"77",
          3019 => x"e9",
          3020 => x"05",
          3021 => x"72",
          3022 => x"9c",
          3023 => x"85",
          3024 => x"d7",
          3025 => x"0c",
          3026 => x"02",
          3027 => x"f6",
          3028 => x"f6",
          3029 => x"74",
          3030 => x"56",
          3031 => x"78",
          3032 => x"04",
          3033 => x"73",
          3034 => x"70",
          3035 => x"2a",
          3036 => x"c4",
          3037 => x"2e",
          3038 => x"7b",
          3039 => x"76",
          3040 => x"85",
          3041 => x"f8",
          3042 => x"71",
          3043 => x"83",
          3044 => x"79",
          3045 => x"83",
          3046 => x"74",
          3047 => x"54",
          3048 => x"0b",
          3049 => x"98",
          3050 => x"38",
          3051 => x"83",
          3052 => x"81",
          3053 => x"27",
          3054 => x"14",
          3055 => x"8e",
          3056 => x"2e",
          3057 => x"86",
          3058 => x"34",
          3059 => x"ff",
          3060 => x"a2",
          3061 => x"83",
          3062 => x"81",
          3063 => x"ff",
          3064 => x"98",
          3065 => x"75",
          3066 => x"06",
          3067 => x"06",
          3068 => x"e7",
          3069 => x"73",
          3070 => x"85",
          3071 => x"34",
          3072 => x"f6",
          3073 => x"83",
          3074 => x"5d",
          3075 => x"f6",
          3076 => x"2e",
          3077 => x"54",
          3078 => x"f6",
          3079 => x"2e",
          3080 => x"54",
          3081 => x"06",
          3082 => x"83",
          3083 => x"2e",
          3084 => x"53",
          3085 => x"83",
          3086 => x"27",
          3087 => x"87",
          3088 => x"54",
          3089 => x"81",
          3090 => x"f6",
          3091 => x"ff",
          3092 => x"f6",
          3093 => x"83",
          3094 => x"72",
          3095 => x"10",
          3096 => x"04",
          3097 => x"2e",
          3098 => x"98",
          3099 => x"fc",
          3100 => x"33",
          3101 => x"74",
          3102 => x"c0",
          3103 => x"73",
          3104 => x"94",
          3105 => x"84",
          3106 => x"f0",
          3107 => x"08",
          3108 => x"72",
          3109 => x"76",
          3110 => x"80",
          3111 => x"57",
          3112 => x"79",
          3113 => x"38",
          3114 => x"81",
          3115 => x"06",
          3116 => x"54",
          3117 => x"80",
          3118 => x"ff",
          3119 => x"72",
          3120 => x"58",
          3121 => x"10",
          3122 => x"83",
          3123 => x"70",
          3124 => x"98",
          3125 => x"fd",
          3126 => x"ff",
          3127 => x"ff",
          3128 => x"78",
          3129 => x"84",
          3130 => x"2e",
          3131 => x"30",
          3132 => x"56",
          3133 => x"81",
          3134 => x"f9",
          3135 => x"10",
          3136 => x"54",
          3137 => x"13",
          3138 => x"73",
          3139 => x"53",
          3140 => x"b6",
          3141 => x"78",
          3142 => x"d4",
          3143 => x"3d",
          3144 => x"54",
          3145 => x"92",
          3146 => x"05",
          3147 => x"fa",
          3148 => x"15",
          3149 => x"34",
          3150 => x"fa",
          3151 => x"72",
          3152 => x"f6",
          3153 => x"fc",
          3154 => x"73",
          3155 => x"38",
          3156 => x"87",
          3157 => x"73",
          3158 => x"9c",
          3159 => x"ff",
          3160 => x"83",
          3161 => x"72",
          3162 => x"06",
          3163 => x"f6",
          3164 => x"33",
          3165 => x"33",
          3166 => x"bf",
          3167 => x"56",
          3168 => x"81",
          3169 => x"81",
          3170 => x"09",
          3171 => x"39",
          3172 => x"98",
          3173 => x"57",
          3174 => x"84",
          3175 => x"39",
          3176 => x"54",
          3177 => x"b6",
          3178 => x"81",
          3179 => x"f7",
          3180 => x"0c",
          3181 => x"70",
          3182 => x"54",
          3183 => x"74",
          3184 => x"06",
          3185 => x"83",
          3186 => x"34",
          3187 => x"06",
          3188 => x"83",
          3189 => x"34",
          3190 => x"83",
          3191 => x"f6",
          3192 => x"84",
          3193 => x"fe",
          3194 => x"e8",
          3195 => x"bb",
          3196 => x"ac",
          3197 => x"0d",
          3198 => x"57",
          3199 => x"83",
          3200 => x"34",
          3201 => x"56",
          3202 => x"86",
          3203 => x"9c",
          3204 => x"ce",
          3205 => x"08",
          3206 => x"70",
          3207 => x"87",
          3208 => x"73",
          3209 => x"db",
          3210 => x"ff",
          3211 => x"71",
          3212 => x"87",
          3213 => x"05",
          3214 => x"87",
          3215 => x"2e",
          3216 => x"98",
          3217 => x"87",
          3218 => x"87",
          3219 => x"26",
          3220 => x"16",
          3221 => x"80",
          3222 => x"52",
          3223 => x"8a",
          3224 => x"3d",
          3225 => x"0c",
          3226 => x"79",
          3227 => x"52",
          3228 => x"88",
          3229 => x"75",
          3230 => x"71",
          3231 => x"70",
          3232 => x"75",
          3233 => x"83",
          3234 => x"34",
          3235 => x"71",
          3236 => x"55",
          3237 => x"0b",
          3238 => x"98",
          3239 => x"80",
          3240 => x"9c",
          3241 => x"51",
          3242 => x"33",
          3243 => x"74",
          3244 => x"2e",
          3245 => x"51",
          3246 => x"38",
          3247 => x"38",
          3248 => x"90",
          3249 => x"52",
          3250 => x"72",
          3251 => x"c0",
          3252 => x"27",
          3253 => x"38",
          3254 => x"75",
          3255 => x"ff",
          3256 => x"75",
          3257 => x"ff",
          3258 => x"51",
          3259 => x"38",
          3260 => x"55",
          3261 => x"71",
          3262 => x"81",
          3263 => x"38",
          3264 => x"0d",
          3265 => x"88",
          3266 => x"fa",
          3267 => x"05",
          3268 => x"f0",
          3269 => x"80",
          3270 => x"55",
          3271 => x"90",
          3272 => x"90",
          3273 => x"86",
          3274 => x"80",
          3275 => x"55",
          3276 => x"70",
          3277 => x"05",
          3278 => x"83",
          3279 => x"34",
          3280 => x"75",
          3281 => x"55",
          3282 => x"0b",
          3283 => x"98",
          3284 => x"80",
          3285 => x"9c",
          3286 => x"51",
          3287 => x"33",
          3288 => x"74",
          3289 => x"2e",
          3290 => x"51",
          3291 => x"38",
          3292 => x"38",
          3293 => x"90",
          3294 => x"52",
          3295 => x"72",
          3296 => x"c0",
          3297 => x"27",
          3298 => x"38",
          3299 => x"75",
          3300 => x"ff",
          3301 => x"75",
          3302 => x"06",
          3303 => x"70",
          3304 => x"83",
          3305 => x"0c",
          3306 => x"39",
          3307 => x"51",
          3308 => x"f2",
          3309 => x"16",
          3310 => x"34",
          3311 => x"f0",
          3312 => x"87",
          3313 => x"98",
          3314 => x"38",
          3315 => x"08",
          3316 => x"71",
          3317 => x"98",
          3318 => x"27",
          3319 => x"2e",
          3320 => x"08",
          3321 => x"98",
          3322 => x"08",
          3323 => x"15",
          3324 => x"52",
          3325 => x"ff",
          3326 => x"08",
          3327 => x"52",
          3328 => x"06",
          3329 => x"72",
          3330 => x"38",
          3331 => x"e8",
          3332 => x"0d",
          3333 => x"08",
          3334 => x"ff",
          3335 => x"70",
          3336 => x"71",
          3337 => x"81",
          3338 => x"2b",
          3339 => x"57",
          3340 => x"24",
          3341 => x"33",
          3342 => x"83",
          3343 => x"12",
          3344 => x"07",
          3345 => x"80",
          3346 => x"33",
          3347 => x"83",
          3348 => x"52",
          3349 => x"73",
          3350 => x"34",
          3351 => x"12",
          3352 => x"07",
          3353 => x"51",
          3354 => x"34",
          3355 => x"0b",
          3356 => x"34",
          3357 => x"14",
          3358 => x"d4",
          3359 => x"71",
          3360 => x"70",
          3361 => x"72",
          3362 => x"0d",
          3363 => x"71",
          3364 => x"11",
          3365 => x"88",
          3366 => x"54",
          3367 => x"34",
          3368 => x"08",
          3369 => x"33",
          3370 => x"56",
          3371 => x"33",
          3372 => x"70",
          3373 => x"86",
          3374 => x"b8",
          3375 => x"33",
          3376 => x"06",
          3377 => x"76",
          3378 => x"b8",
          3379 => x"12",
          3380 => x"07",
          3381 => x"71",
          3382 => x"ff",
          3383 => x"54",
          3384 => x"52",
          3385 => x"34",
          3386 => x"33",
          3387 => x"83",
          3388 => x"12",
          3389 => x"ff",
          3390 => x"55",
          3391 => x"70",
          3392 => x"70",
          3393 => x"71",
          3394 => x"05",
          3395 => x"2b",
          3396 => x"52",
          3397 => x"fc",
          3398 => x"71",
          3399 => x"70",
          3400 => x"34",
          3401 => x"08",
          3402 => x"71",
          3403 => x"05",
          3404 => x"88",
          3405 => x"5c",
          3406 => x"15",
          3407 => x"0d",
          3408 => x"d4",
          3409 => x"38",
          3410 => x"fb",
          3411 => x"ff",
          3412 => x"80",
          3413 => x"80",
          3414 => x"fe",
          3415 => x"55",
          3416 => x"34",
          3417 => x"15",
          3418 => x"b8",
          3419 => x"81",
          3420 => x"08",
          3421 => x"80",
          3422 => x"70",
          3423 => x"88",
          3424 => x"b8",
          3425 => x"b8",
          3426 => x"76",
          3427 => x"34",
          3428 => x"52",
          3429 => x"8e",
          3430 => x"70",
          3431 => x"83",
          3432 => x"84",
          3433 => x"2b",
          3434 => x"81",
          3435 => x"cc",
          3436 => x"33",
          3437 => x"70",
          3438 => x"83",
          3439 => x"53",
          3440 => x"8a",
          3441 => x"73",
          3442 => x"33",
          3443 => x"c1",
          3444 => x"38",
          3445 => x"2b",
          3446 => x"71",
          3447 => x"06",
          3448 => x"79",
          3449 => x"74",
          3450 => x"78",
          3451 => x"2e",
          3452 => x"2b",
          3453 => x"70",
          3454 => x"76",
          3455 => x"b8",
          3456 => x"53",
          3457 => x"34",
          3458 => x"33",
          3459 => x"70",
          3460 => x"05",
          3461 => x"2a",
          3462 => x"75",
          3463 => x"53",
          3464 => x"08",
          3465 => x"15",
          3466 => x"86",
          3467 => x"2b",
          3468 => x"5c",
          3469 => x"72",
          3470 => x"70",
          3471 => x"87",
          3472 => x"88",
          3473 => x"15",
          3474 => x"d4",
          3475 => x"12",
          3476 => x"07",
          3477 => x"75",
          3478 => x"84",
          3479 => x"05",
          3480 => x"88",
          3481 => x"57",
          3482 => x"15",
          3483 => x"05",
          3484 => x"3d",
          3485 => x"33",
          3486 => x"79",
          3487 => x"71",
          3488 => x"5b",
          3489 => x"34",
          3490 => x"08",
          3491 => x"33",
          3492 => x"74",
          3493 => x"71",
          3494 => x"5d",
          3495 => x"86",
          3496 => x"b8",
          3497 => x"33",
          3498 => x"06",
          3499 => x"75",
          3500 => x"b8",
          3501 => x"f1",
          3502 => x"d4",
          3503 => x"38",
          3504 => x"b8",
          3505 => x"51",
          3506 => x"84",
          3507 => x"84",
          3508 => x"a0",
          3509 => x"80",
          3510 => x"51",
          3511 => x"08",
          3512 => x"16",
          3513 => x"84",
          3514 => x"84",
          3515 => x"34",
          3516 => x"d4",
          3517 => x"fe",
          3518 => x"06",
          3519 => x"74",
          3520 => x"84",
          3521 => x"84",
          3522 => x"55",
          3523 => x"15",
          3524 => x"dd",
          3525 => x"65",
          3526 => x"d4",
          3527 => x"84",
          3528 => x"38",
          3529 => x"54",
          3530 => x"05",
          3531 => x"ff",
          3532 => x"06",
          3533 => x"ff",
          3534 => x"70",
          3535 => x"07",
          3536 => x"06",
          3537 => x"83",
          3538 => x"33",
          3539 => x"70",
          3540 => x"53",
          3541 => x"5e",
          3542 => x"38",
          3543 => x"88",
          3544 => x"70",
          3545 => x"71",
          3546 => x"56",
          3547 => x"7a",
          3548 => x"58",
          3549 => x"80",
          3550 => x"77",
          3551 => x"59",
          3552 => x"1e",
          3553 => x"2b",
          3554 => x"33",
          3555 => x"90",
          3556 => x"57",
          3557 => x"38",
          3558 => x"33",
          3559 => x"7a",
          3560 => x"71",
          3561 => x"05",
          3562 => x"88",
          3563 => x"48",
          3564 => x"56",
          3565 => x"34",
          3566 => x"11",
          3567 => x"71",
          3568 => x"33",
          3569 => x"70",
          3570 => x"57",
          3571 => x"87",
          3572 => x"70",
          3573 => x"07",
          3574 => x"5a",
          3575 => x"81",
          3576 => x"1f",
          3577 => x"8b",
          3578 => x"73",
          3579 => x"07",
          3580 => x"5f",
          3581 => x"81",
          3582 => x"1f",
          3583 => x"2b",
          3584 => x"14",
          3585 => x"07",
          3586 => x"5f",
          3587 => x"75",
          3588 => x"70",
          3589 => x"71",
          3590 => x"70",
          3591 => x"05",
          3592 => x"84",
          3593 => x"65",
          3594 => x"5d",
          3595 => x"38",
          3596 => x"95",
          3597 => x"84",
          3598 => x"b8",
          3599 => x"52",
          3600 => x"3f",
          3601 => x"34",
          3602 => x"d4",
          3603 => x"0b",
          3604 => x"5c",
          3605 => x"1d",
          3606 => x"d0",
          3607 => x"70",
          3608 => x"5c",
          3609 => x"77",
          3610 => x"70",
          3611 => x"05",
          3612 => x"34",
          3613 => x"d4",
          3614 => x"80",
          3615 => x"80",
          3616 => x"9b",
          3617 => x"e4",
          3618 => x"84",
          3619 => x"11",
          3620 => x"12",
          3621 => x"ff",
          3622 => x"5e",
          3623 => x"34",
          3624 => x"88",
          3625 => x"7b",
          3626 => x"70",
          3627 => x"88",
          3628 => x"f8",
          3629 => x"06",
          3630 => x"5e",
          3631 => x"76",
          3632 => x"05",
          3633 => x"63",
          3634 => x"84",
          3635 => x"ed",
          3636 => x"7b",
          3637 => x"42",
          3638 => x"ff",
          3639 => x"06",
          3640 => x"88",
          3641 => x"70",
          3642 => x"71",
          3643 => x"58",
          3644 => x"f7",
          3645 => x"fa",
          3646 => x"38",
          3647 => x"7b",
          3648 => x"84",
          3649 => x"a0",
          3650 => x"80",
          3651 => x"51",
          3652 => x"08",
          3653 => x"1b",
          3654 => x"84",
          3655 => x"84",
          3656 => x"34",
          3657 => x"d4",
          3658 => x"fe",
          3659 => x"06",
          3660 => x"74",
          3661 => x"05",
          3662 => x"10",
          3663 => x"05",
          3664 => x"81",
          3665 => x"80",
          3666 => x"ff",
          3667 => x"c0",
          3668 => x"82",
          3669 => x"7f",
          3670 => x"3d",
          3671 => x"83",
          3672 => x"2b",
          3673 => x"12",
          3674 => x"07",
          3675 => x"33",
          3676 => x"43",
          3677 => x"5c",
          3678 => x"7a",
          3679 => x"08",
          3680 => x"33",
          3681 => x"74",
          3682 => x"71",
          3683 => x"41",
          3684 => x"64",
          3685 => x"34",
          3686 => x"81",
          3687 => x"ff",
          3688 => x"5a",
          3689 => x"34",
          3690 => x"11",
          3691 => x"71",
          3692 => x"81",
          3693 => x"88",
          3694 => x"45",
          3695 => x"34",
          3696 => x"33",
          3697 => x"83",
          3698 => x"83",
          3699 => x"88",
          3700 => x"55",
          3701 => x"18",
          3702 => x"82",
          3703 => x"2b",
          3704 => x"2b",
          3705 => x"05",
          3706 => x"d4",
          3707 => x"ff",
          3708 => x"ff",
          3709 => x"80",
          3710 => x"80",
          3711 => x"fe",
          3712 => x"56",
          3713 => x"34",
          3714 => x"16",
          3715 => x"b8",
          3716 => x"81",
          3717 => x"08",
          3718 => x"80",
          3719 => x"70",
          3720 => x"88",
          3721 => x"b8",
          3722 => x"b8",
          3723 => x"7f",
          3724 => x"34",
          3725 => x"fc",
          3726 => x"33",
          3727 => x"79",
          3728 => x"71",
          3729 => x"48",
          3730 => x"05",
          3731 => x"b8",
          3732 => x"85",
          3733 => x"2b",
          3734 => x"15",
          3735 => x"2a",
          3736 => x"40",
          3737 => x"87",
          3738 => x"70",
          3739 => x"07",
          3740 => x"59",
          3741 => x"81",
          3742 => x"1f",
          3743 => x"2b",
          3744 => x"33",
          3745 => x"70",
          3746 => x"05",
          3747 => x"5d",
          3748 => x"34",
          3749 => x"08",
          3750 => x"71",
          3751 => x"05",
          3752 => x"2b",
          3753 => x"2a",
          3754 => x"5b",
          3755 => x"34",
          3756 => x"b3",
          3757 => x"71",
          3758 => x"05",
          3759 => x"88",
          3760 => x"5a",
          3761 => x"79",
          3762 => x"70",
          3763 => x"71",
          3764 => x"05",
          3765 => x"88",
          3766 => x"5e",
          3767 => x"86",
          3768 => x"84",
          3769 => x"12",
          3770 => x"ff",
          3771 => x"55",
          3772 => x"84",
          3773 => x"81",
          3774 => x"2b",
          3775 => x"33",
          3776 => x"8f",
          3777 => x"2a",
          3778 => x"5e",
          3779 => x"17",
          3780 => x"70",
          3781 => x"71",
          3782 => x"81",
          3783 => x"ff",
          3784 => x"5e",
          3785 => x"34",
          3786 => x"08",
          3787 => x"33",
          3788 => x"74",
          3789 => x"71",
          3790 => x"05",
          3791 => x"88",
          3792 => x"49",
          3793 => x"57",
          3794 => x"1d",
          3795 => x"84",
          3796 => x"2b",
          3797 => x"14",
          3798 => x"07",
          3799 => x"40",
          3800 => x"7b",
          3801 => x"16",
          3802 => x"2b",
          3803 => x"2a",
          3804 => x"79",
          3805 => x"70",
          3806 => x"71",
          3807 => x"05",
          3808 => x"2b",
          3809 => x"5d",
          3810 => x"75",
          3811 => x"70",
          3812 => x"8b",
          3813 => x"82",
          3814 => x"2b",
          3815 => x"5d",
          3816 => x"34",
          3817 => x"08",
          3818 => x"33",
          3819 => x"56",
          3820 => x"7e",
          3821 => x"3f",
          3822 => x"61",
          3823 => x"06",
          3824 => x"19",
          3825 => x"71",
          3826 => x"33",
          3827 => x"70",
          3828 => x"55",
          3829 => x"85",
          3830 => x"1e",
          3831 => x"8b",
          3832 => x"86",
          3833 => x"2b",
          3834 => x"48",
          3835 => x"05",
          3836 => x"b8",
          3837 => x"33",
          3838 => x"06",
          3839 => x"78",
          3840 => x"b8",
          3841 => x"12",
          3842 => x"07",
          3843 => x"71",
          3844 => x"ff",
          3845 => x"5d",
          3846 => x"40",
          3847 => x"34",
          3848 => x"33",
          3849 => x"83",
          3850 => x"12",
          3851 => x"ff",
          3852 => x"58",
          3853 => x"78",
          3854 => x"06",
          3855 => x"54",
          3856 => x"5f",
          3857 => x"38",
          3858 => x"08",
          3859 => x"df",
          3860 => x"ef",
          3861 => x"0d",
          3862 => x"58",
          3863 => x"54",
          3864 => x"0c",
          3865 => x"d3",
          3866 => x"b8",
          3867 => x"53",
          3868 => x"fe",
          3869 => x"0c",
          3870 => x"0b",
          3871 => x"84",
          3872 => x"76",
          3873 => x"f0",
          3874 => x"75",
          3875 => x"b8",
          3876 => x"81",
          3877 => x"08",
          3878 => x"87",
          3879 => x"b8",
          3880 => x"07",
          3881 => x"2a",
          3882 => x"34",
          3883 => x"22",
          3884 => x"08",
          3885 => x"15",
          3886 => x"54",
          3887 => x"cc",
          3888 => x"33",
          3889 => x"38",
          3890 => x"84",
          3891 => x"fe",
          3892 => x"83",
          3893 => x"51",
          3894 => x"81",
          3895 => x"84",
          3896 => x"12",
          3897 => x"84",
          3898 => x"7e",
          3899 => x"5a",
          3900 => x"26",
          3901 => x"54",
          3902 => x"bd",
          3903 => x"98",
          3904 => x"51",
          3905 => x"81",
          3906 => x"38",
          3907 => x"e2",
          3908 => x"fc",
          3909 => x"83",
          3910 => x"b8",
          3911 => x"80",
          3912 => x"5a",
          3913 => x"38",
          3914 => x"60",
          3915 => x"5c",
          3916 => x"87",
          3917 => x"73",
          3918 => x"38",
          3919 => x"8c",
          3920 => x"d7",
          3921 => x"ff",
          3922 => x"87",
          3923 => x"38",
          3924 => x"80",
          3925 => x"38",
          3926 => x"e4",
          3927 => x"16",
          3928 => x"55",
          3929 => x"d5",
          3930 => x"05",
          3931 => x"05",
          3932 => x"73",
          3933 => x"33",
          3934 => x"73",
          3935 => x"8c",
          3936 => x"38",
          3937 => x"2e",
          3938 => x"e4",
          3939 => x"0a",
          3940 => x"86",
          3941 => x"80",
          3942 => x"0d",
          3943 => x"8c",
          3944 => x"08",
          3945 => x"70",
          3946 => x"8c",
          3947 => x"98",
          3948 => x"72",
          3949 => x"71",
          3950 => x"ff",
          3951 => x"73",
          3952 => x"0d",
          3953 => x"71",
          3954 => x"81",
          3955 => x"83",
          3956 => x"52",
          3957 => x"84",
          3958 => x"81",
          3959 => x"3d",
          3960 => x"53",
          3961 => x"52",
          3962 => x"b8",
          3963 => x"d9",
          3964 => x"34",
          3965 => x"31",
          3966 => x"5c",
          3967 => x"9b",
          3968 => x"2e",
          3969 => x"54",
          3970 => x"33",
          3971 => x"57",
          3972 => x"fe",
          3973 => x"81",
          3974 => x"b8",
          3975 => x"80",
          3976 => x"17",
          3977 => x"84",
          3978 => x"b7",
          3979 => x"d2",
          3980 => x"ba",
          3981 => x"34",
          3982 => x"80",
          3983 => x"c1",
          3984 => x"0b",
          3985 => x"55",
          3986 => x"2a",
          3987 => x"90",
          3988 => x"74",
          3989 => x"34",
          3990 => x"19",
          3991 => x"a5",
          3992 => x"84",
          3993 => x"74",
          3994 => x"81",
          3995 => x"54",
          3996 => x"51",
          3997 => x"80",
          3998 => x"fb",
          3999 => x"2e",
          4000 => x"3d",
          4001 => x"56",
          4002 => x"08",
          4003 => x"84",
          4004 => x"ff",
          4005 => x"81",
          4006 => x"38",
          4007 => x"38",
          4008 => x"a8",
          4009 => x"b4",
          4010 => x"17",
          4011 => x"06",
          4012 => x"b8",
          4013 => x"e3",
          4014 => x"85",
          4015 => x"18",
          4016 => x"ff",
          4017 => x"70",
          4018 => x"5d",
          4019 => x"b5",
          4020 => x"5c",
          4021 => x"06",
          4022 => x"b8",
          4023 => x"93",
          4024 => x"85",
          4025 => x"18",
          4026 => x"ff",
          4027 => x"2b",
          4028 => x"2a",
          4029 => x"ae",
          4030 => x"e4",
          4031 => x"2a",
          4032 => x"08",
          4033 => x"18",
          4034 => x"2e",
          4035 => x"54",
          4036 => x"33",
          4037 => x"08",
          4038 => x"5a",
          4039 => x"38",
          4040 => x"b8",
          4041 => x"88",
          4042 => x"5b",
          4043 => x"09",
          4044 => x"2a",
          4045 => x"08",
          4046 => x"18",
          4047 => x"2e",
          4048 => x"54",
          4049 => x"33",
          4050 => x"08",
          4051 => x"5a",
          4052 => x"38",
          4053 => x"05",
          4054 => x"33",
          4055 => x"81",
          4056 => x"75",
          4057 => x"06",
          4058 => x"5e",
          4059 => x"81",
          4060 => x"70",
          4061 => x"e2",
          4062 => x"7b",
          4063 => x"84",
          4064 => x"17",
          4065 => x"e4",
          4066 => x"27",
          4067 => x"74",
          4068 => x"38",
          4069 => x"08",
          4070 => x"51",
          4071 => x"39",
          4072 => x"17",
          4073 => x"f6",
          4074 => x"2e",
          4075 => x"b8",
          4076 => x"08",
          4077 => x"18",
          4078 => x"5e",
          4079 => x"b8",
          4080 => x"54",
          4081 => x"53",
          4082 => x"3f",
          4083 => x"2e",
          4084 => x"b8",
          4085 => x"08",
          4086 => x"08",
          4087 => x"fd",
          4088 => x"82",
          4089 => x"81",
          4090 => x"05",
          4091 => x"f4",
          4092 => x"81",
          4093 => x"70",
          4094 => x"da",
          4095 => x"7d",
          4096 => x"84",
          4097 => x"17",
          4098 => x"e4",
          4099 => x"27",
          4100 => x"74",
          4101 => x"38",
          4102 => x"08",
          4103 => x"51",
          4104 => x"39",
          4105 => x"08",
          4106 => x"51",
          4107 => x"5b",
          4108 => x"f2",
          4109 => x"59",
          4110 => x"75",
          4111 => x"33",
          4112 => x"78",
          4113 => x"82",
          4114 => x"90",
          4115 => x"1a",
          4116 => x"08",
          4117 => x"38",
          4118 => x"7c",
          4119 => x"81",
          4120 => x"19",
          4121 => x"e4",
          4122 => x"81",
          4123 => x"79",
          4124 => x"06",
          4125 => x"58",
          4126 => x"2a",
          4127 => x"83",
          4128 => x"90",
          4129 => x"81",
          4130 => x"a8",
          4131 => x"1a",
          4132 => x"e1",
          4133 => x"7c",
          4134 => x"38",
          4135 => x"81",
          4136 => x"b8",
          4137 => x"58",
          4138 => x"58",
          4139 => x"83",
          4140 => x"11",
          4141 => x"7e",
          4142 => x"5c",
          4143 => x"75",
          4144 => x"79",
          4145 => x"7a",
          4146 => x"34",
          4147 => x"70",
          4148 => x"1b",
          4149 => x"b7",
          4150 => x"5e",
          4151 => x"06",
          4152 => x"b8",
          4153 => x"83",
          4154 => x"85",
          4155 => x"1a",
          4156 => x"79",
          4157 => x"1b",
          4158 => x"55",
          4159 => x"2b",
          4160 => x"71",
          4161 => x"0b",
          4162 => x"1a",
          4163 => x"08",
          4164 => x"38",
          4165 => x"53",
          4166 => x"3f",
          4167 => x"2e",
          4168 => x"b8",
          4169 => x"08",
          4170 => x"08",
          4171 => x"5c",
          4172 => x"33",
          4173 => x"81",
          4174 => x"33",
          4175 => x"08",
          4176 => x"58",
          4177 => x"38",
          4178 => x"7b",
          4179 => x"7a",
          4180 => x"71",
          4181 => x"34",
          4182 => x"39",
          4183 => x"53",
          4184 => x"3f",
          4185 => x"2e",
          4186 => x"b8",
          4187 => x"08",
          4188 => x"08",
          4189 => x"5e",
          4190 => x"19",
          4191 => x"06",
          4192 => x"53",
          4193 => x"c2",
          4194 => x"54",
          4195 => x"1a",
          4196 => x"5c",
          4197 => x"81",
          4198 => x"08",
          4199 => x"a8",
          4200 => x"b8",
          4201 => x"7e",
          4202 => x"55",
          4203 => x"e3",
          4204 => x"52",
          4205 => x"7c",
          4206 => x"53",
          4207 => x"52",
          4208 => x"b8",
          4209 => x"fb",
          4210 => x"1a",
          4211 => x"08",
          4212 => x"08",
          4213 => x"fb",
          4214 => x"82",
          4215 => x"81",
          4216 => x"19",
          4217 => x"fa",
          4218 => x"76",
          4219 => x"3f",
          4220 => x"10",
          4221 => x"ff",
          4222 => x"1f",
          4223 => x"1f",
          4224 => x"88",
          4225 => x"06",
          4226 => x"70",
          4227 => x"0a",
          4228 => x"7d",
          4229 => x"b9",
          4230 => x"ba",
          4231 => x"bb",
          4232 => x"0d",
          4233 => x"7a",
          4234 => x"76",
          4235 => x"1a",
          4236 => x"08",
          4237 => x"d7",
          4238 => x"76",
          4239 => x"76",
          4240 => x"26",
          4241 => x"f0",
          4242 => x"2e",
          4243 => x"e4",
          4244 => x"e4",
          4245 => x"80",
          4246 => x"55",
          4247 => x"09",
          4248 => x"74",
          4249 => x"04",
          4250 => x"e4",
          4251 => x"51",
          4252 => x"b8",
          4253 => x"e4",
          4254 => x"2e",
          4255 => x"e4",
          4256 => x"dd",
          4257 => x"76",
          4258 => x"79",
          4259 => x"b8",
          4260 => x"84",
          4261 => x"72",
          4262 => x"b8",
          4263 => x"73",
          4264 => x"80",
          4265 => x"81",
          4266 => x"1a",
          4267 => x"57",
          4268 => x"fe",
          4269 => x"51",
          4270 => x"84",
          4271 => x"e4",
          4272 => x"7a",
          4273 => x"75",
          4274 => x"05",
          4275 => x"26",
          4276 => x"84",
          4277 => x"1a",
          4278 => x"0c",
          4279 => x"b8",
          4280 => x"b8",
          4281 => x"80",
          4282 => x"52",
          4283 => x"e4",
          4284 => x"e4",
          4285 => x"0d",
          4286 => x"b9",
          4287 => x"3d",
          4288 => x"58",
          4289 => x"38",
          4290 => x"38",
          4291 => x"55",
          4292 => x"75",
          4293 => x"2a",
          4294 => x"56",
          4295 => x"08",
          4296 => x"98",
          4297 => x"2e",
          4298 => x"19",
          4299 => x"05",
          4300 => x"b8",
          4301 => x"0b",
          4302 => x"04",
          4303 => x"ff",
          4304 => x"2b",
          4305 => x"9c",
          4306 => x"54",
          4307 => x"38",
          4308 => x"19",
          4309 => x"0c",
          4310 => x"ec",
          4311 => x"84",
          4312 => x"81",
          4313 => x"9e",
          4314 => x"e4",
          4315 => x"76",
          4316 => x"ff",
          4317 => x"0c",
          4318 => x"7f",
          4319 => x"5c",
          4320 => x"86",
          4321 => x"17",
          4322 => x"b2",
          4323 => x"9d",
          4324 => x"58",
          4325 => x"1a",
          4326 => x"f5",
          4327 => x"18",
          4328 => x"0c",
          4329 => x"8f",
          4330 => x"8a",
          4331 => x"06",
          4332 => x"51",
          4333 => x"5d",
          4334 => x"08",
          4335 => x"e4",
          4336 => x"08",
          4337 => x"38",
          4338 => x"17",
          4339 => x"84",
          4340 => x"b8",
          4341 => x"82",
          4342 => x"ff",
          4343 => x"08",
          4344 => x"e4",
          4345 => x"80",
          4346 => x"fe",
          4347 => x"27",
          4348 => x"29",
          4349 => x"b4",
          4350 => x"78",
          4351 => x"58",
          4352 => x"74",
          4353 => x"27",
          4354 => x"53",
          4355 => x"b2",
          4356 => x"38",
          4357 => x"18",
          4358 => x"8f",
          4359 => x"08",
          4360 => x"33",
          4361 => x"e4",
          4362 => x"08",
          4363 => x"1a",
          4364 => x"27",
          4365 => x"7b",
          4366 => x"38",
          4367 => x"08",
          4368 => x"51",
          4369 => x"19",
          4370 => x"55",
          4371 => x"38",
          4372 => x"1a",
          4373 => x"75",
          4374 => x"22",
          4375 => x"98",
          4376 => x"0b",
          4377 => x"04",
          4378 => x"84",
          4379 => x"98",
          4380 => x"2e",
          4381 => x"5a",
          4382 => x"82",
          4383 => x"55",
          4384 => x"94",
          4385 => x"52",
          4386 => x"84",
          4387 => x"ff",
          4388 => x"76",
          4389 => x"08",
          4390 => x"82",
          4391 => x"70",
          4392 => x"1d",
          4393 => x"78",
          4394 => x"71",
          4395 => x"55",
          4396 => x"43",
          4397 => x"75",
          4398 => x"5d",
          4399 => x"84",
          4400 => x"08",
          4401 => x"75",
          4402 => x"0c",
          4403 => x"19",
          4404 => x"51",
          4405 => x"e4",
          4406 => x"ef",
          4407 => x"34",
          4408 => x"84",
          4409 => x"1a",
          4410 => x"33",
          4411 => x"fe",
          4412 => x"a0",
          4413 => x"19",
          4414 => x"fe",
          4415 => x"06",
          4416 => x"06",
          4417 => x"18",
          4418 => x"1f",
          4419 => x"5e",
          4420 => x"55",
          4421 => x"75",
          4422 => x"38",
          4423 => x"1d",
          4424 => x"3d",
          4425 => x"8d",
          4426 => x"81",
          4427 => x"19",
          4428 => x"07",
          4429 => x"77",
          4430 => x"f3",
          4431 => x"83",
          4432 => x"11",
          4433 => x"52",
          4434 => x"38",
          4435 => x"79",
          4436 => x"62",
          4437 => x"8c",
          4438 => x"86",
          4439 => x"2e",
          4440 => x"dd",
          4441 => x"63",
          4442 => x"5e",
          4443 => x"ff",
          4444 => x"c0",
          4445 => x"57",
          4446 => x"05",
          4447 => x"7f",
          4448 => x"59",
          4449 => x"2e",
          4450 => x"0c",
          4451 => x"0d",
          4452 => x"5c",
          4453 => x"3f",
          4454 => x"e4",
          4455 => x"40",
          4456 => x"1b",
          4457 => x"b4",
          4458 => x"83",
          4459 => x"2e",
          4460 => x"54",
          4461 => x"33",
          4462 => x"08",
          4463 => x"57",
          4464 => x"81",
          4465 => x"58",
          4466 => x"8b",
          4467 => x"06",
          4468 => x"81",
          4469 => x"2a",
          4470 => x"ef",
          4471 => x"2e",
          4472 => x"7d",
          4473 => x"75",
          4474 => x"05",
          4475 => x"ff",
          4476 => x"e4",
          4477 => x"ab",
          4478 => x"38",
          4479 => x"70",
          4480 => x"05",
          4481 => x"5a",
          4482 => x"dc",
          4483 => x"ff",
          4484 => x"52",
          4485 => x"e4",
          4486 => x"2e",
          4487 => x"0c",
          4488 => x"1b",
          4489 => x"51",
          4490 => x"e4",
          4491 => x"a4",
          4492 => x"34",
          4493 => x"84",
          4494 => x"1c",
          4495 => x"33",
          4496 => x"fd",
          4497 => x"a0",
          4498 => x"1b",
          4499 => x"fd",
          4500 => x"ab",
          4501 => x"42",
          4502 => x"2a",
          4503 => x"38",
          4504 => x"70",
          4505 => x"59",
          4506 => x"81",
          4507 => x"51",
          4508 => x"5a",
          4509 => x"d9",
          4510 => x"fe",
          4511 => x"ac",
          4512 => x"33",
          4513 => x"c7",
          4514 => x"9a",
          4515 => x"42",
          4516 => x"70",
          4517 => x"55",
          4518 => x"18",
          4519 => x"33",
          4520 => x"75",
          4521 => x"fe",
          4522 => x"a1",
          4523 => x"10",
          4524 => x"1b",
          4525 => x"84",
          4526 => x"fe",
          4527 => x"8c",
          4528 => x"70",
          4529 => x"80",
          4530 => x"38",
          4531 => x"41",
          4532 => x"81",
          4533 => x"84",
          4534 => x"0d",
          4535 => x"bc",
          4536 => x"ea",
          4537 => x"13",
          4538 => x"5e",
          4539 => x"8c",
          4540 => x"74",
          4541 => x"10",
          4542 => x"f4",
          4543 => x"8c",
          4544 => x"81",
          4545 => x"59",
          4546 => x"02",
          4547 => x"58",
          4548 => x"80",
          4549 => x"94",
          4550 => x"58",
          4551 => x"77",
          4552 => x"81",
          4553 => x"ef",
          4554 => x"7a",
          4555 => x"b8",
          4556 => x"58",
          4557 => x"81",
          4558 => x"90",
          4559 => x"60",
          4560 => x"a1",
          4561 => x"25",
          4562 => x"38",
          4563 => x"57",
          4564 => x"b9",
          4565 => x"74",
          4566 => x"84",
          4567 => x"77",
          4568 => x"7a",
          4569 => x"79",
          4570 => x"81",
          4571 => x"38",
          4572 => x"a0",
          4573 => x"16",
          4574 => x"38",
          4575 => x"19",
          4576 => x"34",
          4577 => x"51",
          4578 => x"8b",
          4579 => x"27",
          4580 => x"e4",
          4581 => x"08",
          4582 => x"09",
          4583 => x"db",
          4584 => x"02",
          4585 => x"58",
          4586 => x"5b",
          4587 => x"8c",
          4588 => x"b8",
          4589 => x"51",
          4590 => x"56",
          4591 => x"84",
          4592 => x"98",
          4593 => x"08",
          4594 => x"33",
          4595 => x"82",
          4596 => x"18",
          4597 => x"3f",
          4598 => x"38",
          4599 => x"0c",
          4600 => x"08",
          4601 => x"2e",
          4602 => x"25",
          4603 => x"81",
          4604 => x"2e",
          4605 => x"ee",
          4606 => x"84",
          4607 => x"38",
          4608 => x"38",
          4609 => x"1b",
          4610 => x"08",
          4611 => x"38",
          4612 => x"84",
          4613 => x"1c",
          4614 => x"3f",
          4615 => x"38",
          4616 => x"0c",
          4617 => x"0b",
          4618 => x"70",
          4619 => x"74",
          4620 => x"7b",
          4621 => x"57",
          4622 => x"ff",
          4623 => x"08",
          4624 => x"7c",
          4625 => x"34",
          4626 => x"98",
          4627 => x"80",
          4628 => x"fe",
          4629 => x"51",
          4630 => x"56",
          4631 => x"c7",
          4632 => x"18",
          4633 => x"51",
          4634 => x"77",
          4635 => x"84",
          4636 => x"18",
          4637 => x"a0",
          4638 => x"33",
          4639 => x"84",
          4640 => x"7f",
          4641 => x"53",
          4642 => x"b8",
          4643 => x"fe",
          4644 => x"56",
          4645 => x"81",
          4646 => x"5a",
          4647 => x"06",
          4648 => x"38",
          4649 => x"41",
          4650 => x"1c",
          4651 => x"33",
          4652 => x"82",
          4653 => x"1c",
          4654 => x"3f",
          4655 => x"38",
          4656 => x"0c",
          4657 => x"1c",
          4658 => x"06",
          4659 => x"8f",
          4660 => x"34",
          4661 => x"34",
          4662 => x"5a",
          4663 => x"8b",
          4664 => x"1b",
          4665 => x"33",
          4666 => x"05",
          4667 => x"75",
          4668 => x"57",
          4669 => x"38",
          4670 => x"38",
          4671 => x"76",
          4672 => x"34",
          4673 => x"7d",
          4674 => x"08",
          4675 => x"38",
          4676 => x"38",
          4677 => x"08",
          4678 => x"33",
          4679 => x"84",
          4680 => x"b8",
          4681 => x"08",
          4682 => x"08",
          4683 => x"fb",
          4684 => x"82",
          4685 => x"81",
          4686 => x"05",
          4687 => x"cf",
          4688 => x"76",
          4689 => x"56",
          4690 => x"fa",
          4691 => x"57",
          4692 => x"fa",
          4693 => x"fe",
          4694 => x"53",
          4695 => x"92",
          4696 => x"09",
          4697 => x"08",
          4698 => x"1d",
          4699 => x"27",
          4700 => x"82",
          4701 => x"56",
          4702 => x"58",
          4703 => x"87",
          4704 => x"81",
          4705 => x"fe",
          4706 => x"1c",
          4707 => x"52",
          4708 => x"fc",
          4709 => x"a0",
          4710 => x"18",
          4711 => x"39",
          4712 => x"40",
          4713 => x"98",
          4714 => x"ac",
          4715 => x"80",
          4716 => x"22",
          4717 => x"2e",
          4718 => x"22",
          4719 => x"95",
          4720 => x"ff",
          4721 => x"26",
          4722 => x"11",
          4723 => x"d4",
          4724 => x"30",
          4725 => x"94",
          4726 => x"80",
          4727 => x"1c",
          4728 => x"56",
          4729 => x"85",
          4730 => x"70",
          4731 => x"5b",
          4732 => x"80",
          4733 => x"05",
          4734 => x"70",
          4735 => x"8a",
          4736 => x"88",
          4737 => x"96",
          4738 => x"81",
          4739 => x"81",
          4740 => x"0b",
          4741 => x"11",
          4742 => x"89",
          4743 => x"13",
          4744 => x"9c",
          4745 => x"71",
          4746 => x"14",
          4747 => x"33",
          4748 => x"33",
          4749 => x"5f",
          4750 => x"77",
          4751 => x"16",
          4752 => x"7b",
          4753 => x"81",
          4754 => x"96",
          4755 => x"57",
          4756 => x"07",
          4757 => x"e4",
          4758 => x"ff",
          4759 => x"81",
          4760 => x"7a",
          4761 => x"05",
          4762 => x"5b",
          4763 => x"57",
          4764 => x"39",
          4765 => x"80",
          4766 => x"57",
          4767 => x"81",
          4768 => x"08",
          4769 => x"1f",
          4770 => x"fe",
          4771 => x"59",
          4772 => x"5a",
          4773 => x"1c",
          4774 => x"76",
          4775 => x"72",
          4776 => x"38",
          4777 => x"55",
          4778 => x"34",
          4779 => x"89",
          4780 => x"79",
          4781 => x"83",
          4782 => x"70",
          4783 => x"5d",
          4784 => x"0d",
          4785 => x"80",
          4786 => x"af",
          4787 => x"dc",
          4788 => x"81",
          4789 => x"0c",
          4790 => x"42",
          4791 => x"73",
          4792 => x"61",
          4793 => x"53",
          4794 => x"73",
          4795 => x"ff",
          4796 => x"56",
          4797 => x"83",
          4798 => x"30",
          4799 => x"57",
          4800 => x"74",
          4801 => x"80",
          4802 => x"0b",
          4803 => x"06",
          4804 => x"ab",
          4805 => x"16",
          4806 => x"54",
          4807 => x"06",
          4808 => x"fe",
          4809 => x"5d",
          4810 => x"70",
          4811 => x"73",
          4812 => x"39",
          4813 => x"70",
          4814 => x"55",
          4815 => x"70",
          4816 => x"72",
          4817 => x"32",
          4818 => x"51",
          4819 => x"1d",
          4820 => x"41",
          4821 => x"38",
          4822 => x"81",
          4823 => x"83",
          4824 => x"38",
          4825 => x"93",
          4826 => x"70",
          4827 => x"2e",
          4828 => x"0b",
          4829 => x"de",
          4830 => x"b8",
          4831 => x"73",
          4832 => x"25",
          4833 => x"80",
          4834 => x"62",
          4835 => x"2e",
          4836 => x"30",
          4837 => x"59",
          4838 => x"75",
          4839 => x"84",
          4840 => x"38",
          4841 => x"38",
          4842 => x"22",
          4843 => x"2a",
          4844 => x"ae",
          4845 => x"17",
          4846 => x"19",
          4847 => x"fe",
          4848 => x"ff",
          4849 => x"7a",
          4850 => x"ff",
          4851 => x"f1",
          4852 => x"19",
          4853 => x"ae",
          4854 => x"05",
          4855 => x"8f",
          4856 => x"7c",
          4857 => x"8b",
          4858 => x"70",
          4859 => x"72",
          4860 => x"78",
          4861 => x"54",
          4862 => x"74",
          4863 => x"32",
          4864 => x"54",
          4865 => x"83",
          4866 => x"83",
          4867 => x"30",
          4868 => x"07",
          4869 => x"83",
          4870 => x"38",
          4871 => x"07",
          4872 => x"56",
          4873 => x"fc",
          4874 => x"15",
          4875 => x"74",
          4876 => x"76",
          4877 => x"88",
          4878 => x"58",
          4879 => x"83",
          4880 => x"38",
          4881 => x"9d",
          4882 => x"2e",
          4883 => x"82",
          4884 => x"85",
          4885 => x"1d",
          4886 => x"b8",
          4887 => x"84",
          4888 => x"38",
          4889 => x"81",
          4890 => x"81",
          4891 => x"38",
          4892 => x"82",
          4893 => x"73",
          4894 => x"f9",
          4895 => x"11",
          4896 => x"a0",
          4897 => x"85",
          4898 => x"39",
          4899 => x"09",
          4900 => x"54",
          4901 => x"a0",
          4902 => x"23",
          4903 => x"54",
          4904 => x"73",
          4905 => x"13",
          4906 => x"a0",
          4907 => x"51",
          4908 => x"ab",
          4909 => x"08",
          4910 => x"06",
          4911 => x"33",
          4912 => x"74",
          4913 => x"08",
          4914 => x"11",
          4915 => x"2b",
          4916 => x"7d",
          4917 => x"1d",
          4918 => x"b7",
          4919 => x"fe",
          4920 => x"88",
          4921 => x"76",
          4922 => x"82",
          4923 => x"59",
          4924 => x"fd",
          4925 => x"98",
          4926 => x"88",
          4927 => x"d6",
          4928 => x"80",
          4929 => x"0d",
          4930 => x"81",
          4931 => x"1d",
          4932 => x"79",
          4933 => x"5a",
          4934 => x"83",
          4935 => x"3f",
          4936 => x"06",
          4937 => x"78",
          4938 => x"06",
          4939 => x"74",
          4940 => x"80",
          4941 => x"0b",
          4942 => x"06",
          4943 => x"e0",
          4944 => x"19",
          4945 => x"54",
          4946 => x"06",
          4947 => x"15",
          4948 => x"82",
          4949 => x"ff",
          4950 => x"38",
          4951 => x"e0",
          4952 => x"56",
          4953 => x"74",
          4954 => x"55",
          4955 => x"39",
          4956 => x"06",
          4957 => x"38",
          4958 => x"a0",
          4959 => x"81",
          4960 => x"33",
          4961 => x"71",
          4962 => x"0c",
          4963 => x"a0",
          4964 => x"74",
          4965 => x"5a",
          4966 => x"ff",
          4967 => x"33",
          4968 => x"81",
          4969 => x"74",
          4970 => x"f2",
          4971 => x"93",
          4972 => x"69",
          4973 => x"42",
          4974 => x"08",
          4975 => x"85",
          4976 => x"33",
          4977 => x"2e",
          4978 => x"ba",
          4979 => x"33",
          4980 => x"75",
          4981 => x"08",
          4982 => x"85",
          4983 => x"fe",
          4984 => x"2e",
          4985 => x"bb",
          4986 => x"ff",
          4987 => x"80",
          4988 => x"75",
          4989 => x"81",
          4990 => x"51",
          4991 => x"08",
          4992 => x"56",
          4993 => x"80",
          4994 => x"06",
          4995 => x"80",
          4996 => x"b4",
          4997 => x"54",
          4998 => x"18",
          4999 => x"84",
          5000 => x"ff",
          5001 => x"84",
          5002 => x"33",
          5003 => x"07",
          5004 => x"d5",
          5005 => x"8b",
          5006 => x"61",
          5007 => x"2e",
          5008 => x"26",
          5009 => x"80",
          5010 => x"5e",
          5011 => x"06",
          5012 => x"80",
          5013 => x"57",
          5014 => x"83",
          5015 => x"2b",
          5016 => x"70",
          5017 => x"07",
          5018 => x"75",
          5019 => x"82",
          5020 => x"11",
          5021 => x"8d",
          5022 => x"78",
          5023 => x"c5",
          5024 => x"18",
          5025 => x"c4",
          5026 => x"87",
          5027 => x"c9",
          5028 => x"40",
          5029 => x"06",
          5030 => x"38",
          5031 => x"33",
          5032 => x"a4",
          5033 => x"82",
          5034 => x"2b",
          5035 => x"88",
          5036 => x"5a",
          5037 => x"33",
          5038 => x"07",
          5039 => x"81",
          5040 => x"05",
          5041 => x"78",
          5042 => x"8e",
          5043 => x"b8",
          5044 => x"84",
          5045 => x"f5",
          5046 => x"ff",
          5047 => x"9f",
          5048 => x"82",
          5049 => x"19",
          5050 => x"7b",
          5051 => x"83",
          5052 => x"5c",
          5053 => x"38",
          5054 => x"55",
          5055 => x"19",
          5056 => x"56",
          5057 => x"8d",
          5058 => x"38",
          5059 => x"90",
          5060 => x"34",
          5061 => x"77",
          5062 => x"5d",
          5063 => x"18",
          5064 => x"0c",
          5065 => x"77",
          5066 => x"04",
          5067 => x"3d",
          5068 => x"81",
          5069 => x"26",
          5070 => x"06",
          5071 => x"87",
          5072 => x"d4",
          5073 => x"5b",
          5074 => x"70",
          5075 => x"5a",
          5076 => x"e0",
          5077 => x"ff",
          5078 => x"38",
          5079 => x"55",
          5080 => x"75",
          5081 => x"77",
          5082 => x"30",
          5083 => x"5d",
          5084 => x"38",
          5085 => x"7c",
          5086 => x"a9",
          5087 => x"77",
          5088 => x"7d",
          5089 => x"39",
          5090 => x"e9",
          5091 => x"59",
          5092 => x"80",
          5093 => x"83",
          5094 => x"a6",
          5095 => x"59",
          5096 => x"7a",
          5097 => x"33",
          5098 => x"71",
          5099 => x"70",
          5100 => x"33",
          5101 => x"40",
          5102 => x"ff",
          5103 => x"25",
          5104 => x"33",
          5105 => x"31",
          5106 => x"05",
          5107 => x"5b",
          5108 => x"80",
          5109 => x"18",
          5110 => x"55",
          5111 => x"81",
          5112 => x"17",
          5113 => x"b8",
          5114 => x"55",
          5115 => x"58",
          5116 => x"33",
          5117 => x"58",
          5118 => x"06",
          5119 => x"57",
          5120 => x"38",
          5121 => x"80",
          5122 => x"bc",
          5123 => x"82",
          5124 => x"0b",
          5125 => x"7b",
          5126 => x"81",
          5127 => x"77",
          5128 => x"84",
          5129 => x"d1",
          5130 => x"ee",
          5131 => x"7b",
          5132 => x"81",
          5133 => x"1b",
          5134 => x"80",
          5135 => x"85",
          5136 => x"40",
          5137 => x"33",
          5138 => x"71",
          5139 => x"77",
          5140 => x"2e",
          5141 => x"8d",
          5142 => x"b8",
          5143 => x"58",
          5144 => x"0b",
          5145 => x"5d",
          5146 => x"b8",
          5147 => x"0b",
          5148 => x"5a",
          5149 => x"7a",
          5150 => x"31",
          5151 => x"80",
          5152 => x"e1",
          5153 => x"e4",
          5154 => x"05",
          5155 => x"33",
          5156 => x"42",
          5157 => x"75",
          5158 => x"57",
          5159 => x"58",
          5160 => x"80",
          5161 => x"57",
          5162 => x"f9",
          5163 => x"b4",
          5164 => x"17",
          5165 => x"06",
          5166 => x"b8",
          5167 => x"b0",
          5168 => x"2e",
          5169 => x"b4",
          5170 => x"84",
          5171 => x"b6",
          5172 => x"5e",
          5173 => x"06",
          5174 => x"33",
          5175 => x"88",
          5176 => x"07",
          5177 => x"41",
          5178 => x"8b",
          5179 => x"f8",
          5180 => x"33",
          5181 => x"88",
          5182 => x"07",
          5183 => x"44",
          5184 => x"8a",
          5185 => x"f8",
          5186 => x"33",
          5187 => x"88",
          5188 => x"07",
          5189 => x"1e",
          5190 => x"33",
          5191 => x"88",
          5192 => x"07",
          5193 => x"90",
          5194 => x"45",
          5195 => x"34",
          5196 => x"7c",
          5197 => x"23",
          5198 => x"80",
          5199 => x"7b",
          5200 => x"7f",
          5201 => x"b4",
          5202 => x"81",
          5203 => x"3f",
          5204 => x"81",
          5205 => x"08",
          5206 => x"18",
          5207 => x"27",
          5208 => x"82",
          5209 => x"08",
          5210 => x"80",
          5211 => x"8a",
          5212 => x"fc",
          5213 => x"e2",
          5214 => x"5a",
          5215 => x"17",
          5216 => x"e4",
          5217 => x"71",
          5218 => x"14",
          5219 => x"33",
          5220 => x"82",
          5221 => x"f5",
          5222 => x"f9",
          5223 => x"75",
          5224 => x"77",
          5225 => x"75",
          5226 => x"39",
          5227 => x"08",
          5228 => x"51",
          5229 => x"f0",
          5230 => x"64",
          5231 => x"ff",
          5232 => x"e9",
          5233 => x"70",
          5234 => x"80",
          5235 => x"2e",
          5236 => x"54",
          5237 => x"10",
          5238 => x"55",
          5239 => x"74",
          5240 => x"38",
          5241 => x"0c",
          5242 => x"80",
          5243 => x"51",
          5244 => x"54",
          5245 => x"0d",
          5246 => x"92",
          5247 => x"70",
          5248 => x"89",
          5249 => x"ff",
          5250 => x"2e",
          5251 => x"e4",
          5252 => x"59",
          5253 => x"78",
          5254 => x"12",
          5255 => x"38",
          5256 => x"54",
          5257 => x"89",
          5258 => x"57",
          5259 => x"54",
          5260 => x"38",
          5261 => x"70",
          5262 => x"07",
          5263 => x"38",
          5264 => x"7b",
          5265 => x"98",
          5266 => x"79",
          5267 => x"3d",
          5268 => x"05",
          5269 => x"2e",
          5270 => x"9d",
          5271 => x"05",
          5272 => x"e4",
          5273 => x"2e",
          5274 => x"75",
          5275 => x"04",
          5276 => x"52",
          5277 => x"08",
          5278 => x"81",
          5279 => x"80",
          5280 => x"83",
          5281 => x"38",
          5282 => x"38",
          5283 => x"80",
          5284 => x"33",
          5285 => x"61",
          5286 => x"7d",
          5287 => x"8e",
          5288 => x"a1",
          5289 => x"91",
          5290 => x"17",
          5291 => x"9a",
          5292 => x"7d",
          5293 => x"38",
          5294 => x"80",
          5295 => x"1c",
          5296 => x"55",
          5297 => x"2e",
          5298 => x"7d",
          5299 => x"7c",
          5300 => x"26",
          5301 => x"0c",
          5302 => x"33",
          5303 => x"25",
          5304 => x"5e",
          5305 => x"82",
          5306 => x"84",
          5307 => x"91",
          5308 => x"7d",
          5309 => x"5a",
          5310 => x"81",
          5311 => x"77",
          5312 => x"08",
          5313 => x"67",
          5314 => x"88",
          5315 => x"57",
          5316 => x"7a",
          5317 => x"33",
          5318 => x"88",
          5319 => x"07",
          5320 => x"60",
          5321 => x"52",
          5322 => x"22",
          5323 => x"80",
          5324 => x"1a",
          5325 => x"74",
          5326 => x"2e",
          5327 => x"8a",
          5328 => x"5b",
          5329 => x"25",
          5330 => x"38",
          5331 => x"80",
          5332 => x"51",
          5333 => x"08",
          5334 => x"83",
          5335 => x"ff",
          5336 => x"56",
          5337 => x"91",
          5338 => x"2a",
          5339 => x"b8",
          5340 => x"ed",
          5341 => x"e5",
          5342 => x"dd",
          5343 => x"b8",
          5344 => x"76",
          5345 => x"76",
          5346 => x"95",
          5347 => x"2b",
          5348 => x"5e",
          5349 => x"7b",
          5350 => x"51",
          5351 => x"08",
          5352 => x"81",
          5353 => x"2e",
          5354 => x"ff",
          5355 => x"52",
          5356 => x"b8",
          5357 => x"08",
          5358 => x"5b",
          5359 => x"16",
          5360 => x"07",
          5361 => x"7a",
          5362 => x"39",
          5363 => x"95",
          5364 => x"33",
          5365 => x"90",
          5366 => x"80",
          5367 => x"17",
          5368 => x"cc",
          5369 => x"0b",
          5370 => x"80",
          5371 => x"17",
          5372 => x"09",
          5373 => x"39",
          5374 => x"5d",
          5375 => x"83",
          5376 => x"81",
          5377 => x"b8",
          5378 => x"a3",
          5379 => x"2e",
          5380 => x"b4",
          5381 => x"90",
          5382 => x"bc",
          5383 => x"81",
          5384 => x"70",
          5385 => x"a4",
          5386 => x"2e",
          5387 => x"b8",
          5388 => x"08",
          5389 => x"08",
          5390 => x"ff",
          5391 => x"82",
          5392 => x"81",
          5393 => x"05",
          5394 => x"ff",
          5395 => x"39",
          5396 => x"af",
          5397 => x"a2",
          5398 => x"80",
          5399 => x"9c",
          5400 => x"77",
          5401 => x"22",
          5402 => x"56",
          5403 => x"75",
          5404 => x"56",
          5405 => x"76",
          5406 => x"79",
          5407 => x"08",
          5408 => x"81",
          5409 => x"3d",
          5410 => x"5d",
          5411 => x"80",
          5412 => x"80",
          5413 => x"80",
          5414 => x"1b",
          5415 => x"b7",
          5416 => x"76",
          5417 => x"74",
          5418 => x"06",
          5419 => x"ed",
          5420 => x"71",
          5421 => x"ef",
          5422 => x"60",
          5423 => x"81",
          5424 => x"76",
          5425 => x"75",
          5426 => x"81",
          5427 => x"2e",
          5428 => x"60",
          5429 => x"1a",
          5430 => x"27",
          5431 => x"78",
          5432 => x"74",
          5433 => x"7c",
          5434 => x"83",
          5435 => x"27",
          5436 => x"54",
          5437 => x"51",
          5438 => x"08",
          5439 => x"57",
          5440 => x"19",
          5441 => x"9e",
          5442 => x"b8",
          5443 => x"05",
          5444 => x"34",
          5445 => x"89",
          5446 => x"19",
          5447 => x"1a",
          5448 => x"7b",
          5449 => x"b8",
          5450 => x"84",
          5451 => x"74",
          5452 => x"57",
          5453 => x"31",
          5454 => x"7b",
          5455 => x"2e",
          5456 => x"71",
          5457 => x"81",
          5458 => x"53",
          5459 => x"ff",
          5460 => x"80",
          5461 => x"75",
          5462 => x"60",
          5463 => x"79",
          5464 => x"77",
          5465 => x"81",
          5466 => x"59",
          5467 => x"fe",
          5468 => x"33",
          5469 => x"16",
          5470 => x"81",
          5471 => x"70",
          5472 => x"9e",
          5473 => x"08",
          5474 => x"38",
          5475 => x"b4",
          5476 => x"b8",
          5477 => x"08",
          5478 => x"55",
          5479 => x"d4",
          5480 => x"1a",
          5481 => x"33",
          5482 => x"fe",
          5483 => x"1a",
          5484 => x"08",
          5485 => x"84",
          5486 => x"81",
          5487 => x"84",
          5488 => x"fb",
          5489 => x"fb",
          5490 => x"81",
          5491 => x"0d",
          5492 => x"0b",
          5493 => x"04",
          5494 => x"40",
          5495 => x"57",
          5496 => x"56",
          5497 => x"55",
          5498 => x"22",
          5499 => x"2e",
          5500 => x"76",
          5501 => x"33",
          5502 => x"33",
          5503 => x"87",
          5504 => x"94",
          5505 => x"77",
          5506 => x"80",
          5507 => x"06",
          5508 => x"11",
          5509 => x"5a",
          5510 => x"38",
          5511 => x"84",
          5512 => x"38",
          5513 => x"98",
          5514 => x"74",
          5515 => x"08",
          5516 => x"98",
          5517 => x"fe",
          5518 => x"f0",
          5519 => x"b0",
          5520 => x"2e",
          5521 => x"2a",
          5522 => x"38",
          5523 => x"38",
          5524 => x"53",
          5525 => x"9b",
          5526 => x"a1",
          5527 => x"56",
          5528 => x"80",
          5529 => x"57",
          5530 => x"33",
          5531 => x"16",
          5532 => x"83",
          5533 => x"79",
          5534 => x"1e",
          5535 => x"1f",
          5536 => x"5e",
          5537 => x"56",
          5538 => x"38",
          5539 => x"07",
          5540 => x"75",
          5541 => x"04",
          5542 => x"0d",
          5543 => x"c8",
          5544 => x"9c",
          5545 => x"06",
          5546 => x"79",
          5547 => x"b4",
          5548 => x"0b",
          5549 => x"7f",
          5550 => x"38",
          5551 => x"81",
          5552 => x"84",
          5553 => x"ff",
          5554 => x"7b",
          5555 => x"83",
          5556 => x"7e",
          5557 => x"38",
          5558 => x"70",
          5559 => x"75",
          5560 => x"19",
          5561 => x"16",
          5562 => x"17",
          5563 => x"81",
          5564 => x"09",
          5565 => x"e4",
          5566 => x"a8",
          5567 => x"5d",
          5568 => x"f0",
          5569 => x"2e",
          5570 => x"54",
          5571 => x"53",
          5572 => x"98",
          5573 => x"94",
          5574 => x"26",
          5575 => x"81",
          5576 => x"94",
          5577 => x"1c",
          5578 => x"08",
          5579 => x"84",
          5580 => x"08",
          5581 => x"fd",
          5582 => x"ab",
          5583 => x"84",
          5584 => x"39",
          5585 => x"16",
          5586 => x"ff",
          5587 => x"81",
          5588 => x"17",
          5589 => x"31",
          5590 => x"89",
          5591 => x"2e",
          5592 => x"54",
          5593 => x"53",
          5594 => x"96",
          5595 => x"81",
          5596 => x"84",
          5597 => x"f9",
          5598 => x"f9",
          5599 => x"53",
          5600 => x"52",
          5601 => x"e4",
          5602 => x"08",
          5603 => x"17",
          5604 => x"27",
          5605 => x"77",
          5606 => x"38",
          5607 => x"08",
          5608 => x"51",
          5609 => x"12",
          5610 => x"f4",
          5611 => x"0b",
          5612 => x"04",
          5613 => x"84",
          5614 => x"f5",
          5615 => x"80",
          5616 => x"80",
          5617 => x"80",
          5618 => x"19",
          5619 => x"b5",
          5620 => x"79",
          5621 => x"86",
          5622 => x"2e",
          5623 => x"5a",
          5624 => x"38",
          5625 => x"38",
          5626 => x"81",
          5627 => x"84",
          5628 => x"ff",
          5629 => x"75",
          5630 => x"11",
          5631 => x"18",
          5632 => x"83",
          5633 => x"9a",
          5634 => x"9b",
          5635 => x"19",
          5636 => x"c1",
          5637 => x"34",
          5638 => x"34",
          5639 => x"34",
          5640 => x"34",
          5641 => x"34",
          5642 => x"0b",
          5643 => x"34",
          5644 => x"81",
          5645 => x"96",
          5646 => x"19",
          5647 => x"90",
          5648 => x"8d",
          5649 => x"08",
          5650 => x"33",
          5651 => x"56",
          5652 => x"84",
          5653 => x"17",
          5654 => x"e4",
          5655 => x"27",
          5656 => x"74",
          5657 => x"38",
          5658 => x"08",
          5659 => x"51",
          5660 => x"e8",
          5661 => x"18",
          5662 => x"18",
          5663 => x"34",
          5664 => x"34",
          5665 => x"34",
          5666 => x"34",
          5667 => x"34",
          5668 => x"0b",
          5669 => x"34",
          5670 => x"81",
          5671 => x"94",
          5672 => x"19",
          5673 => x"90",
          5674 => x"33",
          5675 => x"e4",
          5676 => x"38",
          5677 => x"39",
          5678 => x"fb",
          5679 => x"84",
          5680 => x"74",
          5681 => x"72",
          5682 => x"71",
          5683 => x"84",
          5684 => x"96",
          5685 => x"75",
          5686 => x"b8",
          5687 => x"13",
          5688 => x"b8",
          5689 => x"38",
          5690 => x"f6",
          5691 => x"5b",
          5692 => x"81",
          5693 => x"52",
          5694 => x"38",
          5695 => x"c0",
          5696 => x"70",
          5697 => x"b8",
          5698 => x"0b",
          5699 => x"04",
          5700 => x"06",
          5701 => x"38",
          5702 => x"05",
          5703 => x"38",
          5704 => x"79",
          5705 => x"05",
          5706 => x"33",
          5707 => x"99",
          5708 => x"ff",
          5709 => x"70",
          5710 => x"81",
          5711 => x"9f",
          5712 => x"81",
          5713 => x"74",
          5714 => x"9f",
          5715 => x"80",
          5716 => x"5b",
          5717 => x"7a",
          5718 => x"f7",
          5719 => x"39",
          5720 => x"cc",
          5721 => x"3f",
          5722 => x"e4",
          5723 => x"b8",
          5724 => x"5c",
          5725 => x"c5",
          5726 => x"84",
          5727 => x"80",
          5728 => x"5a",
          5729 => x"b2",
          5730 => x"57",
          5731 => x"63",
          5732 => x"88",
          5733 => x"57",
          5734 => x"98",
          5735 => x"98",
          5736 => x"84",
          5737 => x"85",
          5738 => x"0d",
          5739 => x"71",
          5740 => x"07",
          5741 => x"7a",
          5742 => x"b8",
          5743 => x"9e",
          5744 => x"e6",
          5745 => x"80",
          5746 => x"52",
          5747 => x"84",
          5748 => x"08",
          5749 => x"0c",
          5750 => x"3d",
          5751 => x"58",
          5752 => x"d8",
          5753 => x"7a",
          5754 => x"e4",
          5755 => x"92",
          5756 => x"56",
          5757 => x"84",
          5758 => x"5d",
          5759 => x"53",
          5760 => x"ff",
          5761 => x"80",
          5762 => x"76",
          5763 => x"80",
          5764 => x"12",
          5765 => x"33",
          5766 => x"2e",
          5767 => x"0c",
          5768 => x"3f",
          5769 => x"e4",
          5770 => x"51",
          5771 => x"08",
          5772 => x"80",
          5773 => x"12",
          5774 => x"33",
          5775 => x"2e",
          5776 => x"38",
          5777 => x"ff",
          5778 => x"59",
          5779 => x"b4",
          5780 => x"78",
          5781 => x"b8",
          5782 => x"3f",
          5783 => x"79",
          5784 => x"81",
          5785 => x"57",
          5786 => x"78",
          5787 => x"9c",
          5788 => x"18",
          5789 => x"ff",
          5790 => x"75",
          5791 => x"e6",
          5792 => x"34",
          5793 => x"bd",
          5794 => x"80",
          5795 => x"10",
          5796 => x"33",
          5797 => x"2e",
          5798 => x"33",
          5799 => x"1a",
          5800 => x"57",
          5801 => x"5f",
          5802 => x"34",
          5803 => x"38",
          5804 => x"76",
          5805 => x"38",
          5806 => x"b8",
          5807 => x"95",
          5808 => x"2b",
          5809 => x"56",
          5810 => x"94",
          5811 => x"2b",
          5812 => x"5a",
          5813 => x"ce",
          5814 => x"b8",
          5815 => x"ff",
          5816 => x"53",
          5817 => x"52",
          5818 => x"84",
          5819 => x"b8",
          5820 => x"08",
          5821 => x"08",
          5822 => x"fc",
          5823 => x"82",
          5824 => x"81",
          5825 => x"05",
          5826 => x"ff",
          5827 => x"39",
          5828 => x"5c",
          5829 => x"d0",
          5830 => x"d4",
          5831 => x"59",
          5832 => x"06",
          5833 => x"e5",
          5834 => x"79",
          5835 => x"77",
          5836 => x"3d",
          5837 => x"33",
          5838 => x"78",
          5839 => x"59",
          5840 => x"0c",
          5841 => x"0d",
          5842 => x"80",
          5843 => x"80",
          5844 => x"80",
          5845 => x"16",
          5846 => x"a0",
          5847 => x"75",
          5848 => x"72",
          5849 => x"76",
          5850 => x"08",
          5851 => x"cc",
          5852 => x"2b",
          5853 => x"f7",
          5854 => x"bb",
          5855 => x"15",
          5856 => x"bb",
          5857 => x"26",
          5858 => x"70",
          5859 => x"17",
          5860 => x"82",
          5861 => x"38",
          5862 => x"94",
          5863 => x"2a",
          5864 => x"2e",
          5865 => x"ff",
          5866 => x"54",
          5867 => x"a3",
          5868 => x"74",
          5869 => x"9c",
          5870 => x"98",
          5871 => x"91",
          5872 => x"e4",
          5873 => x"33",
          5874 => x"73",
          5875 => x"55",
          5876 => x"81",
          5877 => x"0c",
          5878 => x"90",
          5879 => x"33",
          5880 => x"34",
          5881 => x"2e",
          5882 => x"85",
          5883 => x"84",
          5884 => x"80",
          5885 => x"54",
          5886 => x"98",
          5887 => x"38",
          5888 => x"57",
          5889 => x"76",
          5890 => x"a9",
          5891 => x"fe",
          5892 => x"80",
          5893 => x"29",
          5894 => x"11",
          5895 => x"df",
          5896 => x"39",
          5897 => x"3f",
          5898 => x"39",
          5899 => x"3f",
          5900 => x"72",
          5901 => x"56",
          5902 => x"ff",
          5903 => x"54",
          5904 => x"38",
          5905 => x"ed",
          5906 => x"0c",
          5907 => x"82",
          5908 => x"b8",
          5909 => x"3d",
          5910 => x"2e",
          5911 => x"05",
          5912 => x"9b",
          5913 => x"b8",
          5914 => x"76",
          5915 => x"0c",
          5916 => x"7d",
          5917 => x"84",
          5918 => x"08",
          5919 => x"98",
          5920 => x"38",
          5921 => x"06",
          5922 => x"38",
          5923 => x"12",
          5924 => x"33",
          5925 => x"2e",
          5926 => x"58",
          5927 => x"52",
          5928 => x"b8",
          5929 => x"38",
          5930 => x"76",
          5931 => x"76",
          5932 => x"94",
          5933 => x"2b",
          5934 => x"5a",
          5935 => x"55",
          5936 => x"74",
          5937 => x"72",
          5938 => x"86",
          5939 => x"71",
          5940 => x"57",
          5941 => x"84",
          5942 => x"81",
          5943 => x"84",
          5944 => x"dc",
          5945 => x"39",
          5946 => x"89",
          5947 => x"08",
          5948 => x"33",
          5949 => x"14",
          5950 => x"78",
          5951 => x"59",
          5952 => x"80",
          5953 => x"51",
          5954 => x"08",
          5955 => x"b5",
          5956 => x"76",
          5957 => x"72",
          5958 => x"84",
          5959 => x"70",
          5960 => x"08",
          5961 => x"e4",
          5962 => x"53",
          5963 => x"72",
          5964 => x"84",
          5965 => x"70",
          5966 => x"08",
          5967 => x"52",
          5968 => x"b8",
          5969 => x"3d",
          5970 => x"fd",
          5971 => x"06",
          5972 => x"08",
          5973 => x"0d",
          5974 => x"53",
          5975 => x"84",
          5976 => x"08",
          5977 => x"e4",
          5978 => x"75",
          5979 => x"e4",
          5980 => x"38",
          5981 => x"2b",
          5982 => x"76",
          5983 => x"51",
          5984 => x"e4",
          5985 => x"84",
          5986 => x"ed",
          5987 => x"53",
          5988 => x"51",
          5989 => x"5a",
          5990 => x"75",
          5991 => x"11",
          5992 => x"75",
          5993 => x"79",
          5994 => x"04",
          5995 => x"5b",
          5996 => x"a8",
          5997 => x"5d",
          5998 => x"1d",
          5999 => x"76",
          6000 => x"78",
          6001 => x"54",
          6002 => x"33",
          6003 => x"e4",
          6004 => x"81",
          6005 => x"5b",
          6006 => x"5e",
          6007 => x"17",
          6008 => x"33",
          6009 => x"81",
          6010 => x"75",
          6011 => x"06",
          6012 => x"05",
          6013 => x"ff",
          6014 => x"53",
          6015 => x"38",
          6016 => x"84",
          6017 => x"18",
          6018 => x"3d",
          6019 => x"53",
          6020 => x"52",
          6021 => x"84",
          6022 => x"b8",
          6023 => x"08",
          6024 => x"08",
          6025 => x"fe",
          6026 => x"82",
          6027 => x"81",
          6028 => x"05",
          6029 => x"fe",
          6030 => x"39",
          6031 => x"75",
          6032 => x"84",
          6033 => x"38",
          6034 => x"f7",
          6035 => x"84",
          6036 => x"05",
          6037 => x"9c",
          6038 => x"7f",
          6039 => x"33",
          6040 => x"fe",
          6041 => x"11",
          6042 => x"70",
          6043 => x"83",
          6044 => x"59",
          6045 => x"fe",
          6046 => x"81",
          6047 => x"94",
          6048 => x"58",
          6049 => x"82",
          6050 => x"0d",
          6051 => x"9f",
          6052 => x"97",
          6053 => x"8f",
          6054 => x"59",
          6055 => x"80",
          6056 => x"91",
          6057 => x"90",
          6058 => x"55",
          6059 => x"c4",
          6060 => x"18",
          6061 => x"38",
          6062 => x"81",
          6063 => x"74",
          6064 => x"88",
          6065 => x"0c",
          6066 => x"18",
          6067 => x"91",
          6068 => x"e4",
          6069 => x"78",
          6070 => x"76",
          6071 => x"e4",
          6072 => x"2e",
          6073 => x"81",
          6074 => x"08",
          6075 => x"73",
          6076 => x"84",
          6077 => x"16",
          6078 => x"55",
          6079 => x"81",
          6080 => x"81",
          6081 => x"54",
          6082 => x"39",
          6083 => x"3f",
          6084 => x"73",
          6085 => x"56",
          6086 => x"33",
          6087 => x"18",
          6088 => x"52",
          6089 => x"b8",
          6090 => x"84",
          6091 => x"38",
          6092 => x"b8",
          6093 => x"a1",
          6094 => x"08",
          6095 => x"84",
          6096 => x"84",
          6097 => x"81",
          6098 => x"ff",
          6099 => x"c7",
          6100 => x"b8",
          6101 => x"76",
          6102 => x"e4",
          6103 => x"2e",
          6104 => x"81",
          6105 => x"08",
          6106 => x"73",
          6107 => x"84",
          6108 => x"16",
          6109 => x"55",
          6110 => x"15",
          6111 => x"07",
          6112 => x"77",
          6113 => x"74",
          6114 => x"39",
          6115 => x"90",
          6116 => x"82",
          6117 => x"33",
          6118 => x"e4",
          6119 => x"fa",
          6120 => x"54",
          6121 => x"56",
          6122 => x"db",
          6123 => x"9c",
          6124 => x"fb",
          6125 => x"b8",
          6126 => x"84",
          6127 => x"7d",
          6128 => x"70",
          6129 => x"b8",
          6130 => x"de",
          6131 => x"85",
          6132 => x"77",
          6133 => x"7b",
          6134 => x"33",
          6135 => x"7b",
          6136 => x"9b",
          6137 => x"2b",
          6138 => x"58",
          6139 => x"84",
          6140 => x"80",
          6141 => x"7b",
          6142 => x"41",
          6143 => x"70",
          6144 => x"b8",
          6145 => x"fe",
          6146 => x"74",
          6147 => x"e4",
          6148 => x"38",
          6149 => x"3d",
          6150 => x"33",
          6151 => x"7d",
          6152 => x"84",
          6153 => x"84",
          6154 => x"08",
          6155 => x"74",
          6156 => x"78",
          6157 => x"e4",
          6158 => x"2e",
          6159 => x"80",
          6160 => x"38",
          6161 => x"08",
          6162 => x"9c",
          6163 => x"82",
          6164 => x"fe",
          6165 => x"84",
          6166 => x"b8",
          6167 => x"5a",
          6168 => x"38",
          6169 => x"7a",
          6170 => x"81",
          6171 => x"17",
          6172 => x"b8",
          6173 => x"56",
          6174 => x"56",
          6175 => x"e5",
          6176 => x"90",
          6177 => x"80",
          6178 => x"84",
          6179 => x"08",
          6180 => x"2e",
          6181 => x"56",
          6182 => x"08",
          6183 => x"fe",
          6184 => x"e4",
          6185 => x"a6",
          6186 => x"34",
          6187 => x"84",
          6188 => x"18",
          6189 => x"33",
          6190 => x"fe",
          6191 => x"a0",
          6192 => x"17",
          6193 => x"58",
          6194 => x"27",
          6195 => x"fe",
          6196 => x"5a",
          6197 => x"cb",
          6198 => x"fd",
          6199 => x"2e",
          6200 => x"76",
          6201 => x"e4",
          6202 => x"11",
          6203 => x"7b",
          6204 => x"18",
          6205 => x"7b",
          6206 => x"26",
          6207 => x"39",
          6208 => x"e4",
          6209 => x"fd",
          6210 => x"9f",
          6211 => x"51",
          6212 => x"08",
          6213 => x"8a",
          6214 => x"3d",
          6215 => x"3d",
          6216 => x"84",
          6217 => x"08",
          6218 => x"0c",
          6219 => x"08",
          6220 => x"02",
          6221 => x"81",
          6222 => x"b9",
          6223 => x"70",
          6224 => x"b8",
          6225 => x"e4",
          6226 => x"e4",
          6227 => x"b8",
          6228 => x"75",
          6229 => x"08",
          6230 => x"80",
          6231 => x"fe",
          6232 => x"27",
          6233 => x"29",
          6234 => x"b4",
          6235 => x"79",
          6236 => x"58",
          6237 => x"74",
          6238 => x"27",
          6239 => x"53",
          6240 => x"ee",
          6241 => x"df",
          6242 => x"56",
          6243 => x"08",
          6244 => x"33",
          6245 => x"56",
          6246 => x"b8",
          6247 => x"08",
          6248 => x"18",
          6249 => x"33",
          6250 => x"fe",
          6251 => x"a0",
          6252 => x"17",
          6253 => x"ca",
          6254 => x"55",
          6255 => x"9c",
          6256 => x"52",
          6257 => x"b8",
          6258 => x"80",
          6259 => x"08",
          6260 => x"e4",
          6261 => x"53",
          6262 => x"3f",
          6263 => x"9c",
          6264 => x"5a",
          6265 => x"81",
          6266 => x"81",
          6267 => x"55",
          6268 => x"84",
          6269 => x"8a",
          6270 => x"06",
          6271 => x"81",
          6272 => x"1f",
          6273 => x"57",
          6274 => x"7d",
          6275 => x"58",
          6276 => x"59",
          6277 => x"cf",
          6278 => x"34",
          6279 => x"7d",
          6280 => x"77",
          6281 => x"5b",
          6282 => x"55",
          6283 => x"59",
          6284 => x"57",
          6285 => x"33",
          6286 => x"16",
          6287 => x"0b",
          6288 => x"83",
          6289 => x"80",
          6290 => x"7a",
          6291 => x"74",
          6292 => x"81",
          6293 => x"92",
          6294 => x"84",
          6295 => x"56",
          6296 => x"84",
          6297 => x"0b",
          6298 => x"17",
          6299 => x"18",
          6300 => x"18",
          6301 => x"80",
          6302 => x"16",
          6303 => x"34",
          6304 => x"b8",
          6305 => x"0c",
          6306 => x"55",
          6307 => x"2a",
          6308 => x"fd",
          6309 => x"cc",
          6310 => x"80",
          6311 => x"80",
          6312 => x"fe",
          6313 => x"94",
          6314 => x"95",
          6315 => x"16",
          6316 => x"34",
          6317 => x"b8",
          6318 => x"3d",
          6319 => x"59",
          6320 => x"79",
          6321 => x"26",
          6322 => x"38",
          6323 => x"af",
          6324 => x"05",
          6325 => x"3f",
          6326 => x"e4",
          6327 => x"b8",
          6328 => x"a6",
          6329 => x"3d",
          6330 => x"84",
          6331 => x"08",
          6332 => x"81",
          6333 => x"38",
          6334 => x"58",
          6335 => x"33",
          6336 => x"15",
          6337 => x"b0",
          6338 => x"81",
          6339 => x"59",
          6340 => x"b3",
          6341 => x"d5",
          6342 => x"b8",
          6343 => x"3d",
          6344 => x"84",
          6345 => x"76",
          6346 => x"57",
          6347 => x"82",
          6348 => x"5d",
          6349 => x"80",
          6350 => x"72",
          6351 => x"81",
          6352 => x"5b",
          6353 => x"77",
          6354 => x"81",
          6355 => x"58",
          6356 => x"70",
          6357 => x"70",
          6358 => x"09",
          6359 => x"38",
          6360 => x"07",
          6361 => x"7a",
          6362 => x"1e",
          6363 => x"38",
          6364 => x"39",
          6365 => x"7f",
          6366 => x"05",
          6367 => x"3f",
          6368 => x"e4",
          6369 => x"6c",
          6370 => x"fe",
          6371 => x"3f",
          6372 => x"e4",
          6373 => x"0b",
          6374 => x"05",
          6375 => x"57",
          6376 => x"ff",
          6377 => x"cb",
          6378 => x"33",
          6379 => x"7e",
          6380 => x"8b",
          6381 => x"1e",
          6382 => x"81",
          6383 => x"c5",
          6384 => x"bd",
          6385 => x"33",
          6386 => x"58",
          6387 => x"38",
          6388 => x"5e",
          6389 => x"8a",
          6390 => x"08",
          6391 => x"b5",
          6392 => x"08",
          6393 => x"5f",
          6394 => x"53",
          6395 => x"fe",
          6396 => x"80",
          6397 => x"77",
          6398 => x"d8",
          6399 => x"81",
          6400 => x"81",
          6401 => x"ff",
          6402 => x"34",
          6403 => x"18",
          6404 => x"09",
          6405 => x"5e",
          6406 => x"2a",
          6407 => x"57",
          6408 => x"aa",
          6409 => x"56",
          6410 => x"78",
          6411 => x"e4",
          6412 => x"f5",
          6413 => x"57",
          6414 => x"b4",
          6415 => x"7e",
          6416 => x"38",
          6417 => x"81",
          6418 => x"84",
          6419 => x"ff",
          6420 => x"77",
          6421 => x"5a",
          6422 => x"34",
          6423 => x"80",
          6424 => x"84",
          6425 => x"08",
          6426 => x"74",
          6427 => x"74",
          6428 => x"9d",
          6429 => x"e4",
          6430 => x"84",
          6431 => x"95",
          6432 => x"2b",
          6433 => x"56",
          6434 => x"08",
          6435 => x"e4",
          6436 => x"84",
          6437 => x"81",
          6438 => x"81",
          6439 => x"81",
          6440 => x"09",
          6441 => x"e4",
          6442 => x"a8",
          6443 => x"59",
          6444 => x"a0",
          6445 => x"2e",
          6446 => x"54",
          6447 => x"53",
          6448 => x"e1",
          6449 => x"81",
          6450 => x"70",
          6451 => x"e1",
          6452 => x"08",
          6453 => x"83",
          6454 => x"08",
          6455 => x"74",
          6456 => x"82",
          6457 => x"81",
          6458 => x"17",
          6459 => x"52",
          6460 => x"3f",
          6461 => x"0d",
          6462 => x"05",
          6463 => x"53",
          6464 => x"51",
          6465 => x"08",
          6466 => x"8a",
          6467 => x"3d",
          6468 => x"3d",
          6469 => x"84",
          6470 => x"08",
          6471 => x"81",
          6472 => x"38",
          6473 => x"12",
          6474 => x"51",
          6475 => x"78",
          6476 => x"51",
          6477 => x"08",
          6478 => x"04",
          6479 => x"96",
          6480 => x"ff",
          6481 => x"55",
          6482 => x"38",
          6483 => x"0d",
          6484 => x"d0",
          6485 => x"b8",
          6486 => x"e0",
          6487 => x"a0",
          6488 => x"60",
          6489 => x"90",
          6490 => x"17",
          6491 => x"17",
          6492 => x"17",
          6493 => x"17",
          6494 => x"34",
          6495 => x"b8",
          6496 => x"3d",
          6497 => x"5d",
          6498 => x"52",
          6499 => x"84",
          6500 => x"30",
          6501 => x"25",
          6502 => x"38",
          6503 => x"81",
          6504 => x"80",
          6505 => x"8c",
          6506 => x"78",
          6507 => x"11",
          6508 => x"08",
          6509 => x"33",
          6510 => x"81",
          6511 => x"53",
          6512 => x"fe",
          6513 => x"80",
          6514 => x"76",
          6515 => x"38",
          6516 => x"56",
          6517 => x"56",
          6518 => x"75",
          6519 => x"12",
          6520 => x"07",
          6521 => x"2b",
          6522 => x"5d",
          6523 => x"e4",
          6524 => x"80",
          6525 => x"55",
          6526 => x"08",
          6527 => x"81",
          6528 => x"06",
          6529 => x"57",
          6530 => x"08",
          6531 => x"33",
          6532 => x"59",
          6533 => x"81",
          6534 => x"08",
          6535 => x"17",
          6536 => x"55",
          6537 => x"38",
          6538 => x"09",
          6539 => x"b4",
          6540 => x"7a",
          6541 => x"e2",
          6542 => x"b8",
          6543 => x"da",
          6544 => x"2e",
          6545 => x"52",
          6546 => x"b8",
          6547 => x"fe",
          6548 => x"b8",
          6549 => x"18",
          6550 => x"75",
          6551 => x"78",
          6552 => x"58",
          6553 => x"f2",
          6554 => x"5c",
          6555 => x"fc",
          6556 => x"e1",
          6557 => x"b4",
          6558 => x"eb",
          6559 => x"b8",
          6560 => x"5d",
          6561 => x"81",
          6562 => x"f4",
          6563 => x"70",
          6564 => x"9f",
          6565 => x"90",
          6566 => x"81",
          6567 => x"75",
          6568 => x"81",
          6569 => x"83",
          6570 => x"9f",
          6571 => x"ff",
          6572 => x"e0",
          6573 => x"f4",
          6574 => x"58",
          6575 => x"56",
          6576 => x"70",
          6577 => x"58",
          6578 => x"2e",
          6579 => x"ff",
          6580 => x"ff",
          6581 => x"26",
          6582 => x"8f",
          6583 => x"70",
          6584 => x"76",
          6585 => x"1a",
          6586 => x"ff",
          6587 => x"26",
          6588 => x"86",
          6589 => x"79",
          6590 => x"56",
          6591 => x"a0",
          6592 => x"1a",
          6593 => x"47",
          6594 => x"fe",
          6595 => x"55",
          6596 => x"38",
          6597 => x"a1",
          6598 => x"51",
          6599 => x"83",
          6600 => x"38",
          6601 => x"a1",
          6602 => x"56",
          6603 => x"fe",
          6604 => x"55",
          6605 => x"79",
          6606 => x"7e",
          6607 => x"58",
          6608 => x"ff",
          6609 => x"81",
          6610 => x"d9",
          6611 => x"74",
          6612 => x"fe",
          6613 => x"84",
          6614 => x"06",
          6615 => x"2e",
          6616 => x"76",
          6617 => x"b8",
          6618 => x"75",
          6619 => x"84",
          6620 => x"98",
          6621 => x"08",
          6622 => x"55",
          6623 => x"d7",
          6624 => x"52",
          6625 => x"3f",
          6626 => x"38",
          6627 => x"0c",
          6628 => x"17",
          6629 => x"81",
          6630 => x"70",
          6631 => x"80",
          6632 => x"79",
          6633 => x"51",
          6634 => x"08",
          6635 => x"ff",
          6636 => x"fd",
          6637 => x"38",
          6638 => x"81",
          6639 => x"f4",
          6640 => x"34",
          6641 => x"70",
          6642 => x"05",
          6643 => x"2e",
          6644 => x"58",
          6645 => x"ff",
          6646 => x"39",
          6647 => x"81",
          6648 => x"d7",
          6649 => x"fd",
          6650 => x"81",
          6651 => x"81",
          6652 => x"84",
          6653 => x"06",
          6654 => x"83",
          6655 => x"08",
          6656 => x"8a",
          6657 => x"2e",
          6658 => x"fd",
          6659 => x"51",
          6660 => x"08",
          6661 => x"fd",
          6662 => x"58",
          6663 => x"fe",
          6664 => x"a0",
          6665 => x"18",
          6666 => x"a9",
          6667 => x"88",
          6668 => x"57",
          6669 => x"76",
          6670 => x"74",
          6671 => x"86",
          6672 => x"78",
          6673 => x"73",
          6674 => x"33",
          6675 => x"2e",
          6676 => x"9c",
          6677 => x"81",
          6678 => x"8c",
          6679 => x"2b",
          6680 => x"fd",
          6681 => x"70",
          6682 => x"b8",
          6683 => x"42",
          6684 => x"88",
          6685 => x"38",
          6686 => x"59",
          6687 => x"3f",
          6688 => x"08",
          6689 => x"b8",
          6690 => x"84",
          6691 => x"38",
          6692 => x"81",
          6693 => x"74",
          6694 => x"87",
          6695 => x"0c",
          6696 => x"b8",
          6697 => x"15",
          6698 => x"b8",
          6699 => x"ad",
          6700 => x"a7",
          6701 => x"7a",
          6702 => x"38",
          6703 => x"e6",
          6704 => x"fe",
          6705 => x"56",
          6706 => x"77",
          6707 => x"74",
          6708 => x"55",
          6709 => x"88",
          6710 => x"17",
          6711 => x"18",
          6712 => x"16",
          6713 => x"e9",
          6714 => x"84",
          6715 => x"16",
          6716 => x"54",
          6717 => x"fe",
          6718 => x"81",
          6719 => x"ff",
          6720 => x"3d",
          6721 => x"02",
          6722 => x"42",
          6723 => x"5f",
          6724 => x"38",
          6725 => x"9f",
          6726 => x"9b",
          6727 => x"85",
          6728 => x"80",
          6729 => x"10",
          6730 => x"5a",
          6731 => x"34",
          6732 => x"84",
          6733 => x"81",
          6734 => x"84",
          6735 => x"81",
          6736 => x"ab",
          6737 => x"8a",
          6738 => x"fc",
          6739 => x"d0",
          6740 => x"98",
          6741 => x"90",
          6742 => x"88",
          6743 => x"83",
          6744 => x"84",
          6745 => x"81",
          6746 => x"1f",
          6747 => x"7e",
          6748 => x"70",
          6749 => x"60",
          6750 => x"70",
          6751 => x"57",
          6752 => x"84",
          6753 => x"52",
          6754 => x"57",
          6755 => x"60",
          6756 => x"05",
          6757 => x"8e",
          6758 => x"81",
          6759 => x"61",
          6760 => x"62",
          6761 => x"18",
          6762 => x"90",
          6763 => x"33",
          6764 => x"71",
          6765 => x"82",
          6766 => x"2b",
          6767 => x"88",
          6768 => x"3d",
          6769 => x"0c",
          6770 => x"5a",
          6771 => x"79",
          6772 => x"81",
          6773 => x"2a",
          6774 => x"2e",
          6775 => x"64",
          6776 => x"47",
          6777 => x"30",
          6778 => x"2e",
          6779 => x"8c",
          6780 => x"22",
          6781 => x"74",
          6782 => x"56",
          6783 => x"57",
          6784 => x"75",
          6785 => x"fd",
          6786 => x"10",
          6787 => x"9f",
          6788 => x"b8",
          6789 => x"05",
          6790 => x"4c",
          6791 => x"81",
          6792 => x"68",
          6793 => x"06",
          6794 => x"83",
          6795 => x"77",
          6796 => x"57",
          6797 => x"7c",
          6798 => x"31",
          6799 => x"b8",
          6800 => x"f6",
          6801 => x"82",
          6802 => x"b8",
          6803 => x"89",
          6804 => x"c0",
          6805 => x"a3",
          6806 => x"0c",
          6807 => x"04",
          6808 => x"84",
          6809 => x"b8",
          6810 => x"70",
          6811 => x"89",
          6812 => x"ff",
          6813 => x"2e",
          6814 => x"d4",
          6815 => x"7a",
          6816 => x"81",
          6817 => x"59",
          6818 => x"17",
          6819 => x"9f",
          6820 => x"e0",
          6821 => x"76",
          6822 => x"78",
          6823 => x"ff",
          6824 => x"70",
          6825 => x"4a",
          6826 => x"81",
          6827 => x"25",
          6828 => x"39",
          6829 => x"79",
          6830 => x"84",
          6831 => x"83",
          6832 => x"40",
          6833 => x"55",
          6834 => x"38",
          6835 => x"81",
          6836 => x"ff",
          6837 => x"56",
          6838 => x"93",
          6839 => x"82",
          6840 => x"8b",
          6841 => x"26",
          6842 => x"5b",
          6843 => x"8e",
          6844 => x"3d",
          6845 => x"55",
          6846 => x"f5",
          6847 => x"5b",
          6848 => x"80",
          6849 => x"05",
          6850 => x"38",
          6851 => x"55",
          6852 => x"70",
          6853 => x"74",
          6854 => x"65",
          6855 => x"61",
          6856 => x"06",
          6857 => x"88",
          6858 => x"81",
          6859 => x"70",
          6860 => x"34",
          6861 => x"61",
          6862 => x"ff",
          6863 => x"ff",
          6864 => x"34",
          6865 => x"05",
          6866 => x"61",
          6867 => x"34",
          6868 => x"9b",
          6869 => x"7e",
          6870 => x"34",
          6871 => x"05",
          6872 => x"0c",
          6873 => x"34",
          6874 => x"61",
          6875 => x"34",
          6876 => x"61",
          6877 => x"06",
          6878 => x"88",
          6879 => x"ff",
          6880 => x"a6",
          6881 => x"e4",
          6882 => x"05",
          6883 => x"34",
          6884 => x"83",
          6885 => x"60",
          6886 => x"34",
          6887 => x"51",
          6888 => x"b8",
          6889 => x"5c",
          6890 => x"61",
          6891 => x"58",
          6892 => x"63",
          6893 => x"c0",
          6894 => x"81",
          6895 => x"34",
          6896 => x"64",
          6897 => x"2a",
          6898 => x"34",
          6899 => x"7c",
          6900 => x"38",
          6901 => x"52",
          6902 => x"b8",
          6903 => x"61",
          6904 => x"58",
          6905 => x"78",
          6906 => x"c9",
          6907 => x"2e",
          6908 => x"2e",
          6909 => x"66",
          6910 => x"7a",
          6911 => x"d2",
          6912 => x"38",
          6913 => x"75",
          6914 => x"93",
          6915 => x"26",
          6916 => x"83",
          6917 => x"61",
          6918 => x"b3",
          6919 => x"75",
          6920 => x"59",
          6921 => x"ff",
          6922 => x"47",
          6923 => x"34",
          6924 => x"83",
          6925 => x"6c",
          6926 => x"51",
          6927 => x"05",
          6928 => x"bf",
          6929 => x"84",
          6930 => x"7e",
          6931 => x"83",
          6932 => x"05",
          6933 => x"c9",
          6934 => x"34",
          6935 => x"cb",
          6936 => x"61",
          6937 => x"5f",
          6938 => x"54",
          6939 => x"c2",
          6940 => x"08",
          6941 => x"79",
          6942 => x"84",
          6943 => x"b8",
          6944 => x"3d",
          6945 => x"55",
          6946 => x"45",
          6947 => x"78",
          6948 => x"98",
          6949 => x"38",
          6950 => x"98",
          6951 => x"57",
          6952 => x"76",
          6953 => x"51",
          6954 => x"08",
          6955 => x"2a",
          6956 => x"b8",
          6957 => x"47",
          6958 => x"cb",
          6959 => x"b8",
          6960 => x"e6",
          6961 => x"2a",
          6962 => x"f8",
          6963 => x"80",
          6964 => x"ab",
          6965 => x"88",
          6966 => x"75",
          6967 => x"34",
          6968 => x"05",
          6969 => x"c3",
          6970 => x"34",
          6971 => x"cc",
          6972 => x"a4",
          6973 => x"61",
          6974 => x"78",
          6975 => x"56",
          6976 => x"ac",
          6977 => x"80",
          6978 => x"05",
          6979 => x"61",
          6980 => x"34",
          6981 => x"61",
          6982 => x"c2",
          6983 => x"83",
          6984 => x"81",
          6985 => x"58",
          6986 => x"f9",
          6987 => x"33",
          6988 => x"15",
          6989 => x"81",
          6990 => x"fe",
          6991 => x"e4",
          6992 => x"61",
          6993 => x"34",
          6994 => x"60",
          6995 => x"fc",
          6996 => x"0c",
          6997 => x"04",
          6998 => x"70",
          6999 => x"81",
          7000 => x"61",
          7001 => x"34",
          7002 => x"87",
          7003 => x"ff",
          7004 => x"05",
          7005 => x"b1",
          7006 => x"52",
          7007 => x"80",
          7008 => x"05",
          7009 => x"38",
          7010 => x"05",
          7011 => x"70",
          7012 => x"70",
          7013 => x"34",
          7014 => x"80",
          7015 => x"c1",
          7016 => x"61",
          7017 => x"5b",
          7018 => x"88",
          7019 => x"34",
          7020 => x"ea",
          7021 => x"61",
          7022 => x"ec",
          7023 => x"34",
          7024 => x"61",
          7025 => x"34",
          7026 => x"1f",
          7027 => x"b2",
          7028 => x"52",
          7029 => x"61",
          7030 => x"0d",
          7031 => x"ff",
          7032 => x"b8",
          7033 => x"05",
          7034 => x"ff",
          7035 => x"81",
          7036 => x"74",
          7037 => x"81",
          7038 => x"8a",
          7039 => x"38",
          7040 => x"38",
          7041 => x"8e",
          7042 => x"02",
          7043 => x"77",
          7044 => x"08",
          7045 => x"17",
          7046 => x"77",
          7047 => x"24",
          7048 => x"19",
          7049 => x"8b",
          7050 => x"17",
          7051 => x"3f",
          7052 => x"07",
          7053 => x"81",
          7054 => x"d3",
          7055 => x"3f",
          7056 => x"80",
          7057 => x"80",
          7058 => x"81",
          7059 => x"f4",
          7060 => x"8a",
          7061 => x"76",
          7062 => x"8c",
          7063 => x"16",
          7064 => x"84",
          7065 => x"7c",
          7066 => x"3d",
          7067 => x"05",
          7068 => x"3f",
          7069 => x"7a",
          7070 => x"e4",
          7071 => x"ff",
          7072 => x"52",
          7073 => x"74",
          7074 => x"9f",
          7075 => x"ff",
          7076 => x"eb",
          7077 => x"e4",
          7078 => x"0d",
          7079 => x"52",
          7080 => x"90",
          7081 => x"71",
          7082 => x"04",
          7083 => x"83",
          7084 => x"73",
          7085 => x"22",
          7086 => x"12",
          7087 => x"71",
          7088 => x"83",
          7089 => x"e1",
          7090 => x"06",
          7091 => x"0d",
          7092 => x"22",
          7093 => x"51",
          7094 => x"38",
          7095 => x"84",
          7096 => x"09",
          7097 => x"26",
          7098 => x"05",
          7099 => x"84",
          7100 => x"51",
          7101 => x"38",
          7102 => x"a8",
          7103 => x"d9",
          7104 => x"75",
          7105 => x"26",
          7106 => x"38",
          7107 => x"71",
          7108 => x"70",
          7109 => x"38",
          7110 => x"70",
          7111 => x"70",
          7112 => x"55",
          7113 => x"51",
          7114 => x"0d",
          7115 => x"39",
          7116 => x"10",
          7117 => x"04",
          7118 => x"06",
          7119 => x"b0",
          7120 => x"51",
          7121 => x"ff",
          7122 => x"70",
          7123 => x"39",
          7124 => x"57",
          7125 => x"ff",
          7126 => x"16",
          7127 => x"ff",
          7128 => x"76",
          7129 => x"58",
          7130 => x"31",
          7131 => x"fe",
          7132 => x"ff",
          7133 => x"00",
          7134 => x"19",
          7135 => x"19",
          7136 => x"19",
          7137 => x"19",
          7138 => x"19",
          7139 => x"19",
          7140 => x"19",
          7141 => x"18",
          7142 => x"18",
          7143 => x"18",
          7144 => x"1e",
          7145 => x"1f",
          7146 => x"1f",
          7147 => x"1f",
          7148 => x"1f",
          7149 => x"1f",
          7150 => x"1f",
          7151 => x"1f",
          7152 => x"1f",
          7153 => x"1f",
          7154 => x"1f",
          7155 => x"1f",
          7156 => x"1f",
          7157 => x"1f",
          7158 => x"1f",
          7159 => x"1f",
          7160 => x"1f",
          7161 => x"1f",
          7162 => x"1f",
          7163 => x"1f",
          7164 => x"1f",
          7165 => x"1f",
          7166 => x"1f",
          7167 => x"1f",
          7168 => x"1f",
          7169 => x"1f",
          7170 => x"1f",
          7171 => x"1f",
          7172 => x"1f",
          7173 => x"1f",
          7174 => x"24",
          7175 => x"1f",
          7176 => x"24",
          7177 => x"22",
          7178 => x"1f",
          7179 => x"1f",
          7180 => x"1f",
          7181 => x"1f",
          7182 => x"1f",
          7183 => x"1f",
          7184 => x"1f",
          7185 => x"1f",
          7186 => x"1f",
          7187 => x"1f",
          7188 => x"1f",
          7189 => x"1f",
          7190 => x"1f",
          7191 => x"1f",
          7192 => x"1f",
          7193 => x"1f",
          7194 => x"1f",
          7195 => x"1f",
          7196 => x"1f",
          7197 => x"1f",
          7198 => x"1f",
          7199 => x"1f",
          7200 => x"1f",
          7201 => x"1f",
          7202 => x"1f",
          7203 => x"1f",
          7204 => x"21",
          7205 => x"1f",
          7206 => x"1f",
          7207 => x"1f",
          7208 => x"1f",
          7209 => x"21",
          7210 => x"1f",
          7211 => x"1f",
          7212 => x"21",
          7213 => x"32",
          7214 => x"32",
          7215 => x"32",
          7216 => x"3b",
          7217 => x"38",
          7218 => x"3a",
          7219 => x"37",
          7220 => x"39",
          7221 => x"37",
          7222 => x"34",
          7223 => x"37",
          7224 => x"34",
          7225 => x"37",
          7226 => x"36",
          7227 => x"46",
          7228 => x"46",
          7229 => x"46",
          7230 => x"46",
          7231 => x"47",
          7232 => x"47",
          7233 => x"47",
          7234 => x"47",
          7235 => x"47",
          7236 => x"47",
          7237 => x"47",
          7238 => x"47",
          7239 => x"47",
          7240 => x"47",
          7241 => x"47",
          7242 => x"47",
          7243 => x"47",
          7244 => x"47",
          7245 => x"47",
          7246 => x"48",
          7247 => x"48",
          7248 => x"48",
          7249 => x"47",
          7250 => x"47",
          7251 => x"48",
          7252 => x"47",
          7253 => x"47",
          7254 => x"47",
          7255 => x"47",
          7256 => x"55",
          7257 => x"54",
          7258 => x"54",
          7259 => x"55",
          7260 => x"55",
          7261 => x"52",
          7262 => x"52",
          7263 => x"52",
          7264 => x"55",
          7265 => x"56",
          7266 => x"52",
          7267 => x"52",
          7268 => x"52",
          7269 => x"52",
          7270 => x"52",
          7271 => x"52",
          7272 => x"52",
          7273 => x"52",
          7274 => x"52",
          7275 => x"55",
          7276 => x"52",
          7277 => x"54",
          7278 => x"53",
          7279 => x"52",
          7280 => x"52",
          7281 => x"52",
          7282 => x"59",
          7283 => x"59",
          7284 => x"59",
          7285 => x"59",
          7286 => x"59",
          7287 => x"59",
          7288 => x"59",
          7289 => x"59",
          7290 => x"59",
          7291 => x"59",
          7292 => x"59",
          7293 => x"59",
          7294 => x"59",
          7295 => x"59",
          7296 => x"59",
          7297 => x"59",
          7298 => x"59",
          7299 => x"59",
          7300 => x"5a",
          7301 => x"59",
          7302 => x"5a",
          7303 => x"5a",
          7304 => x"59",
          7305 => x"59",
          7306 => x"59",
          7307 => x"63",
          7308 => x"61",
          7309 => x"61",
          7310 => x"61",
          7311 => x"61",
          7312 => x"61",
          7313 => x"61",
          7314 => x"5e",
          7315 => x"61",
          7316 => x"61",
          7317 => x"61",
          7318 => x"61",
          7319 => x"63",
          7320 => x"63",
          7321 => x"63",
          7322 => x"de",
          7323 => x"de",
          7324 => x"de",
          7325 => x"de",
          7326 => x"0e",
          7327 => x"0b",
          7328 => x"0b",
          7329 => x"0b",
          7330 => x"0b",
          7331 => x"0b",
          7332 => x"0b",
          7333 => x"0f",
          7334 => x"0b",
          7335 => x"0b",
          7336 => x"0b",
          7337 => x"0b",
          7338 => x"0b",
          7339 => x"0b",
          7340 => x"0b",
          7341 => x"0b",
          7342 => x"0b",
          7343 => x"0b",
          7344 => x"0b",
          7345 => x"0b",
          7346 => x"0b",
          7347 => x"0b",
          7348 => x"0b",
          7349 => x"0b",
          7350 => x"0b",
          7351 => x"0b",
          7352 => x"0b",
          7353 => x"0b",
          7354 => x"0e",
          7355 => x"0b",
          7356 => x"0b",
          7357 => x"0b",
          7358 => x"0b",
          7359 => x"0b",
          7360 => x"0e",
          7361 => x"0e",
          7362 => x"0b",
          7363 => x"0b",
          7364 => x"0e",
          7365 => x"0b",
          7366 => x"0e",
          7367 => x"0b",
          7368 => x"0b",
          7369 => x"0b",
          7370 => x"0e",
          7371 => x"00",
          7372 => x"00",
          7373 => x"00",
          7374 => x"00",
          7375 => x"00",
          7376 => x"00",
          7377 => x"00",
          7378 => x"00",
          7379 => x"00",
          7380 => x"68",
          7381 => x"64",
          7382 => x"64",
          7383 => x"6c",
          7384 => x"70",
          7385 => x"74",
          7386 => x"00",
          7387 => x"00",
          7388 => x"00",
          7389 => x"30",
          7390 => x"00",
          7391 => x"00",
          7392 => x"00",
          7393 => x"6b",
          7394 => x"72",
          7395 => x"72",
          7396 => x"20",
          7397 => x"63",
          7398 => x"6f",
          7399 => x"70",
          7400 => x"73",
          7401 => x"73",
          7402 => x"6e",
          7403 => x"79",
          7404 => x"6c",
          7405 => x"63",
          7406 => x"6d",
          7407 => x"70",
          7408 => x"20",
          7409 => x"65",
          7410 => x"72",
          7411 => x"72",
          7412 => x"20",
          7413 => x"62",
          7414 => x"73",
          7415 => x"6f",
          7416 => x"64",
          7417 => x"73",
          7418 => x"6e",
          7419 => x"00",
          7420 => x"6e",
          7421 => x"73",
          7422 => x"64",
          7423 => x"20",
          7424 => x"65",
          7425 => x"74",
          7426 => x"6c",
          7427 => x"65",
          7428 => x"64",
          7429 => x"6c",
          7430 => x"64",
          7431 => x"73",
          7432 => x"63",
          7433 => x"69",
          7434 => x"76",
          7435 => x"6c",
          7436 => x"00",
          7437 => x"68",
          7438 => x"00",
          7439 => x"65",
          7440 => x"00",
          7441 => x"6f",
          7442 => x"2e",
          7443 => x"61",
          7444 => x"2e",
          7445 => x"72",
          7446 => x"63",
          7447 => x"00",
          7448 => x"79",
          7449 => x"61",
          7450 => x"79",
          7451 => x"2e",
          7452 => x"61",
          7453 => x"38",
          7454 => x"20",
          7455 => x"00",
          7456 => x"00",
          7457 => x"34",
          7458 => x"20",
          7459 => x"00",
          7460 => x"20",
          7461 => x"2f",
          7462 => x"00",
          7463 => x"00",
          7464 => x"72",
          7465 => x"29",
          7466 => x"2a",
          7467 => x"55",
          7468 => x"75",
          7469 => x"6c",
          7470 => x"52",
          7471 => x"6e",
          7472 => x"00",
          7473 => x"52",
          7474 => x"72",
          7475 => x"52",
          7476 => x"6e",
          7477 => x"00",
          7478 => x"52",
          7479 => x"72",
          7480 => x"43",
          7481 => x"6e",
          7482 => x"00",
          7483 => x"52",
          7484 => x"72",
          7485 => x"32",
          7486 => x"75",
          7487 => x"6d",
          7488 => x"72",
          7489 => x"74",
          7490 => x"20",
          7491 => x"2e",
          7492 => x"6e",
          7493 => x"2e",
          7494 => x"74",
          7495 => x"61",
          7496 => x"53",
          7497 => x"74",
          7498 => x"20",
          7499 => x"69",
          7500 => x"64",
          7501 => x"2c",
          7502 => x"20",
          7503 => x"6e",
          7504 => x"00",
          7505 => x"3a",
          7506 => x"00",
          7507 => x"6d",
          7508 => x"00",
          7509 => x"6e",
          7510 => x"5c",
          7511 => x"00",
          7512 => x"65",
          7513 => x"2e",
          7514 => x"73",
          7515 => x"20",
          7516 => x"74",
          7517 => x"00",
          7518 => x"67",
          7519 => x"20",
          7520 => x"2e",
          7521 => x"6c",
          7522 => x"6e",
          7523 => x"20",
          7524 => x"00",
          7525 => x"69",
          7526 => x"20",
          7527 => x"20",
          7528 => x"38",
          7529 => x"58",
          7530 => x"38",
          7531 => x"2d",
          7532 => x"69",
          7533 => x"00",
          7534 => x"25",
          7535 => x"30",
          7536 => x"78",
          7537 => x"70",
          7538 => x"00",
          7539 => x"25",
          7540 => x"65",
          7541 => x"2e",
          7542 => x"6d",
          7543 => x"79",
          7544 => x"65",
          7545 => x"3a",
          7546 => x"00",
          7547 => x"20",
          7548 => x"65",
          7549 => x"6f",
          7550 => x"73",
          7551 => x"6e",
          7552 => x"3f",
          7553 => x"25",
          7554 => x"3a",
          7555 => x"0a",
          7556 => x"6e",
          7557 => x"69",
          7558 => x"44",
          7559 => x"69",
          7560 => x"74",
          7561 => x"64",
          7562 => x"00",
          7563 => x"55",
          7564 => x"56",
          7565 => x"64",
          7566 => x"20",
          7567 => x"00",
          7568 => x"55",
          7569 => x"20",
          7570 => x"64",
          7571 => x"20",
          7572 => x"00",
          7573 => x"61",
          7574 => x"74",
          7575 => x"73",
          7576 => x"20",
          7577 => x"00",
          7578 => x"00",
          7579 => x"55",
          7580 => x"20",
          7581 => x"20",
          7582 => x"20",
          7583 => x"00",
          7584 => x"73",
          7585 => x"63",
          7586 => x"20",
          7587 => x"20",
          7588 => x"4d",
          7589 => x"20",
          7590 => x"6e",
          7591 => x"20",
          7592 => x"72",
          7593 => x"25",
          7594 => x"00",
          7595 => x"52",
          7596 => x"6b",
          7597 => x"20",
          7598 => x"20",
          7599 => x"4d",
          7600 => x"20",
          7601 => x"20",
          7602 => x"20",
          7603 => x"00",
          7604 => x"20",
          7605 => x"20",
          7606 => x"4e",
          7607 => x"00",
          7608 => x"54",
          7609 => x"28",
          7610 => x"73",
          7611 => x"0a",
          7612 => x"4d",
          7613 => x"28",
          7614 => x"20",
          7615 => x"0a",
          7616 => x"20",
          7617 => x"28",
          7618 => x"20",
          7619 => x"0a",
          7620 => x"4d",
          7621 => x"28",
          7622 => x"38",
          7623 => x"20",
          7624 => x"20",
          7625 => x"58",
          7626 => x"0a",
          7627 => x"53",
          7628 => x"28",
          7629 => x"38",
          7630 => x"20",
          7631 => x"20",
          7632 => x"58",
          7633 => x"0a",
          7634 => x"20",
          7635 => x"28",
          7636 => x"38",
          7637 => x"66",
          7638 => x"20",
          7639 => x"00",
          7640 => x"6e",
          7641 => x"00",
          7642 => x"00",
          7643 => x"00",
          7644 => x"00",
          7645 => x"f0",
          7646 => x"00",
          7647 => x"00",
          7648 => x"f0",
          7649 => x"00",
          7650 => x"00",
          7651 => x"f0",
          7652 => x"00",
          7653 => x"00",
          7654 => x"f0",
          7655 => x"00",
          7656 => x"00",
          7657 => x"f0",
          7658 => x"00",
          7659 => x"00",
          7660 => x"f0",
          7661 => x"00",
          7662 => x"00",
          7663 => x"f0",
          7664 => x"00",
          7665 => x"00",
          7666 => x"f0",
          7667 => x"00",
          7668 => x"00",
          7669 => x"f0",
          7670 => x"00",
          7671 => x"00",
          7672 => x"f0",
          7673 => x"00",
          7674 => x"00",
          7675 => x"ef",
          7676 => x"00",
          7677 => x"00",
          7678 => x"44",
          7679 => x"42",
          7680 => x"36",
          7681 => x"34",
          7682 => x"33",
          7683 => x"31",
          7684 => x"00",
          7685 => x"00",
          7686 => x"00",
          7687 => x"00",
          7688 => x"00",
          7689 => x"6e",
          7690 => x"6e",
          7691 => x"20",
          7692 => x"20",
          7693 => x"69",
          7694 => x"2e",
          7695 => x"79",
          7696 => x"00",
          7697 => x"36",
          7698 => x"00",
          7699 => x"20",
          7700 => x"74",
          7701 => x"73",
          7702 => x"6c",
          7703 => x"46",
          7704 => x"73",
          7705 => x"31",
          7706 => x"41",
          7707 => x"43",
          7708 => x"31",
          7709 => x"31",
          7710 => x"31",
          7711 => x"31",
          7712 => x"31",
          7713 => x"31",
          7714 => x"31",
          7715 => x"31",
          7716 => x"31",
          7717 => x"32",
          7718 => x"32",
          7719 => x"33",
          7720 => x"46",
          7721 => x"00",
          7722 => x"00",
          7723 => x"64",
          7724 => x"25",
          7725 => x"32",
          7726 => x"25",
          7727 => x"3a",
          7728 => x"64",
          7729 => x"2c",
          7730 => x"00",
          7731 => x"00",
          7732 => x"25",
          7733 => x"70",
          7734 => x"73",
          7735 => x"3a",
          7736 => x"32",
          7737 => x"3a",
          7738 => x"32",
          7739 => x"3a",
          7740 => x"00",
          7741 => x"74",
          7742 => x"64",
          7743 => x"00",
          7744 => x"7c",
          7745 => x"3b",
          7746 => x"54",
          7747 => x"00",
          7748 => x"4f",
          7749 => x"20",
          7750 => x"20",
          7751 => x"20",
          7752 => x"45",
          7753 => x"33",
          7754 => x"f1",
          7755 => x"00",
          7756 => x"05",
          7757 => x"18",
          7758 => x"45",
          7759 => x"45",
          7760 => x"92",
          7761 => x"9a",
          7762 => x"4f",
          7763 => x"aa",
          7764 => x"b2",
          7765 => x"ba",
          7766 => x"c2",
          7767 => x"ca",
          7768 => x"d2",
          7769 => x"da",
          7770 => x"e2",
          7771 => x"ea",
          7772 => x"f2",
          7773 => x"fa",
          7774 => x"2c",
          7775 => x"2a",
          7776 => x"00",
          7777 => x"00",
          7778 => x"00",
          7779 => x"00",
          7780 => x"00",
          7781 => x"00",
          7782 => x"00",
          7783 => x"00",
          7784 => x"00",
          7785 => x"00",
          7786 => x"00",
          7787 => x"00",
          7788 => x"01",
          7789 => x"00",
          7790 => x"00",
          7791 => x"00",
          7792 => x"00",
          7793 => x"25",
          7794 => x"25",
          7795 => x"25",
          7796 => x"25",
          7797 => x"25",
          7798 => x"25",
          7799 => x"25",
          7800 => x"25",
          7801 => x"25",
          7802 => x"25",
          7803 => x"25",
          7804 => x"25",
          7805 => x"03",
          7806 => x"03",
          7807 => x"03",
          7808 => x"22",
          7809 => x"22",
          7810 => x"22",
          7811 => x"22",
          7812 => x"00",
          7813 => x"03",
          7814 => x"00",
          7815 => x"01",
          7816 => x"01",
          7817 => x"01",
          7818 => x"01",
          7819 => x"01",
          7820 => x"01",
          7821 => x"01",
          7822 => x"01",
          7823 => x"01",
          7824 => x"02",
          7825 => x"02",
          7826 => x"01",
          7827 => x"01",
          7828 => x"01",
          7829 => x"01",
          7830 => x"01",
          7831 => x"01",
          7832 => x"01",
          7833 => x"01",
          7834 => x"01",
          7835 => x"01",
          7836 => x"01",
          7837 => x"01",
          7838 => x"01",
          7839 => x"01",
          7840 => x"01",
          7841 => x"00",
          7842 => x"02",
          7843 => x"02",
          7844 => x"02",
          7845 => x"02",
          7846 => x"01",
          7847 => x"02",
          7848 => x"02",
          7849 => x"02",
          7850 => x"01",
          7851 => x"02",
          7852 => x"02",
          7853 => x"01",
          7854 => x"02",
          7855 => x"2c",
          7856 => x"02",
          7857 => x"02",
          7858 => x"02",
          7859 => x"02",
          7860 => x"02",
          7861 => x"03",
          7862 => x"00",
          7863 => x"03",
          7864 => x"00",
          7865 => x"03",
          7866 => x"03",
          7867 => x"03",
          7868 => x"03",
          7869 => x"03",
          7870 => x"04",
          7871 => x"04",
          7872 => x"04",
          7873 => x"04",
          7874 => x"04",
          7875 => x"00",
          7876 => x"1e",
          7877 => x"1f",
          7878 => x"1f",
          7879 => x"1f",
          7880 => x"1f",
          7881 => x"1f",
          7882 => x"00",
          7883 => x"1f",
          7884 => x"1f",
          7885 => x"1f",
          7886 => x"06",
          7887 => x"06",
          7888 => x"1f",
          7889 => x"00",
          7890 => x"1f",
          7891 => x"1f",
          7892 => x"21",
          7893 => x"02",
          7894 => x"24",
          7895 => x"2c",
          7896 => x"2c",
          7897 => x"2d",
          7898 => x"00",
          7899 => x"e6",
          7900 => x"00",
          7901 => x"e6",
          7902 => x"00",
          7903 => x"e6",
          7904 => x"00",
          7905 => x"e6",
          7906 => x"00",
          7907 => x"e6",
          7908 => x"00",
          7909 => x"e6",
          7910 => x"00",
          7911 => x"e6",
          7912 => x"00",
          7913 => x"e6",
          7914 => x"00",
          7915 => x"e6",
          7916 => x"00",
          7917 => x"e6",
          7918 => x"00",
          7919 => x"e6",
          7920 => x"00",
          7921 => x"e6",
          7922 => x"00",
          7923 => x"e6",
          7924 => x"00",
          7925 => x"e6",
          7926 => x"00",
          7927 => x"e6",
          7928 => x"00",
          7929 => x"e6",
          7930 => x"00",
          7931 => x"e6",
          7932 => x"00",
          7933 => x"e6",
          7934 => x"00",
          7935 => x"e6",
          7936 => x"00",
          7937 => x"e6",
          7938 => x"00",
          7939 => x"e6",
          7940 => x"00",
          7941 => x"e6",
          7942 => x"00",
          7943 => x"e6",
          7944 => x"00",
          7945 => x"e6",
          7946 => x"00",
          7947 => x"e6",
          7948 => x"00",
          7949 => x"e6",
          7950 => x"00",
          7951 => x"e7",
          7952 => x"00",
          7953 => x"e7",
          7954 => x"00",
          7955 => x"00",
          7956 => x"7f",
          7957 => x"7f",
          7958 => x"7f",
          7959 => x"00",
          7960 => x"ff",
          7961 => x"00",
          7962 => x"00",
          7963 => x"e1",
          7964 => x"00",
          7965 => x"01",
          7966 => x"00",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"5f",
          7983 => x"40",
          7984 => x"73",
          7985 => x"6b",
          7986 => x"63",
          7987 => x"33",
          7988 => x"2d",
          7989 => x"f3",
          7990 => x"f0",
          7991 => x"82",
          7992 => x"58",
          7993 => x"40",
          7994 => x"53",
          7995 => x"4b",
          7996 => x"43",
          7997 => x"33",
          7998 => x"2d",
          7999 => x"f3",
          8000 => x"f0",
          8001 => x"82",
          8002 => x"58",
          8003 => x"60",
          8004 => x"53",
          8005 => x"4b",
          8006 => x"43",
          8007 => x"23",
          8008 => x"3d",
          8009 => x"e0",
          8010 => x"f0",
          8011 => x"87",
          8012 => x"1e",
          8013 => x"00",
          8014 => x"13",
          8015 => x"0b",
          8016 => x"03",
          8017 => x"f0",
          8018 => x"f0",
          8019 => x"f0",
          8020 => x"f0",
          8021 => x"82",
          8022 => x"cf",
          8023 => x"d7",
          8024 => x"41",
          8025 => x"6c",
          8026 => x"d9",
          8027 => x"7e",
          8028 => x"d1",
          8029 => x"c2",
          8030 => x"f0",
          8031 => x"82",
          8032 => x"00",
          8033 => x"00",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"00",
          8045 => x"00",
          8046 => x"f0",
          8047 => x"f0",
          8048 => x"f0",
          8049 => x"f0",
          8050 => x"f0",
          8051 => x"f0",
          8052 => x"f0",
          8053 => x"f0",
          8054 => x"f0",
          8055 => x"f1",
          8056 => x"f1",
          8057 => x"f1",
          8058 => x"f1",
          8059 => x"f1",
          8060 => x"f1",
          8061 => x"f1",
          8062 => x"f1",
          8063 => x"f1",
          8064 => x"f1",
          8065 => x"f1",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"32",
          9067 => x"00",
          9068 => x"f6",
          9069 => x"fe",
          9070 => x"c6",
          9071 => x"ef",
          9072 => x"66",
          9073 => x"2e",
          9074 => x"26",
          9075 => x"57",
          9076 => x"06",
          9077 => x"0e",
          9078 => x"16",
          9079 => x"be",
          9080 => x"86",
          9081 => x"8e",
          9082 => x"96",
          9083 => x"a5",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"01",
          9100 => x"01",
        others => X"00"
    );

    shared variable RAM6 : ramArray :=
    (
             0 => x"0d",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"83",
             9 => x"2b",
            10 => x"00",
            11 => x"00",
            12 => x"ff",
            13 => x"82",
            14 => x"83",
            15 => x"a5",
            16 => x"05",
            17 => x"09",
            18 => x"51",
            19 => x"00",
            20 => x"2e",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"10",
            26 => x"0a",
            27 => x"00",
            28 => x"2e",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"04",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"53",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"81",
            45 => x"04",
            46 => x"00",
            47 => x"00",
            48 => x"9f",
            49 => x"06",
            50 => x"00",
            51 => x"00",
            52 => x"06",
            53 => x"05",
            54 => x"06",
            55 => x"00",
            56 => x"05",
            57 => x"81",
            58 => x"00",
            59 => x"00",
            60 => x"05",
            61 => x"09",
            62 => x"00",
            63 => x"00",
            64 => x"04",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"05",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"73",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"83",
            77 => x"10",
            78 => x"00",
            79 => x"00",
            80 => x"0b",
            81 => x"10",
            82 => x"b5",
            83 => x"00",
            84 => x"08",
            85 => x"2d",
            86 => x"8c",
            87 => x"00",
            88 => x"08",
            89 => x"2d",
            90 => x"8c",
            91 => x"00",
            92 => x"09",
            93 => x"54",
            94 => x"ff",
            95 => x"00",
            96 => x"09",
            97 => x"70",
            98 => x"05",
            99 => x"04",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"10",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"04",
           133 => x"0b",
           134 => x"8c",
           135 => x"04",
           136 => x"0b",
           137 => x"8c",
           138 => x"04",
           139 => x"0b",
           140 => x"8d",
           141 => x"04",
           142 => x"0b",
           143 => x"8d",
           144 => x"04",
           145 => x"0b",
           146 => x"8e",
           147 => x"04",
           148 => x"0b",
           149 => x"8e",
           150 => x"04",
           151 => x"0b",
           152 => x"8f",
           153 => x"04",
           154 => x"0b",
           155 => x"8f",
           156 => x"04",
           157 => x"0b",
           158 => x"90",
           159 => x"04",
           160 => x"0b",
           161 => x"91",
           162 => x"04",
           163 => x"0b",
           164 => x"91",
           165 => x"04",
           166 => x"0b",
           167 => x"92",
           168 => x"04",
           169 => x"0b",
           170 => x"92",
           171 => x"04",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"84",
           193 => x"84",
           194 => x"04",
           195 => x"84",
           196 => x"04",
           197 => x"84",
           198 => x"04",
           199 => x"84",
           200 => x"04",
           201 => x"84",
           202 => x"04",
           203 => x"84",
           204 => x"04",
           205 => x"84",
           206 => x"04",
           207 => x"84",
           208 => x"04",
           209 => x"84",
           210 => x"04",
           211 => x"84",
           212 => x"04",
           213 => x"84",
           214 => x"04",
           215 => x"84",
           216 => x"04",
           217 => x"2d",
           218 => x"90",
           219 => x"b6",
           220 => x"80",
           221 => x"d2",
           222 => x"c0",
           223 => x"80",
           224 => x"80",
           225 => x"0c",
           226 => x"08",
           227 => x"f0",
           228 => x"f0",
           229 => x"b8",
           230 => x"b8",
           231 => x"84",
           232 => x"84",
           233 => x"04",
           234 => x"2d",
           235 => x"90",
           236 => x"94",
           237 => x"80",
           238 => x"de",
           239 => x"c0",
           240 => x"82",
           241 => x"80",
           242 => x"0c",
           243 => x"08",
           244 => x"f0",
           245 => x"f0",
           246 => x"b8",
           247 => x"b8",
           248 => x"84",
           249 => x"84",
           250 => x"04",
           251 => x"2d",
           252 => x"90",
           253 => x"ac",
           254 => x"80",
           255 => x"93",
           256 => x"c0",
           257 => x"83",
           258 => x"80",
           259 => x"0c",
           260 => x"08",
           261 => x"f0",
           262 => x"f0",
           263 => x"b8",
           264 => x"b8",
           265 => x"84",
           266 => x"84",
           267 => x"04",
           268 => x"2d",
           269 => x"90",
           270 => x"e6",
           271 => x"80",
           272 => x"a0",
           273 => x"c0",
           274 => x"82",
           275 => x"80",
           276 => x"0c",
           277 => x"08",
           278 => x"f0",
           279 => x"f0",
           280 => x"b8",
           281 => x"b8",
           282 => x"84",
           283 => x"84",
           284 => x"04",
           285 => x"2d",
           286 => x"90",
           287 => x"d0",
           288 => x"80",
           289 => x"d0",
           290 => x"c0",
           291 => x"80",
           292 => x"80",
           293 => x"0c",
           294 => x"08",
           295 => x"f0",
           296 => x"08",
           297 => x"f0",
           298 => x"f0",
           299 => x"b8",
           300 => x"b8",
           301 => x"84",
           302 => x"84",
           303 => x"04",
           304 => x"2d",
           305 => x"90",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"73",
           311 => x"81",
           312 => x"07",
           313 => x"72",
           314 => x"09",
           315 => x"0a",
           316 => x"51",
           317 => x"84",
           318 => x"70",
           319 => x"93",
           320 => x"ba",
           321 => x"70",
           322 => x"74",
           323 => x"c5",
           324 => x"0d",
           325 => x"32",
           326 => x"58",
           327 => x"09",
           328 => x"77",
           329 => x"07",
           330 => x"80",
           331 => x"b2",
           332 => x"b8",
           333 => x"ff",
           334 => x"75",
           335 => x"73",
           336 => x"9f",
           337 => x"24",
           338 => x"71",
           339 => x"04",
           340 => x"3d",
           341 => x"86",
           342 => x"56",
           343 => x"53",
           344 => x"9d",
           345 => x"8d",
           346 => x"3d",
           347 => x"85",
           348 => x"0d",
           349 => x"70",
           350 => x"81",
           351 => x"5b",
           352 => x"06",
           353 => x"7b",
           354 => x"81",
           355 => x"81",
           356 => x"81",
           357 => x"70",
           358 => x"38",
           359 => x"2a",
           360 => x"7e",
           361 => x"07",
           362 => x"38",
           363 => x"e4",
           364 => x"2a",
           365 => x"05",
           366 => x"70",
           367 => x"70",
           368 => x"80",
           369 => x"06",
           370 => x"33",
           371 => x"b8",
           372 => x"93",
           373 => x"8a",
           374 => x"38",
           375 => x"8b",
           376 => x"cc",
           377 => x"70",
           378 => x"81",
           379 => x"38",
           380 => x"97",
           381 => x"05",
           382 => x"54",
           383 => x"7c",
           384 => x"7c",
           385 => x"fe",
           386 => x"39",
           387 => x"08",
           388 => x"41",
           389 => x"75",
           390 => x"08",
           391 => x"18",
           392 => x"88",
           393 => x"55",
           394 => x"79",
           395 => x"b8",
           396 => x"c5",
           397 => x"2b",
           398 => x"2e",
           399 => x"fc",
           400 => x"55",
           401 => x"5f",
           402 => x"80",
           403 => x"79",
           404 => x"80",
           405 => x"90",
           406 => x"06",
           407 => x"75",
           408 => x"54",
           409 => x"83",
           410 => x"86",
           411 => x"54",
           412 => x"79",
           413 => x"83",
           414 => x"2e",
           415 => x"06",
           416 => x"2a",
           417 => x"7a",
           418 => x"97",
           419 => x"8f",
           420 => x"7e",
           421 => x"80",
           422 => x"90",
           423 => x"9d",
           424 => x"3f",
           425 => x"80",
           426 => x"54",
           427 => x"06",
           428 => x"79",
           429 => x"05",
           430 => x"75",
           431 => x"87",
           432 => x"29",
           433 => x"5b",
           434 => x"7a",
           435 => x"7a",
           436 => x"e3",
           437 => x"2e",
           438 => x"81",
           439 => x"96",
           440 => x"52",
           441 => x"f4",
           442 => x"81",
           443 => x"38",
           444 => x"80",
           445 => x"55",
           446 => x"52",
           447 => x"7a",
           448 => x"33",
           449 => x"c8",
           450 => x"f8",
           451 => x"08",
           452 => x"42",
           453 => x"84",
           454 => x"13",
           455 => x"84",
           456 => x"70",
           457 => x"41",
           458 => x"5c",
           459 => x"84",
           460 => x"70",
           461 => x"25",
           462 => x"85",
           463 => x"83",
           464 => x"ff",
           465 => x"75",
           466 => x"d8",
           467 => x"ff",
           468 => x"ff",
           469 => x"70",
           470 => x"3f",
           471 => x"fc",
           472 => x"fc",
           473 => x"58",
           474 => x"81",
           475 => x"38",
           476 => x"71",
           477 => x"7e",
           478 => x"bf",
           479 => x"ad",
           480 => x"5b",
           481 => x"7a",
           482 => x"59",
           483 => x"7f",
           484 => x"06",
           485 => x"38",
           486 => x"e4",
           487 => x"31",
           488 => x"58",
           489 => x"7c",
           490 => x"f7",
           491 => x"08",
           492 => x"79",
           493 => x"3f",
           494 => x"06",
           495 => x"c4",
           496 => x"58",
           497 => x"39",
           498 => x"80",
           499 => x"54",
           500 => x"52",
           501 => x"7c",
           502 => x"90",
           503 => x"7c",
           504 => x"88",
           505 => x"fb",
           506 => x"2c",
           507 => x"2c",
           508 => x"53",
           509 => x"7c",
           510 => x"81",
           511 => x"38",
           512 => x"2a",
           513 => x"5b",
           514 => x"c8",
           515 => x"98",
           516 => x"52",
           517 => x"7c",
           518 => x"be",
           519 => x"3f",
           520 => x"06",
           521 => x"fd",
           522 => x"71",
           523 => x"fd",
           524 => x"c4",
           525 => x"b5",
           526 => x"0d",
           527 => x"08",
           528 => x"32",
           529 => x"57",
           530 => x"06",
           531 => x"56",
           532 => x"84",
           533 => x"14",
           534 => x"08",
           535 => x"70",
           536 => x"2e",
           537 => x"d7",
           538 => x"d4",
           539 => x"08",
           540 => x"80",
           541 => x"75",
           542 => x"04",
           543 => x"80",
           544 => x"81",
           545 => x"57",
           546 => x"06",
           547 => x"33",
           548 => x"98",
           549 => x"0c",
           550 => x"05",
           551 => x"38",
           552 => x"53",
           553 => x"2e",
           554 => x"56",
           555 => x"39",
           556 => x"52",
           557 => x"04",
           558 => x"33",
           559 => x"56",
           560 => x"38",
           561 => x"80",
           562 => x"72",
           563 => x"08",
           564 => x"05",
           565 => x"13",
           566 => x"b8",
           567 => x"52",
           568 => x"08",
           569 => x"e4",
           570 => x"05",
           571 => x"fb",
           572 => x"81",
           573 => x"55",
           574 => x"38",
           575 => x"b3",
           576 => x"71",
           577 => x"70",
           578 => x"f0",
           579 => x"08",
           580 => x"ff",
           581 => x"87",
           582 => x"53",
           583 => x"81",
           584 => x"84",
           585 => x"75",
           586 => x"84",
           587 => x"08",
           588 => x"33",
           589 => x"e4",
           590 => x"07",
           591 => x"73",
           592 => x"04",
           593 => x"34",
           594 => x"75",
           595 => x"81",
           596 => x"ff",
           597 => x"33",
           598 => x"34",
           599 => x"0c",
           600 => x"76",
           601 => x"70",
           602 => x"a1",
           603 => x"70",
           604 => x"05",
           605 => x"38",
           606 => x"0d",
           607 => x"d9",
           608 => x"13",
           609 => x"34",
           610 => x"38",
           611 => x"33",
           612 => x"38",
           613 => x"53",
           614 => x"51",
           615 => x"31",
           616 => x"0d",
           617 => x"54",
           618 => x"33",
           619 => x"34",
           620 => x"0c",
           621 => x"75",
           622 => x"70",
           623 => x"05",
           624 => x"34",
           625 => x"84",
           626 => x"fc",
           627 => x"54",
           628 => x"75",
           629 => x"71",
           630 => x"81",
           631 => x"ff",
           632 => x"70",
           633 => x"04",
           634 => x"53",
           635 => x"ff",
           636 => x"2e",
           637 => x"e4",
           638 => x"b8",
           639 => x"3d",
           640 => x"80",
           641 => x"b8",
           642 => x"b2",
           643 => x"84",
           644 => x"84",
           645 => x"34",
           646 => x"08",
           647 => x"08",
           648 => x"3d",
           649 => x"71",
           650 => x"2e",
           651 => x"33",
           652 => x"12",
           653 => x"ea",
           654 => x"52",
           655 => x"0d",
           656 => x"72",
           657 => x"8e",
           658 => x"34",
           659 => x"84",
           660 => x"fa",
           661 => x"52",
           662 => x"80",
           663 => x"e0",
           664 => x"73",
           665 => x"e4",
           666 => x"26",
           667 => x"2e",
           668 => x"2a",
           669 => x"54",
           670 => x"a8",
           671 => x"74",
           672 => x"11",
           673 => x"06",
           674 => x"52",
           675 => x"38",
           676 => x"b8",
           677 => x"3d",
           678 => x"70",
           679 => x"84",
           680 => x"70",
           681 => x"80",
           682 => x"71",
           683 => x"70",
           684 => x"74",
           685 => x"73",
           686 => x"10",
           687 => x"81",
           688 => x"30",
           689 => x"84",
           690 => x"51",
           691 => x"51",
           692 => x"54",
           693 => x"0d",
           694 => x"54",
           695 => x"73",
           696 => x"0c",
           697 => x"0d",
           698 => x"80",
           699 => x"3f",
           700 => x"52",
           701 => x"fe",
           702 => x"31",
           703 => x"c5",
           704 => x"38",
           705 => x"31",
           706 => x"80",
           707 => x"10",
           708 => x"07",
           709 => x"70",
           710 => x"31",
           711 => x"58",
           712 => x"b8",
           713 => x"3d",
           714 => x"7a",
           715 => x"7d",
           716 => x"57",
           717 => x"55",
           718 => x"08",
           719 => x"0c",
           720 => x"7b",
           721 => x"77",
           722 => x"a0",
           723 => x"15",
           724 => x"73",
           725 => x"80",
           726 => x"38",
           727 => x"26",
           728 => x"a0",
           729 => x"74",
           730 => x"ff",
           731 => x"ff",
           732 => x"38",
           733 => x"54",
           734 => x"78",
           735 => x"13",
           736 => x"56",
           737 => x"38",
           738 => x"56",
           739 => x"b8",
           740 => x"70",
           741 => x"56",
           742 => x"fe",
           743 => x"70",
           744 => x"a6",
           745 => x"a0",
           746 => x"38",
           747 => x"89",
           748 => x"b8",
           749 => x"58",
           750 => x"55",
           751 => x"0b",
           752 => x"04",
           753 => x"80",
           754 => x"56",
           755 => x"06",
           756 => x"70",
           757 => x"38",
           758 => x"b0",
           759 => x"80",
           760 => x"8a",
           761 => x"c4",
           762 => x"e0",
           763 => x"d0",
           764 => x"90",
           765 => x"81",
           766 => x"81",
           767 => x"38",
           768 => x"79",
           769 => x"a0",
           770 => x"84",
           771 => x"81",
           772 => x"3d",
           773 => x"0c",
           774 => x"2e",
           775 => x"15",
           776 => x"73",
           777 => x"73",
           778 => x"a0",
           779 => x"80",
           780 => x"e1",
           781 => x"3d",
           782 => x"78",
           783 => x"fe",
           784 => x"0c",
           785 => x"3f",
           786 => x"84",
           787 => x"73",
           788 => x"10",
           789 => x"08",
           790 => x"3f",
           791 => x"51",
           792 => x"83",
           793 => x"3d",
           794 => x"9d",
           795 => x"e4",
           796 => x"04",
           797 => x"83",
           798 => x"ee",
           799 => x"cf",
           800 => x"0d",
           801 => x"3f",
           802 => x"51",
           803 => x"83",
           804 => x"3d",
           805 => x"c5",
           806 => x"ac",
           807 => x"04",
           808 => x"83",
           809 => x"ee",
           810 => x"d0",
           811 => x"0d",
           812 => x"3f",
           813 => x"51",
           814 => x"83",
           815 => x"3d",
           816 => x"ed",
           817 => x"b4",
           818 => x"04",
           819 => x"80",
           820 => x"79",
           821 => x"57",
           822 => x"26",
           823 => x"70",
           824 => x"74",
           825 => x"8c",
           826 => x"3f",
           827 => x"e4",
           828 => x"51",
           829 => x"78",
           830 => x"2a",
           831 => x"80",
           832 => x"08",
           833 => x"38",
           834 => x"f5",
           835 => x"83",
           836 => x"c0",
           837 => x"e4",
           838 => x"e4",
           839 => x"b8",
           840 => x"54",
           841 => x"82",
           842 => x"57",
           843 => x"7a",
           844 => x"74",
           845 => x"87",
           846 => x"84",
           847 => x"a7",
           848 => x"d1",
           849 => x"51",
           850 => x"3d",
           851 => x"33",
           852 => x"52",
           853 => x"e4",
           854 => x"38",
           855 => x"b8",
           856 => x"04",
           857 => x"54",
           858 => x"51",
           859 => x"b8",
           860 => x"3d",
           861 => x"80",
           862 => x"41",
           863 => x"80",
           864 => x"d1",
           865 => x"f4",
           866 => x"79",
           867 => x"ed",
           868 => x"73",
           869 => x"38",
           870 => x"dd",
           871 => x"08",
           872 => x"78",
           873 => x"51",
           874 => x"27",
           875 => x"55",
           876 => x"38",
           877 => x"83",
           878 => x"81",
           879 => x"88",
           880 => x"38",
           881 => x"eb",
           882 => x"26",
           883 => x"d5",
           884 => x"80",
           885 => x"08",
           886 => x"76",
           887 => x"2e",
           888 => x"78",
           889 => x"b8",
           890 => x"d2",
           891 => x"84",
           892 => x"eb",
           893 => x"38",
           894 => x"dc",
           895 => x"08",
           896 => x"73",
           897 => x"53",
           898 => x"52",
           899 => x"82",
           900 => x"a0",
           901 => x"dd",
           902 => x"51",
           903 => x"c8",
           904 => x"3f",
           905 => x"18",
           906 => x"08",
           907 => x"3f",
           908 => x"54",
           909 => x"26",
           910 => x"c8",
           911 => x"81",
           912 => x"d8",
           913 => x"06",
           914 => x"ec",
           915 => x"09",
           916 => x"fc",
           917 => x"84",
           918 => x"2c",
           919 => x"32",
           920 => x"07",
           921 => x"53",
           922 => x"51",
           923 => x"98",
           924 => x"70",
           925 => x"72",
           926 => x"58",
           927 => x"ff",
           928 => x"84",
           929 => x"fe",
           930 => x"53",
           931 => x"3f",
           932 => x"80",
           933 => x"70",
           934 => x"38",
           935 => x"52",
           936 => x"70",
           937 => x"38",
           938 => x"52",
           939 => x"70",
           940 => x"38",
           941 => x"52",
           942 => x"70",
           943 => x"72",
           944 => x"38",
           945 => x"81",
           946 => x"51",
           947 => x"3f",
           948 => x"81",
           949 => x"51",
           950 => x"3f",
           951 => x"80",
           952 => x"9b",
           953 => x"d4",
           954 => x"87",
           955 => x"80",
           956 => x"51",
           957 => x"9b",
           958 => x"72",
           959 => x"71",
           960 => x"39",
           961 => x"c4",
           962 => x"f4",
           963 => x"51",
           964 => x"ff",
           965 => x"83",
           966 => x"51",
           967 => x"81",
           968 => x"94",
           969 => x"bc",
           970 => x"3f",
           971 => x"2a",
           972 => x"2e",
           973 => x"51",
           974 => x"9a",
           975 => x"72",
           976 => x"71",
           977 => x"39",
           978 => x"ff",
           979 => x"52",
           980 => x"b8",
           981 => x"40",
           982 => x"83",
           983 => x"3d",
           984 => x"3f",
           985 => x"7e",
           986 => x"ed",
           987 => x"59",
           988 => x"81",
           989 => x"06",
           990 => x"67",
           991 => x"dc",
           992 => x"09",
           993 => x"33",
           994 => x"80",
           995 => x"90",
           996 => x"52",
           997 => x"08",
           998 => x"7b",
           999 => x"b8",
          1000 => x"5e",
          1001 => x"1c",
          1002 => x"7c",
          1003 => x"7b",
          1004 => x"52",
          1005 => x"e4",
          1006 => x"2e",
          1007 => x"48",
          1008 => x"89",
          1009 => x"06",
          1010 => x"38",
          1011 => x"3f",
          1012 => x"f3",
          1013 => x"7a",
          1014 => x"24",
          1015 => x"e4",
          1016 => x"8c",
          1017 => x"f1",
          1018 => x"56",
          1019 => x"53",
          1020 => x"ae",
          1021 => x"e4",
          1022 => x"80",
          1023 => x"7a",
          1024 => x"7a",
          1025 => x"81",
          1026 => x"7a",
          1027 => x"81",
          1028 => x"61",
          1029 => x"81",
          1030 => x"d3",
          1031 => x"80",
          1032 => x"0b",
          1033 => x"06",
          1034 => x"53",
          1035 => x"51",
          1036 => x"08",
          1037 => x"83",
          1038 => x"80",
          1039 => x"3f",
          1040 => x"38",
          1041 => x"3f",
          1042 => x"81",
          1043 => x"09",
          1044 => x"84",
          1045 => x"82",
          1046 => x"83",
          1047 => x"51",
          1048 => x"79",
          1049 => x"63",
          1050 => x"89",
          1051 => x"83",
          1052 => x"83",
          1053 => x"e4",
          1054 => x"ba",
          1055 => x"b8",
          1056 => x"fb",
          1057 => x"41",
          1058 => x"51",
          1059 => x"e2",
          1060 => x"56",
          1061 => x"53",
          1062 => x"f2",
          1063 => x"3f",
          1064 => x"f9",
          1065 => x"3f",
          1066 => x"fa",
          1067 => x"95",
          1068 => x"d4",
          1069 => x"fa",
          1070 => x"53",
          1071 => x"84",
          1072 => x"38",
          1073 => x"fa",
          1074 => x"e4",
          1075 => x"b8",
          1076 => x"d0",
          1077 => x"ff",
          1078 => x"eb",
          1079 => x"2e",
          1080 => x"a8",
          1081 => x"04",
          1082 => x"80",
          1083 => x"e4",
          1084 => x"3d",
          1085 => x"51",
          1086 => x"86",
          1087 => x"78",
          1088 => x"3f",
          1089 => x"52",
          1090 => x"7e",
          1091 => x"38",
          1092 => x"84",
          1093 => x"3d",
          1094 => x"51",
          1095 => x"80",
          1096 => x"f0",
          1097 => x"b4",
          1098 => x"38",
          1099 => x"83",
          1100 => x"d4",
          1101 => x"51",
          1102 => x"59",
          1103 => x"9f",
          1104 => x"70",
          1105 => x"84",
          1106 => x"f0",
          1107 => x"f8",
          1108 => x"53",
          1109 => x"84",
          1110 => x"38",
          1111 => x"80",
          1112 => x"e4",
          1113 => x"d6",
          1114 => x"5d",
          1115 => x"65",
          1116 => x"7a",
          1117 => x"54",
          1118 => x"f0",
          1119 => x"5c",
          1120 => x"39",
          1121 => x"80",
          1122 => x"e4",
          1123 => x"3d",
          1124 => x"51",
          1125 => x"80",
          1126 => x"f8",
          1127 => x"c8",
          1128 => x"f6",
          1129 => x"ba",
          1130 => x"93",
          1131 => x"5b",
          1132 => x"eb",
          1133 => x"ff",
          1134 => x"b8",
          1135 => x"b8",
          1136 => x"05",
          1137 => x"08",
          1138 => x"83",
          1139 => x"d4",
          1140 => x"51",
          1141 => x"59",
          1142 => x"9f",
          1143 => x"49",
          1144 => x"05",
          1145 => x"b8",
          1146 => x"05",
          1147 => x"08",
          1148 => x"02",
          1149 => x"81",
          1150 => x"53",
          1151 => x"84",
          1152 => x"b9",
          1153 => x"ff",
          1154 => x"b8",
          1155 => x"b8",
          1156 => x"05",
          1157 => x"08",
          1158 => x"fe",
          1159 => x"e6",
          1160 => x"38",
          1161 => x"a4",
          1162 => x"59",
          1163 => x"7a",
          1164 => x"79",
          1165 => x"3f",
          1166 => x"05",
          1167 => x"08",
          1168 => x"88",
          1169 => x"08",
          1170 => x"b8",
          1171 => x"84",
          1172 => x"f4",
          1173 => x"53",
          1174 => x"84",
          1175 => x"e8",
          1176 => x"38",
          1177 => x"fe",
          1178 => x"e5",
          1179 => x"38",
          1180 => x"2e",
          1181 => x"47",
          1182 => x"80",
          1183 => x"e4",
          1184 => x"5c",
          1185 => x"5c",
          1186 => x"07",
          1187 => x"79",
          1188 => x"83",
          1189 => x"d6",
          1190 => x"53",
          1191 => x"83",
          1192 => x"f9",
          1193 => x"84",
          1194 => x"53",
          1195 => x"84",
          1196 => x"38",
          1197 => x"05",
          1198 => x"ff",
          1199 => x"b8",
          1200 => x"64",
          1201 => x"70",
          1202 => x"3d",
          1203 => x"51",
          1204 => x"80",
          1205 => x"80",
          1206 => x"40",
          1207 => x"11",
          1208 => x"3f",
          1209 => x"f1",
          1210 => x"53",
          1211 => x"84",
          1212 => x"38",
          1213 => x"7c",
          1214 => x"39",
          1215 => x"80",
          1216 => x"e4",
          1217 => x"64",
          1218 => x"46",
          1219 => x"09",
          1220 => x"83",
          1221 => x"cc",
          1222 => x"96",
          1223 => x"3f",
          1224 => x"d4",
          1225 => x"fe",
          1226 => x"e0",
          1227 => x"2e",
          1228 => x"05",
          1229 => x"78",
          1230 => x"33",
          1231 => x"83",
          1232 => x"83",
          1233 => x"a1",
          1234 => x"b5",
          1235 => x"3f",
          1236 => x"84",
          1237 => x"cc",
          1238 => x"80",
          1239 => x"49",
          1240 => x"d3",
          1241 => x"ea",
          1242 => x"83",
          1243 => x"83",
          1244 => x"9b",
          1245 => x"dd",
          1246 => x"80",
          1247 => x"47",
          1248 => x"5d",
          1249 => x"c0",
          1250 => x"e6",
          1251 => x"83",
          1252 => x"83",
          1253 => x"fb",
          1254 => x"05",
          1255 => x"80",
          1256 => x"94",
          1257 => x"80",
          1258 => x"b8",
          1259 => x"55",
          1260 => x"bf",
          1261 => x"77",
          1262 => x"56",
          1263 => x"da",
          1264 => x"2b",
          1265 => x"52",
          1266 => x"b8",
          1267 => x"83",
          1268 => x"80",
          1269 => x"81",
          1270 => x"83",
          1271 => x"5e",
          1272 => x"88",
          1273 => x"c8",
          1274 => x"3f",
          1275 => x"fc",
          1276 => x"a4",
          1277 => x"70",
          1278 => x"d2",
          1279 => x"15",
          1280 => x"82",
          1281 => x"80",
          1282 => x"56",
          1283 => x"2e",
          1284 => x"ff",
          1285 => x"81",
          1286 => x"70",
          1287 => x"a0",
          1288 => x"54",
          1289 => x"52",
          1290 => x"72",
          1291 => x"54",
          1292 => x"70",
          1293 => x"86",
          1294 => x"73",
          1295 => x"2e",
          1296 => x"70",
          1297 => x"76",
          1298 => x"88",
          1299 => x"34",
          1300 => x"b8",
          1301 => x"80",
          1302 => x"be",
          1303 => x"70",
          1304 => x"a2",
          1305 => x"81",
          1306 => x"81",
          1307 => x"dc",
          1308 => x"08",
          1309 => x"0c",
          1310 => x"05",
          1311 => x"b8",
          1312 => x"84",
          1313 => x"fc",
          1314 => x"05",
          1315 => x"81",
          1316 => x"54",
          1317 => x"38",
          1318 => x"97",
          1319 => x"54",
          1320 => x"38",
          1321 => x"bb",
          1322 => x"55",
          1323 => x"d9",
          1324 => x"73",
          1325 => x"0b",
          1326 => x"87",
          1327 => x"87",
          1328 => x"87",
          1329 => x"87",
          1330 => x"87",
          1331 => x"87",
          1332 => x"98",
          1333 => x"0c",
          1334 => x"80",
          1335 => x"3d",
          1336 => x"87",
          1337 => x"87",
          1338 => x"23",
          1339 => x"82",
          1340 => x"5a",
          1341 => x"b0",
          1342 => x"c0",
          1343 => x"34",
          1344 => x"86",
          1345 => x"5c",
          1346 => x"a0",
          1347 => x"7d",
          1348 => x"7b",
          1349 => x"33",
          1350 => x"33",
          1351 => x"33",
          1352 => x"83",
          1353 => x"8f",
          1354 => x"93",
          1355 => x"38",
          1356 => x"b8",
          1357 => x"51",
          1358 => x"86",
          1359 => x"84",
          1360 => x"72",
          1361 => x"e4",
          1362 => x"52",
          1363 => x"38",
          1364 => x"b8",
          1365 => x"51",
          1366 => x"39",
          1367 => x"71",
          1368 => x"cd",
          1369 => x"70",
          1370 => x"eb",
          1371 => x"52",
          1372 => x"b8",
          1373 => x"3d",
          1374 => x"9c",
          1375 => x"55",
          1376 => x"c0",
          1377 => x"81",
          1378 => x"8c",
          1379 => x"51",
          1380 => x"81",
          1381 => x"71",
          1382 => x"38",
          1383 => x"94",
          1384 => x"87",
          1385 => x"74",
          1386 => x"04",
          1387 => x"51",
          1388 => x"06",
          1389 => x"93",
          1390 => x"c0",
          1391 => x"96",
          1392 => x"70",
          1393 => x"02",
          1394 => x"2a",
          1395 => x"34",
          1396 => x"78",
          1397 => x"57",
          1398 => x"15",
          1399 => x"06",
          1400 => x"ff",
          1401 => x"96",
          1402 => x"70",
          1403 => x"70",
          1404 => x"72",
          1405 => x"2e",
          1406 => x"52",
          1407 => x"51",
          1408 => x"2e",
          1409 => x"73",
          1410 => x"57",
          1411 => x"e4",
          1412 => x"2a",
          1413 => x"38",
          1414 => x"80",
          1415 => x"06",
          1416 => x"87",
          1417 => x"70",
          1418 => x"38",
          1419 => x"9e",
          1420 => x"52",
          1421 => x"87",
          1422 => x"0c",
          1423 => x"a4",
          1424 => x"f1",
          1425 => x"83",
          1426 => x"08",
          1427 => x"a0",
          1428 => x"9e",
          1429 => x"c0",
          1430 => x"87",
          1431 => x"0c",
          1432 => x"c4",
          1433 => x"f1",
          1434 => x"83",
          1435 => x"08",
          1436 => x"80",
          1437 => x"87",
          1438 => x"0c",
          1439 => x"dc",
          1440 => x"f1",
          1441 => x"34",
          1442 => x"70",
          1443 => x"70",
          1444 => x"34",
          1445 => x"70",
          1446 => x"70",
          1447 => x"83",
          1448 => x"9e",
          1449 => x"51",
          1450 => x"81",
          1451 => x"0b",
          1452 => x"80",
          1453 => x"2e",
          1454 => x"e8",
          1455 => x"08",
          1456 => x"52",
          1457 => x"71",
          1458 => x"c0",
          1459 => x"06",
          1460 => x"38",
          1461 => x"80",
          1462 => x"84",
          1463 => x"80",
          1464 => x"f1",
          1465 => x"90",
          1466 => x"52",
          1467 => x"52",
          1468 => x"87",
          1469 => x"80",
          1470 => x"83",
          1471 => x"34",
          1472 => x"70",
          1473 => x"70",
          1474 => x"83",
          1475 => x"9e",
          1476 => x"52",
          1477 => x"52",
          1478 => x"9e",
          1479 => x"2a",
          1480 => x"80",
          1481 => x"84",
          1482 => x"2e",
          1483 => x"f1",
          1484 => x"f0",
          1485 => x"83",
          1486 => x"9e",
          1487 => x"52",
          1488 => x"71",
          1489 => x"90",
          1490 => x"f4",
          1491 => x"fd",
          1492 => x"a0",
          1493 => x"e4",
          1494 => x"d8",
          1495 => x"e6",
          1496 => x"f1",
          1497 => x"83",
          1498 => x"38",
          1499 => x"ff",
          1500 => x"84",
          1501 => x"75",
          1502 => x"54",
          1503 => x"33",
          1504 => x"e5",
          1505 => x"f1",
          1506 => x"83",
          1507 => x"38",
          1508 => x"f4",
          1509 => x"81",
          1510 => x"bd",
          1511 => x"d8",
          1512 => x"f1",
          1513 => x"ff",
          1514 => x"52",
          1515 => x"3f",
          1516 => x"83",
          1517 => x"51",
          1518 => x"08",
          1519 => x"ca",
          1520 => x"84",
          1521 => x"84",
          1522 => x"51",
          1523 => x"33",
          1524 => x"e6",
          1525 => x"c3",
          1526 => x"f1",
          1527 => x"75",
          1528 => x"08",
          1529 => x"54",
          1530 => x"da",
          1531 => x"51",
          1532 => x"83",
          1533 => x"52",
          1534 => x"e4",
          1535 => x"31",
          1536 => x"83",
          1537 => x"83",
          1538 => x"ff",
          1539 => x"84",
          1540 => x"51",
          1541 => x"52",
          1542 => x"3f",
          1543 => x"80",
          1544 => x"d0",
          1545 => x"b3",
          1546 => x"9d",
          1547 => x"d9",
          1548 => x"f1",
          1549 => x"75",
          1550 => x"08",
          1551 => x"54",
          1552 => x"da",
          1553 => x"f1",
          1554 => x"8d",
          1555 => x"51",
          1556 => x"33",
          1557 => x"fe",
          1558 => x"bf",
          1559 => x"75",
          1560 => x"83",
          1561 => x"83",
          1562 => x"fc",
          1563 => x"51",
          1564 => x"33",
          1565 => x"d7",
          1566 => x"db",
          1567 => x"f1",
          1568 => x"86",
          1569 => x"52",
          1570 => x"3f",
          1571 => x"2e",
          1572 => x"f0",
          1573 => x"b1",
          1574 => x"73",
          1575 => x"83",
          1576 => x"11",
          1577 => x"b1",
          1578 => x"75",
          1579 => x"83",
          1580 => x"11",
          1581 => x"b1",
          1582 => x"73",
          1583 => x"83",
          1584 => x"11",
          1585 => x"b0",
          1586 => x"74",
          1587 => x"83",
          1588 => x"11",
          1589 => x"b0",
          1590 => x"75",
          1591 => x"83",
          1592 => x"11",
          1593 => x"b0",
          1594 => x"73",
          1595 => x"83",
          1596 => x"83",
          1597 => x"83",
          1598 => x"f9",
          1599 => x"02",
          1600 => x"8c",
          1601 => x"05",
          1602 => x"51",
          1603 => x"04",
          1604 => x"3f",
          1605 => x"51",
          1606 => x"04",
          1607 => x"3f",
          1608 => x"51",
          1609 => x"04",
          1610 => x"3f",
          1611 => x"0c",
          1612 => x"0c",
          1613 => x"96",
          1614 => x"3d",
          1615 => x"70",
          1616 => x"08",
          1617 => x"e4",
          1618 => x"ff",
          1619 => x"80",
          1620 => x"3f",
          1621 => x"38",
          1622 => x"e4",
          1623 => x"84",
          1624 => x"b8",
          1625 => x"55",
          1626 => x"70",
          1627 => x"78",
          1628 => x"38",
          1629 => x"53",
          1630 => x"e4",
          1631 => x"38",
          1632 => x"0d",
          1633 => x"fa",
          1634 => x"e8",
          1635 => x"3f",
          1636 => x"08",
          1637 => x"76",
          1638 => x"d2",
          1639 => x"a9",
          1640 => x"3d",
          1641 => x"72",
          1642 => x"2e",
          1643 => x"59",
          1644 => x"d8",
          1645 => x"ba",
          1646 => x"52",
          1647 => x"b8",
          1648 => x"54",
          1649 => x"82",
          1650 => x"ff",
          1651 => x"38",
          1652 => x"aa",
          1653 => x"3d",
          1654 => x"51",
          1655 => x"80",
          1656 => x"52",
          1657 => x"e4",
          1658 => x"2e",
          1659 => x"06",
          1660 => x"38",
          1661 => x"56",
          1662 => x"15",
          1663 => x"a0",
          1664 => x"75",
          1665 => x"3d",
          1666 => x"b8",
          1667 => x"52",
          1668 => x"e4",
          1669 => x"08",
          1670 => x"ce",
          1671 => x"2e",
          1672 => x"3f",
          1673 => x"84",
          1674 => x"b8",
          1675 => x"55",
          1676 => x"81",
          1677 => x"ab",
          1678 => x"06",
          1679 => x"e4",
          1680 => x"0d",
          1681 => x"3d",
          1682 => x"3d",
          1683 => x"d0",
          1684 => x"83",
          1685 => x"2e",
          1686 => x"8d",
          1687 => x"78",
          1688 => x"fd",
          1689 => x"80",
          1690 => x"08",
          1691 => x"79",
          1692 => x"06",
          1693 => x"70",
          1694 => x"98",
          1695 => x"05",
          1696 => x"70",
          1697 => x"5d",
          1698 => x"57",
          1699 => x"75",
          1700 => x"0a",
          1701 => x"2c",
          1702 => x"38",
          1703 => x"57",
          1704 => x"42",
          1705 => x"dd",
          1706 => x"41",
          1707 => x"80",
          1708 => x"34",
          1709 => x"38",
          1710 => x"2c",
          1711 => x"70",
          1712 => x"82",
          1713 => x"53",
          1714 => x"78",
          1715 => x"a0",
          1716 => x"ff",
          1717 => x"81",
          1718 => x"81",
          1719 => x"26",
          1720 => x"82",
          1721 => x"f0",
          1722 => x"ce",
          1723 => x"70",
          1724 => x"bc",
          1725 => x"fe",
          1726 => x"fe",
          1727 => x"fd",
          1728 => x"38",
          1729 => x"d0",
          1730 => x"0c",
          1731 => x"38",
          1732 => x"57",
          1733 => x"08",
          1734 => x"34",
          1735 => x"39",
          1736 => x"2e",
          1737 => x"52",
          1738 => x"d0",
          1739 => x"d0",
          1740 => x"a8",
          1741 => x"a4",
          1742 => x"fc",
          1743 => x"81",
          1744 => x"7b",
          1745 => x"e0",
          1746 => x"8b",
          1747 => x"80",
          1748 => x"83",
          1749 => x"7c",
          1750 => x"a8",
          1751 => x"38",
          1752 => x"ff",
          1753 => x"52",
          1754 => x"d4",
          1755 => x"90",
          1756 => x"5b",
          1757 => x"ff",
          1758 => x"ff",
          1759 => x"34",
          1760 => x"f2",
          1761 => x"7c",
          1762 => x"11",
          1763 => x"74",
          1764 => x"38",
          1765 => x"b8",
          1766 => x"b8",
          1767 => x"53",
          1768 => x"3f",
          1769 => x"33",
          1770 => x"38",
          1771 => x"ff",
          1772 => x"52",
          1773 => x"d4",
          1774 => x"f8",
          1775 => x"55",
          1776 => x"ff",
          1777 => x"33",
          1778 => x"33",
          1779 => x"af",
          1780 => x"15",
          1781 => x"16",
          1782 => x"3f",
          1783 => x"06",
          1784 => x"75",
          1785 => x"c8",
          1786 => x"d0",
          1787 => x"55",
          1788 => x"33",
          1789 => x"33",
          1790 => x"a9",
          1791 => x"33",
          1792 => x"76",
          1793 => x"7a",
          1794 => x"70",
          1795 => x"57",
          1796 => x"84",
          1797 => x"b2",
          1798 => x"98",
          1799 => x"33",
          1800 => x"f9",
          1801 => x"88",
          1802 => x"80",
          1803 => x"98",
          1804 => x"5a",
          1805 => x"d4",
          1806 => x"f8",
          1807 => x"80",
          1808 => x"a4",
          1809 => x"ff",
          1810 => x"58",
          1811 => x"c8",
          1812 => x"c8",
          1813 => x"80",
          1814 => x"a4",
          1815 => x"fe",
          1816 => x"33",
          1817 => x"77",
          1818 => x"81",
          1819 => x"70",
          1820 => x"57",
          1821 => x"fe",
          1822 => x"74",
          1823 => x"c8",
          1824 => x"3f",
          1825 => x"76",
          1826 => x"06",
          1827 => x"7c",
          1828 => x"c8",
          1829 => x"3f",
          1830 => x"8b",
          1831 => x"06",
          1832 => x"a4",
          1833 => x"38",
          1834 => x"83",
          1835 => x"56",
          1836 => x"87",
          1837 => x"18",
          1838 => x"3f",
          1839 => x"f2",
          1840 => x"fc",
          1841 => x"8b",
          1842 => x"75",
          1843 => x"33",
          1844 => x"80",
          1845 => x"84",
          1846 => x"0c",
          1847 => x"33",
          1848 => x"d4",
          1849 => x"a0",
          1850 => x"51",
          1851 => x"08",
          1852 => x"84",
          1853 => x"84",
          1854 => x"55",
          1855 => x"ff",
          1856 => x"a8",
          1857 => x"f5",
          1858 => x"81",
          1859 => x"74",
          1860 => x"08",
          1861 => x"84",
          1862 => x"ae",
          1863 => x"88",
          1864 => x"a8",
          1865 => x"a8",
          1866 => x"cc",
          1867 => x"aa",
          1868 => x"80",
          1869 => x"b8",
          1870 => x"d0",
          1871 => x"56",
          1872 => x"d0",
          1873 => x"d0",
          1874 => x"d0",
          1875 => x"88",
          1876 => x"a8",
          1877 => x"84",
          1878 => x"76",
          1879 => x"c8",
          1880 => x"3f",
          1881 => x"70",
          1882 => x"57",
          1883 => x"38",
          1884 => x"ff",
          1885 => x"29",
          1886 => x"84",
          1887 => x"79",
          1888 => x"08",
          1889 => x"74",
          1890 => x"05",
          1891 => x"5b",
          1892 => x"38",
          1893 => x"17",
          1894 => x"52",
          1895 => x"75",
          1896 => x"05",
          1897 => x"43",
          1898 => x"38",
          1899 => x"34",
          1900 => x"51",
          1901 => x"0a",
          1902 => x"2c",
          1903 => x"60",
          1904 => x"39",
          1905 => x"06",
          1906 => x"38",
          1907 => x"27",
          1908 => x"2c",
          1909 => x"7b",
          1910 => x"75",
          1911 => x"05",
          1912 => x"52",
          1913 => x"81",
          1914 => x"77",
          1915 => x"3d",
          1916 => x"57",
          1917 => x"56",
          1918 => x"84",
          1919 => x"29",
          1920 => x"79",
          1921 => x"60",
          1922 => x"2b",
          1923 => x"5c",
          1924 => x"38",
          1925 => x"ff",
          1926 => x"29",
          1927 => x"84",
          1928 => x"75",
          1929 => x"08",
          1930 => x"75",
          1931 => x"05",
          1932 => x"57",
          1933 => x"38",
          1934 => x"56",
          1935 => x"51",
          1936 => x"08",
          1937 => x"08",
          1938 => x"52",
          1939 => x"d0",
          1940 => x"56",
          1941 => x"d4",
          1942 => x"b8",
          1943 => x"51",
          1944 => x"08",
          1945 => x"84",
          1946 => x"84",
          1947 => x"55",
          1948 => x"3f",
          1949 => x"0c",
          1950 => x"76",
          1951 => x"38",
          1952 => x"52",
          1953 => x"a8",
          1954 => x"81",
          1955 => x"d0",
          1956 => x"24",
          1957 => x"98",
          1958 => x"06",
          1959 => x"ef",
          1960 => x"d0",
          1961 => x"f1",
          1962 => x"74",
          1963 => x"56",
          1964 => x"83",
          1965 => x"55",
          1966 => x"51",
          1967 => x"08",
          1968 => x"83",
          1969 => x"5f",
          1970 => x"d9",
          1971 => x"84",
          1972 => x"ac",
          1973 => x"aa",
          1974 => x"d0",
          1975 => x"ff",
          1976 => x"51",
          1977 => x"d0",
          1978 => x"57",
          1979 => x"84",
          1980 => x"a7",
          1981 => x"a0",
          1982 => x"c8",
          1983 => x"3f",
          1984 => x"79",
          1985 => x"06",
          1986 => x"0b",
          1987 => x"d0",
          1988 => x"b4",
          1989 => x"fa",
          1990 => x"a4",
          1991 => x"06",
          1992 => x"ff",
          1993 => x"ff",
          1994 => x"a8",
          1995 => x"2e",
          1996 => x"52",
          1997 => x"d4",
          1998 => x"f8",
          1999 => x"51",
          2000 => x"33",
          2001 => x"34",
          2002 => x"75",
          2003 => x"e4",
          2004 => x"e4",
          2005 => x"75",
          2006 => x"ff",
          2007 => x"a4",
          2008 => x"5e",
          2009 => x"84",
          2010 => x"a5",
          2011 => x"a0",
          2012 => x"c8",
          2013 => x"3f",
          2014 => x"60",
          2015 => x"06",
          2016 => x"fa",
          2017 => x"2b",
          2018 => x"81",
          2019 => x"dc",
          2020 => x"0c",
          2021 => x"83",
          2022 => x"41",
          2023 => x"53",
          2024 => x"3f",
          2025 => x"81",
          2026 => x"82",
          2027 => x"f4",
          2028 => x"54",
          2029 => x"d8",
          2030 => x"8a",
          2031 => x"d0",
          2032 => x"0b",
          2033 => x"d0",
          2034 => x"b4",
          2035 => x"84",
          2036 => x"3f",
          2037 => x"84",
          2038 => x"83",
          2039 => x"7a",
          2040 => x"e4",
          2041 => x"2e",
          2042 => x"b8",
          2043 => x"84",
          2044 => x"b8",
          2045 => x"b8",
          2046 => x"56",
          2047 => x"83",
          2048 => x"f1",
          2049 => x"59",
          2050 => x"87",
          2051 => x"1a",
          2052 => x"3f",
          2053 => x"f2",
          2054 => x"fc",
          2055 => x"a0",
          2056 => x"5e",
          2057 => x"5d",
          2058 => x"df",
          2059 => x"39",
          2060 => x"a6",
          2061 => x"05",
          2062 => x"7a",
          2063 => x"f2",
          2064 => x"80",
          2065 => x"70",
          2066 => x"fc",
          2067 => x"57",
          2068 => x"08",
          2069 => x"10",
          2070 => x"57",
          2071 => x"38",
          2072 => x"34",
          2073 => x"34",
          2074 => x"ff",
          2075 => x"f8",
          2076 => x"c3",
          2077 => x"05",
          2078 => x"8d",
          2079 => x"81",
          2080 => x"2e",
          2081 => x"59",
          2082 => x"80",
          2083 => x"90",
          2084 => x"83",
          2085 => x"23",
          2086 => x"71",
          2087 => x"71",
          2088 => x"78",
          2089 => x"84",
          2090 => x"05",
          2091 => x"75",
          2092 => x"33",
          2093 => x"55",
          2094 => x"34",
          2095 => x"ff",
          2096 => x"0d",
          2097 => x"f8",
          2098 => x"f8",
          2099 => x"05",
          2100 => x"b0",
          2101 => x"81",
          2102 => x"81",
          2103 => x"83",
          2104 => x"59",
          2105 => x"73",
          2106 => x"29",
          2107 => x"ff",
          2108 => x"ff",
          2109 => x"75",
          2110 => x"5c",
          2111 => x"94",
          2112 => x"29",
          2113 => x"7b",
          2114 => x"55",
          2115 => x"80",
          2116 => x"f8",
          2117 => x"34",
          2118 => x"86",
          2119 => x"33",
          2120 => x"33",
          2121 => x"22",
          2122 => x"5e",
          2123 => x"df",
          2124 => x"ff",
          2125 => x"54",
          2126 => x"0b",
          2127 => x"f8",
          2128 => x"98",
          2129 => x"2b",
          2130 => x"56",
          2131 => x"fd",
          2132 => x"f8",
          2133 => x"10",
          2134 => x"90",
          2135 => x"5e",
          2136 => x"b0",
          2137 => x"70",
          2138 => x"70",
          2139 => x"70",
          2140 => x"60",
          2141 => x"40",
          2142 => x"72",
          2143 => x"57",
          2144 => x"ff",
          2145 => x"ff",
          2146 => x"29",
          2147 => x"78",
          2148 => x"79",
          2149 => x"58",
          2150 => x"5c",
          2151 => x"74",
          2152 => x"39",
          2153 => x"53",
          2154 => x"85",
          2155 => x"80",
          2156 => x"b0",
          2157 => x"80",
          2158 => x"80",
          2159 => x"34",
          2160 => x"51",
          2161 => x"70",
          2162 => x"a0",
          2163 => x"54",
          2164 => x"80",
          2165 => x"72",
          2166 => x"70",
          2167 => x"86",
          2168 => x"f7",
          2169 => x"80",
          2170 => x"0b",
          2171 => x"04",
          2172 => x"0c",
          2173 => x"33",
          2174 => x"b6",
          2175 => x"75",
          2176 => x"d8",
          2177 => x"94",
          2178 => x"a0",
          2179 => x"51",
          2180 => x"83",
          2181 => x"53",
          2182 => x"c4",
          2183 => x"55",
          2184 => x"94",
          2185 => x"7a",
          2186 => x"7a",
          2187 => x"72",
          2188 => x"22",
          2189 => x"d6",
          2190 => x"82",
          2191 => x"71",
          2192 => x"9f",
          2193 => x"14",
          2194 => x"e0",
          2195 => x"33",
          2196 => x"14",
          2197 => x"38",
          2198 => x"f8",
          2199 => x"55",
          2200 => x"73",
          2201 => x"54",
          2202 => x"b6",
          2203 => x"f8",
          2204 => x"06",
          2205 => x"73",
          2206 => x"31",
          2207 => x"71",
          2208 => x"a7",
          2209 => x"79",
          2210 => x"71",
          2211 => x"75",
          2212 => x"16",
          2213 => x"b6",
          2214 => x"5a",
          2215 => x"77",
          2216 => x"84",
          2217 => x"71",
          2218 => x"72",
          2219 => x"84",
          2220 => x"74",
          2221 => x"22",
          2222 => x"d6",
          2223 => x"fd",
          2224 => x"38",
          2225 => x"f8",
          2226 => x"09",
          2227 => x"31",
          2228 => x"71",
          2229 => x"59",
          2230 => x"83",
          2231 => x"74",
          2232 => x"e0",
          2233 => x"05",
          2234 => x"2e",
          2235 => x"16",
          2236 => x"34",
          2237 => x"f4",
          2238 => x"55",
          2239 => x"15",
          2240 => x"74",
          2241 => x"a9",
          2242 => x"05",
          2243 => x"26",
          2244 => x"dc",
          2245 => x"d8",
          2246 => x"71",
          2247 => x"b8",
          2248 => x"0b",
          2249 => x"33",
          2250 => x"80",
          2251 => x"83",
          2252 => x"e4",
          2253 => x"94",
          2254 => x"9f",
          2255 => x"70",
          2256 => x"f8",
          2257 => x"33",
          2258 => x"25",
          2259 => x"94",
          2260 => x"86",
          2261 => x"70",
          2262 => x"72",
          2263 => x"f8",
          2264 => x"0c",
          2265 => x"33",
          2266 => x"11",
          2267 => x"38",
          2268 => x"80",
          2269 => x"0d",
          2270 => x"83",
          2271 => x"ff",
          2272 => x"b4",
          2273 => x"94",
          2274 => x"02",
          2275 => x"b3",
          2276 => x"05",
          2277 => x"33",
          2278 => x"80",
          2279 => x"51",
          2280 => x"09",
          2281 => x"83",
          2282 => x"e4",
          2283 => x"90",
          2284 => x"70",
          2285 => x"b8",
          2286 => x"f8",
          2287 => x"83",
          2288 => x"90",
          2289 => x"70",
          2290 => x"f1",
          2291 => x"84",
          2292 => x"83",
          2293 => x"07",
          2294 => x"b4",
          2295 => x"51",
          2296 => x"39",
          2297 => x"85",
          2298 => x"ff",
          2299 => x"fb",
          2300 => x"90",
          2301 => x"33",
          2302 => x"83",
          2303 => x"f8",
          2304 => x"83",
          2305 => x"f8",
          2306 => x"07",
          2307 => x"cc",
          2308 => x"06",
          2309 => x"34",
          2310 => x"81",
          2311 => x"83",
          2312 => x"f8",
          2313 => x"07",
          2314 => x"94",
          2315 => x"06",
          2316 => x"34",
          2317 => x"81",
          2318 => x"34",
          2319 => x"81",
          2320 => x"f8",
          2321 => x"0d",
          2322 => x"80",
          2323 => x"83",
          2324 => x"84",
          2325 => x"5b",
          2326 => x"78",
          2327 => x"81",
          2328 => x"80",
          2329 => x"f8",
          2330 => x"7c",
          2331 => x"04",
          2332 => x"38",
          2333 => x"0b",
          2334 => x"f8",
          2335 => x"34",
          2336 => x"58",
          2337 => x"d7",
          2338 => x"7b",
          2339 => x"d8",
          2340 => x"b6",
          2341 => x"34",
          2342 => x"f8",
          2343 => x"8f",
          2344 => x"da",
          2345 => x"80",
          2346 => x"83",
          2347 => x"92",
          2348 => x"b7",
          2349 => x"56",
          2350 => x"52",
          2351 => x"3f",
          2352 => x"5a",
          2353 => x"84",
          2354 => x"83",
          2355 => x"81",
          2356 => x"e5",
          2357 => x"dd",
          2358 => x"d2",
          2359 => x"0b",
          2360 => x"94",
          2361 => x"83",
          2362 => x"80",
          2363 => x"84",
          2364 => x"94",
          2365 => x"81",
          2366 => x"c8",
          2367 => x"e4",
          2368 => x"80",
          2369 => x"51",
          2370 => x"e4",
          2371 => x"c8",
          2372 => x"fe",
          2373 => x"ff",
          2374 => x"0d",
          2375 => x"84",
          2376 => x"83",
          2377 => x"86",
          2378 => x"22",
          2379 => x"05",
          2380 => x"ea",
          2381 => x"72",
          2382 => x"2e",
          2383 => x"b9",
          2384 => x"75",
          2385 => x"d8",
          2386 => x"95",
          2387 => x"54",
          2388 => x"a0",
          2389 => x"83",
          2390 => x"72",
          2391 => x"75",
          2392 => x"94",
          2393 => x"83",
          2394 => x"18",
          2395 => x"ff",
          2396 => x"95",
          2397 => x"57",
          2398 => x"97",
          2399 => x"ff",
          2400 => x"99",
          2401 => x"81",
          2402 => x"f8",
          2403 => x"72",
          2404 => x"33",
          2405 => x"80",
          2406 => x"0d",
          2407 => x"8d",
          2408 => x"09",
          2409 => x"81",
          2410 => x"f8",
          2411 => x"96",
          2412 => x"33",
          2413 => x"06",
          2414 => x"a0",
          2415 => x"81",
          2416 => x"ff",
          2417 => x"a5",
          2418 => x"54",
          2419 => x"fa",
          2420 => x"f2",
          2421 => x"3f",
          2422 => x"3d",
          2423 => x"81",
          2424 => x"33",
          2425 => x"53",
          2426 => x"f8",
          2427 => x"d5",
          2428 => x"ff",
          2429 => x"a5",
          2430 => x"34",
          2431 => x"95",
          2432 => x"3f",
          2433 => x"ef",
          2434 => x"0d",
          2435 => x"e0",
          2436 => x"b8",
          2437 => x"78",
          2438 => x"24",
          2439 => x"b9",
          2440 => x"84",
          2441 => x"83",
          2442 => x"58",
          2443 => x"86",
          2444 => x"d8",
          2445 => x"92",
          2446 => x"42",
          2447 => x"83",
          2448 => x"05",
          2449 => x"86",
          2450 => x"d8",
          2451 => x"92",
          2452 => x"29",
          2453 => x"f8",
          2454 => x"81",
          2455 => x"76",
          2456 => x"d9",
          2457 => x"19",
          2458 => x"0b",
          2459 => x"04",
          2460 => x"79",
          2461 => x"9b",
          2462 => x"cc",
          2463 => x"84",
          2464 => x"83",
          2465 => x"5e",
          2466 => x"86",
          2467 => x"d8",
          2468 => x"92",
          2469 => x"59",
          2470 => x"83",
          2471 => x"5b",
          2472 => x"b0",
          2473 => x"70",
          2474 => x"83",
          2475 => x"44",
          2476 => x"33",
          2477 => x"1f",
          2478 => x"77",
          2479 => x"95",
          2480 => x"9c",
          2481 => x"b7",
          2482 => x"78",
          2483 => x"38",
          2484 => x"0b",
          2485 => x"04",
          2486 => x"19",
          2487 => x"84",
          2488 => x"77",
          2489 => x"e8",
          2490 => x"80",
          2491 => x"0b",
          2492 => x"04",
          2493 => x"0b",
          2494 => x"33",
          2495 => x"33",
          2496 => x"84",
          2497 => x"80",
          2498 => x"f8",
          2499 => x"71",
          2500 => x"83",
          2501 => x"33",
          2502 => x"f8",
          2503 => x"34",
          2504 => x"06",
          2505 => x"33",
          2506 => x"58",
          2507 => x"97",
          2508 => x"89",
          2509 => x"3f",
          2510 => x"ae",
          2511 => x"95",
          2512 => x"94",
          2513 => x"a0",
          2514 => x"51",
          2515 => x"ff",
          2516 => x"51",
          2517 => x"a4",
          2518 => x"57",
          2519 => x"75",
          2520 => x"80",
          2521 => x"84",
          2522 => x"e6",
          2523 => x"81",
          2524 => x"84",
          2525 => x"83",
          2526 => x"83",
          2527 => x"83",
          2528 => x"80",
          2529 => x"84",
          2530 => x"78",
          2531 => x"a7",
          2532 => x"d8",
          2533 => x"95",
          2534 => x"29",
          2535 => x"f8",
          2536 => x"05",
          2537 => x"ea",
          2538 => x"5c",
          2539 => x"81",
          2540 => x"83",
          2541 => x"34",
          2542 => x"06",
          2543 => x"05",
          2544 => x"86",
          2545 => x"d8",
          2546 => x"92",
          2547 => x"42",
          2548 => x"34",
          2549 => x"62",
          2550 => x"86",
          2551 => x"d8",
          2552 => x"92",
          2553 => x"29",
          2554 => x"f8",
          2555 => x"34",
          2556 => x"58",
          2557 => x"b6",
          2558 => x"ff",
          2559 => x"83",
          2560 => x"58",
          2561 => x"bb",
          2562 => x"83",
          2563 => x"38",
          2564 => x"f9",
          2565 => x"26",
          2566 => x"c5",
          2567 => x"0b",
          2568 => x"51",
          2569 => x"e4",
          2570 => x"94",
          2571 => x"ff",
          2572 => x"ff",
          2573 => x"a0",
          2574 => x"41",
          2575 => x"ff",
          2576 => x"45",
          2577 => x"82",
          2578 => x"06",
          2579 => x"06",
          2580 => x"84",
          2581 => x"1b",
          2582 => x"95",
          2583 => x"29",
          2584 => x"83",
          2585 => x"33",
          2586 => x"f8",
          2587 => x"34",
          2588 => x"06",
          2589 => x"33",
          2590 => x"40",
          2591 => x"b6",
          2592 => x"ff",
          2593 => x"ac",
          2594 => x"92",
          2595 => x"f8",
          2596 => x"06",
          2597 => x"38",
          2598 => x"33",
          2599 => x"06",
          2600 => x"06",
          2601 => x"5b",
          2602 => x"a7",
          2603 => x"33",
          2604 => x"22",
          2605 => x"56",
          2606 => x"83",
          2607 => x"5a",
          2608 => x"b0",
          2609 => x"70",
          2610 => x"83",
          2611 => x"5b",
          2612 => x"33",
          2613 => x"05",
          2614 => x"7f",
          2615 => x"95",
          2616 => x"b7",
          2617 => x"0c",
          2618 => x"17",
          2619 => x"7a",
          2620 => x"ff",
          2621 => x"39",
          2622 => x"0b",
          2623 => x"04",
          2624 => x"b6",
          2625 => x"94",
          2626 => x"95",
          2627 => x"f4",
          2628 => x"dc",
          2629 => x"d8",
          2630 => x"fb",
          2631 => x"11",
          2632 => x"79",
          2633 => x"ca",
          2634 => x"23",
          2635 => x"33",
          2636 => x"34",
          2637 => x"33",
          2638 => x"f9",
          2639 => x"f8",
          2640 => x"72",
          2641 => x"e0",
          2642 => x"05",
          2643 => x"95",
          2644 => x"29",
          2645 => x"f8",
          2646 => x"76",
          2647 => x"90",
          2648 => x"34",
          2649 => x"06",
          2650 => x"33",
          2651 => x"42",
          2652 => x"b6",
          2653 => x"06",
          2654 => x"38",
          2655 => x"e2",
          2656 => x"95",
          2657 => x"84",
          2658 => x"f3",
          2659 => x"75",
          2660 => x"ea",
          2661 => x"0c",
          2662 => x"33",
          2663 => x"33",
          2664 => x"33",
          2665 => x"b9",
          2666 => x"cc",
          2667 => x"cd",
          2668 => x"ce",
          2669 => x"33",
          2670 => x"84",
          2671 => x"09",
          2672 => x"95",
          2673 => x"33",
          2674 => x"a0",
          2675 => x"ee",
          2676 => x"3f",
          2677 => x"83",
          2678 => x"60",
          2679 => x"83",
          2680 => x"fe",
          2681 => x"33",
          2682 => x"77",
          2683 => x"84",
          2684 => x"41",
          2685 => x"10",
          2686 => x"08",
          2687 => x"80",
          2688 => x"33",
          2689 => x"70",
          2690 => x"42",
          2691 => x"34",
          2692 => x"56",
          2693 => x"b8",
          2694 => x"06",
          2695 => x"75",
          2696 => x"f8",
          2697 => x"83",
          2698 => x"70",
          2699 => x"2e",
          2700 => x"83",
          2701 => x"0b",
          2702 => x"33",
          2703 => x"57",
          2704 => x"17",
          2705 => x"f9",
          2706 => x"80",
          2707 => x"33",
          2708 => x"70",
          2709 => x"41",
          2710 => x"34",
          2711 => x"5b",
          2712 => x"b8",
          2713 => x"81",
          2714 => x"33",
          2715 => x"33",
          2716 => x"80",
          2717 => x"5a",
          2718 => x"ff",
          2719 => x"ff",
          2720 => x"7e",
          2721 => x"80",
          2722 => x"39",
          2723 => x"2e",
          2724 => x"58",
          2725 => x"d9",
          2726 => x"fb",
          2727 => x"75",
          2728 => x"b9",
          2729 => x"05",
          2730 => x"5e",
          2731 => x"57",
          2732 => x"39",
          2733 => x"2e",
          2734 => x"83",
          2735 => x"b6",
          2736 => x"75",
          2737 => x"83",
          2738 => x"e3",
          2739 => x"0b",
          2740 => x"76",
          2741 => x"b8",
          2742 => x"e3",
          2743 => x"17",
          2744 => x"33",
          2745 => x"84",
          2746 => x"2e",
          2747 => x"75",
          2748 => x"52",
          2749 => x"3f",
          2750 => x"57",
          2751 => x"b8",
          2752 => x"06",
          2753 => x"81",
          2754 => x"81",
          2755 => x"5b",
          2756 => x"38",
          2757 => x"76",
          2758 => x"77",
          2759 => x"83",
          2760 => x"ff",
          2761 => x"b4",
          2762 => x"34",
          2763 => x"5f",
          2764 => x"b8",
          2765 => x"5b",
          2766 => x"f8",
          2767 => x"81",
          2768 => x"74",
          2769 => x"83",
          2770 => x"29",
          2771 => x"f6",
          2772 => x"5d",
          2773 => x"83",
          2774 => x"57",
          2775 => x"b6",
          2776 => x"d6",
          2777 => x"92",
          2778 => x"31",
          2779 => x"38",
          2780 => x"27",
          2781 => x"83",
          2782 => x"83",
          2783 => x"76",
          2784 => x"81",
          2785 => x"29",
          2786 => x"a0",
          2787 => x"81",
          2788 => x"71",
          2789 => x"7f",
          2790 => x"1a",
          2791 => x"b6",
          2792 => x"5d",
          2793 => x"7c",
          2794 => x"84",
          2795 => x"71",
          2796 => x"77",
          2797 => x"17",
          2798 => x"7b",
          2799 => x"81",
          2800 => x"5e",
          2801 => x"84",
          2802 => x"43",
          2803 => x"99",
          2804 => x"33",
          2805 => x"80",
          2806 => x"b1",
          2807 => x"b6",
          2808 => x"33",
          2809 => x"94",
          2810 => x"78",
          2811 => x"83",
          2812 => x"06",
          2813 => x"5c",
          2814 => x"b6",
          2815 => x"89",
          2816 => x"76",
          2817 => x"61",
          2818 => x"38",
          2819 => x"62",
          2820 => x"1f",
          2821 => x"79",
          2822 => x"ac",
          2823 => x"a4",
          2824 => x"2b",
          2825 => x"07",
          2826 => x"57",
          2827 => x"70",
          2828 => x"84",
          2829 => x"38",
          2830 => x"33",
          2831 => x"81",
          2832 => x"73",
          2833 => x"77",
          2834 => x"1b",
          2835 => x"75",
          2836 => x"f4",
          2837 => x"97",
          2838 => x"e0",
          2839 => x"5a",
          2840 => x"f4",
          2841 => x"34",
          2842 => x"81",
          2843 => x"f4",
          2844 => x"06",
          2845 => x"90",
          2846 => x"2b",
          2847 => x"58",
          2848 => x"81",
          2849 => x"f8",
          2850 => x"06",
          2851 => x"96",
          2852 => x"33",
          2853 => x"b6",
          2854 => x"b6",
          2855 => x"ee",
          2856 => x"56",
          2857 => x"70",
          2858 => x"39",
          2859 => x"85",
          2860 => x"e5",
          2861 => x"06",
          2862 => x"34",
          2863 => x"f9",
          2864 => x"90",
          2865 => x"81",
          2866 => x"f8",
          2867 => x"0b",
          2868 => x"81",
          2869 => x"83",
          2870 => x"75",
          2871 => x"83",
          2872 => x"07",
          2873 => x"fd",
          2874 => x"06",
          2875 => x"90",
          2876 => x"33",
          2877 => x"75",
          2878 => x"83",
          2879 => x"07",
          2880 => x"c5",
          2881 => x"06",
          2882 => x"34",
          2883 => x"81",
          2884 => x"f8",
          2885 => x"90",
          2886 => x"75",
          2887 => x"83",
          2888 => x"75",
          2889 => x"83",
          2890 => x"75",
          2891 => x"83",
          2892 => x"75",
          2893 => x"83",
          2894 => x"d0",
          2895 => x"fd",
          2896 => x"bf",
          2897 => x"90",
          2898 => x"f8",
          2899 => x"c9",
          2900 => x"33",
          2901 => x"33",
          2902 => x"33",
          2903 => x"0b",
          2904 => x"81",
          2905 => x"84",
          2906 => x"77",
          2907 => x"33",
          2908 => x"56",
          2909 => x"9c",
          2910 => x"fe",
          2911 => x"a1",
          2912 => x"e0",
          2913 => x"80",
          2914 => x"0d",
          2915 => x"e9",
          2916 => x"5c",
          2917 => x"10",
          2918 => x"05",
          2919 => x"0b",
          2920 => x"0b",
          2921 => x"51",
          2922 => x"70",
          2923 => x"e6",
          2924 => x"34",
          2925 => x"ef",
          2926 => x"3f",
          2927 => x"ff",
          2928 => x"06",
          2929 => x"52",
          2930 => x"33",
          2931 => x"75",
          2932 => x"83",
          2933 => x"70",
          2934 => x"f0",
          2935 => x"05",
          2936 => x"59",
          2937 => x"75",
          2938 => x"33",
          2939 => x"77",
          2940 => x"33",
          2941 => x"06",
          2942 => x"11",
          2943 => x"92",
          2944 => x"70",
          2945 => x"33",
          2946 => x"81",
          2947 => x"ff",
          2948 => x"24",
          2949 => x"56",
          2950 => x"16",
          2951 => x"81",
          2952 => x"76",
          2953 => x"33",
          2954 => x"ff",
          2955 => x"7b",
          2956 => x"57",
          2957 => x"38",
          2958 => x"ff",
          2959 => x"79",
          2960 => x"a7",
          2961 => x"81",
          2962 => x"42",
          2963 => x"38",
          2964 => x"17",
          2965 => x"7b",
          2966 => x"81",
          2967 => x"5f",
          2968 => x"84",
          2969 => x"59",
          2970 => x"b1",
          2971 => x"b6",
          2972 => x"5d",
          2973 => x"7d",
          2974 => x"84",
          2975 => x"71",
          2976 => x"75",
          2977 => x"39",
          2978 => x"b6",
          2979 => x"94",
          2980 => x"92",
          2981 => x"5f",
          2982 => x"38",
          2983 => x"06",
          2984 => x"27",
          2985 => x"92",
          2986 => x"58",
          2987 => x"57",
          2988 => x"d8",
          2989 => x"52",
          2990 => x"38",
          2991 => x"eb",
          2992 => x"05",
          2993 => x"40",
          2994 => x"75",
          2995 => x"09",
          2996 => x"95",
          2997 => x"94",
          2998 => x"ff",
          2999 => x"f6",
          3000 => x"f8",
          3001 => x"56",
          3002 => x"39",
          3003 => x"94",
          3004 => x"56",
          3005 => x"76",
          3006 => x"90",
          3007 => x"75",
          3008 => x"70",
          3009 => x"33",
          3010 => x"76",
          3011 => x"7b",
          3012 => x"f1",
          3013 => x"34",
          3014 => x"23",
          3015 => x"92",
          3016 => x"f8",
          3017 => x"96",
          3018 => x"33",
          3019 => x"34",
          3020 => x"97",
          3021 => x"54",
          3022 => x"db",
          3023 => x"0c",
          3024 => x"51",
          3025 => x"e4",
          3026 => x"0d",
          3027 => x"83",
          3028 => x"83",
          3029 => x"59",
          3030 => x"14",
          3031 => x"59",
          3032 => x"0d",
          3033 => x"53",
          3034 => x"32",
          3035 => x"9f",
          3036 => x"f6",
          3037 => x"81",
          3038 => x"54",
          3039 => x"25",
          3040 => x"2e",
          3041 => x"83",
          3042 => x"72",
          3043 => x"05",
          3044 => x"71",
          3045 => x"06",
          3046 => x"58",
          3047 => x"f0",
          3048 => x"80",
          3049 => x"c0",
          3050 => x"f6",
          3051 => x"76",
          3052 => x"70",
          3053 => x"74",
          3054 => x"84",
          3055 => x"f6",
          3056 => x"76",
          3057 => x"2e",
          3058 => x"15",
          3059 => x"81",
          3060 => x"f6",
          3061 => x"33",
          3062 => x"70",
          3063 => x"27",
          3064 => x"70",
          3065 => x"54",
          3066 => x"ff",
          3067 => x"81",
          3068 => x"85",
          3069 => x"34",
          3070 => x"2e",
          3071 => x"be",
          3072 => x"83",
          3073 => x"70",
          3074 => x"33",
          3075 => x"83",
          3076 => x"ff",
          3077 => x"33",
          3078 => x"83",
          3079 => x"ff",
          3080 => x"33",
          3081 => x"ff",
          3082 => x"38",
          3083 => x"81",
          3084 => x"06",
          3085 => x"38",
          3086 => x"74",
          3087 => x"08",
          3088 => x"08",
          3089 => x"38",
          3090 => x"83",
          3091 => x"81",
          3092 => x"fe",
          3093 => x"77",
          3094 => x"53",
          3095 => x"10",
          3096 => x"08",
          3097 => x"80",
          3098 => x"c0",
          3099 => x"27",
          3100 => x"ea",
          3101 => x"38",
          3102 => x"87",
          3103 => x"0c",
          3104 => x"2e",
          3105 => x"54",
          3106 => x"81",
          3107 => x"c4",
          3108 => x"38",
          3109 => x"c3",
          3110 => x"39",
          3111 => x"56",
          3112 => x"38",
          3113 => x"b4",
          3114 => x"79",
          3115 => x"ff",
          3116 => x"2b",
          3117 => x"73",
          3118 => x"81",
          3119 => x"87",
          3120 => x"57",
          3121 => x"78",
          3122 => x"11",
          3123 => x"05",
          3124 => x"c0",
          3125 => x"57",
          3126 => x"2e",
          3127 => x"59",
          3128 => x"39",
          3129 => x"0b",
          3130 => x"81",
          3131 => x"70",
          3132 => x"59",
          3133 => x"09",
          3134 => x"2e",
          3135 => x"10",
          3136 => x"5d",
          3137 => x"81",
          3138 => x"93",
          3139 => x"33",
          3140 => x"84",
          3141 => x"38",
          3142 => x"cc",
          3143 => x"8f",
          3144 => x"f0",
          3145 => x"2e",
          3146 => x"81",
          3147 => x"34",
          3148 => x"ac",
          3149 => x"15",
          3150 => x"34",
          3151 => x"53",
          3152 => x"83",
          3153 => x"27",
          3154 => x"54",
          3155 => x"fc",
          3156 => x"05",
          3157 => x"74",
          3158 => x"98",
          3159 => x"81",
          3160 => x"0b",
          3161 => x"39",
          3162 => x"81",
          3163 => x"83",
          3164 => x"bd",
          3165 => x"be",
          3166 => x"f6",
          3167 => x"5e",
          3168 => x"09",
          3169 => x"7a",
          3170 => x"2e",
          3171 => x"93",
          3172 => x"f8",
          3173 => x"33",
          3174 => x"73",
          3175 => x"ac",
          3176 => x"58",
          3177 => x"84",
          3178 => x"39",
          3179 => x"2e",
          3180 => x"c4",
          3181 => x"33",
          3182 => x"5a",
          3183 => x"55",
          3184 => x"ff",
          3185 => x"27",
          3186 => x"94",
          3187 => x"ff",
          3188 => x"27",
          3189 => x"95",
          3190 => x"52",
          3191 => x"59",
          3192 => x"39",
          3193 => x"51",
          3194 => x"f6",
          3195 => x"fc",
          3196 => x"f5",
          3197 => x"3d",
          3198 => x"53",
          3199 => x"34",
          3200 => x"71",
          3201 => x"55",
          3202 => x"0b",
          3203 => x"98",
          3204 => x"80",
          3205 => x"9c",
          3206 => x"51",
          3207 => x"33",
          3208 => x"74",
          3209 => x"2e",
          3210 => x"51",
          3211 => x"38",
          3212 => x"38",
          3213 => x"90",
          3214 => x"52",
          3215 => x"72",
          3216 => x"c0",
          3217 => x"27",
          3218 => x"38",
          3219 => x"75",
          3220 => x"ff",
          3221 => x"75",
          3222 => x"06",
          3223 => x"2e",
          3224 => x"88",
          3225 => x"e4",
          3226 => x"0d",
          3227 => x"56",
          3228 => x"73",
          3229 => x"70",
          3230 => x"57",
          3231 => x"51",
          3232 => x"56",
          3233 => x"34",
          3234 => x"13",
          3235 => x"e1",
          3236 => x"08",
          3237 => x"80",
          3238 => x"c0",
          3239 => x"55",
          3240 => x"98",
          3241 => x"08",
          3242 => x"14",
          3243 => x"52",
          3244 => x"fe",
          3245 => x"08",
          3246 => x"c8",
          3247 => x"c0",
          3248 => x"ce",
          3249 => x"08",
          3250 => x"74",
          3251 => x"87",
          3252 => x"73",
          3253 => x"db",
          3254 => x"72",
          3255 => x"55",
          3256 => x"53",
          3257 => x"81",
          3258 => x"74",
          3259 => x"aa",
          3260 => x"11",
          3261 => x"38",
          3262 => x"70",
          3263 => x"f0",
          3264 => x"3d",
          3265 => x"0c",
          3266 => x"39",
          3267 => x"a3",
          3268 => x"f2",
          3269 => x"80",
          3270 => x"51",
          3271 => x"72",
          3272 => x"75",
          3273 => x"72",
          3274 => x"08",
          3275 => x"54",
          3276 => x"70",
          3277 => x"81",
          3278 => x"38",
          3279 => x"15",
          3280 => x"e2",
          3281 => x"08",
          3282 => x"80",
          3283 => x"c0",
          3284 => x"55",
          3285 => x"98",
          3286 => x"08",
          3287 => x"14",
          3288 => x"52",
          3289 => x"fe",
          3290 => x"08",
          3291 => x"c8",
          3292 => x"c0",
          3293 => x"ce",
          3294 => x"08",
          3295 => x"74",
          3296 => x"87",
          3297 => x"73",
          3298 => x"db",
          3299 => x"72",
          3300 => x"55",
          3301 => x"53",
          3302 => x"ff",
          3303 => x"51",
          3304 => x"2e",
          3305 => x"e4",
          3306 => x"e8",
          3307 => x"08",
          3308 => x"83",
          3309 => x"81",
          3310 => x"e8",
          3311 => x"f2",
          3312 => x"54",
          3313 => x"c0",
          3314 => x"f6",
          3315 => x"9c",
          3316 => x"38",
          3317 => x"c0",
          3318 => x"74",
          3319 => x"ff",
          3320 => x"9c",
          3321 => x"c0",
          3322 => x"9c",
          3323 => x"81",
          3324 => x"55",
          3325 => x"81",
          3326 => x"a4",
          3327 => x"ff",
          3328 => x"ff",
          3329 => x"38",
          3330 => x"d5",
          3331 => x"e3",
          3332 => x"3d",
          3333 => x"d4",
          3334 => x"83",
          3335 => x"11",
          3336 => x"2b",
          3337 => x"33",
          3338 => x"90",
          3339 => x"5d",
          3340 => x"71",
          3341 => x"11",
          3342 => x"71",
          3343 => x"81",
          3344 => x"2b",
          3345 => x"52",
          3346 => x"13",
          3347 => x"71",
          3348 => x"2a",
          3349 => x"34",
          3350 => x"13",
          3351 => x"84",
          3352 => x"2b",
          3353 => x"54",
          3354 => x"14",
          3355 => x"80",
          3356 => x"13",
          3357 => x"84",
          3358 => x"b8",
          3359 => x"33",
          3360 => x"07",
          3361 => x"74",
          3362 => x"3d",
          3363 => x"33",
          3364 => x"75",
          3365 => x"71",
          3366 => x"58",
          3367 => x"12",
          3368 => x"d4",
          3369 => x"12",
          3370 => x"07",
          3371 => x"12",
          3372 => x"07",
          3373 => x"77",
          3374 => x"84",
          3375 => x"12",
          3376 => x"ff",
          3377 => x"52",
          3378 => x"84",
          3379 => x"81",
          3380 => x"2b",
          3381 => x"33",
          3382 => x"8f",
          3383 => x"2a",
          3384 => x"54",
          3385 => x"14",
          3386 => x"70",
          3387 => x"71",
          3388 => x"81",
          3389 => x"ff",
          3390 => x"53",
          3391 => x"34",
          3392 => x"08",
          3393 => x"33",
          3394 => x"74",
          3395 => x"98",
          3396 => x"5d",
          3397 => x"25",
          3398 => x"33",
          3399 => x"07",
          3400 => x"75",
          3401 => x"d4",
          3402 => x"33",
          3403 => x"74",
          3404 => x"71",
          3405 => x"5c",
          3406 => x"82",
          3407 => x"3d",
          3408 => x"b8",
          3409 => x"8f",
          3410 => x"51",
          3411 => x"84",
          3412 => x"a0",
          3413 => x"80",
          3414 => x"51",
          3415 => x"08",
          3416 => x"16",
          3417 => x"84",
          3418 => x"84",
          3419 => x"34",
          3420 => x"d4",
          3421 => x"fe",
          3422 => x"06",
          3423 => x"74",
          3424 => x"84",
          3425 => x"84",
          3426 => x"55",
          3427 => x"15",
          3428 => x"7b",
          3429 => x"27",
          3430 => x"05",
          3431 => x"70",
          3432 => x"08",
          3433 => x"88",
          3434 => x"55",
          3435 => x"80",
          3436 => x"70",
          3437 => x"07",
          3438 => x"70",
          3439 => x"56",
          3440 => x"27",
          3441 => x"75",
          3442 => x"13",
          3443 => x"75",
          3444 => x"85",
          3445 => x"83",
          3446 => x"33",
          3447 => x"ff",
          3448 => x"70",
          3449 => x"51",
          3450 => x"51",
          3451 => x"75",
          3452 => x"83",
          3453 => x"07",
          3454 => x"5a",
          3455 => x"84",
          3456 => x"53",
          3457 => x"14",
          3458 => x"70",
          3459 => x"07",
          3460 => x"74",
          3461 => x"88",
          3462 => x"52",
          3463 => x"06",
          3464 => x"d4",
          3465 => x"81",
          3466 => x"19",
          3467 => x"8b",
          3468 => x"58",
          3469 => x"34",
          3470 => x"08",
          3471 => x"33",
          3472 => x"70",
          3473 => x"86",
          3474 => x"b8",
          3475 => x"85",
          3476 => x"2b",
          3477 => x"52",
          3478 => x"34",
          3479 => x"78",
          3480 => x"71",
          3481 => x"5c",
          3482 => x"85",
          3483 => x"84",
          3484 => x"8b",
          3485 => x"15",
          3486 => x"07",
          3487 => x"33",
          3488 => x"5a",
          3489 => x"12",
          3490 => x"d4",
          3491 => x"12",
          3492 => x"07",
          3493 => x"33",
          3494 => x"58",
          3495 => x"70",
          3496 => x"84",
          3497 => x"12",
          3498 => x"ff",
          3499 => x"57",
          3500 => x"84",
          3501 => x"fe",
          3502 => x"b8",
          3503 => x"a0",
          3504 => x"84",
          3505 => x"77",
          3506 => x"08",
          3507 => x"04",
          3508 => x"0c",
          3509 => x"82",
          3510 => x"f4",
          3511 => x"d4",
          3512 => x"81",
          3513 => x"76",
          3514 => x"34",
          3515 => x"17",
          3516 => x"b8",
          3517 => x"05",
          3518 => x"ff",
          3519 => x"56",
          3520 => x"34",
          3521 => x"10",
          3522 => x"55",
          3523 => x"83",
          3524 => x"fe",
          3525 => x"0d",
          3526 => x"b8",
          3527 => x"2e",
          3528 => x"af",
          3529 => x"81",
          3530 => x"fb",
          3531 => x"ff",
          3532 => x"ff",
          3533 => x"83",
          3534 => x"11",
          3535 => x"2b",
          3536 => x"ff",
          3537 => x"73",
          3538 => x"12",
          3539 => x"2b",
          3540 => x"44",
          3541 => x"52",
          3542 => x"fd",
          3543 => x"71",
          3544 => x"19",
          3545 => x"2b",
          3546 => x"56",
          3547 => x"38",
          3548 => x"1b",
          3549 => x"60",
          3550 => x"58",
          3551 => x"18",
          3552 => x"76",
          3553 => x"8b",
          3554 => x"70",
          3555 => x"71",
          3556 => x"53",
          3557 => x"ba",
          3558 => x"12",
          3559 => x"07",
          3560 => x"33",
          3561 => x"7e",
          3562 => x"71",
          3563 => x"57",
          3564 => x"59",
          3565 => x"1d",
          3566 => x"84",
          3567 => x"2b",
          3568 => x"14",
          3569 => x"07",
          3570 => x"40",
          3571 => x"7b",
          3572 => x"16",
          3573 => x"2b",
          3574 => x"2a",
          3575 => x"79",
          3576 => x"70",
          3577 => x"71",
          3578 => x"05",
          3579 => x"2b",
          3580 => x"5d",
          3581 => x"75",
          3582 => x"70",
          3583 => x"8b",
          3584 => x"82",
          3585 => x"2b",
          3586 => x"5d",
          3587 => x"34",
          3588 => x"08",
          3589 => x"33",
          3590 => x"56",
          3591 => x"7e",
          3592 => x"3f",
          3593 => x"61",
          3594 => x"06",
          3595 => x"b6",
          3596 => x"0c",
          3597 => x"0b",
          3598 => x"84",
          3599 => x"60",
          3600 => x"f9",
          3601 => x"7e",
          3602 => x"b8",
          3603 => x"81",
          3604 => x"08",
          3605 => x"87",
          3606 => x"b8",
          3607 => x"07",
          3608 => x"2a",
          3609 => x"34",
          3610 => x"22",
          3611 => x"08",
          3612 => x"15",
          3613 => x"b8",
          3614 => x"76",
          3615 => x"7f",
          3616 => x"f4",
          3617 => x"b8",
          3618 => x"1c",
          3619 => x"71",
          3620 => x"81",
          3621 => x"ff",
          3622 => x"5b",
          3623 => x"1c",
          3624 => x"7c",
          3625 => x"34",
          3626 => x"08",
          3627 => x"71",
          3628 => x"ff",
          3629 => x"ff",
          3630 => x"57",
          3631 => x"34",
          3632 => x"83",
          3633 => x"5b",
          3634 => x"61",
          3635 => x"51",
          3636 => x"39",
          3637 => x"06",
          3638 => x"ff",
          3639 => x"ff",
          3640 => x"71",
          3641 => x"1b",
          3642 => x"2b",
          3643 => x"54",
          3644 => x"f9",
          3645 => x"24",
          3646 => x"8f",
          3647 => x"61",
          3648 => x"39",
          3649 => x"0c",
          3650 => x"82",
          3651 => x"f4",
          3652 => x"d4",
          3653 => x"81",
          3654 => x"7e",
          3655 => x"34",
          3656 => x"19",
          3657 => x"b8",
          3658 => x"05",
          3659 => x"ff",
          3660 => x"44",
          3661 => x"89",
          3662 => x"10",
          3663 => x"f8",
          3664 => x"34",
          3665 => x"39",
          3666 => x"83",
          3667 => x"fb",
          3668 => x"2e",
          3669 => x"3f",
          3670 => x"95",
          3671 => x"33",
          3672 => x"83",
          3673 => x"87",
          3674 => x"2b",
          3675 => x"15",
          3676 => x"2a",
          3677 => x"53",
          3678 => x"34",
          3679 => x"d4",
          3680 => x"12",
          3681 => x"07",
          3682 => x"33",
          3683 => x"5b",
          3684 => x"73",
          3685 => x"05",
          3686 => x"33",
          3687 => x"81",
          3688 => x"5c",
          3689 => x"1e",
          3690 => x"82",
          3691 => x"2b",
          3692 => x"33",
          3693 => x"70",
          3694 => x"57",
          3695 => x"1d",
          3696 => x"70",
          3697 => x"71",
          3698 => x"33",
          3699 => x"70",
          3700 => x"5c",
          3701 => x"83",
          3702 => x"1f",
          3703 => x"88",
          3704 => x"83",
          3705 => x"84",
          3706 => x"b8",
          3707 => x"ff",
          3708 => x"84",
          3709 => x"a0",
          3710 => x"80",
          3711 => x"51",
          3712 => x"08",
          3713 => x"17",
          3714 => x"84",
          3715 => x"84",
          3716 => x"34",
          3717 => x"d4",
          3718 => x"fe",
          3719 => x"06",
          3720 => x"61",
          3721 => x"84",
          3722 => x"84",
          3723 => x"5d",
          3724 => x"1c",
          3725 => x"54",
          3726 => x"1a",
          3727 => x"07",
          3728 => x"33",
          3729 => x"5c",
          3730 => x"84",
          3731 => x"84",
          3732 => x"33",
          3733 => x"83",
          3734 => x"87",
          3735 => x"88",
          3736 => x"59",
          3737 => x"64",
          3738 => x"1d",
          3739 => x"2b",
          3740 => x"2a",
          3741 => x"7f",
          3742 => x"70",
          3743 => x"8b",
          3744 => x"70",
          3745 => x"07",
          3746 => x"77",
          3747 => x"5a",
          3748 => x"17",
          3749 => x"d4",
          3750 => x"33",
          3751 => x"74",
          3752 => x"88",
          3753 => x"88",
          3754 => x"41",
          3755 => x"05",
          3756 => x"fa",
          3757 => x"33",
          3758 => x"79",
          3759 => x"71",
          3760 => x"5e",
          3761 => x"34",
          3762 => x"08",
          3763 => x"33",
          3764 => x"74",
          3765 => x"71",
          3766 => x"56",
          3767 => x"60",
          3768 => x"34",
          3769 => x"81",
          3770 => x"ff",
          3771 => x"58",
          3772 => x"34",
          3773 => x"33",
          3774 => x"83",
          3775 => x"12",
          3776 => x"2b",
          3777 => x"88",
          3778 => x"42",
          3779 => x"83",
          3780 => x"1f",
          3781 => x"2b",
          3782 => x"33",
          3783 => x"81",
          3784 => x"54",
          3785 => x"7c",
          3786 => x"d4",
          3787 => x"12",
          3788 => x"07",
          3789 => x"33",
          3790 => x"78",
          3791 => x"71",
          3792 => x"57",
          3793 => x"5a",
          3794 => x"85",
          3795 => x"17",
          3796 => x"8b",
          3797 => x"86",
          3798 => x"2b",
          3799 => x"52",
          3800 => x"34",
          3801 => x"08",
          3802 => x"88",
          3803 => x"88",
          3804 => x"34",
          3805 => x"08",
          3806 => x"33",
          3807 => x"74",
          3808 => x"88",
          3809 => x"45",
          3810 => x"34",
          3811 => x"08",
          3812 => x"71",
          3813 => x"05",
          3814 => x"88",
          3815 => x"45",
          3816 => x"1a",
          3817 => x"d4",
          3818 => x"12",
          3819 => x"62",
          3820 => x"5d",
          3821 => x"d4",
          3822 => x"05",
          3823 => x"ff",
          3824 => x"86",
          3825 => x"2b",
          3826 => x"1c",
          3827 => x"07",
          3828 => x"41",
          3829 => x"61",
          3830 => x"70",
          3831 => x"71",
          3832 => x"05",
          3833 => x"88",
          3834 => x"5f",
          3835 => x"86",
          3836 => x"84",
          3837 => x"12",
          3838 => x"ff",
          3839 => x"55",
          3840 => x"84",
          3841 => x"81",
          3842 => x"2b",
          3843 => x"33",
          3844 => x"8f",
          3845 => x"2a",
          3846 => x"58",
          3847 => x"1e",
          3848 => x"70",
          3849 => x"71",
          3850 => x"81",
          3851 => x"ff",
          3852 => x"49",
          3853 => x"34",
          3854 => x"ff",
          3855 => x"52",
          3856 => x"08",
          3857 => x"93",
          3858 => x"e4",
          3859 => x"51",
          3860 => x"27",
          3861 => x"3d",
          3862 => x"08",
          3863 => x"77",
          3864 => x"e4",
          3865 => x"e4",
          3866 => x"84",
          3867 => x"77",
          3868 => x"51",
          3869 => x"e4",
          3870 => x"f4",
          3871 => x"0b",
          3872 => x"53",
          3873 => x"b6",
          3874 => x"76",
          3875 => x"84",
          3876 => x"34",
          3877 => x"d4",
          3878 => x"0b",
          3879 => x"84",
          3880 => x"80",
          3881 => x"88",
          3882 => x"17",
          3883 => x"d0",
          3884 => x"d4",
          3885 => x"82",
          3886 => x"77",
          3887 => x"fe",
          3888 => x"05",
          3889 => x"87",
          3890 => x"71",
          3891 => x"04",
          3892 => x"52",
          3893 => x"71",
          3894 => x"08",
          3895 => x"72",
          3896 => x"e0",
          3897 => x"0c",
          3898 => x"7c",
          3899 => x"33",
          3900 => x"74",
          3901 => x"33",
          3902 => x"73",
          3903 => x"c0",
          3904 => x"76",
          3905 => x"08",
          3906 => x"a7",
          3907 => x"73",
          3908 => x"74",
          3909 => x"2e",
          3910 => x"84",
          3911 => x"84",
          3912 => x"06",
          3913 => x"ac",
          3914 => x"7e",
          3915 => x"5a",
          3916 => x"26",
          3917 => x"54",
          3918 => x"bd",
          3919 => x"98",
          3920 => x"51",
          3921 => x"81",
          3922 => x"38",
          3923 => x"e2",
          3924 => x"fc",
          3925 => x"83",
          3926 => x"b8",
          3927 => x"80",
          3928 => x"5a",
          3929 => x"38",
          3930 => x"84",
          3931 => x"9f",
          3932 => x"71",
          3933 => x"12",
          3934 => x"53",
          3935 => x"98",
          3936 => x"96",
          3937 => x"83",
          3938 => x"b8",
          3939 => x"80",
          3940 => x"0c",
          3941 => x"0c",
          3942 => x"3d",
          3943 => x"92",
          3944 => x"71",
          3945 => x"51",
          3946 => x"98",
          3947 => x"c0",
          3948 => x"81",
          3949 => x"52",
          3950 => x"2e",
          3951 => x"54",
          3952 => x"3d",
          3953 => x"33",
          3954 => x"09",
          3955 => x"75",
          3956 => x"80",
          3957 => x"3f",
          3958 => x"38",
          3959 => x"8c",
          3960 => x"08",
          3961 => x"33",
          3962 => x"84",
          3963 => x"06",
          3964 => x"19",
          3965 => x"08",
          3966 => x"08",
          3967 => x"ff",
          3968 => x"82",
          3969 => x"81",
          3970 => x"18",
          3971 => x"33",
          3972 => x"06",
          3973 => x"76",
          3974 => x"38",
          3975 => x"57",
          3976 => x"ff",
          3977 => x"0b",
          3978 => x"84",
          3979 => x"80",
          3980 => x"0b",
          3981 => x"19",
          3982 => x"34",
          3983 => x"80",
          3984 => x"e1",
          3985 => x"08",
          3986 => x"88",
          3987 => x"74",
          3988 => x"34",
          3989 => x"19",
          3990 => x"a4",
          3991 => x"84",
          3992 => x"75",
          3993 => x"55",
          3994 => x"08",
          3995 => x"81",
          3996 => x"33",
          3997 => x"34",
          3998 => x"51",
          3999 => x"80",
          4000 => x"f3",
          4001 => x"56",
          4002 => x"17",
          4003 => x"77",
          4004 => x"04",
          4005 => x"2e",
          4006 => x"a5",
          4007 => x"dd",
          4008 => x"2a",
          4009 => x"5b",
          4010 => x"83",
          4011 => x"81",
          4012 => x"53",
          4013 => x"f8",
          4014 => x"2e",
          4015 => x"b4",
          4016 => x"83",
          4017 => x"1c",
          4018 => x"53",
          4019 => x"2e",
          4020 => x"71",
          4021 => x"81",
          4022 => x"53",
          4023 => x"f8",
          4024 => x"2e",
          4025 => x"b4",
          4026 => x"83",
          4027 => x"88",
          4028 => x"84",
          4029 => x"fe",
          4030 => x"b8",
          4031 => x"88",
          4032 => x"17",
          4033 => x"83",
          4034 => x"7b",
          4035 => x"81",
          4036 => x"17",
          4037 => x"e4",
          4038 => x"81",
          4039 => x"df",
          4040 => x"05",
          4041 => x"71",
          4042 => x"57",
          4043 => x"2e",
          4044 => x"87",
          4045 => x"17",
          4046 => x"83",
          4047 => x"7b",
          4048 => x"81",
          4049 => x"17",
          4050 => x"e4",
          4051 => x"81",
          4052 => x"f7",
          4053 => x"77",
          4054 => x"12",
          4055 => x"07",
          4056 => x"2b",
          4057 => x"80",
          4058 => x"5c",
          4059 => x"04",
          4060 => x"17",
          4061 => x"f6",
          4062 => x"08",
          4063 => x"38",
          4064 => x"b4",
          4065 => x"b8",
          4066 => x"08",
          4067 => x"55",
          4068 => x"f7",
          4069 => x"18",
          4070 => x"33",
          4071 => x"df",
          4072 => x"b8",
          4073 => x"5c",
          4074 => x"7b",
          4075 => x"84",
          4076 => x"17",
          4077 => x"a0",
          4078 => x"33",
          4079 => x"84",
          4080 => x"81",
          4081 => x"70",
          4082 => x"bb",
          4083 => x"7b",
          4084 => x"84",
          4085 => x"17",
          4086 => x"e4",
          4087 => x"27",
          4088 => x"74",
          4089 => x"38",
          4090 => x"08",
          4091 => x"51",
          4092 => x"39",
          4093 => x"17",
          4094 => x"f4",
          4095 => x"08",
          4096 => x"38",
          4097 => x"b4",
          4098 => x"b8",
          4099 => x"08",
          4100 => x"55",
          4101 => x"84",
          4102 => x"18",
          4103 => x"33",
          4104 => x"ec",
          4105 => x"18",
          4106 => x"33",
          4107 => x"81",
          4108 => x"39",
          4109 => x"57",
          4110 => x"38",
          4111 => x"78",
          4112 => x"74",
          4113 => x"2e",
          4114 => x"0c",
          4115 => x"a8",
          4116 => x"1a",
          4117 => x"b6",
          4118 => x"7c",
          4119 => x"38",
          4120 => x"81",
          4121 => x"b8",
          4122 => x"58",
          4123 => x"58",
          4124 => x"fe",
          4125 => x"06",
          4126 => x"88",
          4127 => x"0b",
          4128 => x"0c",
          4129 => x"09",
          4130 => x"2a",
          4131 => x"b4",
          4132 => x"85",
          4133 => x"5d",
          4134 => x"bd",
          4135 => x"52",
          4136 => x"84",
          4137 => x"ff",
          4138 => x"79",
          4139 => x"2b",
          4140 => x"83",
          4141 => x"06",
          4142 => x"5e",
          4143 => x"56",
          4144 => x"5a",
          4145 => x"5b",
          4146 => x"1a",
          4147 => x"16",
          4148 => x"b4",
          4149 => x"2e",
          4150 => x"71",
          4151 => x"81",
          4152 => x"53",
          4153 => x"f0",
          4154 => x"2e",
          4155 => x"b4",
          4156 => x"38",
          4157 => x"81",
          4158 => x"7a",
          4159 => x"84",
          4160 => x"06",
          4161 => x"81",
          4162 => x"a8",
          4163 => x"1a",
          4164 => x"dd",
          4165 => x"70",
          4166 => x"9b",
          4167 => x"7f",
          4168 => x"84",
          4169 => x"19",
          4170 => x"1b",
          4171 => x"56",
          4172 => x"19",
          4173 => x"38",
          4174 => x"19",
          4175 => x"e4",
          4176 => x"81",
          4177 => x"83",
          4178 => x"05",
          4179 => x"38",
          4180 => x"06",
          4181 => x"76",
          4182 => x"cb",
          4183 => x"70",
          4184 => x"8b",
          4185 => x"7c",
          4186 => x"84",
          4187 => x"19",
          4188 => x"1b",
          4189 => x"40",
          4190 => x"82",
          4191 => x"81",
          4192 => x"1e",
          4193 => x"ee",
          4194 => x"81",
          4195 => x"81",
          4196 => x"81",
          4197 => x"09",
          4198 => x"e4",
          4199 => x"70",
          4200 => x"84",
          4201 => x"74",
          4202 => x"33",
          4203 => x"fc",
          4204 => x"76",
          4205 => x"3f",
          4206 => x"76",
          4207 => x"33",
          4208 => x"84",
          4209 => x"06",
          4210 => x"83",
          4211 => x"1b",
          4212 => x"e4",
          4213 => x"27",
          4214 => x"74",
          4215 => x"38",
          4216 => x"81",
          4217 => x"5a",
          4218 => x"53",
          4219 => x"f3",
          4220 => x"76",
          4221 => x"83",
          4222 => x"b8",
          4223 => x"b9",
          4224 => x"fd",
          4225 => x"fc",
          4226 => x"33",
          4227 => x"f0",
          4228 => x"58",
          4229 => x"75",
          4230 => x"79",
          4231 => x"7a",
          4232 => x"3d",
          4233 => x"5a",
          4234 => x"57",
          4235 => x"9c",
          4236 => x"19",
          4237 => x"80",
          4238 => x"38",
          4239 => x"08",
          4240 => x"77",
          4241 => x"51",
          4242 => x"80",
          4243 => x"b8",
          4244 => x"b8",
          4245 => x"07",
          4246 => x"55",
          4247 => x"2e",
          4248 => x"55",
          4249 => x"0d",
          4250 => x"b8",
          4251 => x"79",
          4252 => x"84",
          4253 => x"b8",
          4254 => x"ff",
          4255 => x"b8",
          4256 => x"fe",
          4257 => x"08",
          4258 => x"52",
          4259 => x"84",
          4260 => x"38",
          4261 => x"70",
          4262 => x"84",
          4263 => x"55",
          4264 => x"08",
          4265 => x"54",
          4266 => x"9c",
          4267 => x"70",
          4268 => x"2e",
          4269 => x"78",
          4270 => x"08",
          4271 => x"b8",
          4272 => x"55",
          4273 => x"38",
          4274 => x"fe",
          4275 => x"78",
          4276 => x"0c",
          4277 => x"84",
          4278 => x"e4",
          4279 => x"84",
          4280 => x"84",
          4281 => x"73",
          4282 => x"7a",
          4283 => x"b8",
          4284 => x"b8",
          4285 => x"3d",
          4286 => x"ff",
          4287 => x"f8",
          4288 => x"55",
          4289 => x"df",
          4290 => x"d7",
          4291 => x"08",
          4292 => x"56",
          4293 => x"85",
          4294 => x"5a",
          4295 => x"17",
          4296 => x"0c",
          4297 => x"80",
          4298 => x"98",
          4299 => x"b8",
          4300 => x"84",
          4301 => x"82",
          4302 => x"0d",
          4303 => x"2e",
          4304 => x"89",
          4305 => x"38",
          4306 => x"14",
          4307 => x"8d",
          4308 => x"b0",
          4309 => x"19",
          4310 => x"51",
          4311 => x"55",
          4312 => x"38",
          4313 => x"ff",
          4314 => x"b8",
          4315 => x"73",
          4316 => x"38",
          4317 => x"e4",
          4318 => x"0d",
          4319 => x"05",
          4320 => x"27",
          4321 => x"98",
          4322 => x"2e",
          4323 => x"7a",
          4324 => x"57",
          4325 => x"88",
          4326 => x"81",
          4327 => x"90",
          4328 => x"18",
          4329 => x"0c",
          4330 => x"0c",
          4331 => x"2a",
          4332 => x"76",
          4333 => x"08",
          4334 => x"e4",
          4335 => x"b8",
          4336 => x"19",
          4337 => x"91",
          4338 => x"94",
          4339 => x"3f",
          4340 => x"84",
          4341 => x"38",
          4342 => x"2e",
          4343 => x"e4",
          4344 => x"b8",
          4345 => x"7d",
          4346 => x"08",
          4347 => x"78",
          4348 => x"71",
          4349 => x"7b",
          4350 => x"80",
          4351 => x"05",
          4352 => x"38",
          4353 => x"75",
          4354 => x"1c",
          4355 => x"e4",
          4356 => x"e7",
          4357 => x"98",
          4358 => x"0c",
          4359 => x"19",
          4360 => x"1a",
          4361 => x"b8",
          4362 => x"e4",
          4363 => x"a8",
          4364 => x"08",
          4365 => x"5c",
          4366 => x"db",
          4367 => x"1a",
          4368 => x"33",
          4369 => x"8a",
          4370 => x"06",
          4371 => x"a7",
          4372 => x"9c",
          4373 => x"58",
          4374 => x"19",
          4375 => x"05",
          4376 => x"81",
          4377 => x"0d",
          4378 => x"5c",
          4379 => x"70",
          4380 => x"80",
          4381 => x"75",
          4382 => x"2e",
          4383 => x"58",
          4384 => x"81",
          4385 => x"19",
          4386 => x"3f",
          4387 => x"38",
          4388 => x"0c",
          4389 => x"1c",
          4390 => x"2e",
          4391 => x"06",
          4392 => x"86",
          4393 => x"30",
          4394 => x"25",
          4395 => x"57",
          4396 => x"06",
          4397 => x"38",
          4398 => x"ff",
          4399 => x"3f",
          4400 => x"e4",
          4401 => x"56",
          4402 => x"e4",
          4403 => x"b4",
          4404 => x"33",
          4405 => x"b8",
          4406 => x"fe",
          4407 => x"1a",
          4408 => x"31",
          4409 => x"a0",
          4410 => x"19",
          4411 => x"06",
          4412 => x"08",
          4413 => x"81",
          4414 => x"57",
          4415 => x"81",
          4416 => x"81",
          4417 => x"8d",
          4418 => x"90",
          4419 => x"5e",
          4420 => x"ff",
          4421 => x"56",
          4422 => x"be",
          4423 => x"98",
          4424 => x"94",
          4425 => x"39",
          4426 => x"09",
          4427 => x"9b",
          4428 => x"2b",
          4429 => x"38",
          4430 => x"29",
          4431 => x"5b",
          4432 => x"81",
          4433 => x"07",
          4434 => x"c5",
          4435 => x"38",
          4436 => x"75",
          4437 => x"57",
          4438 => x"70",
          4439 => x"80",
          4440 => x"fe",
          4441 => x"80",
          4442 => x"06",
          4443 => x"ff",
          4444 => x"fe",
          4445 => x"8b",
          4446 => x"29",
          4447 => x"40",
          4448 => x"19",
          4449 => x"7e",
          4450 => x"1d",
          4451 => x"3d",
          4452 => x"08",
          4453 => x"cf",
          4454 => x"b8",
          4455 => x"70",
          4456 => x"b8",
          4457 => x"58",
          4458 => x"38",
          4459 => x"78",
          4460 => x"81",
          4461 => x"1b",
          4462 => x"e4",
          4463 => x"81",
          4464 => x"76",
          4465 => x"33",
          4466 => x"38",
          4467 => x"ff",
          4468 => x"76",
          4469 => x"83",
          4470 => x"81",
          4471 => x"8f",
          4472 => x"78",
          4473 => x"2a",
          4474 => x"81",
          4475 => x"81",
          4476 => x"76",
          4477 => x"38",
          4478 => x"a7",
          4479 => x"78",
          4480 => x"81",
          4481 => x"1a",
          4482 => x"81",
          4483 => x"81",
          4484 => x"80",
          4485 => x"b8",
          4486 => x"80",
          4487 => x"e4",
          4488 => x"b4",
          4489 => x"33",
          4490 => x"b8",
          4491 => x"fe",
          4492 => x"1c",
          4493 => x"31",
          4494 => x"a0",
          4495 => x"1b",
          4496 => x"06",
          4497 => x"08",
          4498 => x"81",
          4499 => x"57",
          4500 => x"39",
          4501 => x"06",
          4502 => x"86",
          4503 => x"93",
          4504 => x"06",
          4505 => x"0c",
          4506 => x"38",
          4507 => x"7b",
          4508 => x"08",
          4509 => x"fc",
          4510 => x"2e",
          4511 => x"0b",
          4512 => x"19",
          4513 => x"06",
          4514 => x"33",
          4515 => x"59",
          4516 => x"33",
          4517 => x"5b",
          4518 => x"e4",
          4519 => x"71",
          4520 => x"57",
          4521 => x"81",
          4522 => x"81",
          4523 => x"7a",
          4524 => x"81",
          4525 => x"75",
          4526 => x"06",
          4527 => x"58",
          4528 => x"33",
          4529 => x"75",
          4530 => x"8d",
          4531 => x"41",
          4532 => x"70",
          4533 => x"39",
          4534 => x"3d",
          4535 => x"ff",
          4536 => x"39",
          4537 => x"ab",
          4538 => x"5d",
          4539 => x"74",
          4540 => x"5d",
          4541 => x"70",
          4542 => x"74",
          4543 => x"40",
          4544 => x"70",
          4545 => x"05",
          4546 => x"38",
          4547 => x"06",
          4548 => x"38",
          4549 => x"0b",
          4550 => x"7b",
          4551 => x"55",
          4552 => x"70",
          4553 => x"74",
          4554 => x"38",
          4555 => x"2e",
          4556 => x"8f",
          4557 => x"76",
          4558 => x"72",
          4559 => x"57",
          4560 => x"a0",
          4561 => x"80",
          4562 => x"ca",
          4563 => x"05",
          4564 => x"55",
          4565 => x"55",
          4566 => x"78",
          4567 => x"38",
          4568 => x"76",
          4569 => x"38",
          4570 => x"38",
          4571 => x"a2",
          4572 => x"74",
          4573 => x"81",
          4574 => x"8e",
          4575 => x"81",
          4576 => x"77",
          4577 => x"7d",
          4578 => x"08",
          4579 => x"7b",
          4580 => x"80",
          4581 => x"e4",
          4582 => x"2e",
          4583 => x"80",
          4584 => x"08",
          4585 => x"57",
          4586 => x"81",
          4587 => x"52",
          4588 => x"84",
          4589 => x"7d",
          4590 => x"08",
          4591 => x"38",
          4592 => x"59",
          4593 => x"18",
          4594 => x"18",
          4595 => x"06",
          4596 => x"b8",
          4597 => x"a4",
          4598 => x"85",
          4599 => x"19",
          4600 => x"1e",
          4601 => x"e5",
          4602 => x"80",
          4603 => x"2e",
          4604 => x"7b",
          4605 => x"51",
          4606 => x"56",
          4607 => x"88",
          4608 => x"89",
          4609 => x"ff",
          4610 => x"1e",
          4611 => x"af",
          4612 => x"7f",
          4613 => x"b8",
          4614 => x"9c",
          4615 => x"85",
          4616 => x"1d",
          4617 => x"a0",
          4618 => x"76",
          4619 => x"55",
          4620 => x"08",
          4621 => x"05",
          4622 => x"34",
          4623 => x"1e",
          4624 => x"5a",
          4625 => x"1d",
          4626 => x"0c",
          4627 => x"70",
          4628 => x"74",
          4629 => x"7d",
          4630 => x"08",
          4631 => x"fd",
          4632 => x"b4",
          4633 => x"33",
          4634 => x"08",
          4635 => x"38",
          4636 => x"b4",
          4637 => x"74",
          4638 => x"18",
          4639 => x"38",
          4640 => x"39",
          4641 => x"31",
          4642 => x"84",
          4643 => x"08",
          4644 => x"08",
          4645 => x"75",
          4646 => x"05",
          4647 => x"ff",
          4648 => x"e4",
          4649 => x"43",
          4650 => x"b4",
          4651 => x"1c",
          4652 => x"06",
          4653 => x"b8",
          4654 => x"dc",
          4655 => x"85",
          4656 => x"1d",
          4657 => x"8c",
          4658 => x"ff",
          4659 => x"34",
          4660 => x"1c",
          4661 => x"1c",
          4662 => x"77",
          4663 => x"2e",
          4664 => x"81",
          4665 => x"18",
          4666 => x"81",
          4667 => x"75",
          4668 => x"ff",
          4669 => x"cb",
          4670 => x"b3",
          4671 => x"58",
          4672 => x"7b",
          4673 => x"52",
          4674 => x"e4",
          4675 => x"f1",
          4676 => x"a9",
          4677 => x"1c",
          4678 => x"1d",
          4679 => x"56",
          4680 => x"84",
          4681 => x"1c",
          4682 => x"e4",
          4683 => x"27",
          4684 => x"61",
          4685 => x"38",
          4686 => x"08",
          4687 => x"51",
          4688 => x"39",
          4689 => x"43",
          4690 => x"06",
          4691 => x"70",
          4692 => x"38",
          4693 => x"5d",
          4694 => x"08",
          4695 => x"cf",
          4696 => x"2e",
          4697 => x"e4",
          4698 => x"a8",
          4699 => x"08",
          4700 => x"7e",
          4701 => x"08",
          4702 => x"41",
          4703 => x"fc",
          4704 => x"39",
          4705 => x"fc",
          4706 => x"b4",
          4707 => x"61",
          4708 => x"3f",
          4709 => x"08",
          4710 => x"81",
          4711 => x"e3",
          4712 => x"08",
          4713 => x"34",
          4714 => x"38",
          4715 => x"38",
          4716 => x"70",
          4717 => x"78",
          4718 => x"70",
          4719 => x"82",
          4720 => x"83",
          4721 => x"ff",
          4722 => x"76",
          4723 => x"79",
          4724 => x"70",
          4725 => x"18",
          4726 => x"34",
          4727 => x"9c",
          4728 => x"58",
          4729 => x"74",
          4730 => x"32",
          4731 => x"55",
          4732 => x"72",
          4733 => x"81",
          4734 => x"77",
          4735 => x"58",
          4736 => x"18",
          4737 => x"34",
          4738 => x"77",
          4739 => x"34",
          4740 => x"80",
          4741 => x"8c",
          4742 => x"73",
          4743 => x"8b",
          4744 => x"08",
          4745 => x"33",
          4746 => x"81",
          4747 => x"75",
          4748 => x"16",
          4749 => x"07",
          4750 => x"55",
          4751 => x"98",
          4752 => x"54",
          4753 => x"04",
          4754 => x"1d",
          4755 => x"5b",
          4756 => x"74",
          4757 => x"b8",
          4758 => x"81",
          4759 => x"27",
          4760 => x"73",
          4761 => x"78",
          4762 => x"56",
          4763 => x"5c",
          4764 => x"ba",
          4765 => x"07",
          4766 => x"55",
          4767 => x"34",
          4768 => x"1f",
          4769 => x"89",
          4770 => x"2e",
          4771 => x"57",
          4772 => x"11",
          4773 => x"9c",
          4774 => x"88",
          4775 => x"53",
          4776 => x"8a",
          4777 => x"06",
          4778 => x"5a",
          4779 => x"71",
          4780 => x"56",
          4781 => x"72",
          4782 => x"30",
          4783 => x"53",
          4784 => x"3d",
          4785 => x"5c",
          4786 => x"74",
          4787 => x"80",
          4788 => x"2e",
          4789 => x"1d",
          4790 => x"41",
          4791 => x"38",
          4792 => x"57",
          4793 => x"55",
          4794 => x"0c",
          4795 => x"ff",
          4796 => x"18",
          4797 => x"73",
          4798 => x"70",
          4799 => x"07",
          4800 => x"38",
          4801 => x"74",
          4802 => x"80",
          4803 => x"ff",
          4804 => x"81",
          4805 => x"81",
          4806 => x"56",
          4807 => x"ff",
          4808 => x"81",
          4809 => x"18",
          4810 => x"70",
          4811 => x"57",
          4812 => x"cb",
          4813 => x"30",
          4814 => x"58",
          4815 => x"14",
          4816 => x"55",
          4817 => x"dc",
          4818 => x"07",
          4819 => x"88",
          4820 => x"3d",
          4821 => x"90",
          4822 => x"51",
          4823 => x"08",
          4824 => x"8d",
          4825 => x"0c",
          4826 => x"33",
          4827 => x"80",
          4828 => x"80",
          4829 => x"51",
          4830 => x"84",
          4831 => x"81",
          4832 => x"80",
          4833 => x"7d",
          4834 => x"80",
          4835 => x"af",
          4836 => x"70",
          4837 => x"54",
          4838 => x"9f",
          4839 => x"2e",
          4840 => x"d1",
          4841 => x"a7",
          4842 => x"70",
          4843 => x"9f",
          4844 => x"7c",
          4845 => x"ff",
          4846 => x"77",
          4847 => x"2e",
          4848 => x"83",
          4849 => x"56",
          4850 => x"83",
          4851 => x"82",
          4852 => x"77",
          4853 => x"78",
          4854 => x"fe",
          4855 => x"2e",
          4856 => x"54",
          4857 => x"38",
          4858 => x"74",
          4859 => x"53",
          4860 => x"88",
          4861 => x"57",
          4862 => x"38",
          4863 => x"ae",
          4864 => x"5a",
          4865 => x"72",
          4866 => x"26",
          4867 => x"70",
          4868 => x"7c",
          4869 => x"2e",
          4870 => x"83",
          4871 => x"83",
          4872 => x"76",
          4873 => x"81",
          4874 => x"77",
          4875 => x"53",
          4876 => x"57",
          4877 => x"7c",
          4878 => x"06",
          4879 => x"7d",
          4880 => x"e3",
          4881 => x"75",
          4882 => x"80",
          4883 => x"7d",
          4884 => x"2e",
          4885 => x"ab",
          4886 => x"84",
          4887 => x"54",
          4888 => x"ac",
          4889 => x"09",
          4890 => x"2a",
          4891 => x"f0",
          4892 => x"78",
          4893 => x"56",
          4894 => x"57",
          4895 => x"79",
          4896 => x"7c",
          4897 => x"fd",
          4898 => x"8a",
          4899 => x"2e",
          4900 => x"22",
          4901 => x"fc",
          4902 => x"7b",
          4903 => x"ae",
          4904 => x"54",
          4905 => x"81",
          4906 => x"79",
          4907 => x"7b",
          4908 => x"08",
          4909 => x"e4",
          4910 => x"81",
          4911 => x"1c",
          4912 => x"5d",
          4913 => x"1c",
          4914 => x"d3",
          4915 => x"88",
          4916 => x"54",
          4917 => x"88",
          4918 => x"fe",
          4919 => x"2e",
          4920 => x"fb",
          4921 => x"07",
          4922 => x"7d",
          4923 => x"06",
          4924 => x"06",
          4925 => x"fd",
          4926 => x"7c",
          4927 => x"38",
          4928 => x"34",
          4929 => x"3d",
          4930 => x"38",
          4931 => x"ff",
          4932 => x"38",
          4933 => x"5c",
          4934 => x"5a",
          4935 => x"f6",
          4936 => x"ff",
          4937 => x"55",
          4938 => x"ff",
          4939 => x"54",
          4940 => x"74",
          4941 => x"8c",
          4942 => x"ff",
          4943 => x"80",
          4944 => x"81",
          4945 => x"56",
          4946 => x"ff",
          4947 => x"bf",
          4948 => x"7d",
          4949 => x"53",
          4950 => x"93",
          4951 => x"06",
          4952 => x"58",
          4953 => x"59",
          4954 => x"16",
          4955 => x"b3",
          4956 => x"ff",
          4957 => x"ae",
          4958 => x"1d",
          4959 => x"34",
          4960 => x"14",
          4961 => x"2b",
          4962 => x"1f",
          4963 => x"1b",
          4964 => x"72",
          4965 => x"05",
          4966 => x"5b",
          4967 => x"1d",
          4968 => x"09",
          4969 => x"39",
          4970 => x"f6",
          4971 => x"0c",
          4972 => x"67",
          4973 => x"33",
          4974 => x"7e",
          4975 => x"2e",
          4976 => x"5b",
          4977 => x"ba",
          4978 => x"75",
          4979 => x"c0",
          4980 => x"38",
          4981 => x"70",
          4982 => x"2e",
          4983 => x"81",
          4984 => x"80",
          4985 => x"ff",
          4986 => x"81",
          4987 => x"7c",
          4988 => x"34",
          4989 => x"33",
          4990 => x"33",
          4991 => x"e4",
          4992 => x"41",
          4993 => x"78",
          4994 => x"81",
          4995 => x"38",
          4996 => x"0b",
          4997 => x"81",
          4998 => x"81",
          4999 => x"3f",
          5000 => x"38",
          5001 => x"0c",
          5002 => x"17",
          5003 => x"2b",
          5004 => x"d4",
          5005 => x"26",
          5006 => x"42",
          5007 => x"84",
          5008 => x"81",
          5009 => x"33",
          5010 => x"07",
          5011 => x"81",
          5012 => x"33",
          5013 => x"07",
          5014 => x"17",
          5015 => x"90",
          5016 => x"33",
          5017 => x"71",
          5018 => x"56",
          5019 => x"33",
          5020 => x"ff",
          5021 => x"59",
          5022 => x"38",
          5023 => x"80",
          5024 => x"8a",
          5025 => x"87",
          5026 => x"61",
          5027 => x"80",
          5028 => x"56",
          5029 => x"8f",
          5030 => x"98",
          5031 => x"18",
          5032 => x"74",
          5033 => x"33",
          5034 => x"88",
          5035 => x"07",
          5036 => x"44",
          5037 => x"17",
          5038 => x"2b",
          5039 => x"2e",
          5040 => x"2a",
          5041 => x"38",
          5042 => x"ee",
          5043 => x"84",
          5044 => x"38",
          5045 => x"ff",
          5046 => x"83",
          5047 => x"75",
          5048 => x"5d",
          5049 => x"a4",
          5050 => x"0c",
          5051 => x"7c",
          5052 => x"22",
          5053 => x"e0",
          5054 => x"19",
          5055 => x"10",
          5056 => x"05",
          5057 => x"59",
          5058 => x"b8",
          5059 => x"0b",
          5060 => x"18",
          5061 => x"7c",
          5062 => x"05",
          5063 => x"86",
          5064 => x"18",
          5065 => x"58",
          5066 => x"0d",
          5067 => x"97",
          5068 => x"70",
          5069 => x"89",
          5070 => x"ff",
          5071 => x"2e",
          5072 => x"e4",
          5073 => x"5a",
          5074 => x"79",
          5075 => x"12",
          5076 => x"38",
          5077 => x"55",
          5078 => x"89",
          5079 => x"58",
          5080 => x"55",
          5081 => x"38",
          5082 => x"70",
          5083 => x"07",
          5084 => x"98",
          5085 => x"83",
          5086 => x"f9",
          5087 => x"38",
          5088 => x"58",
          5089 => x"c0",
          5090 => x"81",
          5091 => x"81",
          5092 => x"70",
          5093 => x"77",
          5094 => x"83",
          5095 => x"83",
          5096 => x"5b",
          5097 => x"16",
          5098 => x"2b",
          5099 => x"33",
          5100 => x"1b",
          5101 => x"40",
          5102 => x"0c",
          5103 => x"80",
          5104 => x"1d",
          5105 => x"71",
          5106 => x"f0",
          5107 => x"43",
          5108 => x"7a",
          5109 => x"83",
          5110 => x"7a",
          5111 => x"38",
          5112 => x"81",
          5113 => x"84",
          5114 => x"ff",
          5115 => x"84",
          5116 => x"7f",
          5117 => x"83",
          5118 => x"81",
          5119 => x"33",
          5120 => x"b7",
          5121 => x"70",
          5122 => x"7f",
          5123 => x"38",
          5124 => x"80",
          5125 => x"58",
          5126 => x"38",
          5127 => x"38",
          5128 => x"1a",
          5129 => x"fe",
          5130 => x"80",
          5131 => x"58",
          5132 => x"70",
          5133 => x"ff",
          5134 => x"2e",
          5135 => x"38",
          5136 => x"98",
          5137 => x"5d",
          5138 => x"71",
          5139 => x"40",
          5140 => x"80",
          5141 => x"39",
          5142 => x"84",
          5143 => x"75",
          5144 => x"85",
          5145 => x"40",
          5146 => x"84",
          5147 => x"83",
          5148 => x"5c",
          5149 => x"33",
          5150 => x"71",
          5151 => x"77",
          5152 => x"2e",
          5153 => x"83",
          5154 => x"81",
          5155 => x"5c",
          5156 => x"58",
          5157 => x"38",
          5158 => x"77",
          5159 => x"81",
          5160 => x"33",
          5161 => x"07",
          5162 => x"06",
          5163 => x"5a",
          5164 => x"83",
          5165 => x"81",
          5166 => x"53",
          5167 => x"ff",
          5168 => x"80",
          5169 => x"77",
          5170 => x"79",
          5171 => x"84",
          5172 => x"57",
          5173 => x"81",
          5174 => x"11",
          5175 => x"71",
          5176 => x"72",
          5177 => x"5e",
          5178 => x"84",
          5179 => x"06",
          5180 => x"11",
          5181 => x"71",
          5182 => x"72",
          5183 => x"47",
          5184 => x"86",
          5185 => x"06",
          5186 => x"11",
          5187 => x"71",
          5188 => x"72",
          5189 => x"94",
          5190 => x"11",
          5191 => x"71",
          5192 => x"72",
          5193 => x"62",
          5194 => x"5c",
          5195 => x"77",
          5196 => x"5d",
          5197 => x"18",
          5198 => x"0c",
          5199 => x"39",
          5200 => x"7a",
          5201 => x"54",
          5202 => x"53",
          5203 => x"b3",
          5204 => x"09",
          5205 => x"e4",
          5206 => x"a8",
          5207 => x"08",
          5208 => x"60",
          5209 => x"e4",
          5210 => x"74",
          5211 => x"81",
          5212 => x"58",
          5213 => x"80",
          5214 => x"5f",
          5215 => x"88",
          5216 => x"80",
          5217 => x"33",
          5218 => x"81",
          5219 => x"75",
          5220 => x"7d",
          5221 => x"40",
          5222 => x"2e",
          5223 => x"39",
          5224 => x"3d",
          5225 => x"39",
          5226 => x"bf",
          5227 => x"18",
          5228 => x"33",
          5229 => x"39",
          5230 => x"33",
          5231 => x"5d",
          5232 => x"80",
          5233 => x"33",
          5234 => x"2e",
          5235 => x"ba",
          5236 => x"33",
          5237 => x"73",
          5238 => x"08",
          5239 => x"80",
          5240 => x"86",
          5241 => x"75",
          5242 => x"38",
          5243 => x"05",
          5244 => x"08",
          5245 => x"3d",
          5246 => x"0c",
          5247 => x"11",
          5248 => x"73",
          5249 => x"81",
          5250 => x"79",
          5251 => x"83",
          5252 => x"7e",
          5253 => x"33",
          5254 => x"9f",
          5255 => x"89",
          5256 => x"56",
          5257 => x"26",
          5258 => x"06",
          5259 => x"58",
          5260 => x"85",
          5261 => x"32",
          5262 => x"79",
          5263 => x"92",
          5264 => x"83",
          5265 => x"fe",
          5266 => x"7a",
          5267 => x"e6",
          5268 => x"fb",
          5269 => x"80",
          5270 => x"54",
          5271 => x"84",
          5272 => x"b8",
          5273 => x"80",
          5274 => x"56",
          5275 => x"0d",
          5276 => x"70",
          5277 => x"e4",
          5278 => x"2e",
          5279 => x"7c",
          5280 => x"2e",
          5281 => x"ea",
          5282 => x"bb",
          5283 => x"7a",
          5284 => x"11",
          5285 => x"07",
          5286 => x"56",
          5287 => x"0b",
          5288 => x"34",
          5289 => x"0b",
          5290 => x"8b",
          5291 => x"0b",
          5292 => x"34",
          5293 => x"a9",
          5294 => x"34",
          5295 => x"9e",
          5296 => x"7e",
          5297 => x"80",
          5298 => x"08",
          5299 => x"81",
          5300 => x"7c",
          5301 => x"79",
          5302 => x"05",
          5303 => x"80",
          5304 => x"06",
          5305 => x"fe",
          5306 => x"70",
          5307 => x"82",
          5308 => x"5e",
          5309 => x"06",
          5310 => x"2a",
          5311 => x"38",
          5312 => x"11",
          5313 => x"0c",
          5314 => x"71",
          5315 => x"40",
          5316 => x"38",
          5317 => x"11",
          5318 => x"71",
          5319 => x"72",
          5320 => x"70",
          5321 => x"51",
          5322 => x"1a",
          5323 => x"34",
          5324 => x"9c",
          5325 => x"55",
          5326 => x"80",
          5327 => x"0c",
          5328 => x"52",
          5329 => x"80",
          5330 => x"92",
          5331 => x"7d",
          5332 => x"78",
          5333 => x"e4",
          5334 => x"26",
          5335 => x"08",
          5336 => x"31",
          5337 => x"33",
          5338 => x"82",
          5339 => x"fc",
          5340 => x"fb",
          5341 => x"fb",
          5342 => x"fb",
          5343 => x"84",
          5344 => x"57",
          5345 => x"7a",
          5346 => x"39",
          5347 => x"98",
          5348 => x"5d",
          5349 => x"7c",
          5350 => x"79",
          5351 => x"e4",
          5352 => x"2e",
          5353 => x"81",
          5354 => x"08",
          5355 => x"74",
          5356 => x"84",
          5357 => x"17",
          5358 => x"56",
          5359 => x"81",
          5360 => x"81",
          5361 => x"55",
          5362 => x"d9",
          5363 => x"0b",
          5364 => x"16",
          5365 => x"71",
          5366 => x"5b",
          5367 => x"8f",
          5368 => x"80",
          5369 => x"a0",
          5370 => x"5e",
          5371 => x"9b",
          5372 => x"2e",
          5373 => x"a9",
          5374 => x"57",
          5375 => x"38",
          5376 => x"09",
          5377 => x"53",
          5378 => x"ff",
          5379 => x"80",
          5380 => x"76",
          5381 => x"1d",
          5382 => x"fb",
          5383 => x"39",
          5384 => x"16",
          5385 => x"ff",
          5386 => x"7d",
          5387 => x"84",
          5388 => x"16",
          5389 => x"e4",
          5390 => x"27",
          5391 => x"74",
          5392 => x"38",
          5393 => x"08",
          5394 => x"51",
          5395 => x"ec",
          5396 => x"f8",
          5397 => x"f8",
          5398 => x"79",
          5399 => x"19",
          5400 => x"5a",
          5401 => x"1a",
          5402 => x"05",
          5403 => x"38",
          5404 => x"76",
          5405 => x"0c",
          5406 => x"80",
          5407 => x"e4",
          5408 => x"39",
          5409 => x"f0",
          5410 => x"40",
          5411 => x"79",
          5412 => x"75",
          5413 => x"74",
          5414 => x"84",
          5415 => x"84",
          5416 => x"55",
          5417 => x"55",
          5418 => x"81",
          5419 => x"81",
          5420 => x"08",
          5421 => x"81",
          5422 => x"38",
          5423 => x"7a",
          5424 => x"05",
          5425 => x"38",
          5426 => x"55",
          5427 => x"ff",
          5428 => x"0c",
          5429 => x"9c",
          5430 => x"60",
          5431 => x"70",
          5432 => x"56",
          5433 => x"15",
          5434 => x"2e",
          5435 => x"75",
          5436 => x"77",
          5437 => x"33",
          5438 => x"e4",
          5439 => x"33",
          5440 => x"b4",
          5441 => x"27",
          5442 => x"1e",
          5443 => x"81",
          5444 => x"59",
          5445 => x"77",
          5446 => x"08",
          5447 => x"08",
          5448 => x"5c",
          5449 => x"84",
          5450 => x"74",
          5451 => x"04",
          5452 => x"08",
          5453 => x"71",
          5454 => x"38",
          5455 => x"77",
          5456 => x"33",
          5457 => x"09",
          5458 => x"76",
          5459 => x"51",
          5460 => x"08",
          5461 => x"5b",
          5462 => x"38",
          5463 => x"11",
          5464 => x"59",
          5465 => x"70",
          5466 => x"05",
          5467 => x"2e",
          5468 => x"56",
          5469 => x"ff",
          5470 => x"39",
          5471 => x"19",
          5472 => x"ff",
          5473 => x"e4",
          5474 => x"9c",
          5475 => x"34",
          5476 => x"84",
          5477 => x"1a",
          5478 => x"33",
          5479 => x"fe",
          5480 => x"a0",
          5481 => x"19",
          5482 => x"5b",
          5483 => x"94",
          5484 => x"1a",
          5485 => x"3f",
          5486 => x"39",
          5487 => x"3f",
          5488 => x"74",
          5489 => x"57",
          5490 => x"34",
          5491 => x"3d",
          5492 => x"82",
          5493 => x"0d",
          5494 => x"66",
          5495 => x"89",
          5496 => x"08",
          5497 => x"33",
          5498 => x"16",
          5499 => x"78",
          5500 => x"41",
          5501 => x"1a",
          5502 => x"1a",
          5503 => x"58",
          5504 => x"38",
          5505 => x"7b",
          5506 => x"7a",
          5507 => x"ff",
          5508 => x"8a",
          5509 => x"06",
          5510 => x"9e",
          5511 => x"2e",
          5512 => x"a1",
          5513 => x"74",
          5514 => x"38",
          5515 => x"16",
          5516 => x"38",
          5517 => x"08",
          5518 => x"85",
          5519 => x"29",
          5520 => x"80",
          5521 => x"89",
          5522 => x"98",
          5523 => x"85",
          5524 => x"7b",
          5525 => x"ff",
          5526 => x"85",
          5527 => x"31",
          5528 => x"84",
          5529 => x"1f",
          5530 => x"56",
          5531 => x"ff",
          5532 => x"75",
          5533 => x"7a",
          5534 => x"79",
          5535 => x"94",
          5536 => x"57",
          5537 => x"74",
          5538 => x"85",
          5539 => x"c0",
          5540 => x"56",
          5541 => x"0d",
          5542 => x"3d",
          5543 => x"82",
          5544 => x"60",
          5545 => x"ff",
          5546 => x"7a",
          5547 => x"57",
          5548 => x"80",
          5549 => x"5f",
          5550 => x"d5",
          5551 => x"52",
          5552 => x"3f",
          5553 => x"38",
          5554 => x"0c",
          5555 => x"08",
          5556 => x"05",
          5557 => x"95",
          5558 => x"75",
          5559 => x"56",
          5560 => x"83",
          5561 => x"b4",
          5562 => x"81",
          5563 => x"3f",
          5564 => x"2e",
          5565 => x"b8",
          5566 => x"08",
          5567 => x"08",
          5568 => x"fe",
          5569 => x"82",
          5570 => x"81",
          5571 => x"05",
          5572 => x"ff",
          5573 => x"39",
          5574 => x"77",
          5575 => x"7f",
          5576 => x"0c",
          5577 => x"9c",
          5578 => x"1a",
          5579 => x"3f",
          5580 => x"e4",
          5581 => x"58",
          5582 => x"ff",
          5583 => x"55",
          5584 => x"e4",
          5585 => x"b8",
          5586 => x"57",
          5587 => x"08",
          5588 => x"83",
          5589 => x"08",
          5590 => x"fd",
          5591 => x"82",
          5592 => x"81",
          5593 => x"05",
          5594 => x"ff",
          5595 => x"39",
          5596 => x"3f",
          5597 => x"74",
          5598 => x"57",
          5599 => x"08",
          5600 => x"33",
          5601 => x"b8",
          5602 => x"e4",
          5603 => x"a8",
          5604 => x"08",
          5605 => x"58",
          5606 => x"8b",
          5607 => x"17",
          5608 => x"33",
          5609 => x"b4",
          5610 => x"fd",
          5611 => x"81",
          5612 => x"0d",
          5613 => x"0b",
          5614 => x"04",
          5615 => x"77",
          5616 => x"75",
          5617 => x"74",
          5618 => x"84",
          5619 => x"83",
          5620 => x"56",
          5621 => x"70",
          5622 => x"80",
          5623 => x"08",
          5624 => x"ac",
          5625 => x"bc",
          5626 => x"52",
          5627 => x"3f",
          5628 => x"38",
          5629 => x"0c",
          5630 => x"8b",
          5631 => x"8b",
          5632 => x"70",
          5633 => x"7a",
          5634 => x"79",
          5635 => x"96",
          5636 => x"81",
          5637 => x"7b",
          5638 => x"18",
          5639 => x"18",
          5640 => x"18",
          5641 => x"18",
          5642 => x"cc",
          5643 => x"18",
          5644 => x"5b",
          5645 => x"ff",
          5646 => x"90",
          5647 => x"79",
          5648 => x"0c",
          5649 => x"17",
          5650 => x"18",
          5651 => x"81",
          5652 => x"38",
          5653 => x"b4",
          5654 => x"b8",
          5655 => x"08",
          5656 => x"55",
          5657 => x"81",
          5658 => x"18",
          5659 => x"33",
          5660 => x"fd",
          5661 => x"94",
          5662 => x"95",
          5663 => x"7b",
          5664 => x"18",
          5665 => x"18",
          5666 => x"18",
          5667 => x"18",
          5668 => x"cc",
          5669 => x"18",
          5670 => x"5b",
          5671 => x"ff",
          5672 => x"90",
          5673 => x"79",
          5674 => x"16",
          5675 => x"b8",
          5676 => x"ba",
          5677 => x"b4",
          5678 => x"55",
          5679 => x"54",
          5680 => x"56",
          5681 => x"53",
          5682 => x"52",
          5683 => x"22",
          5684 => x"2e",
          5685 => x"54",
          5686 => x"84",
          5687 => x"81",
          5688 => x"84",
          5689 => x"da",
          5690 => x"39",
          5691 => x"57",
          5692 => x"70",
          5693 => x"52",
          5694 => x"ee",
          5695 => x"d0",
          5696 => x"38",
          5697 => x"84",
          5698 => x"8b",
          5699 => x"0d",
          5700 => x"ff",
          5701 => x"91",
          5702 => x"d0",
          5703 => x"f5",
          5704 => x"58",
          5705 => x"81",
          5706 => x"57",
          5707 => x"70",
          5708 => x"81",
          5709 => x"51",
          5710 => x"70",
          5711 => x"70",
          5712 => x"09",
          5713 => x"38",
          5714 => x"07",
          5715 => x"76",
          5716 => x"1b",
          5717 => x"38",
          5718 => x"24",
          5719 => x"c3",
          5720 => x"3d",
          5721 => x"94",
          5722 => x"b8",
          5723 => x"84",
          5724 => x"7a",
          5725 => x"51",
          5726 => x"55",
          5727 => x"02",
          5728 => x"58",
          5729 => x"02",
          5730 => x"06",
          5731 => x"7a",
          5732 => x"71",
          5733 => x"5b",
          5734 => x"76",
          5735 => x"0c",
          5736 => x"08",
          5737 => x"38",
          5738 => x"3d",
          5739 => x"33",
          5740 => x"79",
          5741 => x"39",
          5742 => x"84",
          5743 => x"ff",
          5744 => x"80",
          5745 => x"34",
          5746 => x"05",
          5747 => x"3f",
          5748 => x"e4",
          5749 => x"3d",
          5750 => x"dd",
          5751 => x"5b",
          5752 => x"80",
          5753 => x"52",
          5754 => x"b8",
          5755 => x"83",
          5756 => x"58",
          5757 => x"38",
          5758 => x"5f",
          5759 => x"76",
          5760 => x"51",
          5761 => x"08",
          5762 => x"59",
          5763 => x"38",
          5764 => x"9a",
          5765 => x"70",
          5766 => x"83",
          5767 => x"3d",
          5768 => x"b7",
          5769 => x"b8",
          5770 => x"7a",
          5771 => x"e4",
          5772 => x"38",
          5773 => x"9a",
          5774 => x"70",
          5775 => x"83",
          5776 => x"a4",
          5777 => x"51",
          5778 => x"08",
          5779 => x"ff",
          5780 => x"38",
          5781 => x"fd",
          5782 => x"89",
          5783 => x"57",
          5784 => x"56",
          5785 => x"57",
          5786 => x"75",
          5787 => x"2e",
          5788 => x"ff",
          5789 => x"19",
          5790 => x"33",
          5791 => x"80",
          5792 => x"7e",
          5793 => x"fd",
          5794 => x"38",
          5795 => x"10",
          5796 => x"70",
          5797 => x"7a",
          5798 => x"70",
          5799 => x"82",
          5800 => x"80",
          5801 => x"16",
          5802 => x"5e",
          5803 => x"ee",
          5804 => x"34",
          5805 => x"df",
          5806 => x"84",
          5807 => x"04",
          5808 => x"98",
          5809 => x"59",
          5810 => x"33",
          5811 => x"90",
          5812 => x"0c",
          5813 => x"a0",
          5814 => x"84",
          5815 => x"38",
          5816 => x"08",
          5817 => x"33",
          5818 => x"59",
          5819 => x"84",
          5820 => x"16",
          5821 => x"e4",
          5822 => x"27",
          5823 => x"74",
          5824 => x"38",
          5825 => x"08",
          5826 => x"51",
          5827 => x"dd",
          5828 => x"11",
          5829 => x"84",
          5830 => x"e4",
          5831 => x"59",
          5832 => x"81",
          5833 => x"80",
          5834 => x"5a",
          5835 => x"34",
          5836 => x"e5",
          5837 => x"79",
          5838 => x"7f",
          5839 => x"82",
          5840 => x"e4",
          5841 => x"3d",
          5842 => x"74",
          5843 => x"73",
          5844 => x"72",
          5845 => x"84",
          5846 => x"83",
          5847 => x"53",
          5848 => x"53",
          5849 => x"56",
          5850 => x"15",
          5851 => x"81",
          5852 => x"89",
          5853 => x"81",
          5854 => x"fd",
          5855 => x"ff",
          5856 => x"fd",
          5857 => x"73",
          5858 => x"06",
          5859 => x"98",
          5860 => x"2e",
          5861 => x"d9",
          5862 => x"17",
          5863 => x"81",
          5864 => x"80",
          5865 => x"51",
          5866 => x"08",
          5867 => x"81",
          5868 => x"81",
          5869 => x"73",
          5870 => x"73",
          5871 => x"0b",
          5872 => x"b8",
          5873 => x"15",
          5874 => x"58",
          5875 => x"08",
          5876 => x"09",
          5877 => x"16",
          5878 => x"27",
          5879 => x"15",
          5880 => x"16",
          5881 => x"80",
          5882 => x"2e",
          5883 => x"0b",
          5884 => x"04",
          5885 => x"08",
          5886 => x"73",
          5887 => x"c2",
          5888 => x"08",
          5889 => x"0c",
          5890 => x"2e",
          5891 => x"08",
          5892 => x"27",
          5893 => x"71",
          5894 => x"2a",
          5895 => x"80",
          5896 => x"e9",
          5897 => x"b7",
          5898 => x"8a",
          5899 => x"a2",
          5900 => x"53",
          5901 => x"54",
          5902 => x"51",
          5903 => x"08",
          5904 => x"98",
          5905 => x"fd",
          5906 => x"16",
          5907 => x"39",
          5908 => x"84",
          5909 => x"f6",
          5910 => x"80",
          5911 => x"fc",
          5912 => x"c5",
          5913 => x"84",
          5914 => x"80",
          5915 => x"e4",
          5916 => x"0c",
          5917 => x"3f",
          5918 => x"e4",
          5919 => x"70",
          5920 => x"af",
          5921 => x"81",
          5922 => x"c5",
          5923 => x"9a",
          5924 => x"70",
          5925 => x"83",
          5926 => x"7a",
          5927 => x"74",
          5928 => x"84",
          5929 => x"8d",
          5930 => x"80",
          5931 => x"80",
          5932 => x"33",
          5933 => x"90",
          5934 => x"5a",
          5935 => x"78",
          5936 => x"38",
          5937 => x"38",
          5938 => x"38",
          5939 => x"52",
          5940 => x"71",
          5941 => x"73",
          5942 => x"04",
          5943 => x"3f",
          5944 => x"71",
          5945 => x"d7",
          5946 => x"55",
          5947 => x"74",
          5948 => x"73",
          5949 => x"86",
          5950 => x"72",
          5951 => x"72",
          5952 => x"76",
          5953 => x"74",
          5954 => x"e4",
          5955 => x"2e",
          5956 => x"38",
          5957 => x"3f",
          5958 => x"3f",
          5959 => x"30",
          5960 => x"e4",
          5961 => x"b8",
          5962 => x"77",
          5963 => x"3f",
          5964 => x"3f",
          5965 => x"30",
          5966 => x"e4",
          5967 => x"75",
          5968 => x"84",
          5969 => x"8a",
          5970 => x"fe",
          5971 => x"81",
          5972 => x"75",
          5973 => x"3d",
          5974 => x"70",
          5975 => x"3f",
          5976 => x"e4",
          5977 => x"b8",
          5978 => x"52",
          5979 => x"b8",
          5980 => x"e5",
          5981 => x"98",
          5982 => x"38",
          5983 => x"75",
          5984 => x"b8",
          5985 => x"0b",
          5986 => x"04",
          5987 => x"80",
          5988 => x"3d",
          5989 => x"08",
          5990 => x"7f",
          5991 => x"fe",
          5992 => x"57",
          5993 => x"0c",
          5994 => x"0d",
          5995 => x"5a",
          5996 => x"77",
          5997 => x"5a",
          5998 => x"81",
          5999 => x"08",
          6000 => x"33",
          6001 => x"81",
          6002 => x"17",
          6003 => x"b8",
          6004 => x"5a",
          6005 => x"7e",
          6006 => x"33",
          6007 => x"77",
          6008 => x"12",
          6009 => x"07",
          6010 => x"2b",
          6011 => x"80",
          6012 => x"63",
          6013 => x"62",
          6014 => x"52",
          6015 => x"f2",
          6016 => x"0c",
          6017 => x"84",
          6018 => x"95",
          6019 => x"08",
          6020 => x"33",
          6021 => x"5e",
          6022 => x"84",
          6023 => x"17",
          6024 => x"e4",
          6025 => x"27",
          6026 => x"74",
          6027 => x"38",
          6028 => x"08",
          6029 => x"51",
          6030 => x"97",
          6031 => x"56",
          6032 => x"3f",
          6033 => x"e8",
          6034 => x"80",
          6035 => x"70",
          6036 => x"7c",
          6037 => x"5c",
          6038 => x"7a",
          6039 => x"17",
          6040 => x"34",
          6041 => x"81",
          6042 => x"07",
          6043 => x"1d",
          6044 => x"5f",
          6045 => x"38",
          6046 => x"39",
          6047 => x"7a",
          6048 => x"07",
          6049 => x"39",
          6050 => x"3d",
          6051 => x"2e",
          6052 => x"2e",
          6053 => x"2e",
          6054 => x"22",
          6055 => x"38",
          6056 => x"38",
          6057 => x"38",
          6058 => x"06",
          6059 => x"80",
          6060 => x"8c",
          6061 => x"d5",
          6062 => x"54",
          6063 => x"08",
          6064 => x"0b",
          6065 => x"18",
          6066 => x"90",
          6067 => x"75",
          6068 => x"b8",
          6069 => x"54",
          6070 => x"52",
          6071 => x"b8",
          6072 => x"80",
          6073 => x"08",
          6074 => x"e4",
          6075 => x"53",
          6076 => x"3f",
          6077 => x"9c",
          6078 => x"57",
          6079 => x"38",
          6080 => x"33",
          6081 => x"78",
          6082 => x"9c",
          6083 => x"e2",
          6084 => x"54",
          6085 => x"55",
          6086 => x"18",
          6087 => x"88",
          6088 => x"08",
          6089 => x"84",
          6090 => x"38",
          6091 => x"be",
          6092 => x"84",
          6093 => x"81",
          6094 => x"18",
          6095 => x"0b",
          6096 => x"38",
          6097 => x"27",
          6098 => x"38",
          6099 => x"83",
          6100 => x"84",
          6101 => x"52",
          6102 => x"b8",
          6103 => x"80",
          6104 => x"08",
          6105 => x"e4",
          6106 => x"53",
          6107 => x"3f",
          6108 => x"9c",
          6109 => x"57",
          6110 => x"81",
          6111 => x"81",
          6112 => x"54",
          6113 => x"55",
          6114 => x"f3",
          6115 => x"0b",
          6116 => x"39",
          6117 => x"18",
          6118 => x"b8",
          6119 => x"fd",
          6120 => x"59",
          6121 => x"08",
          6122 => x"39",
          6123 => x"ff",
          6124 => x"b7",
          6125 => x"84",
          6126 => x"75",
          6127 => x"04",
          6128 => x"3d",
          6129 => x"84",
          6130 => x"08",
          6131 => x"70",
          6132 => x"56",
          6133 => x"80",
          6134 => x"05",
          6135 => x"56",
          6136 => x"08",
          6137 => x"88",
          6138 => x"57",
          6139 => x"76",
          6140 => x"2e",
          6141 => x"08",
          6142 => x"7a",
          6143 => x"3d",
          6144 => x"84",
          6145 => x"08",
          6146 => x"52",
          6147 => x"b8",
          6148 => x"a0",
          6149 => x"a7",
          6150 => x"17",
          6151 => x"07",
          6152 => x"39",
          6153 => x"38",
          6154 => x"78",
          6155 => x"57",
          6156 => x"52",
          6157 => x"b8",
          6158 => x"80",
          6159 => x"07",
          6160 => x"9a",
          6161 => x"79",
          6162 => x"38",
          6163 => x"38",
          6164 => x"51",
          6165 => x"08",
          6166 => x"04",
          6167 => x"80",
          6168 => x"b9",
          6169 => x"74",
          6170 => x"38",
          6171 => x"81",
          6172 => x"84",
          6173 => x"ff",
          6174 => x"77",
          6175 => x"58",
          6176 => x"34",
          6177 => x"38",
          6178 => x"3f",
          6179 => x"e4",
          6180 => x"84",
          6181 => x"82",
          6182 => x"17",
          6183 => x"51",
          6184 => x"b8",
          6185 => x"ff",
          6186 => x"18",
          6187 => x"31",
          6188 => x"a0",
          6189 => x"17",
          6190 => x"06",
          6191 => x"08",
          6192 => x"81",
          6193 => x"79",
          6194 => x"78",
          6195 => x"51",
          6196 => x"08",
          6197 => x"80",
          6198 => x"2e",
          6199 => x"ff",
          6200 => x"52",
          6201 => x"b8",
          6202 => x"fe",
          6203 => x"75",
          6204 => x"94",
          6205 => x"5c",
          6206 => x"7a",
          6207 => x"a2",
          6208 => x"b8",
          6209 => x"56",
          6210 => x"53",
          6211 => x"3d",
          6212 => x"e4",
          6213 => x"2e",
          6214 => x"9f",
          6215 => x"93",
          6216 => x"3f",
          6217 => x"e4",
          6218 => x"e4",
          6219 => x"e4",
          6220 => x"38",
          6221 => x"2a",
          6222 => x"ff",
          6223 => x"3d",
          6224 => x"84",
          6225 => x"b8",
          6226 => x"b8",
          6227 => x"84",
          6228 => x"38",
          6229 => x"e4",
          6230 => x"7a",
          6231 => x"08",
          6232 => x"79",
          6233 => x"71",
          6234 => x"7a",
          6235 => x"80",
          6236 => x"05",
          6237 => x"38",
          6238 => x"75",
          6239 => x"1b",
          6240 => x"fe",
          6241 => x"81",
          6242 => x"82",
          6243 => x"17",
          6244 => x"18",
          6245 => x"81",
          6246 => x"84",
          6247 => x"17",
          6248 => x"a0",
          6249 => x"17",
          6250 => x"06",
          6251 => x"08",
          6252 => x"81",
          6253 => x"fe",
          6254 => x"58",
          6255 => x"7b",
          6256 => x"74",
          6257 => x"84",
          6258 => x"08",
          6259 => x"e4",
          6260 => x"b8",
          6261 => x"80",
          6262 => x"b0",
          6263 => x"38",
          6264 => x"08",
          6265 => x"38",
          6266 => x"33",
          6267 => x"79",
          6268 => x"75",
          6269 => x"04",
          6270 => x"ff",
          6271 => x"09",
          6272 => x"b8",
          6273 => x"05",
          6274 => x"38",
          6275 => x"7d",
          6276 => x"7d",
          6277 => x"80",
          6278 => x"1a",
          6279 => x"34",
          6280 => x"56",
          6281 => x"2a",
          6282 => x"33",
          6283 => x"7d",
          6284 => x"1b",
          6285 => x"56",
          6286 => x"ff",
          6287 => x"ae",
          6288 => x"71",
          6289 => x"78",
          6290 => x"5b",
          6291 => x"55",
          6292 => x"5b",
          6293 => x"ff",
          6294 => x"56",
          6295 => x"69",
          6296 => x"34",
          6297 => x"a1",
          6298 => x"99",
          6299 => x"9a",
          6300 => x"9b",
          6301 => x"2e",
          6302 => x"8b",
          6303 => x"18",
          6304 => x"84",
          6305 => x"e4",
          6306 => x"2a",
          6307 => x"88",
          6308 => x"fe",
          6309 => x"80",
          6310 => x"74",
          6311 => x"0b",
          6312 => x"56",
          6313 => x"77",
          6314 => x"7b",
          6315 => x"8b",
          6316 => x"18",
          6317 => x"84",
          6318 => x"d1",
          6319 => x"70",
          6320 => x"38",
          6321 => x"9f",
          6322 => x"b8",
          6323 => x"81",
          6324 => x"fc",
          6325 => x"b4",
          6326 => x"b8",
          6327 => x"84",
          6328 => x"7f",
          6329 => x"a5",
          6330 => x"3f",
          6331 => x"e4",
          6332 => x"33",
          6333 => x"ce",
          6334 => x"08",
          6335 => x"57",
          6336 => x"ff",
          6337 => x"58",
          6338 => x"70",
          6339 => x"05",
          6340 => x"38",
          6341 => x"9e",
          6342 => x"84",
          6343 => x"a8",
          6344 => x"0b",
          6345 => x"04",
          6346 => x"06",
          6347 => x"38",
          6348 => x"05",
          6349 => x"38",
          6350 => x"08",
          6351 => x"70",
          6352 => x"05",
          6353 => x"56",
          6354 => x"70",
          6355 => x"17",
          6356 => x"17",
          6357 => x"30",
          6358 => x"2e",
          6359 => x"be",
          6360 => x"72",
          6361 => x"55",
          6362 => x"84",
          6363 => x"c2",
          6364 => x"96",
          6365 => x"79",
          6366 => x"fc",
          6367 => x"e4",
          6368 => x"b8",
          6369 => x"39",
          6370 => x"06",
          6371 => x"a8",
          6372 => x"b8",
          6373 => x"93",
          6374 => x"cd",
          6375 => x"05",
          6376 => x"34",
          6377 => x"80",
          6378 => x"18",
          6379 => x"56",
          6380 => x"76",
          6381 => x"83",
          6382 => x"2a",
          6383 => x"81",
          6384 => x"81",
          6385 => x"1a",
          6386 => x"41",
          6387 => x"e0",
          6388 => x"05",
          6389 => x"38",
          6390 => x"19",
          6391 => x"82",
          6392 => x"17",
          6393 => x"33",
          6394 => x"75",
          6395 => x"51",
          6396 => x"08",
          6397 => x"5c",
          6398 => x"80",
          6399 => x"38",
          6400 => x"09",
          6401 => x"ff",
          6402 => x"18",
          6403 => x"f3",
          6404 => x"2e",
          6405 => x"2a",
          6406 => x"88",
          6407 => x"7f",
          6408 => x"08",
          6409 => x"5c",
          6410 => x"52",
          6411 => x"b8",
          6412 => x"80",
          6413 => x"08",
          6414 => x"2e",
          6415 => x"5f",
          6416 => x"a8",
          6417 => x"52",
          6418 => x"3f",
          6419 => x"38",
          6420 => x"0c",
          6421 => x"08",
          6422 => x"17",
          6423 => x"38",
          6424 => x"3f",
          6425 => x"e4",
          6426 => x"56",
          6427 => x"56",
          6428 => x"e5",
          6429 => x"b8",
          6430 => x"0b",
          6431 => x"04",
          6432 => x"98",
          6433 => x"58",
          6434 => x"e4",
          6435 => x"b8",
          6436 => x"75",
          6437 => x"04",
          6438 => x"52",
          6439 => x"3f",
          6440 => x"2e",
          6441 => x"b8",
          6442 => x"08",
          6443 => x"08",
          6444 => x"fe",
          6445 => x"82",
          6446 => x"81",
          6447 => x"05",
          6448 => x"fe",
          6449 => x"39",
          6450 => x"17",
          6451 => x"fe",
          6452 => x"e4",
          6453 => x"08",
          6454 => x"18",
          6455 => x"55",
          6456 => x"38",
          6457 => x"09",
          6458 => x"b4",
          6459 => x"7a",
          6460 => x"eb",
          6461 => x"3d",
          6462 => x"84",
          6463 => x"82",
          6464 => x"3d",
          6465 => x"e4",
          6466 => x"2e",
          6467 => x"96",
          6468 => x"96",
          6469 => x"3f",
          6470 => x"e4",
          6471 => x"33",
          6472 => x"d2",
          6473 => x"8b",
          6474 => x"07",
          6475 => x"34",
          6476 => x"78",
          6477 => x"e4",
          6478 => x"0d",
          6479 => x"53",
          6480 => x"51",
          6481 => x"08",
          6482 => x"8a",
          6483 => x"3d",
          6484 => x"3d",
          6485 => x"84",
          6486 => x"08",
          6487 => x"81",
          6488 => x"38",
          6489 => x"71",
          6490 => x"96",
          6491 => x"97",
          6492 => x"98",
          6493 => x"99",
          6494 => x"18",
          6495 => x"84",
          6496 => x"96",
          6497 => x"6d",
          6498 => x"05",
          6499 => x"3f",
          6500 => x"08",
          6501 => x"80",
          6502 => x"8b",
          6503 => x"78",
          6504 => x"07",
          6505 => x"81",
          6506 => x"58",
          6507 => x"a4",
          6508 => x"16",
          6509 => x"16",
          6510 => x"09",
          6511 => x"76",
          6512 => x"51",
          6513 => x"08",
          6514 => x"59",
          6515 => x"bd",
          6516 => x"c3",
          6517 => x"e4",
          6518 => x"56",
          6519 => x"82",
          6520 => x"2b",
          6521 => x"88",
          6522 => x"5f",
          6523 => x"b8",
          6524 => x"5e",
          6525 => x"52",
          6526 => x"e4",
          6527 => x"2e",
          6528 => x"81",
          6529 => x"80",
          6530 => x"16",
          6531 => x"17",
          6532 => x"77",
          6533 => x"09",
          6534 => x"e4",
          6535 => x"a8",
          6536 => x"5a",
          6537 => x"ad",
          6538 => x"2e",
          6539 => x"54",
          6540 => x"53",
          6541 => x"db",
          6542 => x"53",
          6543 => x"fe",
          6544 => x"80",
          6545 => x"75",
          6546 => x"84",
          6547 => x"08",
          6548 => x"84",
          6549 => x"79",
          6550 => x"56",
          6551 => x"8a",
          6552 => x"57",
          6553 => x"fc",
          6554 => x"33",
          6555 => x"38",
          6556 => x"39",
          6557 => x"ff",
          6558 => x"9c",
          6559 => x"84",
          6560 => x"3d",
          6561 => x"70",
          6562 => x"74",
          6563 => x"33",
          6564 => x"5a",
          6565 => x"3d",
          6566 => x"06",
          6567 => x"38",
          6568 => x"26",
          6569 => x"3f",
          6570 => x"51",
          6571 => x"83",
          6572 => x"81",
          6573 => x"e5",
          6574 => x"56",
          6575 => x"74",
          6576 => x"18",
          6577 => x"57",
          6578 => x"77",
          6579 => x"81",
          6580 => x"81",
          6581 => x"89",
          6582 => x"27",
          6583 => x"7b",
          6584 => x"5a",
          6585 => x"81",
          6586 => x"81",
          6587 => x"9f",
          6588 => x"57",
          6589 => x"38",
          6590 => x"05",
          6591 => x"7a",
          6592 => x"ff",
          6593 => x"80",
          6594 => x"56",
          6595 => x"08",
          6596 => x"b4",
          6597 => x"0c",
          6598 => x"74",
          6599 => x"08",
          6600 => x"f8",
          6601 => x"0c",
          6602 => x"33",
          6603 => x"51",
          6604 => x"08",
          6605 => x"38",
          6606 => x"6c",
          6607 => x"05",
          6608 => x"34",
          6609 => x"5d",
          6610 => x"fe",
          6611 => x"55",
          6612 => x"27",
          6613 => x"39",
          6614 => x"81",
          6615 => x"75",
          6616 => x"53",
          6617 => x"84",
          6618 => x"08",
          6619 => x"38",
          6620 => x"5a",
          6621 => x"18",
          6622 => x"33",
          6623 => x"81",
          6624 => x"18",
          6625 => x"c4",
          6626 => x"85",
          6627 => x"19",
          6628 => x"9c",
          6629 => x"74",
          6630 => x"30",
          6631 => x"74",
          6632 => x"5a",
          6633 => x"75",
          6634 => x"e4",
          6635 => x"2e",
          6636 => x"2e",
          6637 => x"b9",
          6638 => x"70",
          6639 => x"74",
          6640 => x"17",
          6641 => x"76",
          6642 => x"81",
          6643 => x"80",
          6644 => x"05",
          6645 => x"34",
          6646 => x"d6",
          6647 => x"5d",
          6648 => x"fe",
          6649 => x"55",
          6650 => x"39",
          6651 => x"52",
          6652 => x"3f",
          6653 => x"81",
          6654 => x"08",
          6655 => x"19",
          6656 => x"27",
          6657 => x"82",
          6658 => x"59",
          6659 => x"75",
          6660 => x"e4",
          6661 => x"2e",
          6662 => x"70",
          6663 => x"38",
          6664 => x"08",
          6665 => x"81",
          6666 => x"fd",
          6667 => x"02",
          6668 => x"5b",
          6669 => x"38",
          6670 => x"38",
          6671 => x"38",
          6672 => x"59",
          6673 => x"54",
          6674 => x"17",
          6675 => x"80",
          6676 => x"81",
          6677 => x"2a",
          6678 => x"81",
          6679 => x"89",
          6680 => x"59",
          6681 => x"06",
          6682 => x"84",
          6683 => x"79",
          6684 => x"27",
          6685 => x"83",
          6686 => x"80",
          6687 => x"87",
          6688 => x"14",
          6689 => x"84",
          6690 => x"38",
          6691 => x"d8",
          6692 => x"38",
          6693 => x"38",
          6694 => x"38",
          6695 => x"e4",
          6696 => x"84",
          6697 => x"81",
          6698 => x"84",
          6699 => x"fe",
          6700 => x"fe",
          6701 => x"38",
          6702 => x"ab",
          6703 => x"80",
          6704 => x"51",
          6705 => x"08",
          6706 => x"38",
          6707 => x"5e",
          6708 => x"0c",
          6709 => x"7a",
          6710 => x"90",
          6711 => x"90",
          6712 => x"94",
          6713 => x"fe",
          6714 => x"0c",
          6715 => x"84",
          6716 => x"ff",
          6717 => x"59",
          6718 => x"39",
          6719 => x"5e",
          6720 => x"e3",
          6721 => x"08",
          6722 => x"44",
          6723 => x"70",
          6724 => x"8a",
          6725 => x"70",
          6726 => x"85",
          6727 => x"2e",
          6728 => x"56",
          6729 => x"10",
          6730 => x"56",
          6731 => x"75",
          6732 => x"33",
          6733 => x"5d",
          6734 => x"3f",
          6735 => x"70",
          6736 => x"84",
          6737 => x"40",
          6738 => x"3d",
          6739 => x"fe",
          6740 => x"84",
          6741 => x"84",
          6742 => x"84",
          6743 => x"74",
          6744 => x"38",
          6745 => x"7e",
          6746 => x"ff",
          6747 => x"38",
          6748 => x"2a",
          6749 => x"5b",
          6750 => x"30",
          6751 => x"91",
          6752 => x"2e",
          6753 => x"60",
          6754 => x"81",
          6755 => x"38",
          6756 => x"fe",
          6757 => x"56",
          6758 => x"09",
          6759 => x"29",
          6760 => x"58",
          6761 => x"b6",
          6762 => x"71",
          6763 => x"14",
          6764 => x"33",
          6765 => x"33",
          6766 => x"88",
          6767 => x"07",
          6768 => x"a2",
          6769 => x"3d",
          6770 => x"41",
          6771 => x"ff",
          6772 => x"7a",
          6773 => x"81",
          6774 => x"80",
          6775 => x"45",
          6776 => x"06",
          6777 => x"70",
          6778 => x"83",
          6779 => x"78",
          6780 => x"88",
          6781 => x"38",
          6782 => x"88",
          6783 => x"57",
          6784 => x"76",
          6785 => x"51",
          6786 => x"08",
          6787 => x"08",
          6788 => x"84",
          6789 => x"08",
          6790 => x"57",
          6791 => x"5d",
          6792 => x"11",
          6793 => x"6b",
          6794 => x"62",
          6795 => x"5d",
          6796 => x"56",
          6797 => x"78",
          6798 => x"68",
          6799 => x"84",
          6800 => x"89",
          6801 => x"06",
          6802 => x"84",
          6803 => x"7a",
          6804 => x"80",
          6805 => x"fe",
          6806 => x"e4",
          6807 => x"0c",
          6808 => x"0b",
          6809 => x"84",
          6810 => x"11",
          6811 => x"74",
          6812 => x"81",
          6813 => x"7a",
          6814 => x"e4",
          6815 => x"5b",
          6816 => x"70",
          6817 => x"45",
          6818 => x"e0",
          6819 => x"ff",
          6820 => x"38",
          6821 => x"46",
          6822 => x"76",
          6823 => x"78",
          6824 => x"30",
          6825 => x"5d",
          6826 => x"38",
          6827 => x"7c",
          6828 => x"e0",
          6829 => x"52",
          6830 => x"57",
          6831 => x"61",
          6832 => x"08",
          6833 => x"6c",
          6834 => x"9c",
          6835 => x"39",
          6836 => x"24",
          6837 => x"0c",
          6838 => x"48",
          6839 => x"38",
          6840 => x"fc",
          6841 => x"f5",
          6842 => x"18",
          6843 => x"38",
          6844 => x"9f",
          6845 => x"80",
          6846 => x"9f",
          6847 => x"06",
          6848 => x"84",
          6849 => x"81",
          6850 => x"f4",
          6851 => x"57",
          6852 => x"76",
          6853 => x"55",
          6854 => x"74",
          6855 => x"77",
          6856 => x"ff",
          6857 => x"6a",
          6858 => x"34",
          6859 => x"32",
          6860 => x"05",
          6861 => x"68",
          6862 => x"83",
          6863 => x"83",
          6864 => x"05",
          6865 => x"94",
          6866 => x"bf",
          6867 => x"05",
          6868 => x"61",
          6869 => x"34",
          6870 => x"05",
          6871 => x"9e",
          6872 => x"f0",
          6873 => x"05",
          6874 => x"80",
          6875 => x"05",
          6876 => x"cc",
          6877 => x"ff",
          6878 => x"74",
          6879 => x"34",
          6880 => x"61",
          6881 => x"83",
          6882 => x"81",
          6883 => x"58",
          6884 => x"60",
          6885 => x"34",
          6886 => x"6b",
          6887 => x"79",
          6888 => x"84",
          6889 => x"17",
          6890 => x"69",
          6891 => x"05",
          6892 => x"38",
          6893 => x"86",
          6894 => x"62",
          6895 => x"61",
          6896 => x"74",
          6897 => x"90",
          6898 => x"46",
          6899 => x"34",
          6900 => x"83",
          6901 => x"60",
          6902 => x"84",
          6903 => x"80",
          6904 => x"05",
          6905 => x"38",
          6906 => x"76",
          6907 => x"80",
          6908 => x"83",
          6909 => x"75",
          6910 => x"54",
          6911 => x"c4",
          6912 => x"9b",
          6913 => x"5b",
          6914 => x"2e",
          6915 => x"ff",
          6916 => x"2e",
          6917 => x"38",
          6918 => x"81",
          6919 => x"80",
          6920 => x"19",
          6921 => x"34",
          6922 => x"05",
          6923 => x"05",
          6924 => x"67",
          6925 => x"34",
          6926 => x"1f",
          6927 => x"85",
          6928 => x"2a",
          6929 => x"34",
          6930 => x"34",
          6931 => x"61",
          6932 => x"c8",
          6933 => x"83",
          6934 => x"05",
          6935 => x"83",
          6936 => x"77",
          6937 => x"2a",
          6938 => x"81",
          6939 => x"fe",
          6940 => x"e4",
          6941 => x"52",
          6942 => x"57",
          6943 => x"84",
          6944 => x"9f",
          6945 => x"62",
          6946 => x"16",
          6947 => x"38",
          6948 => x"e6",
          6949 => x"9d",
          6950 => x"e6",
          6951 => x"22",
          6952 => x"38",
          6953 => x"78",
          6954 => x"e4",
          6955 => x"89",
          6956 => x"84",
          6957 => x"58",
          6958 => x"f5",
          6959 => x"84",
          6960 => x"f8",
          6961 => x"81",
          6962 => x"57",
          6963 => x"63",
          6964 => x"f4",
          6965 => x"75",
          6966 => x"34",
          6967 => x"05",
          6968 => x"a3",
          6969 => x"80",
          6970 => x"05",
          6971 => x"80",
          6972 => x"61",
          6973 => x"7b",
          6974 => x"59",
          6975 => x"2a",
          6976 => x"61",
          6977 => x"34",
          6978 => x"af",
          6979 => x"80",
          6980 => x"05",
          6981 => x"80",
          6982 => x"80",
          6983 => x"05",
          6984 => x"70",
          6985 => x"05",
          6986 => x"2e",
          6987 => x"58",
          6988 => x"ff",
          6989 => x"39",
          6990 => x"51",
          6991 => x"b8",
          6992 => x"29",
          6993 => x"05",
          6994 => x"53",
          6995 => x"3f",
          6996 => x"e4",
          6997 => x"0c",
          6998 => x"6a",
          6999 => x"70",
          7000 => x"ff",
          7001 => x"05",
          7002 => x"61",
          7003 => x"34",
          7004 => x"8a",
          7005 => x"f9",
          7006 => x"60",
          7007 => x"84",
          7008 => x"81",
          7009 => x"f4",
          7010 => x"81",
          7011 => x"75",
          7012 => x"75",
          7013 => x"75",
          7014 => x"34",
          7015 => x"80",
          7016 => x"e1",
          7017 => x"05",
          7018 => x"7a",
          7019 => x"05",
          7020 => x"83",
          7021 => x"7f",
          7022 => x"83",
          7023 => x"05",
          7024 => x"76",
          7025 => x"69",
          7026 => x"87",
          7027 => x"bd",
          7028 => x"60",
          7029 => x"69",
          7030 => x"3d",
          7031 => x"61",
          7032 => x"25",
          7033 => x"f8",
          7034 => x"51",
          7035 => x"09",
          7036 => x"55",
          7037 => x"70",
          7038 => x"74",
          7039 => x"cd",
          7040 => x"83",
          7041 => x"0c",
          7042 => x"7b",
          7043 => x"57",
          7044 => x"17",
          7045 => x"88",
          7046 => x"59",
          7047 => x"bb",
          7048 => x"81",
          7049 => x"04",
          7050 => x"8c",
          7051 => x"d1",
          7052 => x"72",
          7053 => x"0c",
          7054 => x"56",
          7055 => x"94",
          7056 => x"02",
          7057 => x"58",
          7058 => x"70",
          7059 => x"74",
          7060 => x"77",
          7061 => x"80",
          7062 => x"17",
          7063 => x"81",
          7064 => x"74",
          7065 => x"0c",
          7066 => x"9f",
          7067 => x"c0",
          7068 => x"c9",
          7069 => x"7c",
          7070 => x"b8",
          7071 => x"3d",
          7072 => x"05",
          7073 => x"3f",
          7074 => x"07",
          7075 => x"56",
          7076 => x"fd",
          7077 => x"b8",
          7078 => x"3d",
          7079 => x"22",
          7080 => x"26",
          7081 => x"52",
          7082 => x"0d",
          7083 => x"70",
          7084 => x"38",
          7085 => x"a8",
          7086 => x"81",
          7087 => x"54",
          7088 => x"10",
          7089 => x"51",
          7090 => x"ff",
          7091 => x"3d",
          7092 => x"05",
          7093 => x"53",
          7094 => x"8c",
          7095 => x"0c",
          7096 => x"2e",
          7097 => x"ff",
          7098 => x"a8",
          7099 => x"51",
          7100 => x"77",
          7101 => x"e1",
          7102 => x"e8",
          7103 => x"80",
          7104 => x"22",
          7105 => x"7a",
          7106 => x"b7",
          7107 => x"72",
          7108 => x"06",
          7109 => x"b1",
          7110 => x"70",
          7111 => x"30",
          7112 => x"53",
          7113 => x"75",
          7114 => x"3d",
          7115 => x"a2",
          7116 => x"10",
          7117 => x"08",
          7118 => x"ff",
          7119 => x"ff",
          7120 => x"57",
          7121 => x"ff",
          7122 => x"16",
          7123 => x"db",
          7124 => x"06",
          7125 => x"83",
          7126 => x"f0",
          7127 => x"51",
          7128 => x"06",
          7129 => x"06",
          7130 => x"73",
          7131 => x"52",
          7132 => x"ff",
          7133 => x"ff",
          7134 => x"00",
          7135 => x"00",
          7136 => x"00",
          7137 => x"00",
          7138 => x"00",
          7139 => x"00",
          7140 => x"00",
          7141 => x"00",
          7142 => x"00",
          7143 => x"00",
          7144 => x"00",
          7145 => x"00",
          7146 => x"00",
          7147 => x"00",
          7148 => x"00",
          7149 => x"00",
          7150 => x"00",
          7151 => x"00",
          7152 => x"00",
          7153 => x"00",
          7154 => x"00",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"00",
          7372 => x"6c",
          7373 => x"00",
          7374 => x"00",
          7375 => x"00",
          7376 => x"72",
          7377 => x"00",
          7378 => x"00",
          7379 => x"00",
          7380 => x"65",
          7381 => x"69",
          7382 => x"66",
          7383 => x"61",
          7384 => x"6d",
          7385 => x"72",
          7386 => x"00",
          7387 => x"00",
          7388 => x"00",
          7389 => x"38",
          7390 => x"63",
          7391 => x"63",
          7392 => x"00",
          7393 => x"6e",
          7394 => x"72",
          7395 => x"61",
          7396 => x"73",
          7397 => x"65",
          7398 => x"6f",
          7399 => x"6f",
          7400 => x"65",
          7401 => x"6e",
          7402 => x"65",
          7403 => x"72",
          7404 => x"69",
          7405 => x"6f",
          7406 => x"69",
          7407 => x"6f",
          7408 => x"6e",
          7409 => x"6c",
          7410 => x"6f",
          7411 => x"6f",
          7412 => x"6f",
          7413 => x"69",
          7414 => x"65",
          7415 => x"66",
          7416 => x"20",
          7417 => x"69",
          7418 => x"65",
          7419 => x"00",
          7420 => x"20",
          7421 => x"69",
          7422 => x"69",
          7423 => x"44",
          7424 => x"74",
          7425 => x"63",
          7426 => x"69",
          7427 => x"6c",
          7428 => x"69",
          7429 => x"69",
          7430 => x"61",
          7431 => x"74",
          7432 => x"63",
          7433 => x"6e",
          7434 => x"6e",
          7435 => x"69",
          7436 => x"00",
          7437 => x"74",
          7438 => x"2e",
          7439 => x"6c",
          7440 => x"2e",
          7441 => x"6e",
          7442 => x"79",
          7443 => x"6e",
          7444 => x"72",
          7445 => x"45",
          7446 => x"75",
          7447 => x"00",
          7448 => x"62",
          7449 => x"20",
          7450 => x"62",
          7451 => x"63",
          7452 => x"65",
          7453 => x"30",
          7454 => x"20",
          7455 => x"00",
          7456 => x"00",
          7457 => x"30",
          7458 => x"20",
          7459 => x"00",
          7460 => x"2a",
          7461 => x"36",
          7462 => x"31",
          7463 => x"00",
          7464 => x"20",
          7465 => x"78",
          7466 => x"20",
          7467 => x"50",
          7468 => x"72",
          7469 => x"64",
          7470 => x"41",
          7471 => x"69",
          7472 => x"74",
          7473 => x"20",
          7474 => x"72",
          7475 => x"41",
          7476 => x"69",
          7477 => x"74",
          7478 => x"20",
          7479 => x"72",
          7480 => x"4f",
          7481 => x"69",
          7482 => x"74",
          7483 => x"20",
          7484 => x"72",
          7485 => x"53",
          7486 => x"72",
          7487 => x"69",
          7488 => x"65",
          7489 => x"65",
          7490 => x"70",
          7491 => x"2e",
          7492 => x"69",
          7493 => x"72",
          7494 => x"75",
          7495 => x"62",
          7496 => x"4f",
          7497 => x"73",
          7498 => x"64",
          7499 => x"74",
          7500 => x"73",
          7501 => x"30",
          7502 => x"65",
          7503 => x"61",
          7504 => x"00",
          7505 => x"64",
          7506 => x"3a",
          7507 => x"6f",
          7508 => x"00",
          7509 => x"69",
          7510 => x"73",
          7511 => x"00",
          7512 => x"72",
          7513 => x"67",
          7514 => x"65",
          7515 => x"67",
          7516 => x"61",
          7517 => x"00",
          7518 => x"6e",
          7519 => x"40",
          7520 => x"2e",
          7521 => x"61",
          7522 => x"72",
          7523 => x"65",
          7524 => x"00",
          7525 => x"74",
          7526 => x"65",
          7527 => x"78",
          7528 => x"30",
          7529 => x"6c",
          7530 => x"30",
          7531 => x"58",
          7532 => x"72",
          7533 => x"00",
          7534 => x"28",
          7535 => x"25",
          7536 => x"38",
          7537 => x"6f",
          7538 => x"2e",
          7539 => x"20",
          7540 => x"6c",
          7541 => x"2e",
          7542 => x"75",
          7543 => x"72",
          7544 => x"6c",
          7545 => x"64",
          7546 => x"00",
          7547 => x"79",
          7548 => x"74",
          7549 => x"6e",
          7550 => x"65",
          7551 => x"61",
          7552 => x"3f",
          7553 => x"2f",
          7554 => x"64",
          7555 => x"64",
          7556 => x"6f",
          7557 => x"74",
          7558 => x"0a",
          7559 => x"20",
          7560 => x"6e",
          7561 => x"64",
          7562 => x"3a",
          7563 => x"50",
          7564 => x"20",
          7565 => x"41",
          7566 => x"3d",
          7567 => x"00",
          7568 => x"50",
          7569 => x"79",
          7570 => x"41",
          7571 => x"3d",
          7572 => x"00",
          7573 => x"74",
          7574 => x"72",
          7575 => x"73",
          7576 => x"3d",
          7577 => x"00",
          7578 => x"00",
          7579 => x"50",
          7580 => x"20",
          7581 => x"20",
          7582 => x"3d",
          7583 => x"00",
          7584 => x"79",
          7585 => x"6f",
          7586 => x"20",
          7587 => x"3d",
          7588 => x"64",
          7589 => x"20",
          7590 => x"6f",
          7591 => x"4d",
          7592 => x"46",
          7593 => x"2e",
          7594 => x"0a",
          7595 => x"44",
          7596 => x"63",
          7597 => x"20",
          7598 => x"3d",
          7599 => x"64",
          7600 => x"20",
          7601 => x"20",
          7602 => x"20",
          7603 => x"00",
          7604 => x"42",
          7605 => x"20",
          7606 => x"4f",
          7607 => x"00",
          7608 => x"4e",
          7609 => x"20",
          7610 => x"6c",
          7611 => x"2e",
          7612 => x"49",
          7613 => x"20",
          7614 => x"20",
          7615 => x"2e",
          7616 => x"44",
          7617 => x"20",
          7618 => x"73",
          7619 => x"2e",
          7620 => x"41",
          7621 => x"20",
          7622 => x"30",
          7623 => x"20",
          7624 => x"20",
          7625 => x"38",
          7626 => x"2e",
          7627 => x"4e",
          7628 => x"20",
          7629 => x"30",
          7630 => x"20",
          7631 => x"20",
          7632 => x"38",
          7633 => x"2e",
          7634 => x"42",
          7635 => x"20",
          7636 => x"30",
          7637 => x"28",
          7638 => x"43",
          7639 => x"29",
          7640 => x"77",
          7641 => x"00",
          7642 => x"00",
          7643 => x"6d",
          7644 => x"00",
          7645 => x"00",
          7646 => x"00",
          7647 => x"00",
          7648 => x"00",
          7649 => x"00",
          7650 => x"00",
          7651 => x"00",
          7652 => x"00",
          7653 => x"00",
          7654 => x"00",
          7655 => x"00",
          7656 => x"00",
          7657 => x"00",
          7658 => x"00",
          7659 => x"00",
          7660 => x"00",
          7661 => x"00",
          7662 => x"00",
          7663 => x"00",
          7664 => x"00",
          7665 => x"00",
          7666 => x"00",
          7667 => x"00",
          7668 => x"00",
          7669 => x"00",
          7670 => x"00",
          7671 => x"00",
          7672 => x"00",
          7673 => x"00",
          7674 => x"00",
          7675 => x"00",
          7676 => x"00",
          7677 => x"00",
          7678 => x"5b",
          7679 => x"5b",
          7680 => x"5b",
          7681 => x"5b",
          7682 => x"5b",
          7683 => x"5b",
          7684 => x"00",
          7685 => x"00",
          7686 => x"00",
          7687 => x"00",
          7688 => x"00",
          7689 => x"61",
          7690 => x"65",
          7691 => x"65",
          7692 => x"79",
          7693 => x"64",
          7694 => x"67",
          7695 => x"72",
          7696 => x"00",
          7697 => x"30",
          7698 => x"0a",
          7699 => x"64",
          7700 => x"65",
          7701 => x"69",
          7702 => x"69",
          7703 => x"4f",
          7704 => x"25",
          7705 => x"5b",
          7706 => x"5b",
          7707 => x"5b",
          7708 => x"5b",
          7709 => x"5b",
          7710 => x"5b",
          7711 => x"5b",
          7712 => x"5b",
          7713 => x"5b",
          7714 => x"5b",
          7715 => x"5b",
          7716 => x"5b",
          7717 => x"5b",
          7718 => x"5b",
          7719 => x"5b",
          7720 => x"5b",
          7721 => x"00",
          7722 => x"00",
          7723 => x"25",
          7724 => x"2c",
          7725 => x"30",
          7726 => x"3a",
          7727 => x"64",
          7728 => x"25",
          7729 => x"64",
          7730 => x"00",
          7731 => x"00",
          7732 => x"3b",
          7733 => x"65",
          7734 => x"72",
          7735 => x"70",
          7736 => x"30",
          7737 => x"77",
          7738 => x"30",
          7739 => x"64",
          7740 => x"00",
          7741 => x"73",
          7742 => x"65",
          7743 => x"44",
          7744 => x"3f",
          7745 => x"2c",
          7746 => x"41",
          7747 => x"00",
          7748 => x"44",
          7749 => x"4f",
          7750 => x"20",
          7751 => x"20",
          7752 => x"4d",
          7753 => x"54",
          7754 => x"00",
          7755 => x"00",
          7756 => x"03",
          7757 => x"16",
          7758 => x"9a",
          7759 => x"45",
          7760 => x"92",
          7761 => x"99",
          7762 => x"49",
          7763 => x"a9",
          7764 => x"b1",
          7765 => x"b9",
          7766 => x"c1",
          7767 => x"c9",
          7768 => x"d1",
          7769 => x"d9",
          7770 => x"e1",
          7771 => x"e9",
          7772 => x"f1",
          7773 => x"f9",
          7774 => x"2e",
          7775 => x"22",
          7776 => x"00",
          7777 => x"10",
          7778 => x"00",
          7779 => x"04",
          7780 => x"00",
          7781 => x"e9",
          7782 => x"e5",
          7783 => x"e8",
          7784 => x"c4",
          7785 => x"c6",
          7786 => x"fb",
          7787 => x"dc",
          7788 => x"a7",
          7789 => x"f3",
          7790 => x"aa",
          7791 => x"ac",
          7792 => x"ab",
          7793 => x"93",
          7794 => x"62",
          7795 => x"51",
          7796 => x"5b",
          7797 => x"2c",
          7798 => x"5e",
          7799 => x"69",
          7800 => x"6c",
          7801 => x"65",
          7802 => x"53",
          7803 => x"0c",
          7804 => x"90",
          7805 => x"93",
          7806 => x"b5",
          7807 => x"a9",
          7808 => x"b5",
          7809 => x"65",
          7810 => x"f7",
          7811 => x"b7",
          7812 => x"a0",
          7813 => x"e0",
          7814 => x"ff",
          7815 => x"30",
          7816 => x"10",
          7817 => x"06",
          7818 => x"81",
          7819 => x"84",
          7820 => x"89",
          7821 => x"8d",
          7822 => x"91",
          7823 => x"f6",
          7824 => x"98",
          7825 => x"9d",
          7826 => x"a0",
          7827 => x"a4",
          7828 => x"a9",
          7829 => x"ac",
          7830 => x"b1",
          7831 => x"b5",
          7832 => x"b8",
          7833 => x"bc",
          7834 => x"c1",
          7835 => x"c5",
          7836 => x"c7",
          7837 => x"cd",
          7838 => x"8e",
          7839 => x"03",
          7840 => x"f8",
          7841 => x"3a",
          7842 => x"3b",
          7843 => x"40",
          7844 => x"0a",
          7845 => x"86",
          7846 => x"58",
          7847 => x"5c",
          7848 => x"93",
          7849 => x"64",
          7850 => x"97",
          7851 => x"6c",
          7852 => x"70",
          7853 => x"74",
          7854 => x"78",
          7855 => x"7c",
          7856 => x"a6",
          7857 => x"84",
          7858 => x"ae",
          7859 => x"45",
          7860 => x"90",
          7861 => x"03",
          7862 => x"ac",
          7863 => x"89",
          7864 => x"c2",
          7865 => x"c4",
          7866 => x"8c",
          7867 => x"18",
          7868 => x"f3",
          7869 => x"f7",
          7870 => x"fa",
          7871 => x"10",
          7872 => x"36",
          7873 => x"01",
          7874 => x"61",
          7875 => x"7d",
          7876 => x"96",
          7877 => x"08",
          7878 => x"08",
          7879 => x"06",
          7880 => x"52",
          7881 => x"56",
          7882 => x"70",
          7883 => x"c8",
          7884 => x"da",
          7885 => x"ea",
          7886 => x"80",
          7887 => x"a0",
          7888 => x"b8",
          7889 => x"cc",
          7890 => x"02",
          7891 => x"01",
          7892 => x"fc",
          7893 => x"70",
          7894 => x"83",
          7895 => x"2f",
          7896 => x"06",
          7897 => x"64",
          7898 => x"1a",
          7899 => x"00",
          7900 => x"00",
          7901 => x"00",
          7902 => x"00",
          7903 => x"00",
          7904 => x"00",
          7905 => x"00",
          7906 => x"00",
          7907 => x"00",
          7908 => x"00",
          7909 => x"00",
          7910 => x"00",
          7911 => x"00",
          7912 => x"00",
          7913 => x"00",
          7914 => x"00",
          7915 => x"00",
          7916 => x"00",
          7917 => x"00",
          7918 => x"00",
          7919 => x"00",
          7920 => x"00",
          7921 => x"00",
          7922 => x"00",
          7923 => x"00",
          7924 => x"00",
          7925 => x"00",
          7926 => x"00",
          7927 => x"00",
          7928 => x"00",
          7929 => x"00",
          7930 => x"00",
          7931 => x"00",
          7932 => x"00",
          7933 => x"00",
          7934 => x"00",
          7935 => x"00",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"00",
          7940 => x"00",
          7941 => x"00",
          7942 => x"00",
          7943 => x"00",
          7944 => x"00",
          7945 => x"00",
          7946 => x"00",
          7947 => x"00",
          7948 => x"00",
          7949 => x"00",
          7950 => x"00",
          7951 => x"00",
          7952 => x"00",
          7953 => x"00",
          7954 => x"00",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"00",
          7959 => x"81",
          7960 => x"7f",
          7961 => x"00",
          7962 => x"00",
          7963 => x"f5",
          7964 => x"00",
          7965 => x"01",
          7966 => x"00",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"00",
          7980 => x"00",
          7981 => x"00",
          7982 => x"fc",
          7983 => x"7a",
          7984 => x"72",
          7985 => x"6a",
          7986 => x"62",
          7987 => x"32",
          7988 => x"f3",
          7989 => x"7f",
          7990 => x"f0",
          7991 => x"81",
          7992 => x"fc",
          7993 => x"5a",
          7994 => x"52",
          7995 => x"4a",
          7996 => x"42",
          7997 => x"32",
          7998 => x"f3",
          7999 => x"7f",
          8000 => x"f0",
          8001 => x"81",
          8002 => x"fc",
          8003 => x"5a",
          8004 => x"52",
          8005 => x"4a",
          8006 => x"42",
          8007 => x"22",
          8008 => x"7e",
          8009 => x"e2",
          8010 => x"f0",
          8011 => x"86",
          8012 => x"fe",
          8013 => x"1a",
          8014 => x"12",
          8015 => x"0a",
          8016 => x"02",
          8017 => x"f0",
          8018 => x"1e",
          8019 => x"f0",
          8020 => x"f0",
          8021 => x"81",
          8022 => x"f0",
          8023 => x"77",
          8024 => x"70",
          8025 => x"5d",
          8026 => x"6e",
          8027 => x"36",
          8028 => x"9f",
          8029 => x"c5",
          8030 => x"f0",
          8031 => x"81",
          8032 => x"00",
          8033 => x"00",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"00",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"cf",
          9069 => x"fd",
          9070 => x"c5",
          9071 => x"ee",
          9072 => x"65",
          9073 => x"2a",
          9074 => x"25",
          9075 => x"2b",
          9076 => x"05",
          9077 => x"0d",
          9078 => x"15",
          9079 => x"54",
          9080 => x"85",
          9081 => x"8d",
          9082 => x"95",
          9083 => x"40",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"04",
          9100 => x"04",
        others => X"00"
    );

    shared variable RAM7 : ramArray :=
    (
             0 => x"f8",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"90",
             5 => x"8c",
             6 => x"00",
             7 => x"00",
             8 => x"72",
             9 => x"83",
            10 => x"04",
            11 => x"00",
            12 => x"83",
            13 => x"05",
            14 => x"73",
            15 => x"83",
            16 => x"72",
            17 => x"73",
            18 => x"53",
            19 => x"00",
            20 => x"73",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"0a",
            26 => x"05",
            27 => x"04",
            28 => x"73",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"cd",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"0a",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"09",
            45 => x"05",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"81",
            50 => x"04",
            51 => x"00",
            52 => x"04",
            53 => x"82",
            54 => x"fc",
            55 => x"00",
            56 => x"72",
            57 => x"0a",
            58 => x"00",
            59 => x"00",
            60 => x"72",
            61 => x"0a",
            62 => x"00",
            63 => x"00",
            64 => x"52",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"05",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"73",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"72",
            77 => x"10",
            78 => x"04",
            79 => x"00",
            80 => x"0b",
            81 => x"10",
            82 => x"93",
            83 => x"00",
            84 => x"90",
            85 => x"cc",
            86 => x"0c",
            87 => x"00",
            88 => x"90",
            89 => x"ab",
            90 => x"0c",
            91 => x"00",
            92 => x"05",
            93 => x"70",
            94 => x"05",
            95 => x"04",
            96 => x"05",
            97 => x"05",
            98 => x"74",
            99 => x"51",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"04",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"10",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"05",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"81",
           133 => x"0b",
           134 => x"0b",
           135 => x"b6",
           136 => x"0b",
           137 => x"0b",
           138 => x"f6",
           139 => x"0b",
           140 => x"0b",
           141 => x"b6",
           142 => x"0b",
           143 => x"0b",
           144 => x"f9",
           145 => x"0b",
           146 => x"0b",
           147 => x"bd",
           148 => x"0b",
           149 => x"0b",
           150 => x"81",
           151 => x"0b",
           152 => x"0b",
           153 => x"c5",
           154 => x"0b",
           155 => x"0b",
           156 => x"89",
           157 => x"0b",
           158 => x"0b",
           159 => x"cd",
           160 => x"0b",
           161 => x"0b",
           162 => x"91",
           163 => x"0b",
           164 => x"0b",
           165 => x"d5",
           166 => x"0b",
           167 => x"0b",
           168 => x"99",
           169 => x"0b",
           170 => x"0b",
           171 => x"dc",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"04",
           193 => x"2d",
           194 => x"90",
           195 => x"2d",
           196 => x"90",
           197 => x"2d",
           198 => x"90",
           199 => x"2d",
           200 => x"90",
           201 => x"2d",
           202 => x"90",
           203 => x"2d",
           204 => x"90",
           205 => x"2d",
           206 => x"90",
           207 => x"2d",
           208 => x"90",
           209 => x"2d",
           210 => x"90",
           211 => x"2d",
           212 => x"90",
           213 => x"2d",
           214 => x"90",
           215 => x"2d",
           216 => x"90",
           217 => x"d1",
           218 => x"80",
           219 => x"d5",
           220 => x"c0",
           221 => x"80",
           222 => x"80",
           223 => x"0c",
           224 => x"08",
           225 => x"f0",
           226 => x"f0",
           227 => x"b8",
           228 => x"b8",
           229 => x"84",
           230 => x"84",
           231 => x"04",
           232 => x"2d",
           233 => x"90",
           234 => x"8c",
           235 => x"80",
           236 => x"fa",
           237 => x"c0",
           238 => x"82",
           239 => x"80",
           240 => x"0c",
           241 => x"08",
           242 => x"f0",
           243 => x"f0",
           244 => x"b8",
           245 => x"b8",
           246 => x"84",
           247 => x"84",
           248 => x"04",
           249 => x"2d",
           250 => x"90",
           251 => x"f5",
           252 => x"80",
           253 => x"f5",
           254 => x"c0",
           255 => x"83",
           256 => x"80",
           257 => x"0c",
           258 => x"08",
           259 => x"f0",
           260 => x"f0",
           261 => x"b8",
           262 => x"b8",
           263 => x"84",
           264 => x"84",
           265 => x"04",
           266 => x"2d",
           267 => x"90",
           268 => x"89",
           269 => x"80",
           270 => x"99",
           271 => x"c0",
           272 => x"83",
           273 => x"80",
           274 => x"0c",
           275 => x"08",
           276 => x"f0",
           277 => x"f0",
           278 => x"b8",
           279 => x"b8",
           280 => x"84",
           281 => x"84",
           282 => x"04",
           283 => x"2d",
           284 => x"90",
           285 => x"d1",
           286 => x"80",
           287 => x"f5",
           288 => x"c0",
           289 => x"80",
           290 => x"80",
           291 => x"0c",
           292 => x"08",
           293 => x"f0",
           294 => x"f0",
           295 => x"b8",
           296 => x"f0",
           297 => x"b8",
           298 => x"b8",
           299 => x"84",
           300 => x"84",
           301 => x"04",
           302 => x"2d",
           303 => x"90",
           304 => x"80",
           305 => x"80",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"00",
           311 => x"09",
           312 => x"2b",
           313 => x"04",
           314 => x"05",
           315 => x"72",
           316 => x"51",
           317 => x"70",
           318 => x"71",
           319 => x"0b",
           320 => x"ce",
           321 => x"3d",
           322 => x"53",
           323 => x"81",
           324 => x"3d",
           325 => x"81",
           326 => x"56",
           327 => x"2e",
           328 => x"14",
           329 => x"72",
           330 => x"54",
           331 => x"2e",
           332 => x"84",
           333 => x"08",
           334 => x"08",
           335 => x"14",
           336 => x"07",
           337 => x"80",
           338 => x"52",
           339 => x"0d",
           340 => x"88",
           341 => x"54",
           342 => x"73",
           343 => x"05",
           344 => x"51",
           345 => x"34",
           346 => x"86",
           347 => x"51",
           348 => x"3d",
           349 => x"80",
           350 => x"70",
           351 => x"55",
           352 => x"81",
           353 => x"76",
           354 => x"7b",
           355 => x"81",
           356 => x"26",
           357 => x"30",
           358 => x"ae",
           359 => x"83",
           360 => x"54",
           361 => x"80",
           362 => x"bd",
           363 => x"b8",
           364 => x"83",
           365 => x"10",
           366 => x"19",
           367 => x"05",
           368 => x"5f",
           369 => x"81",
           370 => x"7c",
           371 => x"ff",
           372 => x"06",
           373 => x"5b",
           374 => x"dd",
           375 => x"51",
           376 => x"fe",
           377 => x"2a",
           378 => x"38",
           379 => x"95",
           380 => x"26",
           381 => x"f4",
           382 => x"18",
           383 => x"38",
           384 => x"80",
           385 => x"38",
           386 => x"f6",
           387 => x"71",
           388 => x"58",
           389 => x"52",
           390 => x"e4",
           391 => x"08",
           392 => x"26",
           393 => x"05",
           394 => x"34",
           395 => x"84",
           396 => x"08",
           397 => x"98",
           398 => x"80",
           399 => x"29",
           400 => x"59",
           401 => x"55",
           402 => x"84",
           403 => x"53",
           404 => x"80",
           405 => x"72",
           406 => x"81",
           407 => x"38",
           408 => x"54",
           409 => x"7a",
           410 => x"71",
           411 => x"06",
           412 => x"77",
           413 => x"7c",
           414 => x"80",
           415 => x"81",
           416 => x"84",
           417 => x"38",
           418 => x"86",
           419 => x"85",
           420 => x"5f",
           421 => x"84",
           422 => x"70",
           423 => x"25",
           424 => x"a9",
           425 => x"fc",
           426 => x"40",
           427 => x"81",
           428 => x"78",
           429 => x"0a",
           430 => x"80",
           431 => x"51",
           432 => x"0a",
           433 => x"2c",
           434 => x"38",
           435 => x"55",
           436 => x"80",
           437 => x"f3",
           438 => x"2e",
           439 => x"2e",
           440 => x"33",
           441 => x"b8",
           442 => x"74",
           443 => x"a7",
           444 => x"fc",
           445 => x"40",
           446 => x"7c",
           447 => x"39",
           448 => x"7c",
           449 => x"fa",
           450 => x"80",
           451 => x"71",
           452 => x"59",
           453 => x"60",
           454 => x"83",
           455 => x"7c",
           456 => x"05",
           457 => x"57",
           458 => x"06",
           459 => x"78",
           460 => x"05",
           461 => x"7f",
           462 => x"51",
           463 => x"70",
           464 => x"83",
           465 => x"52",
           466 => x"85",
           467 => x"83",
           468 => x"ff",
           469 => x"75",
           470 => x"b9",
           471 => x"81",
           472 => x"29",
           473 => x"5a",
           474 => x"70",
           475 => x"c6",
           476 => x"05",
           477 => x"80",
           478 => x"ff",
           479 => x"fa",
           480 => x"58",
           481 => x"39",
           482 => x"58",
           483 => x"39",
           484 => x"81",
           485 => x"8a",
           486 => x"b8",
           487 => x"71",
           488 => x"2c",
           489 => x"07",
           490 => x"38",
           491 => x"71",
           492 => x"54",
           493 => x"bb",
           494 => x"ff",
           495 => x"5a",
           496 => x"33",
           497 => x"c9",
           498 => x"fc",
           499 => x"54",
           500 => x"7c",
           501 => x"39",
           502 => x"79",
           503 => x"38",
           504 => x"7a",
           505 => x"2e",
           506 => x"98",
           507 => x"90",
           508 => x"51",
           509 => x"39",
           510 => x"7e",
           511 => x"a2",
           512 => x"98",
           513 => x"06",
           514 => x"fb",
           515 => x"70",
           516 => x"7c",
           517 => x"39",
           518 => x"ff",
           519 => x"8b",
           520 => x"ff",
           521 => x"5a",
           522 => x"30",
           523 => x"5b",
           524 => x"d4",
           525 => x"f3",
           526 => x"3d",
           527 => x"c8",
           528 => x"81",
           529 => x"55",
           530 => x"81",
           531 => x"05",
           532 => x"38",
           533 => x"90",
           534 => x"e4",
           535 => x"74",
           536 => x"80",
           537 => x"54",
           538 => x"84",
           539 => x"14",
           540 => x"08",
           541 => x"56",
           542 => x"0d",
           543 => x"54",
           544 => x"2a",
           545 => x"57",
           546 => x"81",
           547 => x"55",
           548 => x"06",
           549 => x"e4",
           550 => x"81",
           551 => x"ea",
           552 => x"08",
           553 => x"80",
           554 => x"05",
           555 => x"ca",
           556 => x"08",
           557 => x"0d",
           558 => x"11",
           559 => x"06",
           560 => x"ae",
           561 => x"73",
           562 => x"53",
           563 => x"74",
           564 => x"81",
           565 => x"81",
           566 => x"84",
           567 => x"74",
           568 => x"15",
           569 => x"b8",
           570 => x"81",
           571 => x"39",
           572 => x"70",
           573 => x"06",
           574 => x"b3",
           575 => x"71",
           576 => x"52",
           577 => x"08",
           578 => x"80",
           579 => x"16",
           580 => x"81",
           581 => x"0c",
           582 => x"06",
           583 => x"08",
           584 => x"33",
           585 => x"04",
           586 => x"2d",
           587 => x"e4",
           588 => x"16",
           589 => x"b8",
           590 => x"a0",
           591 => x"54",
           592 => x"0d",
           593 => x"17",
           594 => x"0d",
           595 => x"70",
           596 => x"38",
           597 => x"54",
           598 => x"54",
           599 => x"e4",
           600 => x"0d",
           601 => x"54",
           602 => x"27",
           603 => x"71",
           604 => x"81",
           605 => x"ef",
           606 => x"3d",
           607 => x"27",
           608 => x"ff",
           609 => x"73",
           610 => x"d9",
           611 => x"71",
           612 => x"df",
           613 => x"70",
           614 => x"33",
           615 => x"74",
           616 => x"3d",
           617 => x"71",
           618 => x"54",
           619 => x"54",
           620 => x"e4",
           621 => x"0d",
           622 => x"54",
           623 => x"81",
           624 => x"55",
           625 => x"73",
           626 => x"04",
           627 => x"56",
           628 => x"33",
           629 => x"52",
           630 => x"38",
           631 => x"38",
           632 => x"51",
           633 => x"0d",
           634 => x"33",
           635 => x"38",
           636 => x"80",
           637 => x"b8",
           638 => x"84",
           639 => x"fb",
           640 => x"56",
           641 => x"84",
           642 => x"81",
           643 => x"54",
           644 => x"38",
           645 => x"74",
           646 => x"e4",
           647 => x"e4",
           648 => x"87",
           649 => x"77",
           650 => x"80",
           651 => x"54",
           652 => x"ff",
           653 => x"06",
           654 => x"52",
           655 => x"3d",
           656 => x"79",
           657 => x"2e",
           658 => x"54",
           659 => x"73",
           660 => x"04",
           661 => x"a0",
           662 => x"51",
           663 => x"52",
           664 => x"38",
           665 => x"b8",
           666 => x"9f",
           667 => x"9f",
           668 => x"71",
           669 => x"57",
           670 => x"2e",
           671 => x"07",
           672 => x"ff",
           673 => x"72",
           674 => x"56",
           675 => x"da",
           676 => x"84",
           677 => x"fc",
           678 => x"06",
           679 => x"70",
           680 => x"2a",
           681 => x"70",
           682 => x"74",
           683 => x"30",
           684 => x"31",
           685 => x"05",
           686 => x"25",
           687 => x"70",
           688 => x"70",
           689 => x"05",
           690 => x"55",
           691 => x"55",
           692 => x"56",
           693 => x"3d",
           694 => x"54",
           695 => x"08",
           696 => x"e4",
           697 => x"3d",
           698 => x"76",
           699 => x"cf",
           700 => x"13",
           701 => x"51",
           702 => x"08",
           703 => x"80",
           704 => x"be",
           705 => x"72",
           706 => x"55",
           707 => x"72",
           708 => x"77",
           709 => x"2c",
           710 => x"71",
           711 => x"55",
           712 => x"84",
           713 => x"fa",
           714 => x"2c",
           715 => x"2c",
           716 => x"31",
           717 => x"59",
           718 => x"e4",
           719 => x"e4",
           720 => x"0d",
           721 => x"0c",
           722 => x"73",
           723 => x"81",
           724 => x"55",
           725 => x"2e",
           726 => x"83",
           727 => x"89",
           728 => x"56",
           729 => x"e0",
           730 => x"81",
           731 => x"81",
           732 => x"8f",
           733 => x"54",
           734 => x"72",
           735 => x"29",
           736 => x"33",
           737 => x"be",
           738 => x"30",
           739 => x"84",
           740 => x"81",
           741 => x"56",
           742 => x"06",
           743 => x"0c",
           744 => x"2e",
           745 => x"2e",
           746 => x"c6",
           747 => x"58",
           748 => x"84",
           749 => x"82",
           750 => x"33",
           751 => x"80",
           752 => x"0d",
           753 => x"57",
           754 => x"33",
           755 => x"81",
           756 => x"0c",
           757 => x"f3",
           758 => x"73",
           759 => x"58",
           760 => x"38",
           761 => x"80",
           762 => x"38",
           763 => x"53",
           764 => x"53",
           765 => x"70",
           766 => x"27",
           767 => x"83",
           768 => x"70",
           769 => x"73",
           770 => x"2e",
           771 => x"0c",
           772 => x"8b",
           773 => x"79",
           774 => x"b0",
           775 => x"81",
           776 => x"55",
           777 => x"58",
           778 => x"56",
           779 => x"53",
           780 => x"fe",
           781 => x"8b",
           782 => x"70",
           783 => x"56",
           784 => x"e4",
           785 => x"d1",
           786 => x"06",
           787 => x"0d",
           788 => x"71",
           789 => x"71",
           790 => x"be",
           791 => x"9c",
           792 => x"04",
           793 => x"83",
           794 => x"ef",
           795 => x"ce",
           796 => x"0d",
           797 => x"3f",
           798 => x"51",
           799 => x"83",
           800 => x"3d",
           801 => x"e6",
           802 => x"e0",
           803 => x"04",
           804 => x"83",
           805 => x"ee",
           806 => x"d0",
           807 => x"0d",
           808 => x"3f",
           809 => x"51",
           810 => x"83",
           811 => x"3d",
           812 => x"8e",
           813 => x"88",
           814 => x"04",
           815 => x"83",
           816 => x"ed",
           817 => x"d1",
           818 => x"0d",
           819 => x"05",
           820 => x"68",
           821 => x"51",
           822 => x"ff",
           823 => x"07",
           824 => x"57",
           825 => x"52",
           826 => x"c8",
           827 => x"b8",
           828 => x"77",
           829 => x"70",
           830 => x"9f",
           831 => x"77",
           832 => x"88",
           833 => x"e0",
           834 => x"51",
           835 => x"54",
           836 => x"d1",
           837 => x"b8",
           838 => x"b8",
           839 => x"84",
           840 => x"05",
           841 => x"51",
           842 => x"08",
           843 => x"38",
           844 => x"38",
           845 => x"39",
           846 => x"3f",
           847 => x"f4",
           848 => x"83",
           849 => x"c0",
           850 => x"f8",
           851 => x"05",
           852 => x"7b",
           853 => x"b8",
           854 => x"91",
           855 => x"84",
           856 => x"78",
           857 => x"60",
           858 => x"7e",
           859 => x"84",
           860 => x"f3",
           861 => x"05",
           862 => x"68",
           863 => x"78",
           864 => x"83",
           865 => x"d1",
           866 => x"73",
           867 => x"81",
           868 => x"38",
           869 => x"a7",
           870 => x"51",
           871 => x"c8",
           872 => x"3f",
           873 => x"80",
           874 => x"79",
           875 => x"33",
           876 => x"83",
           877 => x"27",
           878 => x"70",
           879 => x"2e",
           880 => x"ee",
           881 => x"51",
           882 => x"76",
           883 => x"e9",
           884 => x"58",
           885 => x"e4",
           886 => x"54",
           887 => x"9b",
           888 => x"76",
           889 => x"84",
           890 => x"83",
           891 => x"14",
           892 => x"51",
           893 => x"b8",
           894 => x"51",
           895 => x"c8",
           896 => x"3f",
           897 => x"18",
           898 => x"22",
           899 => x"3f",
           900 => x"54",
           901 => x"26",
           902 => x"94",
           903 => x"d4",
           904 => x"a9",
           905 => x"73",
           906 => x"72",
           907 => x"ab",
           908 => x"53",
           909 => x"74",
           910 => x"d4",
           911 => x"3f",
           912 => x"ce",
           913 => x"ff",
           914 => x"fc",
           915 => x"2e",
           916 => x"59",
           917 => x"3f",
           918 => x"98",
           919 => x"9b",
           920 => x"75",
           921 => x"58",
           922 => x"80",
           923 => x"08",
           924 => x"32",
           925 => x"70",
           926 => x"55",
           927 => x"24",
           928 => x"0b",
           929 => x"04",
           930 => x"08",
           931 => x"ed",
           932 => x"3f",
           933 => x"2a",
           934 => x"b7",
           935 => x"51",
           936 => x"2a",
           937 => x"db",
           938 => x"51",
           939 => x"2a",
           940 => x"ff",
           941 => x"51",
           942 => x"2a",
           943 => x"38",
           944 => x"88",
           945 => x"04",
           946 => x"f4",
           947 => x"ed",
           948 => x"04",
           949 => x"88",
           950 => x"d5",
           951 => x"72",
           952 => x"51",
           953 => x"9b",
           954 => x"72",
           955 => x"71",
           956 => x"81",
           957 => x"51",
           958 => x"3f",
           959 => x"52",
           960 => x"be",
           961 => x"d3",
           962 => x"9a",
           963 => x"06",
           964 => x"38",
           965 => x"3f",
           966 => x"80",
           967 => x"70",
           968 => x"fe",
           969 => x"9a",
           970 => x"cd",
           971 => x"83",
           972 => x"80",
           973 => x"81",
           974 => x"51",
           975 => x"3f",
           976 => x"52",
           977 => x"bd",
           978 => x"41",
           979 => x"81",
           980 => x"84",
           981 => x"3d",
           982 => x"38",
           983 => x"98",
           984 => x"c3",
           985 => x"52",
           986 => x"83",
           987 => x"5b",
           988 => x"79",
           989 => x"ff",
           990 => x"38",
           991 => x"83",
           992 => x"2e",
           993 => x"70",
           994 => x"38",
           995 => x"7b",
           996 => x"08",
           997 => x"e4",
           998 => x"53",
           999 => x"84",
          1000 => x"33",
          1001 => x"81",
          1002 => x"9b",
          1003 => x"5c",
          1004 => x"f8",
          1005 => x"b8",
          1006 => x"80",
          1007 => x"08",
          1008 => x"91",
          1009 => x"62",
          1010 => x"84",
          1011 => x"8b",
          1012 => x"80",
          1013 => x"5b",
          1014 => x"82",
          1015 => x"82",
          1016 => x"d5",
          1017 => x"83",
          1018 => x"7d",
          1019 => x"0a",
          1020 => x"f5",
          1021 => x"b8",
          1022 => x"07",
          1023 => x"5a",
          1024 => x"78",
          1025 => x"38",
          1026 => x"5a",
          1027 => x"61",
          1028 => x"38",
          1029 => x"51",
          1030 => x"51",
          1031 => x"53",
          1032 => x"0b",
          1033 => x"ff",
          1034 => x"81",
          1035 => x"f4",
          1036 => x"e4",
          1037 => x"0b",
          1038 => x"53",
          1039 => x"b7",
          1040 => x"a0",
          1041 => x"e6",
          1042 => x"70",
          1043 => x"2e",
          1044 => x"39",
          1045 => x"3f",
          1046 => x"34",
          1047 => x"7e",
          1048 => x"5a",
          1049 => x"1a",
          1050 => x"81",
          1051 => x"10",
          1052 => x"04",
          1053 => x"51",
          1054 => x"84",
          1055 => x"84",
          1056 => x"06",
          1057 => x"45",
          1058 => x"98",
          1059 => x"92",
          1060 => x"a8",
          1061 => x"80",
          1062 => x"d2",
          1063 => x"9a",
          1064 => x"fa",
          1065 => x"93",
          1066 => x"3f",
          1067 => x"de",
          1068 => x"d5",
          1069 => x"3f",
          1070 => x"11",
          1071 => x"3f",
          1072 => x"ba",
          1073 => x"d0",
          1074 => x"b8",
          1075 => x"84",
          1076 => x"51",
          1077 => x"3d",
          1078 => x"51",
          1079 => x"80",
          1080 => x"d6",
          1081 => x"78",
          1082 => x"ff",
          1083 => x"b8",
          1084 => x"b8",
          1085 => x"05",
          1086 => x"08",
          1087 => x"53",
          1088 => x"83",
          1089 => x"f8",
          1090 => x"48",
          1091 => x"a2",
          1092 => x"64",
          1093 => x"b8",
          1094 => x"05",
          1095 => x"08",
          1096 => x"fe",
          1097 => x"e8",
          1098 => x"b0",
          1099 => x"52",
          1100 => x"84",
          1101 => x"7e",
          1102 => x"33",
          1103 => x"78",
          1104 => x"05",
          1105 => x"ff",
          1106 => x"e9",
          1107 => x"2e",
          1108 => x"11",
          1109 => x"3f",
          1110 => x"8a",
          1111 => x"ff",
          1112 => x"b8",
          1113 => x"83",
          1114 => x"67",
          1115 => x"38",
          1116 => x"5a",
          1117 => x"79",
          1118 => x"d6",
          1119 => x"5b",
          1120 => x"d2",
          1121 => x"ff",
          1122 => x"b8",
          1123 => x"b8",
          1124 => x"05",
          1125 => x"08",
          1126 => x"fe",
          1127 => x"e8",
          1128 => x"2e",
          1129 => x"cd",
          1130 => x"82",
          1131 => x"05",
          1132 => x"46",
          1133 => x"53",
          1134 => x"84",
          1135 => x"38",
          1136 => x"80",
          1137 => x"e4",
          1138 => x"52",
          1139 => x"84",
          1140 => x"7e",
          1141 => x"33",
          1142 => x"78",
          1143 => x"05",
          1144 => x"db",
          1145 => x"49",
          1146 => x"80",
          1147 => x"e4",
          1148 => x"59",
          1149 => x"68",
          1150 => x"11",
          1151 => x"3f",
          1152 => x"f5",
          1153 => x"53",
          1154 => x"84",
          1155 => x"38",
          1156 => x"80",
          1157 => x"e4",
          1158 => x"3d",
          1159 => x"51",
          1160 => x"86",
          1161 => x"d7",
          1162 => x"5b",
          1163 => x"5b",
          1164 => x"79",
          1165 => x"f1",
          1166 => x"80",
          1167 => x"e4",
          1168 => x"59",
          1169 => x"e4",
          1170 => x"84",
          1171 => x"38",
          1172 => x"3f",
          1173 => x"11",
          1174 => x"3f",
          1175 => x"f1",
          1176 => x"c0",
          1177 => x"3d",
          1178 => x"51",
          1179 => x"91",
          1180 => x"80",
          1181 => x"08",
          1182 => x"ff",
          1183 => x"b8",
          1184 => x"66",
          1185 => x"81",
          1186 => x"72",
          1187 => x"5d",
          1188 => x"2e",
          1189 => x"51",
          1190 => x"65",
          1191 => x"3f",
          1192 => x"f2",
          1193 => x"64",
          1194 => x"11",
          1195 => x"3f",
          1196 => x"da",
          1197 => x"84",
          1198 => x"53",
          1199 => x"84",
          1200 => x"39",
          1201 => x"7e",
          1202 => x"b8",
          1203 => x"05",
          1204 => x"08",
          1205 => x"02",
          1206 => x"05",
          1207 => x"f0",
          1208 => x"bd",
          1209 => x"38",
          1210 => x"11",
          1211 => x"3f",
          1212 => x"dc",
          1213 => x"33",
          1214 => x"9b",
          1215 => x"ff",
          1216 => x"b8",
          1217 => x"64",
          1218 => x"70",
          1219 => x"2e",
          1220 => x"55",
          1221 => x"d7",
          1222 => x"f3",
          1223 => x"8a",
          1224 => x"51",
          1225 => x"3d",
          1226 => x"51",
          1227 => x"80",
          1228 => x"ce",
          1229 => x"23",
          1230 => x"e9",
          1231 => x"38",
          1232 => x"39",
          1233 => x"2e",
          1234 => x"fc",
          1235 => x"d6",
          1236 => x"d8",
          1237 => x"f6",
          1238 => x"78",
          1239 => x"08",
          1240 => x"51",
          1241 => x"f1",
          1242 => x"38",
          1243 => x"39",
          1244 => x"2e",
          1245 => x"fb",
          1246 => x"7d",
          1247 => x"08",
          1248 => x"33",
          1249 => x"f1",
          1250 => x"f1",
          1251 => x"38",
          1252 => x"39",
          1253 => x"49",
          1254 => x"88",
          1255 => x"0d",
          1256 => x"c0",
          1257 => x"84",
          1258 => x"84",
          1259 => x"57",
          1260 => x"da",
          1261 => x"07",
          1262 => x"08",
          1263 => x"51",
          1264 => x"90",
          1265 => x"80",
          1266 => x"84",
          1267 => x"80",
          1268 => x"8c",
          1269 => x"0c",
          1270 => x"5d",
          1271 => x"80",
          1272 => x"70",
          1273 => x"d4",
          1274 => x"83",
          1275 => x"94",
          1276 => x"d2",
          1277 => x"d4",
          1278 => x"83",
          1279 => x"81",
          1280 => x"c4",
          1281 => x"3f",
          1282 => x"08",
          1283 => x"73",
          1284 => x"81",
          1285 => x"09",
          1286 => x"33",
          1287 => x"70",
          1288 => x"06",
          1289 => x"74",
          1290 => x"80",
          1291 => x"54",
          1292 => x"54",
          1293 => x"2e",
          1294 => x"80",
          1295 => x"a0",
          1296 => x"54",
          1297 => x"25",
          1298 => x"2e",
          1299 => x"54",
          1300 => x"84",
          1301 => x"70",
          1302 => x"ff",
          1303 => x"33",
          1304 => x"70",
          1305 => x"39",
          1306 => x"72",
          1307 => x"38",
          1308 => x"72",
          1309 => x"e4",
          1310 => x"fc",
          1311 => x"84",
          1312 => x"74",
          1313 => x"04",
          1314 => x"ff",
          1315 => x"26",
          1316 => x"05",
          1317 => x"8a",
          1318 => x"70",
          1319 => x"33",
          1320 => x"f2",
          1321 => x"74",
          1322 => x"22",
          1323 => x"80",
          1324 => x"52",
          1325 => x"81",
          1326 => x"22",
          1327 => x"33",
          1328 => x"33",
          1329 => x"33",
          1330 => x"33",
          1331 => x"33",
          1332 => x"c0",
          1333 => x"a0",
          1334 => x"0c",
          1335 => x"86",
          1336 => x"5b",
          1337 => x"0c",
          1338 => x"7b",
          1339 => x"7b",
          1340 => x"08",
          1341 => x"98",
          1342 => x"87",
          1343 => x"1c",
          1344 => x"7b",
          1345 => x"08",
          1346 => x"98",
          1347 => x"80",
          1348 => x"59",
          1349 => x"1b",
          1350 => x"1b",
          1351 => x"1b",
          1352 => x"52",
          1353 => x"3f",
          1354 => x"02",
          1355 => x"a8",
          1356 => x"84",
          1357 => x"2c",
          1358 => x"06",
          1359 => x"71",
          1360 => x"04",
          1361 => x"b8",
          1362 => x"51",
          1363 => x"df",
          1364 => x"84",
          1365 => x"2c",
          1366 => x"c7",
          1367 => x"52",
          1368 => x"e7",
          1369 => x"2b",
          1370 => x"2e",
          1371 => x"54",
          1372 => x"84",
          1373 => x"fc",
          1374 => x"f1",
          1375 => x"55",
          1376 => x"87",
          1377 => x"70",
          1378 => x"2e",
          1379 => x"06",
          1380 => x"32",
          1381 => x"38",
          1382 => x"cf",
          1383 => x"c0",
          1384 => x"38",
          1385 => x"0c",
          1386 => x"0d",
          1387 => x"51",
          1388 => x"81",
          1389 => x"71",
          1390 => x"2e",
          1391 => x"70",
          1392 => x"52",
          1393 => x"0d",
          1394 => x"9f",
          1395 => x"9c",
          1396 => x"0d",
          1397 => x"52",
          1398 => x"81",
          1399 => x"ff",
          1400 => x"80",
          1401 => x"70",
          1402 => x"52",
          1403 => x"2a",
          1404 => x"38",
          1405 => x"80",
          1406 => x"06",
          1407 => x"06",
          1408 => x"80",
          1409 => x"52",
          1410 => x"55",
          1411 => x"b8",
          1412 => x"91",
          1413 => x"98",
          1414 => x"72",
          1415 => x"81",
          1416 => x"38",
          1417 => x"2a",
          1418 => x"ce",
          1419 => x"c0",
          1420 => x"06",
          1421 => x"38",
          1422 => x"a0",
          1423 => x"f1",
          1424 => x"83",
          1425 => x"08",
          1426 => x"9c",
          1427 => x"9e",
          1428 => x"c0",
          1429 => x"87",
          1430 => x"0c",
          1431 => x"c0",
          1432 => x"f1",
          1433 => x"83",
          1434 => x"08",
          1435 => x"c4",
          1436 => x"9e",
          1437 => x"23",
          1438 => x"d8",
          1439 => x"f1",
          1440 => x"83",
          1441 => x"e4",
          1442 => x"08",
          1443 => x"52",
          1444 => x"e5",
          1445 => x"08",
          1446 => x"52",
          1447 => x"71",
          1448 => x"c0",
          1449 => x"06",
          1450 => x"38",
          1451 => x"80",
          1452 => x"88",
          1453 => x"80",
          1454 => x"f1",
          1455 => x"90",
          1456 => x"52",
          1457 => x"52",
          1458 => x"87",
          1459 => x"80",
          1460 => x"83",
          1461 => x"34",
          1462 => x"70",
          1463 => x"70",
          1464 => x"83",
          1465 => x"9e",
          1466 => x"51",
          1467 => x"81",
          1468 => x"0b",
          1469 => x"80",
          1470 => x"2e",
          1471 => x"ed",
          1472 => x"08",
          1473 => x"52",
          1474 => x"71",
          1475 => x"c0",
          1476 => x"51",
          1477 => x"81",
          1478 => x"c0",
          1479 => x"8a",
          1480 => x"34",
          1481 => x"70",
          1482 => x"80",
          1483 => x"f1",
          1484 => x"83",
          1485 => x"71",
          1486 => x"c0",
          1487 => x"52",
          1488 => x"52",
          1489 => x"9e",
          1490 => x"f1",
          1491 => x"52",
          1492 => x"d8",
          1493 => x"f1",
          1494 => x"83",
          1495 => x"f1",
          1496 => x"83",
          1497 => x"38",
          1498 => x"a8",
          1499 => x"84",
          1500 => x"73",
          1501 => x"56",
          1502 => x"33",
          1503 => x"f1",
          1504 => x"f1",
          1505 => x"83",
          1506 => x"38",
          1507 => x"93",
          1508 => x"82",
          1509 => x"73",
          1510 => x"c2",
          1511 => x"83",
          1512 => x"83",
          1513 => x"51",
          1514 => x"08",
          1515 => x"ab",
          1516 => x"3f",
          1517 => x"d8",
          1518 => x"d8",
          1519 => x"51",
          1520 => x"bd",
          1521 => x"54",
          1522 => x"80",
          1523 => x"eb",
          1524 => x"f1",
          1525 => x"51",
          1526 => x"83",
          1527 => x"52",
          1528 => x"e4",
          1529 => x"31",
          1530 => x"83",
          1531 => x"8a",
          1532 => x"04",
          1533 => x"c0",
          1534 => x"b8",
          1535 => x"71",
          1536 => x"52",
          1537 => x"3f",
          1538 => x"2e",
          1539 => x"db",
          1540 => x"cc",
          1541 => x"08",
          1542 => x"d3",
          1543 => x"d9",
          1544 => x"f1",
          1545 => x"ff",
          1546 => x"c0",
          1547 => x"83",
          1548 => x"83",
          1549 => x"52",
          1550 => x"e4",
          1551 => x"31",
          1552 => x"83",
          1553 => x"83",
          1554 => x"fe",
          1555 => x"8c",
          1556 => x"ee",
          1557 => x"38",
          1558 => x"ff",
          1559 => x"56",
          1560 => x"39",
          1561 => x"3f",
          1562 => x"2e",
          1563 => x"ac",
          1564 => x"e7",
          1565 => x"38",
          1566 => x"83",
          1567 => x"83",
          1568 => x"fc",
          1569 => x"33",
          1570 => x"f3",
          1571 => x"80",
          1572 => x"f1",
          1573 => x"ff",
          1574 => x"54",
          1575 => x"39",
          1576 => x"08",
          1577 => x"ff",
          1578 => x"56",
          1579 => x"39",
          1580 => x"08",
          1581 => x"ff",
          1582 => x"54",
          1583 => x"39",
          1584 => x"08",
          1585 => x"ff",
          1586 => x"55",
          1587 => x"39",
          1588 => x"08",
          1589 => x"ff",
          1590 => x"56",
          1591 => x"39",
          1592 => x"08",
          1593 => x"ff",
          1594 => x"54",
          1595 => x"39",
          1596 => x"3f",
          1597 => x"3f",
          1598 => x"2e",
          1599 => x"0d",
          1600 => x"26",
          1601 => x"ec",
          1602 => x"c0",
          1603 => x"0d",
          1604 => x"e3",
          1605 => x"d0",
          1606 => x"0d",
          1607 => x"cb",
          1608 => x"e0",
          1609 => x"0d",
          1610 => x"b3",
          1611 => x"80",
          1612 => x"84",
          1613 => x"c0",
          1614 => x"aa",
          1615 => x"81",
          1616 => x"d0",
          1617 => x"b8",
          1618 => x"57",
          1619 => x"55",
          1620 => x"8f",
          1621 => x"a4",
          1622 => x"b8",
          1623 => x"0b",
          1624 => x"84",
          1625 => x"55",
          1626 => x"30",
          1627 => x"55",
          1628 => x"b0",
          1629 => x"08",
          1630 => x"b8",
          1631 => x"9a",
          1632 => x"3d",
          1633 => x"ad",
          1634 => x"06",
          1635 => x"aa",
          1636 => x"3d",
          1637 => x"34",
          1638 => x"ad",
          1639 => x"0c",
          1640 => x"ab",
          1641 => x"5d",
          1642 => x"a0",
          1643 => x"3d",
          1644 => x"f2",
          1645 => x"bf",
          1646 => x"79",
          1647 => x"84",
          1648 => x"33",
          1649 => x"73",
          1650 => x"81",
          1651 => x"c2",
          1652 => x"0c",
          1653 => x"aa",
          1654 => x"05",
          1655 => x"08",
          1656 => x"78",
          1657 => x"b8",
          1658 => x"80",
          1659 => x"ff",
          1660 => x"fa",
          1661 => x"05",
          1662 => x"81",
          1663 => x"73",
          1664 => x"38",
          1665 => x"8d",
          1666 => x"84",
          1667 => x"08",
          1668 => x"b8",
          1669 => x"d0",
          1670 => x"82",
          1671 => x"80",
          1672 => x"e3",
          1673 => x"0b",
          1674 => x"84",
          1675 => x"58",
          1676 => x"52",
          1677 => x"ff",
          1678 => x"81",
          1679 => x"b8",
          1680 => x"3d",
          1681 => x"b9",
          1682 => x"b4",
          1683 => x"f2",
          1684 => x"74",
          1685 => x"80",
          1686 => x"91",
          1687 => x"57",
          1688 => x"90",
          1689 => x"5f",
          1690 => x"e4",
          1691 => x"56",
          1692 => x"ff",
          1693 => x"2b",
          1694 => x"70",
          1695 => x"2c",
          1696 => x"05",
          1697 => x"5c",
          1698 => x"81",
          1699 => x"78",
          1700 => x"80",
          1701 => x"98",
          1702 => x"cb",
          1703 => x"56",
          1704 => x"33",
          1705 => x"83",
          1706 => x"56",
          1707 => x"76",
          1708 => x"9c",
          1709 => x"99",
          1710 => x"98",
          1711 => x"2b",
          1712 => x"70",
          1713 => x"5f",
          1714 => x"7a",
          1715 => x"d0",
          1716 => x"76",
          1717 => x"29",
          1718 => x"70",
          1719 => x"95",
          1720 => x"70",
          1721 => x"dd",
          1722 => x"25",
          1723 => x"18",
          1724 => x"ff",
          1725 => x"38",
          1726 => x"2e",
          1727 => x"56",
          1728 => x"e9",
          1729 => x"84",
          1730 => x"7f",
          1731 => x"b0",
          1732 => x"05",
          1733 => x"15",
          1734 => x"a0",
          1735 => x"d9",
          1736 => x"80",
          1737 => x"08",
          1738 => x"84",
          1739 => x"84",
          1740 => x"d0",
          1741 => x"d0",
          1742 => x"27",
          1743 => x"52",
          1744 => x"34",
          1745 => x"b5",
          1746 => x"2e",
          1747 => x"f2",
          1748 => x"8f",
          1749 => x"75",
          1750 => x"d0",
          1751 => x"b6",
          1752 => x"51",
          1753 => x"08",
          1754 => x"84",
          1755 => x"b5",
          1756 => x"05",
          1757 => x"81",
          1758 => x"51",
          1759 => x"a8",
          1760 => x"83",
          1761 => x"38",
          1762 => x"fc",
          1763 => x"38",
          1764 => x"a8",
          1765 => x"84",
          1766 => x"84",
          1767 => x"05",
          1768 => x"a5",
          1769 => x"a8",
          1770 => x"9e",
          1771 => x"51",
          1772 => x"08",
          1773 => x"84",
          1774 => x"b3",
          1775 => x"05",
          1776 => x"81",
          1777 => x"a8",
          1778 => x"a4",
          1779 => x"fa",
          1780 => x"81",
          1781 => x"7b",
          1782 => x"b9",
          1783 => x"ff",
          1784 => x"55",
          1785 => x"d4",
          1786 => x"84",
          1787 => x"52",
          1788 => x"a8",
          1789 => x"a4",
          1790 => x"ff",
          1791 => x"a8",
          1792 => x"74",
          1793 => x"5b",
          1794 => x"2b",
          1795 => x"43",
          1796 => x"38",
          1797 => x"ff",
          1798 => x"70",
          1799 => x"a4",
          1800 => x"24",
          1801 => x"52",
          1802 => x"81",
          1803 => x"70",
          1804 => x"56",
          1805 => x"84",
          1806 => x"b1",
          1807 => x"81",
          1808 => x"d0",
          1809 => x"25",
          1810 => x"16",
          1811 => x"d4",
          1812 => x"b1",
          1813 => x"81",
          1814 => x"d0",
          1815 => x"25",
          1816 => x"18",
          1817 => x"52",
          1818 => x"75",
          1819 => x"05",
          1820 => x"5b",
          1821 => x"38",
          1822 => x"55",
          1823 => x"d4",
          1824 => x"e9",
          1825 => x"57",
          1826 => x"ff",
          1827 => x"33",
          1828 => x"d4",
          1829 => x"c1",
          1830 => x"f4",
          1831 => x"ff",
          1832 => x"d0",
          1833 => x"d8",
          1834 => x"10",
          1835 => x"5e",
          1836 => x"2b",
          1837 => x"81",
          1838 => x"fb",
          1839 => x"83",
          1840 => x"f1",
          1841 => x"74",
          1842 => x"56",
          1843 => x"cc",
          1844 => x"38",
          1845 => x"0b",
          1846 => x"e4",
          1847 => x"a8",
          1848 => x"84",
          1849 => x"af",
          1850 => x"a0",
          1851 => x"c8",
          1852 => x"3f",
          1853 => x"75",
          1854 => x"06",
          1855 => x"51",
          1856 => x"d0",
          1857 => x"34",
          1858 => x"0b",
          1859 => x"55",
          1860 => x"c8",
          1861 => x"3f",
          1862 => x"ff",
          1863 => x"52",
          1864 => x"d0",
          1865 => x"d0",
          1866 => x"74",
          1867 => x"9f",
          1868 => x"34",
          1869 => x"84",
          1870 => x"84",
          1871 => x"5c",
          1872 => x"84",
          1873 => x"84",
          1874 => x"84",
          1875 => x"52",
          1876 => x"d0",
          1877 => x"2c",
          1878 => x"56",
          1879 => x"d4",
          1880 => x"a9",
          1881 => x"2b",
          1882 => x"5d",
          1883 => x"f0",
          1884 => x"51",
          1885 => x"0a",
          1886 => x"2c",
          1887 => x"74",
          1888 => x"c8",
          1889 => x"3f",
          1890 => x"0a",
          1891 => x"33",
          1892 => x"b9",
          1893 => x"81",
          1894 => x"08",
          1895 => x"3f",
          1896 => x"0a",
          1897 => x"33",
          1898 => x"e6",
          1899 => x"77",
          1900 => x"33",
          1901 => x"80",
          1902 => x"98",
          1903 => x"5b",
          1904 => x"b6",
          1905 => x"ff",
          1906 => x"b8",
          1907 => x"75",
          1908 => x"98",
          1909 => x"38",
          1910 => x"34",
          1911 => x"0a",
          1912 => x"33",
          1913 => x"38",
          1914 => x"34",
          1915 => x"b3",
          1916 => x"33",
          1917 => x"17",
          1918 => x"57",
          1919 => x"0a",
          1920 => x"2c",
          1921 => x"58",
          1922 => x"98",
          1923 => x"06",
          1924 => x"a8",
          1925 => x"51",
          1926 => x"0a",
          1927 => x"2c",
          1928 => x"75",
          1929 => x"c8",
          1930 => x"3f",
          1931 => x"0a",
          1932 => x"33",
          1933 => x"b9",
          1934 => x"08",
          1935 => x"75",
          1936 => x"e4",
          1937 => x"e4",
          1938 => x"75",
          1939 => x"84",
          1940 => x"56",
          1941 => x"84",
          1942 => x"a9",
          1943 => x"a0",
          1944 => x"c8",
          1945 => x"3f",
          1946 => x"7a",
          1947 => x"06",
          1948 => x"8b",
          1949 => x"d0",
          1950 => x"38",
          1951 => x"ca",
          1952 => x"08",
          1953 => x"ff",
          1954 => x"29",
          1955 => x"84",
          1956 => x"76",
          1957 => x"70",
          1958 => x"ff",
          1959 => x"25",
          1960 => x"f2",
          1961 => x"83",
          1962 => x"55",
          1963 => x"58",
          1964 => x"0b",
          1965 => x"08",
          1966 => x"74",
          1967 => x"d0",
          1968 => x"0b",
          1969 => x"3d",
          1970 => x"80",
          1971 => x"16",
          1972 => x"ff",
          1973 => x"ff",
          1974 => x"84",
          1975 => x"81",
          1976 => x"7b",
          1977 => x"84",
          1978 => x"57",
          1979 => x"38",
          1980 => x"ff",
          1981 => x"52",
          1982 => x"d4",
          1983 => x"f1",
          1984 => x"5a",
          1985 => x"ff",
          1986 => x"80",
          1987 => x"84",
          1988 => x"0c",
          1989 => x"a9",
          1990 => x"d0",
          1991 => x"ff",
          1992 => x"51",
          1993 => x"81",
          1994 => x"d0",
          1995 => x"80",
          1996 => x"08",
          1997 => x"84",
          1998 => x"a5",
          1999 => x"88",
          2000 => x"a8",
          2001 => x"a8",
          2002 => x"39",
          2003 => x"b8",
          2004 => x"b8",
          2005 => x"53",
          2006 => x"3f",
          2007 => x"d0",
          2008 => x"58",
          2009 => x"38",
          2010 => x"ff",
          2011 => x"52",
          2012 => x"d4",
          2013 => x"81",
          2014 => x"41",
          2015 => x"ff",
          2016 => x"d6",
          2017 => x"82",
          2018 => x"05",
          2019 => x"80",
          2020 => x"7b",
          2021 => x"10",
          2022 => x"41",
          2023 => x"75",
          2024 => x"a5",
          2025 => x"70",
          2026 => x"27",
          2027 => x"34",
          2028 => x"05",
          2029 => x"81",
          2030 => x"52",
          2031 => x"f2",
          2032 => x"80",
          2033 => x"84",
          2034 => x"0c",
          2035 => x"52",
          2036 => x"f8",
          2037 => x"38",
          2038 => x"5d",
          2039 => x"52",
          2040 => x"b8",
          2041 => x"7b",
          2042 => x"84",
          2043 => x"3f",
          2044 => x"84",
          2045 => x"84",
          2046 => x"58",
          2047 => x"06",
          2048 => x"83",
          2049 => x"58",
          2050 => x"2b",
          2051 => x"81",
          2052 => x"cb",
          2053 => x"83",
          2054 => x"f1",
          2055 => x"74",
          2056 => x"06",
          2057 => x"80",
          2058 => x"fe",
          2059 => x"e6",
          2060 => x"ff",
          2061 => x"81",
          2062 => x"93",
          2063 => x"83",
          2064 => x"51",
          2065 => x"33",
          2066 => x"f1",
          2067 => x"56",
          2068 => x"e4",
          2069 => x"70",
          2070 => x"08",
          2071 => x"82",
          2072 => x"d4",
          2073 => x"d4",
          2074 => x"51",
          2075 => x"38",
          2076 => x"80",
          2077 => x"c7",
          2078 => x"81",
          2079 => x"38",
          2080 => x"82",
          2081 => x"80",
          2082 => x"57",
          2083 => x"2e",
          2084 => x"75",
          2085 => x"92",
          2086 => x"2b",
          2087 => x"07",
          2088 => x"5b",
          2089 => x"70",
          2090 => x"84",
          2091 => x"38",
          2092 => x"90",
          2093 => x"31",
          2094 => x"15",
          2095 => x"34",
          2096 => x"3d",
          2097 => x"83",
          2098 => x"83",
          2099 => x"74",
          2100 => x"a7",
          2101 => x"70",
          2102 => x"70",
          2103 => x"70",
          2104 => x"5d",
          2105 => x"73",
          2106 => x"75",
          2107 => x"81",
          2108 => x"83",
          2109 => x"70",
          2110 => x"5b",
          2111 => x"f8",
          2112 => x"7d",
          2113 => x"5c",
          2114 => x"7d",
          2115 => x"38",
          2116 => x"83",
          2117 => x"56",
          2118 => x"59",
          2119 => x"d8",
          2120 => x"d7",
          2121 => x"92",
          2122 => x"57",
          2123 => x"81",
          2124 => x"81",
          2125 => x"54",
          2126 => x"80",
          2127 => x"83",
          2128 => x"70",
          2129 => x"88",
          2130 => x"56",
          2131 => x"38",
          2132 => x"83",
          2133 => x"70",
          2134 => x"71",
          2135 => x"11",
          2136 => x"a7",
          2137 => x"33",
          2138 => x"33",
          2139 => x"22",
          2140 => x"29",
          2141 => x"5f",
          2142 => x"38",
          2143 => x"19",
          2144 => x"81",
          2145 => x"ff",
          2146 => x"75",
          2147 => x"7b",
          2148 => x"53",
          2149 => x"5b",
          2150 => x"06",
          2151 => x"39",
          2152 => x"9a",
          2153 => x"8c",
          2154 => x"34",
          2155 => x"ee",
          2156 => x"ff",
          2157 => x"56",
          2158 => x"ee",
          2159 => x"74",
          2160 => x"83",
          2161 => x"e0",
          2162 => x"86",
          2163 => x"07",
          2164 => x"70",
          2165 => x"53",
          2166 => x"08",
          2167 => x"72",
          2168 => x"81",
          2169 => x"34",
          2170 => x"80",
          2171 => x"0d",
          2172 => x"e4",
          2173 => x"05",
          2174 => x"84",
          2175 => x"53",
          2176 => x"b6",
          2177 => x"f8",
          2178 => x"a7",
          2179 => x"5f",
          2180 => x"70",
          2181 => x"33",
          2182 => x"83",
          2183 => x"05",
          2184 => x"f8",
          2185 => x"06",
          2186 => x"72",
          2187 => x"53",
          2188 => x"92",
          2189 => x"b6",
          2190 => x"26",
          2191 => x"76",
          2192 => x"9f",
          2193 => x"70",
          2194 => x"e0",
          2195 => x"54",
          2196 => x"81",
          2197 => x"e3",
          2198 => x"83",
          2199 => x"54",
          2200 => x"74",
          2201 => x"14",
          2202 => x"84",
          2203 => x"83",
          2204 => x"ff",
          2205 => x"54",
          2206 => x"74",
          2207 => x"71",
          2208 => x"86",
          2209 => x"80",
          2210 => x"06",
          2211 => x"57",
          2212 => x"b6",
          2213 => x"84",
          2214 => x"05",
          2215 => x"33",
          2216 => x"15",
          2217 => x"33",
          2218 => x"55",
          2219 => x"72",
          2220 => x"04",
          2221 => x"92",
          2222 => x"b6",
          2223 => x"27",
          2224 => x"dd",
          2225 => x"83",
          2226 => x"2e",
          2227 => x"76",
          2228 => x"71",
          2229 => x"52",
          2230 => x"38",
          2231 => x"15",
          2232 => x"0b",
          2233 => x"81",
          2234 => x"80",
          2235 => x"e0",
          2236 => x"57",
          2237 => x"fd",
          2238 => x"33",
          2239 => x"96",
          2240 => x"33",
          2241 => x"fc",
          2242 => x"84",
          2243 => x"86",
          2244 => x"c3",
          2245 => x"b6",
          2246 => x"38",
          2247 => x"84",
          2248 => x"80",
          2249 => x"94",
          2250 => x"72",
          2251 => x"70",
          2252 => x"b8",
          2253 => x"f8",
          2254 => x"70",
          2255 => x"54",
          2256 => x"83",
          2257 => x"d7",
          2258 => x"75",
          2259 => x"f8",
          2260 => x"0c",
          2261 => x"33",
          2262 => x"2c",
          2263 => x"83",
          2264 => x"e4",
          2265 => x"95",
          2266 => x"ff",
          2267 => x"83",
          2268 => x"34",
          2269 => x"3d",
          2270 => x"34",
          2271 => x"33",
          2272 => x"fe",
          2273 => x"f8",
          2274 => x"0d",
          2275 => x"26",
          2276 => x"f8",
          2277 => x"90",
          2278 => x"2b",
          2279 => x"07",
          2280 => x"2e",
          2281 => x"0b",
          2282 => x"b8",
          2283 => x"f8",
          2284 => x"51",
          2285 => x"84",
          2286 => x"83",
          2287 => x"70",
          2288 => x"f8",
          2289 => x"51",
          2290 => x"80",
          2291 => x"0b",
          2292 => x"04",
          2293 => x"84",
          2294 => x"ff",
          2295 => x"07",
          2296 => x"a5",
          2297 => x"06",
          2298 => x"34",
          2299 => x"81",
          2300 => x"f8",
          2301 => x"90",
          2302 => x"70",
          2303 => x"83",
          2304 => x"70",
          2305 => x"83",
          2306 => x"d0",
          2307 => x"fe",
          2308 => x"bf",
          2309 => x"90",
          2310 => x"33",
          2311 => x"70",
          2312 => x"83",
          2313 => x"c0",
          2314 => x"fe",
          2315 => x"af",
          2316 => x"90",
          2317 => x"33",
          2318 => x"90",
          2319 => x"33",
          2320 => x"83",
          2321 => x"3d",
          2322 => x"05",
          2323 => x"33",
          2324 => x"33",
          2325 => x"5d",
          2326 => x"38",
          2327 => x"2e",
          2328 => x"34",
          2329 => x"83",
          2330 => x"23",
          2331 => x"0d",
          2332 => x"db",
          2333 => x"81",
          2334 => x"83",
          2335 => x"95",
          2336 => x"79",
          2337 => x"b6",
          2338 => x"55",
          2339 => x"e2",
          2340 => x"84",
          2341 => x"dc",
          2342 => x"83",
          2343 => x"34",
          2344 => x"b6",
          2345 => x"34",
          2346 => x"0b",
          2347 => x"f8",
          2348 => x"84",
          2349 => x"33",
          2350 => x"7a",
          2351 => x"8b",
          2352 => x"5a",
          2353 => x"10",
          2354 => x"59",
          2355 => x"3f",
          2356 => x"b7",
          2357 => x"26",
          2358 => x"80",
          2359 => x"80",
          2360 => x"f8",
          2361 => x"7c",
          2362 => x"04",
          2363 => x"0b",
          2364 => x"f8",
          2365 => x"34",
          2366 => x"f6",
          2367 => x"b8",
          2368 => x"ff",
          2369 => x"c8",
          2370 => x"b8",
          2371 => x"f6",
          2372 => x"51",
          2373 => x"81",
          2374 => x"3d",
          2375 => x"33",
          2376 => x"33",
          2377 => x"12",
          2378 => x"92",
          2379 => x"29",
          2380 => x"f6",
          2381 => x"57",
          2382 => x"89",
          2383 => x"81",
          2384 => x"38",
          2385 => x"b6",
          2386 => x"f8",
          2387 => x"56",
          2388 => x"a7",
          2389 => x"33",
          2390 => x"22",
          2391 => x"53",
          2392 => x"f8",
          2393 => x"54",
          2394 => x"80",
          2395 => x"81",
          2396 => x"f8",
          2397 => x"5b",
          2398 => x"84",
          2399 => x"81",
          2400 => x"81",
          2401 => x"77",
          2402 => x"83",
          2403 => x"53",
          2404 => x"dc",
          2405 => x"38",
          2406 => x"3d",
          2407 => x"75",
          2408 => x"2e",
          2409 => x"52",
          2410 => x"83",
          2411 => x"f8",
          2412 => x"13",
          2413 => x"81",
          2414 => x"52",
          2415 => x"70",
          2416 => x"26",
          2417 => x"fd",
          2418 => x"06",
          2419 => x"fe",
          2420 => x"fe",
          2421 => x"de",
          2422 => x"89",
          2423 => x"09",
          2424 => x"95",
          2425 => x"05",
          2426 => x"83",
          2427 => x"fc",
          2428 => x"81",
          2429 => x"fe",
          2430 => x"95",
          2431 => x"f8",
          2432 => x"e2",
          2433 => x"51",
          2434 => x"3d",
          2435 => x"b7",
          2436 => x"81",
          2437 => x"38",
          2438 => x"8a",
          2439 => x"84",
          2440 => x"38",
          2441 => x"33",
          2442 => x"05",
          2443 => x"33",
          2444 => x"b6",
          2445 => x"f8",
          2446 => x"5a",
          2447 => x"34",
          2448 => x"62",
          2449 => x"7f",
          2450 => x"b6",
          2451 => x"f8",
          2452 => x"72",
          2453 => x"83",
          2454 => x"34",
          2455 => x"58",
          2456 => x"b6",
          2457 => x"ff",
          2458 => x"80",
          2459 => x"0d",
          2460 => x"b7",
          2461 => x"2e",
          2462 => x"89",
          2463 => x"0c",
          2464 => x"33",
          2465 => x"05",
          2466 => x"33",
          2467 => x"b6",
          2468 => x"f8",
          2469 => x"5f",
          2470 => x"34",
          2471 => x"19",
          2472 => x"a7",
          2473 => x"33",
          2474 => x"22",
          2475 => x"11",
          2476 => x"90",
          2477 => x"81",
          2478 => x"60",
          2479 => x"f8",
          2480 => x"0c",
          2481 => x"82",
          2482 => x"38",
          2483 => x"a8",
          2484 => x"80",
          2485 => x"0d",
          2486 => x"d0",
          2487 => x"38",
          2488 => x"57",
          2489 => x"b7",
          2490 => x"59",
          2491 => x"80",
          2492 => x"0d",
          2493 => x"80",
          2494 => x"d8",
          2495 => x"95",
          2496 => x"40",
          2497 => x"a0",
          2498 => x"83",
          2499 => x"72",
          2500 => x"78",
          2501 => x"94",
          2502 => x"83",
          2503 => x"1b",
          2504 => x"ff",
          2505 => x"95",
          2506 => x"43",
          2507 => x"84",
          2508 => x"fe",
          2509 => x"fa",
          2510 => x"fe",
          2511 => x"f8",
          2512 => x"f8",
          2513 => x"a7",
          2514 => x"40",
          2515 => x"83",
          2516 => x"5a",
          2517 => x"86",
          2518 => x"1a",
          2519 => x"56",
          2520 => x"39",
          2521 => x"0b",
          2522 => x"b7",
          2523 => x"34",
          2524 => x"0b",
          2525 => x"04",
          2526 => x"34",
          2527 => x"34",
          2528 => x"34",
          2529 => x"0b",
          2530 => x"04",
          2531 => x"fa",
          2532 => x"b6",
          2533 => x"f8",
          2534 => x"75",
          2535 => x"83",
          2536 => x"29",
          2537 => x"f6",
          2538 => x"5b",
          2539 => x"78",
          2540 => x"75",
          2541 => x"95",
          2542 => x"ff",
          2543 => x"29",
          2544 => x"33",
          2545 => x"b6",
          2546 => x"f8",
          2547 => x"5e",
          2548 => x"18",
          2549 => x"29",
          2550 => x"33",
          2551 => x"b6",
          2552 => x"f8",
          2553 => x"72",
          2554 => x"83",
          2555 => x"05",
          2556 => x"5c",
          2557 => x"84",
          2558 => x"38",
          2559 => x"34",
          2560 => x"06",
          2561 => x"78",
          2562 => x"2e",
          2563 => x"a8",
          2564 => x"83",
          2565 => x"b4",
          2566 => x"83",
          2567 => x"80",
          2568 => x"81",
          2569 => x"b8",
          2570 => x"f8",
          2571 => x"81",
          2572 => x"81",
          2573 => x"a7",
          2574 => x"5c",
          2575 => x"ff",
          2576 => x"53",
          2577 => x"2e",
          2578 => x"ff",
          2579 => x"ff",
          2580 => x"40",
          2581 => x"80",
          2582 => x"f8",
          2583 => x"71",
          2584 => x"0b",
          2585 => x"94",
          2586 => x"83",
          2587 => x"1a",
          2588 => x"ff",
          2589 => x"95",
          2590 => x"5a",
          2591 => x"97",
          2592 => x"81",
          2593 => x"81",
          2594 => x"77",
          2595 => x"83",
          2596 => x"ff",
          2597 => x"a7",
          2598 => x"d8",
          2599 => x"ff",
          2600 => x"ff",
          2601 => x"43",
          2602 => x"86",
          2603 => x"d8",
          2604 => x"92",
          2605 => x"5e",
          2606 => x"34",
          2607 => x"1e",
          2608 => x"a7",
          2609 => x"33",
          2610 => x"22",
          2611 => x"11",
          2612 => x"90",
          2613 => x"81",
          2614 => x"79",
          2615 => x"f8",
          2616 => x"84",
          2617 => x"e4",
          2618 => x"96",
          2619 => x"33",
          2620 => x"81",
          2621 => x"ca",
          2622 => x"80",
          2623 => x"0d",
          2624 => x"84",
          2625 => x"f8",
          2626 => x"f8",
          2627 => x"fc",
          2628 => x"3d",
          2629 => x"8a",
          2630 => x"2e",
          2631 => x"81",
          2632 => x"34",
          2633 => x"80",
          2634 => x"05",
          2635 => x"17",
          2636 => x"7b",
          2637 => x"d8",
          2638 => x"5c",
          2639 => x"83",
          2640 => x"72",
          2641 => x"b6",
          2642 => x"80",
          2643 => x"f8",
          2644 => x"71",
          2645 => x"83",
          2646 => x"33",
          2647 => x"f8",
          2648 => x"05",
          2649 => x"ff",
          2650 => x"95",
          2651 => x"5a",
          2652 => x"97",
          2653 => x"ff",
          2654 => x"a2",
          2655 => x"90",
          2656 => x"f8",
          2657 => x"0c",
          2658 => x"2e",
          2659 => x"56",
          2660 => x"51",
          2661 => x"e4",
          2662 => x"cc",
          2663 => x"cd",
          2664 => x"ce",
          2665 => x"ff",
          2666 => x"b8",
          2667 => x"b8",
          2668 => x"b8",
          2669 => x"e5",
          2670 => x"38",
          2671 => x"2e",
          2672 => x"f8",
          2673 => x"94",
          2674 => x"e3",
          2675 => x"fe",
          2676 => x"83",
          2677 => x"06",
          2678 => x"41",
          2679 => x"52",
          2680 => x"3f",
          2681 => x"e5",
          2682 => x"5b",
          2683 => x"10",
          2684 => x"57",
          2685 => x"75",
          2686 => x"7e",
          2687 => x"7d",
          2688 => x"94",
          2689 => x"31",
          2690 => x"5a",
          2691 => x"94",
          2692 => x"33",
          2693 => x"84",
          2694 => x"ff",
          2695 => x"5f",
          2696 => x"83",
          2697 => x"0b",
          2698 => x"33",
          2699 => x"80",
          2700 => x"75",
          2701 => x"80",
          2702 => x"94",
          2703 => x"57",
          2704 => x"81",
          2705 => x"fc",
          2706 => x"7f",
          2707 => x"95",
          2708 => x"31",
          2709 => x"5a",
          2710 => x"95",
          2711 => x"33",
          2712 => x"84",
          2713 => x"09",
          2714 => x"d8",
          2715 => x"94",
          2716 => x"a0",
          2717 => x"51",
          2718 => x"83",
          2719 => x"87",
          2720 => x"5d",
          2721 => x"38",
          2722 => x"f2",
          2723 => x"80",
          2724 => x"22",
          2725 => x"fb",
          2726 => x"34",
          2727 => x"56",
          2728 => x"b8",
          2729 => x"7c",
          2730 => x"59",
          2731 => x"75",
          2732 => x"a2",
          2733 => x"80",
          2734 => x"33",
          2735 => x"84",
          2736 => x"56",
          2737 => x"76",
          2738 => x"83",
          2739 => x"80",
          2740 => x"76",
          2741 => x"84",
          2742 => x"83",
          2743 => x"81",
          2744 => x"e5",
          2745 => x"0b",
          2746 => x"80",
          2747 => x"56",
          2748 => x"81",
          2749 => x"f3",
          2750 => x"33",
          2751 => x"84",
          2752 => x"ff",
          2753 => x"70",
          2754 => x"70",
          2755 => x"52",
          2756 => x"83",
          2757 => x"23",
          2758 => x"5f",
          2759 => x"76",
          2760 => x"33",
          2761 => x"f9",
          2762 => x"95",
          2763 => x"33",
          2764 => x"84",
          2765 => x"40",
          2766 => x"83",
          2767 => x"70",
          2768 => x"71",
          2769 => x"05",
          2770 => x"7e",
          2771 => x"83",
          2772 => x"5f",
          2773 => x"79",
          2774 => x"5d",
          2775 => x"84",
          2776 => x"8e",
          2777 => x"f8",
          2778 => x"7c",
          2779 => x"e5",
          2780 => x"76",
          2781 => x"75",
          2782 => x"06",
          2783 => x"5a",
          2784 => x"31",
          2785 => x"71",
          2786 => x"a7",
          2787 => x"7f",
          2788 => x"71",
          2789 => x"79",
          2790 => x"b6",
          2791 => x"84",
          2792 => x"05",
          2793 => x"33",
          2794 => x"18",
          2795 => x"33",
          2796 => x"58",
          2797 => x"e0",
          2798 => x"33",
          2799 => x"70",
          2800 => x"05",
          2801 => x"33",
          2802 => x"1d",
          2803 => x"ff",
          2804 => x"e5",
          2805 => x"38",
          2806 => x"d8",
          2807 => x"84",
          2808 => x"e5",
          2809 => x"2e",
          2810 => x"75",
          2811 => x"38",
          2812 => x"ff",
          2813 => x"5c",
          2814 => x"84",
          2815 => x"f6",
          2816 => x"60",
          2817 => x"26",
          2818 => x"f2",
          2819 => x"29",
          2820 => x"70",
          2821 => x"05",
          2822 => x"8b",
          2823 => x"8b",
          2824 => x"98",
          2825 => x"2b",
          2826 => x"5f",
          2827 => x"77",
          2828 => x"70",
          2829 => x"ee",
          2830 => x"d7",
          2831 => x"60",
          2832 => x"7d",
          2833 => x"5a",
          2834 => x"31",
          2835 => x"40",
          2836 => x"26",
          2837 => x"84",
          2838 => x"e0",
          2839 => x"05",
          2840 => x"26",
          2841 => x"19",
          2842 => x"34",
          2843 => x"38",
          2844 => x"ff",
          2845 => x"f8",
          2846 => x"84",
          2847 => x"07",
          2848 => x"09",
          2849 => x"83",
          2850 => x"ff",
          2851 => x"f8",
          2852 => x"1e",
          2853 => x"84",
          2854 => x"84",
          2855 => x"fa",
          2856 => x"07",
          2857 => x"18",
          2858 => x"fb",
          2859 => x"06",
          2860 => x"34",
          2861 => x"fb",
          2862 => x"90",
          2863 => x"81",
          2864 => x"f8",
          2865 => x"33",
          2866 => x"83",
          2867 => x"f1",
          2868 => x"70",
          2869 => x"39",
          2870 => x"56",
          2871 => x"39",
          2872 => x"90",
          2873 => x"fe",
          2874 => x"ef",
          2875 => x"f8",
          2876 => x"90",
          2877 => x"56",
          2878 => x"39",
          2879 => x"a0",
          2880 => x"fe",
          2881 => x"fe",
          2882 => x"90",
          2883 => x"33",
          2884 => x"83",
          2885 => x"f8",
          2886 => x"56",
          2887 => x"39",
          2888 => x"56",
          2889 => x"39",
          2890 => x"56",
          2891 => x"39",
          2892 => x"56",
          2893 => x"39",
          2894 => x"80",
          2895 => x"34",
          2896 => x"81",
          2897 => x"f8",
          2898 => x"83",
          2899 => x"d2",
          2900 => x"cc",
          2901 => x"cd",
          2902 => x"ce",
          2903 => x"80",
          2904 => x"39",
          2905 => x"0b",
          2906 => x"04",
          2907 => x"95",
          2908 => x"05",
          2909 => x"42",
          2910 => x"51",
          2911 => x"08",
          2912 => x"b7",
          2913 => x"34",
          2914 => x"3d",
          2915 => x"ef",
          2916 => x"11",
          2917 => x"7b",
          2918 => x"ca",
          2919 => x"80",
          2920 => x"80",
          2921 => x"81",
          2922 => x"33",
          2923 => x"56",
          2924 => x"95",
          2925 => x"3f",
          2926 => x"e9",
          2927 => x"33",
          2928 => x"72",
          2929 => x"75",
          2930 => x"d8",
          2931 => x"38",
          2932 => x"39",
          2933 => x"09",
          2934 => x"57",
          2935 => x"81",
          2936 => x"59",
          2937 => x"38",
          2938 => x"d7",
          2939 => x"81",
          2940 => x"94",
          2941 => x"ff",
          2942 => x"29",
          2943 => x"f8",
          2944 => x"05",
          2945 => x"ea",
          2946 => x"77",
          2947 => x"ff",
          2948 => x"7b",
          2949 => x"33",
          2950 => x"ff",
          2951 => x"7c",
          2952 => x"80",
          2953 => x"d7",
          2954 => x"38",
          2955 => x"34",
          2956 => x"22",
          2957 => x"90",
          2958 => x"81",
          2959 => x"5f",
          2960 => x"86",
          2961 => x"7f",
          2962 => x"41",
          2963 => x"ea",
          2964 => x"e0",
          2965 => x"33",
          2966 => x"70",
          2967 => x"05",
          2968 => x"33",
          2969 => x"1d",
          2970 => x"ec",
          2971 => x"84",
          2972 => x"05",
          2973 => x"33",
          2974 => x"18",
          2975 => x"33",
          2976 => x"58",
          2977 => x"fa",
          2978 => x"84",
          2979 => x"f8",
          2980 => x"f8",
          2981 => x"5c",
          2982 => x"d2",
          2983 => x"ff",
          2984 => x"61",
          2985 => x"f8",
          2986 => x"19",
          2987 => x"80",
          2988 => x"b6",
          2989 => x"12",
          2990 => x"8d",
          2991 => x"34",
          2992 => x"81",
          2993 => x"59",
          2994 => x"38",
          2995 => x"2e",
          2996 => x"f8",
          2997 => x"f8",
          2998 => x"76",
          2999 => x"38",
          3000 => x"83",
          3001 => x"1a",
          3002 => x"e7",
          3003 => x"f8",
          3004 => x"58",
          3005 => x"80",
          3006 => x"f8",
          3007 => x"34",
          3008 => x"76",
          3009 => x"90",
          3010 => x"79",
          3011 => x"79",
          3012 => x"23",
          3013 => x"94",
          3014 => x"92",
          3015 => x"f8",
          3016 => x"83",
          3017 => x"f8",
          3018 => x"1a",
          3019 => x"e9",
          3020 => x"02",
          3021 => x"54",
          3022 => x"51",
          3023 => x"e4",
          3024 => x"73",
          3025 => x"b8",
          3026 => x"3d",
          3027 => x"0b",
          3028 => x"06",
          3029 => x"55",
          3030 => x"81",
          3031 => x"74",
          3032 => x"3d",
          3033 => x"82",
          3034 => x"73",
          3035 => x"70",
          3036 => x"83",
          3037 => x"7b",
          3038 => x"7b",
          3039 => x"80",
          3040 => x"80",
          3041 => x"33",
          3042 => x"33",
          3043 => x"80",
          3044 => x"5d",
          3045 => x"ff",
          3046 => x"55",
          3047 => x"81",
          3048 => x"34",
          3049 => x"87",
          3050 => x"2e",
          3051 => x"57",
          3052 => x"14",
          3053 => x"f9",
          3054 => x"f6",
          3055 => x"83",
          3056 => x"72",
          3057 => x"ff",
          3058 => x"98",
          3059 => x"79",
          3060 => x"83",
          3061 => x"14",
          3062 => x"14",
          3063 => x"74",
          3064 => x"33",
          3065 => x"56",
          3066 => x"81",
          3067 => x"70",
          3068 => x"2e",
          3069 => x"bd",
          3070 => x"80",
          3071 => x"f6",
          3072 => x"33",
          3073 => x"33",
          3074 => x"bf",
          3075 => x"56",
          3076 => x"81",
          3077 => x"16",
          3078 => x"38",
          3079 => x"81",
          3080 => x"16",
          3081 => x"81",
          3082 => x"8d",
          3083 => x"72",
          3084 => x"ff",
          3085 => x"8c",
          3086 => x"81",
          3087 => x"b8",
          3088 => x"9c",
          3089 => x"ec",
          3090 => x"08",
          3091 => x"70",
          3092 => x"27",
          3093 => x"34",
          3094 => x"19",
          3095 => x"72",
          3096 => x"79",
          3097 => x"73",
          3098 => x"87",
          3099 => x"7d",
          3100 => x"f6",
          3101 => x"83",
          3102 => x"34",
          3103 => x"ec",
          3104 => x"81",
          3105 => x"33",
          3106 => x"34",
          3107 => x"f6",
          3108 => x"9c",
          3109 => x"80",
          3110 => x"8a",
          3111 => x"74",
          3112 => x"9b",
          3113 => x"83",
          3114 => x"38",
          3115 => x"81",
          3116 => x"98",
          3117 => x"38",
          3118 => x"70",
          3119 => x"06",
          3120 => x"53",
          3121 => x"38",
          3122 => x"76",
          3123 => x"f4",
          3124 => x"87",
          3125 => x"0c",
          3126 => x"81",
          3127 => x"06",
          3128 => x"9b",
          3129 => x"80",
          3130 => x"72",
          3131 => x"32",
          3132 => x"40",
          3133 => x"2e",
          3134 => x"ff",
          3135 => x"10",
          3136 => x"33",
          3137 => x"38",
          3138 => x"57",
          3139 => x"db",
          3140 => x"38",
          3141 => x"91",
          3142 => x"51",
          3143 => x"0c",
          3144 => x"81",
          3145 => x"ff",
          3146 => x"33",
          3147 => x"15",
          3148 => x"f6",
          3149 => x"98",
          3150 => x"15",
          3151 => x"06",
          3152 => x"38",
          3153 => x"75",
          3154 => x"06",
          3155 => x"fb",
          3156 => x"fa",
          3157 => x"55",
          3158 => x"c0",
          3159 => x"76",
          3160 => x"ff",
          3161 => x"ca",
          3162 => x"09",
          3163 => x"72",
          3164 => x"f6",
          3165 => x"f6",
          3166 => x"83",
          3167 => x"5c",
          3168 => x"2e",
          3169 => x"59",
          3170 => x"81",
          3171 => x"fd",
          3172 => x"54",
          3173 => x"db",
          3174 => x"54",
          3175 => x"f7",
          3176 => x"33",
          3177 => x"73",
          3178 => x"95",
          3179 => x"84",
          3180 => x"f6",
          3181 => x"d7",
          3182 => x"57",
          3183 => x"80",
          3184 => x"81",
          3185 => x"73",
          3186 => x"f8",
          3187 => x"81",
          3188 => x"75",
          3189 => x"f8",
          3190 => x"81",
          3191 => x"ff",
          3192 => x"95",
          3193 => x"c8",
          3194 => x"83",
          3195 => x"59",
          3196 => x"51",
          3197 => x"fa",
          3198 => x"08",
          3199 => x"13",
          3200 => x"e0",
          3201 => x"08",
          3202 => x"80",
          3203 => x"c0",
          3204 => x"55",
          3205 => x"98",
          3206 => x"08",
          3207 => x"14",
          3208 => x"52",
          3209 => x"fe",
          3210 => x"08",
          3211 => x"c8",
          3212 => x"c0",
          3213 => x"ce",
          3214 => x"08",
          3215 => x"74",
          3216 => x"87",
          3217 => x"73",
          3218 => x"db",
          3219 => x"72",
          3220 => x"55",
          3221 => x"53",
          3222 => x"ff",
          3223 => x"ff",
          3224 => x"0c",
          3225 => x"b8",
          3226 => x"3d",
          3227 => x"33",
          3228 => x"08",
          3229 => x"06",
          3230 => x"55",
          3231 => x"2a",
          3232 => x"2a",
          3233 => x"15",
          3234 => x"82",
          3235 => x"80",
          3236 => x"f0",
          3237 => x"34",
          3238 => x"87",
          3239 => x"08",
          3240 => x"c0",
          3241 => x"9c",
          3242 => x"81",
          3243 => x"56",
          3244 => x"81",
          3245 => x"a4",
          3246 => x"80",
          3247 => x"80",
          3248 => x"80",
          3249 => x"9c",
          3250 => x"55",
          3251 => x"33",
          3252 => x"70",
          3253 => x"2e",
          3254 => x"55",
          3255 => x"71",
          3256 => x"57",
          3257 => x"74",
          3258 => x"38",
          3259 => x"75",
          3260 => x"80",
          3261 => x"92",
          3262 => x"71",
          3263 => x"26",
          3264 => x"88",
          3265 => x"e4",
          3266 => x"c2",
          3267 => x"05",
          3268 => x"83",
          3269 => x"fc",
          3270 => x"07",
          3271 => x"34",
          3272 => x"34",
          3273 => x"34",
          3274 => x"f0",
          3275 => x"56",
          3276 => x"38",
          3277 => x"70",
          3278 => x"f0",
          3279 => x"82",
          3280 => x"80",
          3281 => x"f0",
          3282 => x"34",
          3283 => x"87",
          3284 => x"08",
          3285 => x"c0",
          3286 => x"9c",
          3287 => x"81",
          3288 => x"56",
          3289 => x"81",
          3290 => x"a4",
          3291 => x"80",
          3292 => x"80",
          3293 => x"80",
          3294 => x"9c",
          3295 => x"55",
          3296 => x"33",
          3297 => x"70",
          3298 => x"2e",
          3299 => x"55",
          3300 => x"71",
          3301 => x"57",
          3302 => x"81",
          3303 => x"74",
          3304 => x"80",
          3305 => x"b8",
          3306 => x"51",
          3307 => x"f0",
          3308 => x"0b",
          3309 => x"0b",
          3310 => x"80",
          3311 => x"83",
          3312 => x"05",
          3313 => x"87",
          3314 => x"2e",
          3315 => x"98",
          3316 => x"87",
          3317 => x"87",
          3318 => x"70",
          3319 => x"71",
          3320 => x"98",
          3321 => x"87",
          3322 => x"98",
          3323 => x"38",
          3324 => x"08",
          3325 => x"71",
          3326 => x"98",
          3327 => x"38",
          3328 => x"81",
          3329 => x"8a",
          3330 => x"fe",
          3331 => x"83",
          3332 => x"82",
          3333 => x"b8",
          3334 => x"70",
          3335 => x"73",
          3336 => x"8b",
          3337 => x"70",
          3338 => x"71",
          3339 => x"53",
          3340 => x"80",
          3341 => x"82",
          3342 => x"2b",
          3343 => x"33",
          3344 => x"90",
          3345 => x"56",
          3346 => x"84",
          3347 => x"2b",
          3348 => x"88",
          3349 => x"13",
          3350 => x"87",
          3351 => x"17",
          3352 => x"88",
          3353 => x"59",
          3354 => x"85",
          3355 => x"52",
          3356 => x"87",
          3357 => x"74",
          3358 => x"84",
          3359 => x"12",
          3360 => x"80",
          3361 => x"52",
          3362 => x"89",
          3363 => x"13",
          3364 => x"07",
          3365 => x"33",
          3366 => x"58",
          3367 => x"84",
          3368 => x"b8",
          3369 => x"85",
          3370 => x"2b",
          3371 => x"86",
          3372 => x"2b",
          3373 => x"52",
          3374 => x"34",
          3375 => x"81",
          3376 => x"ff",
          3377 => x"54",
          3378 => x"34",
          3379 => x"33",
          3380 => x"83",
          3381 => x"12",
          3382 => x"2b",
          3383 => x"88",
          3384 => x"57",
          3385 => x"83",
          3386 => x"17",
          3387 => x"2b",
          3388 => x"33",
          3389 => x"81",
          3390 => x"52",
          3391 => x"73",
          3392 => x"d4",
          3393 => x"12",
          3394 => x"07",
          3395 => x"71",
          3396 => x"53",
          3397 => x"80",
          3398 => x"13",
          3399 => x"80",
          3400 => x"76",
          3401 => x"b8",
          3402 => x"12",
          3403 => x"07",
          3404 => x"33",
          3405 => x"57",
          3406 => x"72",
          3407 => x"89",
          3408 => x"84",
          3409 => x"2e",
          3410 => x"77",
          3411 => x"04",
          3412 => x"0c",
          3413 => x"82",
          3414 => x"f4",
          3415 => x"d4",
          3416 => x"81",
          3417 => x"76",
          3418 => x"34",
          3419 => x"17",
          3420 => x"b8",
          3421 => x"05",
          3422 => x"ff",
          3423 => x"56",
          3424 => x"34",
          3425 => x"10",
          3426 => x"55",
          3427 => x"83",
          3428 => x"0d",
          3429 => x"72",
          3430 => x"82",
          3431 => x"51",
          3432 => x"d4",
          3433 => x"71",
          3434 => x"58",
          3435 => x"2e",
          3436 => x"17",
          3437 => x"2b",
          3438 => x"31",
          3439 => x"27",
          3440 => x"74",
          3441 => x"38",
          3442 => x"85",
          3443 => x"5a",
          3444 => x"2e",
          3445 => x"76",
          3446 => x"12",
          3447 => x"ff",
          3448 => x"59",
          3449 => x"80",
          3450 => x"78",
          3451 => x"72",
          3452 => x"70",
          3453 => x"80",
          3454 => x"56",
          3455 => x"34",
          3456 => x"2a",
          3457 => x"83",
          3458 => x"19",
          3459 => x"2b",
          3460 => x"06",
          3461 => x"70",
          3462 => x"52",
          3463 => x"ff",
          3464 => x"b8",
          3465 => x"72",
          3466 => x"70",
          3467 => x"71",
          3468 => x"05",
          3469 => x"15",
          3470 => x"d4",
          3471 => x"11",
          3472 => x"07",
          3473 => x"70",
          3474 => x"84",
          3475 => x"33",
          3476 => x"83",
          3477 => x"5a",
          3478 => x"15",
          3479 => x"55",
          3480 => x"33",
          3481 => x"54",
          3482 => x"79",
          3483 => x"18",
          3484 => x"0c",
          3485 => x"87",
          3486 => x"2b",
          3487 => x"18",
          3488 => x"2a",
          3489 => x"84",
          3490 => x"b8",
          3491 => x"85",
          3492 => x"2b",
          3493 => x"15",
          3494 => x"2a",
          3495 => x"52",
          3496 => x"34",
          3497 => x"81",
          3498 => x"ff",
          3499 => x"54",
          3500 => x"34",
          3501 => x"51",
          3502 => x"84",
          3503 => x"2e",
          3504 => x"73",
          3505 => x"04",
          3506 => x"e4",
          3507 => x"0d",
          3508 => x"d4",
          3509 => x"23",
          3510 => x"ff",
          3511 => x"b8",
          3512 => x"0b",
          3513 => x"54",
          3514 => x"15",
          3515 => x"86",
          3516 => x"84",
          3517 => x"ff",
          3518 => x"ff",
          3519 => x"55",
          3520 => x"17",
          3521 => x"10",
          3522 => x"05",
          3523 => x"0b",
          3524 => x"2e",
          3525 => x"3d",
          3526 => x"84",
          3527 => x"61",
          3528 => x"85",
          3529 => x"38",
          3530 => x"7f",
          3531 => x"83",
          3532 => x"ff",
          3533 => x"70",
          3534 => x"7a",
          3535 => x"88",
          3536 => x"ff",
          3537 => x"05",
          3538 => x"81",
          3539 => x"90",
          3540 => x"46",
          3541 => x"59",
          3542 => x"85",
          3543 => x"33",
          3544 => x"10",
          3545 => x"98",
          3546 => x"53",
          3547 => x"c9",
          3548 => x"63",
          3549 => x"38",
          3550 => x"1b",
          3551 => x"63",
          3552 => x"38",
          3553 => x"71",
          3554 => x"11",
          3555 => x"2b",
          3556 => x"52",
          3557 => x"8c",
          3558 => x"83",
          3559 => x"2b",
          3560 => x"12",
          3561 => x"07",
          3562 => x"33",
          3563 => x"59",
          3564 => x"5c",
          3565 => x"85",
          3566 => x"17",
          3567 => x"8b",
          3568 => x"86",
          3569 => x"2b",
          3570 => x"52",
          3571 => x"34",
          3572 => x"08",
          3573 => x"88",
          3574 => x"88",
          3575 => x"34",
          3576 => x"08",
          3577 => x"33",
          3578 => x"74",
          3579 => x"88",
          3580 => x"45",
          3581 => x"34",
          3582 => x"08",
          3583 => x"71",
          3584 => x"05",
          3585 => x"88",
          3586 => x"45",
          3587 => x"1a",
          3588 => x"d4",
          3589 => x"12",
          3590 => x"62",
          3591 => x"5d",
          3592 => x"fd",
          3593 => x"05",
          3594 => x"ff",
          3595 => x"81",
          3596 => x"e4",
          3597 => x"f4",
          3598 => x"0b",
          3599 => x"53",
          3600 => x"c7",
          3601 => x"60",
          3602 => x"84",
          3603 => x"34",
          3604 => x"d4",
          3605 => x"0b",
          3606 => x"84",
          3607 => x"80",
          3608 => x"88",
          3609 => x"18",
          3610 => x"d0",
          3611 => x"d4",
          3612 => x"82",
          3613 => x"84",
          3614 => x"38",
          3615 => x"54",
          3616 => x"51",
          3617 => x"84",
          3618 => x"61",
          3619 => x"2b",
          3620 => x"33",
          3621 => x"81",
          3622 => x"44",
          3623 => x"81",
          3624 => x"05",
          3625 => x"19",
          3626 => x"d4",
          3627 => x"33",
          3628 => x"8f",
          3629 => x"ff",
          3630 => x"47",
          3631 => x"05",
          3632 => x"63",
          3633 => x"1e",
          3634 => x"34",
          3635 => x"05",
          3636 => x"bc",
          3637 => x"ff",
          3638 => x"81",
          3639 => x"ff",
          3640 => x"33",
          3641 => x"10",
          3642 => x"98",
          3643 => x"53",
          3644 => x"25",
          3645 => x"78",
          3646 => x"8b",
          3647 => x"5b",
          3648 => x"8f",
          3649 => x"d4",
          3650 => x"23",
          3651 => x"ff",
          3652 => x"b8",
          3653 => x"0b",
          3654 => x"59",
          3655 => x"1a",
          3656 => x"86",
          3657 => x"84",
          3658 => x"ff",
          3659 => x"ff",
          3660 => x"57",
          3661 => x"64",
          3662 => x"70",
          3663 => x"05",
          3664 => x"05",
          3665 => x"ee",
          3666 => x"61",
          3667 => x"27",
          3668 => x"80",
          3669 => x"fb",
          3670 => x"0c",
          3671 => x"11",
          3672 => x"71",
          3673 => x"33",
          3674 => x"83",
          3675 => x"85",
          3676 => x"88",
          3677 => x"58",
          3678 => x"05",
          3679 => x"b8",
          3680 => x"85",
          3681 => x"2b",
          3682 => x"15",
          3683 => x"2a",
          3684 => x"41",
          3685 => x"87",
          3686 => x"70",
          3687 => x"07",
          3688 => x"5f",
          3689 => x"81",
          3690 => x"1f",
          3691 => x"8b",
          3692 => x"73",
          3693 => x"07",
          3694 => x"43",
          3695 => x"81",
          3696 => x"1f",
          3697 => x"2b",
          3698 => x"14",
          3699 => x"07",
          3700 => x"40",
          3701 => x"60",
          3702 => x"70",
          3703 => x"71",
          3704 => x"70",
          3705 => x"05",
          3706 => x"84",
          3707 => x"83",
          3708 => x"39",
          3709 => x"0c",
          3710 => x"82",
          3711 => x"f4",
          3712 => x"d4",
          3713 => x"81",
          3714 => x"7f",
          3715 => x"34",
          3716 => x"15",
          3717 => x"b8",
          3718 => x"05",
          3719 => x"ff",
          3720 => x"5e",
          3721 => x"34",
          3722 => x"10",
          3723 => x"5c",
          3724 => x"83",
          3725 => x"7f",
          3726 => x"87",
          3727 => x"2b",
          3728 => x"1d",
          3729 => x"2a",
          3730 => x"61",
          3731 => x"34",
          3732 => x"11",
          3733 => x"71",
          3734 => x"33",
          3735 => x"70",
          3736 => x"56",
          3737 => x"78",
          3738 => x"08",
          3739 => x"88",
          3740 => x"88",
          3741 => x"34",
          3742 => x"08",
          3743 => x"71",
          3744 => x"05",
          3745 => x"2b",
          3746 => x"06",
          3747 => x"5d",
          3748 => x"82",
          3749 => x"b8",
          3750 => x"12",
          3751 => x"07",
          3752 => x"71",
          3753 => x"70",
          3754 => x"5a",
          3755 => x"81",
          3756 => x"5b",
          3757 => x"16",
          3758 => x"07",
          3759 => x"33",
          3760 => x"5e",
          3761 => x"1e",
          3762 => x"d4",
          3763 => x"12",
          3764 => x"07",
          3765 => x"33",
          3766 => x"44",
          3767 => x"7c",
          3768 => x"05",
          3769 => x"33",
          3770 => x"81",
          3771 => x"5b",
          3772 => x"16",
          3773 => x"70",
          3774 => x"71",
          3775 => x"81",
          3776 => x"83",
          3777 => x"63",
          3778 => x"59",
          3779 => x"7b",
          3780 => x"70",
          3781 => x"8b",
          3782 => x"70",
          3783 => x"07",
          3784 => x"5d",
          3785 => x"75",
          3786 => x"b8",
          3787 => x"83",
          3788 => x"2b",
          3789 => x"12",
          3790 => x"07",
          3791 => x"33",
          3792 => x"59",
          3793 => x"5d",
          3794 => x"79",
          3795 => x"70",
          3796 => x"71",
          3797 => x"05",
          3798 => x"88",
          3799 => x"5e",
          3800 => x"16",
          3801 => x"d4",
          3802 => x"71",
          3803 => x"70",
          3804 => x"79",
          3805 => x"d4",
          3806 => x"12",
          3807 => x"07",
          3808 => x"71",
          3809 => x"5c",
          3810 => x"79",
          3811 => x"d4",
          3812 => x"33",
          3813 => x"74",
          3814 => x"71",
          3815 => x"5c",
          3816 => x"82",
          3817 => x"b8",
          3818 => x"83",
          3819 => x"57",
          3820 => x"5a",
          3821 => x"b6",
          3822 => x"84",
          3823 => x"ff",
          3824 => x"39",
          3825 => x"8b",
          3826 => x"84",
          3827 => x"2b",
          3828 => x"43",
          3829 => x"63",
          3830 => x"08",
          3831 => x"33",
          3832 => x"74",
          3833 => x"71",
          3834 => x"41",
          3835 => x"64",
          3836 => x"34",
          3837 => x"81",
          3838 => x"ff",
          3839 => x"42",
          3840 => x"34",
          3841 => x"33",
          3842 => x"83",
          3843 => x"12",
          3844 => x"2b",
          3845 => x"88",
          3846 => x"45",
          3847 => x"83",
          3848 => x"1f",
          3849 => x"2b",
          3850 => x"33",
          3851 => x"81",
          3852 => x"5f",
          3853 => x"7d",
          3854 => x"ff",
          3855 => x"60",
          3856 => x"e4",
          3857 => x"2e",
          3858 => x"b8",
          3859 => x"73",
          3860 => x"7b",
          3861 => x"f9",
          3862 => x"d4",
          3863 => x"38",
          3864 => x"b8",
          3865 => x"51",
          3866 => x"54",
          3867 => x"38",
          3868 => x"08",
          3869 => x"b8",
          3870 => x"ff",
          3871 => x"80",
          3872 => x"80",
          3873 => x"fe",
          3874 => x"55",
          3875 => x"34",
          3876 => x"15",
          3877 => x"b8",
          3878 => x"81",
          3879 => x"08",
          3880 => x"80",
          3881 => x"70",
          3882 => x"88",
          3883 => x"b8",
          3884 => x"b8",
          3885 => x"76",
          3886 => x"34",
          3887 => x"38",
          3888 => x"8f",
          3889 => x"26",
          3890 => x"52",
          3891 => x"0d",
          3892 => x"33",
          3893 => x"38",
          3894 => x"e4",
          3895 => x"38",
          3896 => x"b8",
          3897 => x"e4",
          3898 => x"0d",
          3899 => x"05",
          3900 => x"76",
          3901 => x"17",
          3902 => x"55",
          3903 => x"87",
          3904 => x"52",
          3905 => x"e4",
          3906 => x"2e",
          3907 => x"54",
          3908 => x"38",
          3909 => x"80",
          3910 => x"74",
          3911 => x"04",
          3912 => x"ff",
          3913 => x"ff",
          3914 => x"7c",
          3915 => x"33",
          3916 => x"74",
          3917 => x"33",
          3918 => x"73",
          3919 => x"c0",
          3920 => x"76",
          3921 => x"08",
          3922 => x"a7",
          3923 => x"73",
          3924 => x"74",
          3925 => x"2e",
          3926 => x"84",
          3927 => x"84",
          3928 => x"06",
          3929 => x"ac",
          3930 => x"02",
          3931 => x"05",
          3932 => x"53",
          3933 => x"e0",
          3934 => x"83",
          3935 => x"c0",
          3936 => x"2e",
          3937 => x"70",
          3938 => x"84",
          3939 => x"88",
          3940 => x"e4",
          3941 => x"75",
          3942 => x"86",
          3943 => x"c0",
          3944 => x"38",
          3945 => x"51",
          3946 => x"c0",
          3947 => x"87",
          3948 => x"38",
          3949 => x"14",
          3950 => x"80",
          3951 => x"06",
          3952 => x"f6",
          3953 => x"19",
          3954 => x"2e",
          3955 => x"56",
          3956 => x"53",
          3957 => x"a3",
          3958 => x"83",
          3959 => x"0c",
          3960 => x"18",
          3961 => x"19",
          3962 => x"59",
          3963 => x"81",
          3964 => x"83",
          3965 => x"1a",
          3966 => x"e4",
          3967 => x"27",
          3968 => x"74",
          3969 => x"38",
          3970 => x"81",
          3971 => x"78",
          3972 => x"81",
          3973 => x"57",
          3974 => x"ee",
          3975 => x"56",
          3976 => x"34",
          3977 => x"d5",
          3978 => x"0b",
          3979 => x"34",
          3980 => x"e1",
          3981 => x"bb",
          3982 => x"19",
          3983 => x"34",
          3984 => x"80",
          3985 => x"18",
          3986 => x"74",
          3987 => x"34",
          3988 => x"19",
          3989 => x"a3",
          3990 => x"84",
          3991 => x"74",
          3992 => x"56",
          3993 => x"2a",
          3994 => x"18",
          3995 => x"5b",
          3996 => x"18",
          3997 => x"19",
          3998 => x"33",
          3999 => x"08",
          4000 => x"39",
          4001 => x"59",
          4002 => x"9c",
          4003 => x"58",
          4004 => x"0d",
          4005 => x"82",
          4006 => x"82",
          4007 => x"06",
          4008 => x"89",
          4009 => x"80",
          4010 => x"38",
          4011 => x"09",
          4012 => x"78",
          4013 => x"51",
          4014 => x"80",
          4015 => x"78",
          4016 => x"79",
          4017 => x"81",
          4018 => x"05",
          4019 => x"79",
          4020 => x"33",
          4021 => x"09",
          4022 => x"78",
          4023 => x"51",
          4024 => x"80",
          4025 => x"78",
          4026 => x"7a",
          4027 => x"70",
          4028 => x"71",
          4029 => x"79",
          4030 => x"84",
          4031 => x"75",
          4032 => x"b4",
          4033 => x"0b",
          4034 => x"7b",
          4035 => x"38",
          4036 => x"81",
          4037 => x"b8",
          4038 => x"59",
          4039 => x"fd",
          4040 => x"77",
          4041 => x"33",
          4042 => x"0c",
          4043 => x"83",
          4044 => x"75",
          4045 => x"b4",
          4046 => x"0b",
          4047 => x"7c",
          4048 => x"38",
          4049 => x"81",
          4050 => x"b8",
          4051 => x"59",
          4052 => x"fc",
          4053 => x"06",
          4054 => x"82",
          4055 => x"2b",
          4056 => x"88",
          4057 => x"fe",
          4058 => x"41",
          4059 => x"0d",
          4060 => x"b8",
          4061 => x"5c",
          4062 => x"e4",
          4063 => x"be",
          4064 => x"34",
          4065 => x"84",
          4066 => x"18",
          4067 => x"33",
          4068 => x"fd",
          4069 => x"a0",
          4070 => x"17",
          4071 => x"fd",
          4072 => x"53",
          4073 => x"52",
          4074 => x"08",
          4075 => x"38",
          4076 => x"b4",
          4077 => x"7c",
          4078 => x"17",
          4079 => x"38",
          4080 => x"39",
          4081 => x"17",
          4082 => x"f5",
          4083 => x"08",
          4084 => x"38",
          4085 => x"b4",
          4086 => x"b8",
          4087 => x"08",
          4088 => x"55",
          4089 => x"b8",
          4090 => x"18",
          4091 => x"33",
          4092 => x"a0",
          4093 => x"b8",
          4094 => x"5e",
          4095 => x"e4",
          4096 => x"cb",
          4097 => x"34",
          4098 => x"84",
          4099 => x"18",
          4100 => x"33",
          4101 => x"fb",
          4102 => x"a0",
          4103 => x"17",
          4104 => x"fa",
          4105 => x"a0",
          4106 => x"17",
          4107 => x"39",
          4108 => x"9f",
          4109 => x"5d",
          4110 => x"9c",
          4111 => x"38",
          4112 => x"38",
          4113 => x"81",
          4114 => x"e4",
          4115 => x"2a",
          4116 => x"b4",
          4117 => x"86",
          4118 => x"5d",
          4119 => x"fa",
          4120 => x"52",
          4121 => x"84",
          4122 => x"ff",
          4123 => x"79",
          4124 => x"83",
          4125 => x"ff",
          4126 => x"76",
          4127 => x"81",
          4128 => x"e4",
          4129 => x"2e",
          4130 => x"87",
          4131 => x"0b",
          4132 => x"2e",
          4133 => x"5b",
          4134 => x"84",
          4135 => x"19",
          4136 => x"3f",
          4137 => x"38",
          4138 => x"0c",
          4139 => x"82",
          4140 => x"11",
          4141 => x"0a",
          4142 => x"57",
          4143 => x"2a",
          4144 => x"2a",
          4145 => x"2a",
          4146 => x"83",
          4147 => x"2a",
          4148 => x"05",
          4149 => x"78",
          4150 => x"33",
          4151 => x"09",
          4152 => x"77",
          4153 => x"51",
          4154 => x"80",
          4155 => x"77",
          4156 => x"ac",
          4157 => x"05",
          4158 => x"57",
          4159 => x"7a",
          4160 => x"8f",
          4161 => x"34",
          4162 => x"2a",
          4163 => x"b4",
          4164 => x"83",
          4165 => x"19",
          4166 => x"f0",
          4167 => x"08",
          4168 => x"38",
          4169 => x"b4",
          4170 => x"a0",
          4171 => x"5c",
          4172 => x"82",
          4173 => x"e4",
          4174 => x"81",
          4175 => x"b8",
          4176 => x"56",
          4177 => x"fc",
          4178 => x"b8",
          4179 => x"8f",
          4180 => x"f0",
          4181 => x"74",
          4182 => x"fc",
          4183 => x"19",
          4184 => x"ef",
          4185 => x"08",
          4186 => x"38",
          4187 => x"b4",
          4188 => x"a0",
          4189 => x"59",
          4190 => x"38",
          4191 => x"09",
          4192 => x"76",
          4193 => x"51",
          4194 => x"39",
          4195 => x"53",
          4196 => x"3f",
          4197 => x"2e",
          4198 => x"b8",
          4199 => x"08",
          4200 => x"08",
          4201 => x"5f",
          4202 => x"19",
          4203 => x"06",
          4204 => x"53",
          4205 => x"e4",
          4206 => x"54",
          4207 => x"1a",
          4208 => x"5a",
          4209 => x"81",
          4210 => x"08",
          4211 => x"a8",
          4212 => x"b8",
          4213 => x"7d",
          4214 => x"55",
          4215 => x"fa",
          4216 => x"52",
          4217 => x"7b",
          4218 => x"1c",
          4219 => x"ec",
          4220 => x"7b",
          4221 => x"7c",
          4222 => x"76",
          4223 => x"79",
          4224 => x"58",
          4225 => x"83",
          4226 => x"11",
          4227 => x"7f",
          4228 => x"5d",
          4229 => x"56",
          4230 => x"5a",
          4231 => x"5b",
          4232 => x"f6",
          4233 => x"5c",
          4234 => x"08",
          4235 => x"76",
          4236 => x"94",
          4237 => x"2e",
          4238 => x"93",
          4239 => x"19",
          4240 => x"75",
          4241 => x"79",
          4242 => x"08",
          4243 => x"84",
          4244 => x"84",
          4245 => x"72",
          4246 => x"51",
          4247 => x"77",
          4248 => x"73",
          4249 => x"3d",
          4250 => x"84",
          4251 => x"52",
          4252 => x"74",
          4253 => x"84",
          4254 => x"08",
          4255 => x"84",
          4256 => x"57",
          4257 => x"19",
          4258 => x"75",
          4259 => x"58",
          4260 => x"a0",
          4261 => x"30",
          4262 => x"07",
          4263 => x"55",
          4264 => x"e4",
          4265 => x"08",
          4266 => x"73",
          4267 => x"73",
          4268 => x"80",
          4269 => x"52",
          4270 => x"e4",
          4271 => x"84",
          4272 => x"58",
          4273 => x"e3",
          4274 => x"08",
          4275 => x"74",
          4276 => x"1a",
          4277 => x"79",
          4278 => x"b8",
          4279 => x"0b",
          4280 => x"04",
          4281 => x"39",
          4282 => x"53",
          4283 => x"84",
          4284 => x"84",
          4285 => x"8c",
          4286 => x"2e",
          4287 => x"39",
          4288 => x"59",
          4289 => x"80",
          4290 => x"80",
          4291 => x"18",
          4292 => x"33",
          4293 => x"73",
          4294 => x"22",
          4295 => x"ac",
          4296 => x"19",
          4297 => x"72",
          4298 => x"13",
          4299 => x"17",
          4300 => x"75",
          4301 => x"04",
          4302 => x"3d",
          4303 => x"80",
          4304 => x"70",
          4305 => x"a5",
          4306 => x"fe",
          4307 => x"27",
          4308 => x"29",
          4309 => x"98",
          4310 => x"77",
          4311 => x"08",
          4312 => x"a4",
          4313 => x"27",
          4314 => x"84",
          4315 => x"38",
          4316 => x"cd",
          4317 => x"b8",
          4318 => x"3d",
          4319 => x"a0",
          4320 => x"7a",
          4321 => x"0c",
          4322 => x"80",
          4323 => x"5b",
          4324 => x"08",
          4325 => x"2a",
          4326 => x"27",
          4327 => x"79",
          4328 => x"9c",
          4329 => x"e4",
          4330 => x"18",
          4331 => x"89",
          4332 => x"52",
          4333 => x"e4",
          4334 => x"b8",
          4335 => x"84",
          4336 => x"9c",
          4337 => x"82",
          4338 => x"38",
          4339 => x"a7",
          4340 => x"56",
          4341 => x"9c",
          4342 => x"81",
          4343 => x"b8",
          4344 => x"84",
          4345 => x"58",
          4346 => x"1a",
          4347 => x"75",
          4348 => x"76",
          4349 => x"5e",
          4350 => x"84",
          4351 => x"81",
          4352 => x"f4",
          4353 => x"75",
          4354 => x"75",
          4355 => x"51",
          4356 => x"80",
          4357 => x"7a",
          4358 => x"e4",
          4359 => x"b4",
          4360 => x"81",
          4361 => x"84",
          4362 => x"b8",
          4363 => x"08",
          4364 => x"1a",
          4365 => x"33",
          4366 => x"fe",
          4367 => x"a0",
          4368 => x"19",
          4369 => x"39",
          4370 => x"ff",
          4371 => x"06",
          4372 => x"1d",
          4373 => x"80",
          4374 => x"8a",
          4375 => x"08",
          4376 => x"39",
          4377 => x"3d",
          4378 => x"41",
          4379 => x"ff",
          4380 => x"75",
          4381 => x"5f",
          4382 => x"76",
          4383 => x"78",
          4384 => x"06",
          4385 => x"b8",
          4386 => x"bd",
          4387 => x"85",
          4388 => x"1a",
          4389 => x"9c",
          4390 => x"80",
          4391 => x"bf",
          4392 => x"60",
          4393 => x"70",
          4394 => x"80",
          4395 => x"45",
          4396 => x"df",
          4397 => x"bf",
          4398 => x"81",
          4399 => x"f6",
          4400 => x"b8",
          4401 => x"08",
          4402 => x"b8",
          4403 => x"54",
          4404 => x"19",
          4405 => x"84",
          4406 => x"06",
          4407 => x"83",
          4408 => x"08",
          4409 => x"7a",
          4410 => x"82",
          4411 => x"81",
          4412 => x"19",
          4413 => x"52",
          4414 => x"77",
          4415 => x"09",
          4416 => x"2a",
          4417 => x"38",
          4418 => x"70",
          4419 => x"59",
          4420 => x"81",
          4421 => x"81",
          4422 => x"fe",
          4423 => x"0b",
          4424 => x"0c",
          4425 => x"df",
          4426 => x"2e",
          4427 => x"08",
          4428 => x"88",
          4429 => x"b7",
          4430 => x"8d",
          4431 => x"58",
          4432 => x"05",
          4433 => x"2b",
          4434 => x"80",
          4435 => x"87",
          4436 => x"42",
          4437 => x"17",
          4438 => x"33",
          4439 => x"77",
          4440 => x"26",
          4441 => x"43",
          4442 => x"ff",
          4443 => x"83",
          4444 => x"55",
          4445 => x"55",
          4446 => x"80",
          4447 => x"33",
          4448 => x"ff",
          4449 => x"74",
          4450 => x"ac",
          4451 => x"94",
          4452 => x"70",
          4453 => x"f5",
          4454 => x"84",
          4455 => x"ff",
          4456 => x"0c",
          4457 => x"80",
          4458 => x"cc",
          4459 => x"74",
          4460 => x"38",
          4461 => x"81",
          4462 => x"b8",
          4463 => x"56",
          4464 => x"5a",
          4465 => x"70",
          4466 => x"99",
          4467 => x"81",
          4468 => x"34",
          4469 => x"75",
          4470 => x"2e",
          4471 => x"75",
          4472 => x"38",
          4473 => x"81",
          4474 => x"70",
          4475 => x"70",
          4476 => x"5d",
          4477 => x"cd",
          4478 => x"76",
          4479 => x"57",
          4480 => x"70",
          4481 => x"ff",
          4482 => x"2e",
          4483 => x"38",
          4484 => x"0c",
          4485 => x"84",
          4486 => x"08",
          4487 => x"b8",
          4488 => x"54",
          4489 => x"1b",
          4490 => x"84",
          4491 => x"06",
          4492 => x"83",
          4493 => x"08",
          4494 => x"78",
          4495 => x"82",
          4496 => x"81",
          4497 => x"1b",
          4498 => x"52",
          4499 => x"77",
          4500 => x"e4",
          4501 => x"81",
          4502 => x"76",
          4503 => x"2e",
          4504 => x"bf",
          4505 => x"05",
          4506 => x"af",
          4507 => x"52",
          4508 => x"e4",
          4509 => x"2e",
          4510 => x"80",
          4511 => x"ff",
          4512 => x"8d",
          4513 => x"81",
          4514 => x"1a",
          4515 => x"07",
          4516 => x"78",
          4517 => x"05",
          4518 => x"e4",
          4519 => x"33",
          4520 => x"42",
          4521 => x"79",
          4522 => x"51",
          4523 => x"08",
          4524 => x"43",
          4525 => x"3f",
          4526 => x"81",
          4527 => x"18",
          4528 => x"78",
          4529 => x"59",
          4530 => x"2e",
          4531 => x"22",
          4532 => x"1d",
          4533 => x"ae",
          4534 => x"93",
          4535 => x"2e",
          4536 => x"94",
          4537 => x"70",
          4538 => x"5a",
          4539 => x"38",
          4540 => x"57",
          4541 => x"1d",
          4542 => x"5d",
          4543 => x"5b",
          4544 => x"75",
          4545 => x"81",
          4546 => x"ef",
          4547 => x"81",
          4548 => x"aa",
          4549 => x"81",
          4550 => x"08",
          4551 => x"57",
          4552 => x"76",
          4553 => x"55",
          4554 => x"c2",
          4555 => x"80",
          4556 => x"56",
          4557 => x"07",
          4558 => x"06",
          4559 => x"56",
          4560 => x"84",
          4561 => x"77",
          4562 => x"74",
          4563 => x"cf",
          4564 => x"06",
          4565 => x"15",
          4566 => x"19",
          4567 => x"e3",
          4568 => x"34",
          4569 => x"a0",
          4570 => x"98",
          4571 => x"88",
          4572 => x"57",
          4573 => x"38",
          4574 => x"26",
          4575 => x"05",
          4576 => x"74",
          4577 => x"38",
          4578 => x"e4",
          4579 => x"e3",
          4580 => x"7a",
          4581 => x"b8",
          4582 => x"84",
          4583 => x"02",
          4584 => x"7d",
          4585 => x"33",
          4586 => x"5f",
          4587 => x"8d",
          4588 => x"3f",
          4589 => x"52",
          4590 => x"e4",
          4591 => x"82",
          4592 => x"5e",
          4593 => x"b4",
          4594 => x"83",
          4595 => x"81",
          4596 => x"53",
          4597 => x"d4",
          4598 => x"2e",
          4599 => x"b4",
          4600 => x"9c",
          4601 => x"81",
          4602 => x"70",
          4603 => x"80",
          4604 => x"78",
          4605 => x"7d",
          4606 => x"08",
          4607 => x"ff",
          4608 => x"81",
          4609 => x"38",
          4610 => x"98",
          4611 => x"2e",
          4612 => x"40",
          4613 => x"53",
          4614 => x"d3",
          4615 => x"2e",
          4616 => x"b4",
          4617 => x"38",
          4618 => x"80",
          4619 => x"15",
          4620 => x"1f",
          4621 => x"81",
          4622 => x"59",
          4623 => x"9c",
          4624 => x"5e",
          4625 => x"83",
          4626 => x"e4",
          4627 => x"30",
          4628 => x"57",
          4629 => x"52",
          4630 => x"e4",
          4631 => x"2e",
          4632 => x"54",
          4633 => x"18",
          4634 => x"e4",
          4635 => x"bf",
          4636 => x"34",
          4637 => x"55",
          4638 => x"82",
          4639 => x"ac",
          4640 => x"9c",
          4641 => x"71",
          4642 => x"3f",
          4643 => x"e4",
          4644 => x"e4",
          4645 => x"2a",
          4646 => x"81",
          4647 => x"81",
          4648 => x"76",
          4649 => x"1d",
          4650 => x"56",
          4651 => x"83",
          4652 => x"81",
          4653 => x"53",
          4654 => x"d0",
          4655 => x"2e",
          4656 => x"b4",
          4657 => x"38",
          4658 => x"81",
          4659 => x"1c",
          4660 => x"8c",
          4661 => x"9b",
          4662 => x"76",
          4663 => x"ff",
          4664 => x"22",
          4665 => x"e4",
          4666 => x"70",
          4667 => x"56",
          4668 => x"ff",
          4669 => x"27",
          4670 => x"81",
          4671 => x"58",
          4672 => x"7c",
          4673 => x"80",
          4674 => x"b8",
          4675 => x"fc",
          4676 => x"fe",
          4677 => x"b4",
          4678 => x"81",
          4679 => x"81",
          4680 => x"38",
          4681 => x"b4",
          4682 => x"b8",
          4683 => x"08",
          4684 => x"42",
          4685 => x"bc",
          4686 => x"1d",
          4687 => x"33",
          4688 => x"a4",
          4689 => x"57",
          4690 => x"81",
          4691 => x"81",
          4692 => x"9f",
          4693 => x"07",
          4694 => x"1c",
          4695 => x"51",
          4696 => x"76",
          4697 => x"b8",
          4698 => x"08",
          4699 => x"1d",
          4700 => x"5f",
          4701 => x"e4",
          4702 => x"1c",
          4703 => x"38",
          4704 => x"e8",
          4705 => x"2e",
          4706 => x"54",
          4707 => x"53",
          4708 => x"ac",
          4709 => x"18",
          4710 => x"52",
          4711 => x"f8",
          4712 => x"71",
          4713 => x"1e",
          4714 => x"b5",
          4715 => x"d9",
          4716 => x"08",
          4717 => x"72",
          4718 => x"14",
          4719 => x"7a",
          4720 => x"70",
          4721 => x"8f",
          4722 => x"1a",
          4723 => x"5b",
          4724 => x"25",
          4725 => x"7c",
          4726 => x"18",
          4727 => x"58",
          4728 => x"18",
          4729 => x"38",
          4730 => x"89",
          4731 => x"25",
          4732 => x"38",
          4733 => x"70",
          4734 => x"74",
          4735 => x"18",
          4736 => x"7c",
          4737 => x"16",
          4738 => x"38",
          4739 => x"1e",
          4740 => x"56",
          4741 => x"08",
          4742 => x"38",
          4743 => x"53",
          4744 => x"1c",
          4745 => x"12",
          4746 => x"07",
          4747 => x"2b",
          4748 => x"97",
          4749 => x"2b",
          4750 => x"5b",
          4751 => x"33",
          4752 => x"5d",
          4753 => x"0d",
          4754 => x"77",
          4755 => x"58",
          4756 => x"2b",
          4757 => x"84",
          4758 => x"55",
          4759 => x"76",
          4760 => x"54",
          4761 => x"82",
          4762 => x"08",
          4763 => x"22",
          4764 => x"fd",
          4765 => x"78",
          4766 => x"58",
          4767 => x"7a",
          4768 => x"8c",
          4769 => x"73",
          4770 => x"80",
          4771 => x"7e",
          4772 => x"bf",
          4773 => x"38",
          4774 => x"5b",
          4775 => x"2a",
          4776 => x"2e",
          4777 => x"ff",
          4778 => x"05",
          4779 => x"19",
          4780 => x"56",
          4781 => x"39",
          4782 => x"7b",
          4783 => x"06",
          4784 => x"ef",
          4785 => x"57",
          4786 => x"53",
          4787 => x"74",
          4788 => x"80",
          4789 => x"88",
          4790 => x"3d",
          4791 => x"a7",
          4792 => x"80",
          4793 => x"33",
          4794 => x"7f",
          4795 => x"83",
          4796 => x"10",
          4797 => x"57",
          4798 => x"32",
          4799 => x"25",
          4800 => x"90",
          4801 => x"38",
          4802 => x"e4",
          4803 => x"81",
          4804 => x"2e",
          4805 => x"38",
          4806 => x"06",
          4807 => x"81",
          4808 => x"76",
          4809 => x"10",
          4810 => x"62",
          4811 => x"54",
          4812 => x"80",
          4813 => x"70",
          4814 => x"55",
          4815 => x"81",
          4816 => x"54",
          4817 => x"80",
          4818 => x"77",
          4819 => x"72",
          4820 => x"94",
          4821 => x"fe",
          4822 => x"73",
          4823 => x"e4",
          4824 => x"fe",
          4825 => x"e4",
          4826 => x"80",
          4827 => x"7a",
          4828 => x"ff",
          4829 => x"7b",
          4830 => x"08",
          4831 => x"04",
          4832 => x"70",
          4833 => x"56",
          4834 => x"42",
          4835 => x"72",
          4836 => x"32",
          4837 => x"40",
          4838 => x"0c",
          4839 => x"81",
          4840 => x"83",
          4841 => x"2e",
          4842 => x"05",
          4843 => x"70",
          4844 => x"59",
          4845 => x"38",
          4846 => x"59",
          4847 => x"80",
          4848 => x"70",
          4849 => x"55",
          4850 => x"73",
          4851 => x"2e",
          4852 => x"38",
          4853 => x"54",
          4854 => x"18",
          4855 => x"80",
          4856 => x"5e",
          4857 => x"eb",
          4858 => x"a0",
          4859 => x"13",
          4860 => x"5e",
          4861 => x"59",
          4862 => x"ed",
          4863 => x"74",
          4864 => x"55",
          4865 => x"38",
          4866 => x"7b",
          4867 => x"32",
          4868 => x"70",
          4869 => x"80",
          4870 => x"86",
          4871 => x"79",
          4872 => x"38",
          4873 => x"2b",
          4874 => x"5d",
          4875 => x"56",
          4876 => x"33",
          4877 => x"38",
          4878 => x"8c",
          4879 => x"38",
          4880 => x"82",
          4881 => x"56",
          4882 => x"7c",
          4883 => x"5a",
          4884 => x"80",
          4885 => x"79",
          4886 => x"3f",
          4887 => x"56",
          4888 => x"81",
          4889 => x"2e",
          4890 => x"85",
          4891 => x"84",
          4892 => x"59",
          4893 => x"55",
          4894 => x"80",
          4895 => x"11",
          4896 => x"56",
          4897 => x"2e",
          4898 => x"fd",
          4899 => x"ae",
          4900 => x"77",
          4901 => x"06",
          4902 => x"80",
          4903 => x"53",
          4904 => x"a0",
          4905 => x"34",
          4906 => x"38",
          4907 => x"34",
          4908 => x"e4",
          4909 => x"b8",
          4910 => x"2a",
          4911 => x"86",
          4912 => x"56",
          4913 => x"90",
          4914 => x"80",
          4915 => x"71",
          4916 => x"54",
          4917 => x"74",
          4918 => x"56",
          4919 => x"ae",
          4920 => x"76",
          4921 => x"83",
          4922 => x"39",
          4923 => x"8c",
          4924 => x"81",
          4925 => x"5a",
          4926 => x"34",
          4927 => x"f6",
          4928 => x"1d",
          4929 => x"93",
          4930 => x"9d",
          4931 => x"38",
          4932 => x"f7",
          4933 => x"57",
          4934 => x"07",
          4935 => x"85",
          4936 => x"ff",
          4937 => x"5a",
          4938 => x"80",
          4939 => x"56",
          4940 => x"38",
          4941 => x"e4",
          4942 => x"81",
          4943 => x"2e",
          4944 => x"38",
          4945 => x"06",
          4946 => x"81",
          4947 => x"ff",
          4948 => x"38",
          4949 => x"5f",
          4950 => x"26",
          4951 => x"ff",
          4952 => x"06",
          4953 => x"05",
          4954 => x"75",
          4955 => x"fa",
          4956 => x"81",
          4957 => x"ff",
          4958 => x"7d",
          4959 => x"79",
          4960 => x"cd",
          4961 => x"98",
          4962 => x"88",
          4963 => x"7b",
          4964 => x"54",
          4965 => x"a0",
          4966 => x"1b",
          4967 => x"a0",
          4968 => x"2e",
          4969 => x"a3",
          4970 => x"7b",
          4971 => x"e4",
          4972 => x"0d",
          4973 => x"05",
          4974 => x"ff",
          4975 => x"80",
          4976 => x"05",
          4977 => x"75",
          4978 => x"38",
          4979 => x"d0",
          4980 => x"b2",
          4981 => x"05",
          4982 => x"80",
          4983 => x"7f",
          4984 => x"7b",
          4985 => x"51",
          4986 => x"08",
          4987 => x"58",
          4988 => x"77",
          4989 => x"1d",
          4990 => x"17",
          4991 => x"b8",
          4992 => x"06",
          4993 => x"38",
          4994 => x"2a",
          4995 => x"b1",
          4996 => x"ff",
          4997 => x"55",
          4998 => x"53",
          4999 => x"95",
          5000 => x"85",
          5001 => x"18",
          5002 => x"b7",
          5003 => x"88",
          5004 => x"82",
          5005 => x"81",
          5006 => x"33",
          5007 => x"75",
          5008 => x"75",
          5009 => x"17",
          5010 => x"2b",
          5011 => x"09",
          5012 => x"17",
          5013 => x"2b",
          5014 => x"dc",
          5015 => x"71",
          5016 => x"14",
          5017 => x"33",
          5018 => x"5f",
          5019 => x"17",
          5020 => x"33",
          5021 => x"40",
          5022 => x"d9",
          5023 => x"29",
          5024 => x"77",
          5025 => x"2e",
          5026 => x"42",
          5027 => x"33",
          5028 => x"07",
          5029 => x"75",
          5030 => x"82",
          5031 => x"cb",
          5032 => x"5c",
          5033 => x"11",
          5034 => x"71",
          5035 => x"72",
          5036 => x"53",
          5037 => x"c7",
          5038 => x"88",
          5039 => x"80",
          5040 => x"84",
          5041 => x"c1",
          5042 => x"fd",
          5043 => x"56",
          5044 => x"a9",
          5045 => x"ff",
          5046 => x"75",
          5047 => x"5d",
          5048 => x"81",
          5049 => x"7b",
          5050 => x"1a",
          5051 => x"59",
          5052 => x"17",
          5053 => x"80",
          5054 => x"78",
          5055 => x"78",
          5056 => x"06",
          5057 => x"2a",
          5058 => x"26",
          5059 => x"ff",
          5060 => x"84",
          5061 => x"38",
          5062 => x"81",
          5063 => x"7c",
          5064 => x"8c",
          5065 => x"80",
          5066 => x"3d",
          5067 => x"0c",
          5068 => x"11",
          5069 => x"74",
          5070 => x"81",
          5071 => x"7a",
          5072 => x"83",
          5073 => x"7f",
          5074 => x"33",
          5075 => x"9f",
          5076 => x"89",
          5077 => x"57",
          5078 => x"26",
          5079 => x"06",
          5080 => x"59",
          5081 => x"85",
          5082 => x"32",
          5083 => x"7a",
          5084 => x"87",
          5085 => x"5c",
          5086 => x"56",
          5087 => x"cf",
          5088 => x"8a",
          5089 => x"fe",
          5090 => x"75",
          5091 => x"38",
          5092 => x"30",
          5093 => x"5c",
          5094 => x"2e",
          5095 => x"5a",
          5096 => x"59",
          5097 => x"81",
          5098 => x"90",
          5099 => x"19",
          5100 => x"fe",
          5101 => x"40",
          5102 => x"5c",
          5103 => x"78",
          5104 => x"d9",
          5105 => x"72",
          5106 => x"05",
          5107 => x"52",
          5108 => x"56",
          5109 => x"0b",
          5110 => x"0c",
          5111 => x"a5",
          5112 => x"52",
          5113 => x"3f",
          5114 => x"38",
          5115 => x"0c",
          5116 => x"33",
          5117 => x"5e",
          5118 => x"09",
          5119 => x"18",
          5120 => x"82",
          5121 => x"30",
          5122 => x"42",
          5123 => x"b6",
          5124 => x"56",
          5125 => x"5d",
          5126 => x"83",
          5127 => x"bd",
          5128 => x"81",
          5129 => x"27",
          5130 => x"0b",
          5131 => x"5d",
          5132 => x"7e",
          5133 => x"31",
          5134 => x"80",
          5135 => x"e1",
          5136 => x"e4",
          5137 => x"05",
          5138 => x"33",
          5139 => x"42",
          5140 => x"75",
          5141 => x"f3",
          5142 => x"77",
          5143 => x"04",
          5144 => x"38",
          5145 => x"98",
          5146 => x"0b",
          5147 => x"04",
          5148 => x"94",
          5149 => x"5a",
          5150 => x"71",
          5151 => x"5f",
          5152 => x"80",
          5153 => x"18",
          5154 => x"70",
          5155 => x"05",
          5156 => x"5b",
          5157 => x"91",
          5158 => x"3d",
          5159 => x"39",
          5160 => x"17",
          5161 => x"2b",
          5162 => x"81",
          5163 => x"80",
          5164 => x"38",
          5165 => x"09",
          5166 => x"77",
          5167 => x"51",
          5168 => x"08",
          5169 => x"5a",
          5170 => x"38",
          5171 => x"33",
          5172 => x"07",
          5173 => x"09",
          5174 => x"83",
          5175 => x"2b",
          5176 => x"70",
          5177 => x"07",
          5178 => x"77",
          5179 => x"81",
          5180 => x"83",
          5181 => x"2b",
          5182 => x"70",
          5183 => x"07",
          5184 => x"60",
          5185 => x"81",
          5186 => x"83",
          5187 => x"2b",
          5188 => x"70",
          5189 => x"07",
          5190 => x"83",
          5191 => x"2b",
          5192 => x"70",
          5193 => x"07",
          5194 => x"46",
          5195 => x"7c",
          5196 => x"05",
          5197 => x"86",
          5198 => x"18",
          5199 => x"cf",
          5200 => x"7b",
          5201 => x"75",
          5202 => x"70",
          5203 => x"af",
          5204 => x"2e",
          5205 => x"b8",
          5206 => x"08",
          5207 => x"18",
          5208 => x"41",
          5209 => x"b8",
          5210 => x"56",
          5211 => x"0b",
          5212 => x"5a",
          5213 => x"33",
          5214 => x"07",
          5215 => x"38",
          5216 => x"38",
          5217 => x"12",
          5218 => x"07",
          5219 => x"2b",
          5220 => x"5a",
          5221 => x"59",
          5222 => x"80",
          5223 => x"e3",
          5224 => x"93",
          5225 => x"f2",
          5226 => x"fc",
          5227 => x"a0",
          5228 => x"17",
          5229 => x"85",
          5230 => x"05",
          5231 => x"57",
          5232 => x"2e",
          5233 => x"5a",
          5234 => x"ba",
          5235 => x"74",
          5236 => x"c0",
          5237 => x"38",
          5238 => x"70",
          5239 => x"38",
          5240 => x"2e",
          5241 => x"73",
          5242 => x"92",
          5243 => x"84",
          5244 => x"e4",
          5245 => x"92",
          5246 => x"e4",
          5247 => x"d0",
          5248 => x"57",
          5249 => x"77",
          5250 => x"77",
          5251 => x"08",
          5252 => x"08",
          5253 => x"5b",
          5254 => x"ff",
          5255 => x"26",
          5256 => x"06",
          5257 => x"99",
          5258 => x"ff",
          5259 => x"2a",
          5260 => x"06",
          5261 => x"79",
          5262 => x"2a",
          5263 => x"2e",
          5264 => x"5b",
          5265 => x"54",
          5266 => x"38",
          5267 => x"39",
          5268 => x"80",
          5269 => x"78",
          5270 => x"70",
          5271 => x"3d",
          5272 => x"84",
          5273 => x"08",
          5274 => x"76",
          5275 => x"3d",
          5276 => x"3d",
          5277 => x"b8",
          5278 => x"80",
          5279 => x"5d",
          5280 => x"80",
          5281 => x"83",
          5282 => x"ff",
          5283 => x"5b",
          5284 => x"9b",
          5285 => x"2b",
          5286 => x"5e",
          5287 => x"80",
          5288 => x"17",
          5289 => x"cc",
          5290 => x"0b",
          5291 => x"80",
          5292 => x"17",
          5293 => x"84",
          5294 => x"1c",
          5295 => x"0b",
          5296 => x"34",
          5297 => x"7b",
          5298 => x"11",
          5299 => x"57",
          5300 => x"08",
          5301 => x"80",
          5302 => x"e7",
          5303 => x"7b",
          5304 => x"9c",
          5305 => x"76",
          5306 => x"33",
          5307 => x"7b",
          5308 => x"06",
          5309 => x"81",
          5310 => x"83",
          5311 => x"86",
          5312 => x"b4",
          5313 => x"1b",
          5314 => x"33",
          5315 => x"5e",
          5316 => x"f1",
          5317 => x"83",
          5318 => x"2b",
          5319 => x"70",
          5320 => x"07",
          5321 => x"0c",
          5322 => x"86",
          5323 => x"1a",
          5324 => x"0b",
          5325 => x"06",
          5326 => x"75",
          5327 => x"1a",
          5328 => x"7c",
          5329 => x"07",
          5330 => x"84",
          5331 => x"5b",
          5332 => x"52",
          5333 => x"b8",
          5334 => x"81",
          5335 => x"e4",
          5336 => x"7a",
          5337 => x"05",
          5338 => x"77",
          5339 => x"2e",
          5340 => x"0c",
          5341 => x"0c",
          5342 => x"0c",
          5343 => x"3f",
          5344 => x"59",
          5345 => x"39",
          5346 => x"f3",
          5347 => x"71",
          5348 => x"07",
          5349 => x"55",
          5350 => x"52",
          5351 => x"b8",
          5352 => x"80",
          5353 => x"08",
          5354 => x"e4",
          5355 => x"53",
          5356 => x"3f",
          5357 => x"9c",
          5358 => x"58",
          5359 => x"38",
          5360 => x"33",
          5361 => x"7c",
          5362 => x"80",
          5363 => x"80",
          5364 => x"95",
          5365 => x"2b",
          5366 => x"56",
          5367 => x"0b",
          5368 => x"34",
          5369 => x"56",
          5370 => x"57",
          5371 => x"0b",
          5372 => x"83",
          5373 => x"ff",
          5374 => x"59",
          5375 => x"ae",
          5376 => x"2e",
          5377 => x"7d",
          5378 => x"51",
          5379 => x"08",
          5380 => x"5b",
          5381 => x"ff",
          5382 => x"2e",
          5383 => x"97",
          5384 => x"b8",
          5385 => x"5a",
          5386 => x"08",
          5387 => x"38",
          5388 => x"b4",
          5389 => x"b8",
          5390 => x"08",
          5391 => x"55",
          5392 => x"85",
          5393 => x"17",
          5394 => x"33",
          5395 => x"fe",
          5396 => x"56",
          5397 => x"76",
          5398 => x"5a",
          5399 => x"fe",
          5400 => x"59",
          5401 => x"8a",
          5402 => x"08",
          5403 => x"cd",
          5404 => x"0c",
          5405 => x"1a",
          5406 => x"57",
          5407 => x"b8",
          5408 => x"cf",
          5409 => x"39",
          5410 => x"40",
          5411 => x"57",
          5412 => x"56",
          5413 => x"55",
          5414 => x"22",
          5415 => x"2e",
          5416 => x"76",
          5417 => x"33",
          5418 => x"33",
          5419 => x"2e",
          5420 => x"1b",
          5421 => x"26",
          5422 => x"d5",
          5423 => x"5b",
          5424 => x"ff",
          5425 => x"9b",
          5426 => x"08",
          5427 => x"74",
          5428 => x"1b",
          5429 => x"05",
          5430 => x"76",
          5431 => x"22",
          5432 => x"56",
          5433 => x"7a",
          5434 => x"80",
          5435 => x"75",
          5436 => x"58",
          5437 => x"19",
          5438 => x"b8",
          5439 => x"11",
          5440 => x"38",
          5441 => x"78",
          5442 => x"29",
          5443 => x"70",
          5444 => x"05",
          5445 => x"38",
          5446 => x"7e",
          5447 => x"1c",
          5448 => x"5e",
          5449 => x"75",
          5450 => x"04",
          5451 => x"0d",
          5452 => x"1a",
          5453 => x"80",
          5454 => x"83",
          5455 => x"08",
          5456 => x"1a",
          5457 => x"2e",
          5458 => x"54",
          5459 => x"33",
          5460 => x"e4",
          5461 => x"81",
          5462 => x"dc",
          5463 => x"06",
          5464 => x"56",
          5465 => x"74",
          5466 => x"81",
          5467 => x"80",
          5468 => x"05",
          5469 => x"34",
          5470 => x"bc",
          5471 => x"b8",
          5472 => x"40",
          5473 => x"b8",
          5474 => x"ff",
          5475 => x"1a",
          5476 => x"31",
          5477 => x"a0",
          5478 => x"19",
          5479 => x"06",
          5480 => x"08",
          5481 => x"81",
          5482 => x"7e",
          5483 => x"0c",
          5484 => x"98",
          5485 => x"98",
          5486 => x"a1",
          5487 => x"83",
          5488 => x"55",
          5489 => x"56",
          5490 => x"1b",
          5491 => x"92",
          5492 => x"34",
          5493 => x"3d",
          5494 => x"67",
          5495 => x"0c",
          5496 => x"79",
          5497 => x"75",
          5498 => x"86",
          5499 => x"78",
          5500 => x"74",
          5501 => x"91",
          5502 => x"90",
          5503 => x"58",
          5504 => x"a1",
          5505 => x"57",
          5506 => x"5b",
          5507 => x"83",
          5508 => x"60",
          5509 => x"2a",
          5510 => x"84",
          5511 => x"80",
          5512 => x"86",
          5513 => x"38",
          5514 => x"85",
          5515 => x"b4",
          5516 => x"d3",
          5517 => x"17",
          5518 => x"27",
          5519 => x"79",
          5520 => x"74",
          5521 => x"7b",
          5522 => x"83",
          5523 => x"27",
          5524 => x"54",
          5525 => x"51",
          5526 => x"08",
          5527 => x"7d",
          5528 => x"38",
          5529 => x"29",
          5530 => x"05",
          5531 => x"34",
          5532 => x"59",
          5533 => x"59",
          5534 => x"0c",
          5535 => x"71",
          5536 => x"5a",
          5537 => x"38",
          5538 => x"fe",
          5539 => x"80",
          5540 => x"80",
          5541 => x"3d",
          5542 => x"92",
          5543 => x"74",
          5544 => x"39",
          5545 => x"83",
          5546 => x"5c",
          5547 => x"77",
          5548 => x"38",
          5549 => x"41",
          5550 => x"80",
          5551 => x"16",
          5552 => x"cd",
          5553 => x"85",
          5554 => x"17",
          5555 => x"1b",
          5556 => x"b8",
          5557 => x"2e",
          5558 => x"33",
          5559 => x"16",
          5560 => x"0b",
          5561 => x"54",
          5562 => x"53",
          5563 => x"f4",
          5564 => x"7f",
          5565 => x"84",
          5566 => x"16",
          5567 => x"e4",
          5568 => x"27",
          5569 => x"74",
          5570 => x"38",
          5571 => x"08",
          5572 => x"51",
          5573 => x"ca",
          5574 => x"08",
          5575 => x"40",
          5576 => x"12",
          5577 => x"7c",
          5578 => x"98",
          5579 => x"e7",
          5580 => x"b8",
          5581 => x"33",
          5582 => x"51",
          5583 => x"08",
          5584 => x"38",
          5585 => x"53",
          5586 => x"52",
          5587 => x"e4",
          5588 => x"08",
          5589 => x"17",
          5590 => x"27",
          5591 => x"7b",
          5592 => x"38",
          5593 => x"08",
          5594 => x"51",
          5595 => x"89",
          5596 => x"9b",
          5597 => x"55",
          5598 => x"56",
          5599 => x"16",
          5600 => x"17",
          5601 => x"84",
          5602 => x"b8",
          5603 => x"08",
          5604 => x"17",
          5605 => x"33",
          5606 => x"fe",
          5607 => x"a0",
          5608 => x"16",
          5609 => x"7c",
          5610 => x"56",
          5611 => x"34",
          5612 => x"3d",
          5613 => x"82",
          5614 => x"0d",
          5615 => x"5a",
          5616 => x"56",
          5617 => x"55",
          5618 => x"22",
          5619 => x"2e",
          5620 => x"79",
          5621 => x"33",
          5622 => x"7a",
          5623 => x"19",
          5624 => x"2e",
          5625 => x"81",
          5626 => x"17",
          5627 => x"f5",
          5628 => x"85",
          5629 => x"18",
          5630 => x"08",
          5631 => x"78",
          5632 => x"08",
          5633 => x"56",
          5634 => x"5a",
          5635 => x"33",
          5636 => x"2e",
          5637 => x"74",
          5638 => x"9d",
          5639 => x"9e",
          5640 => x"9f",
          5641 => x"97",
          5642 => x"80",
          5643 => x"92",
          5644 => x"7b",
          5645 => x"51",
          5646 => x"08",
          5647 => x"56",
          5648 => x"e4",
          5649 => x"b4",
          5650 => x"81",
          5651 => x"3f",
          5652 => x"c9",
          5653 => x"34",
          5654 => x"84",
          5655 => x"18",
          5656 => x"33",
          5657 => x"fe",
          5658 => x"a0",
          5659 => x"17",
          5660 => x"56",
          5661 => x"74",
          5662 => x"75",
          5663 => x"74",
          5664 => x"9d",
          5665 => x"9e",
          5666 => x"9f",
          5667 => x"97",
          5668 => x"80",
          5669 => x"92",
          5670 => x"7b",
          5671 => x"51",
          5672 => x"08",
          5673 => x"56",
          5674 => x"81",
          5675 => x"84",
          5676 => x"fc",
          5677 => x"fc",
          5678 => x"52",
          5679 => x"08",
          5680 => x"89",
          5681 => x"08",
          5682 => x"33",
          5683 => x"13",
          5684 => x"77",
          5685 => x"75",
          5686 => x"73",
          5687 => x"04",
          5688 => x"3f",
          5689 => x"72",
          5690 => x"d5",
          5691 => x"5b",
          5692 => x"75",
          5693 => x"26",
          5694 => x"70",
          5695 => x"84",
          5696 => x"90",
          5697 => x"0b",
          5698 => x"04",
          5699 => x"3d",
          5700 => x"81",
          5701 => x"26",
          5702 => x"06",
          5703 => x"80",
          5704 => x"5b",
          5705 => x"70",
          5706 => x"05",
          5707 => x"52",
          5708 => x"70",
          5709 => x"13",
          5710 => x"13",
          5711 => x"30",
          5712 => x"2e",
          5713 => x"be",
          5714 => x"72",
          5715 => x"52",
          5716 => x"84",
          5717 => x"99",
          5718 => x"83",
          5719 => x"fe",
          5720 => x"98",
          5721 => x"d1",
          5722 => x"84",
          5723 => x"74",
          5724 => x"04",
          5725 => x"05",
          5726 => x"08",
          5727 => x"38",
          5728 => x"2b",
          5729 => x"38",
          5730 => x"81",
          5731 => x"38",
          5732 => x"33",
          5733 => x"5a",
          5734 => x"38",
          5735 => x"e4",
          5736 => x"e4",
          5737 => x"8f",
          5738 => x"98",
          5739 => x"17",
          5740 => x"07",
          5741 => x"cc",
          5742 => x"74",
          5743 => x"04",
          5744 => x"08",
          5745 => x"7c",
          5746 => x"b4",
          5747 => x"c5",
          5748 => x"b8",
          5749 => x"d9",
          5750 => x"80",
          5751 => x"08",
          5752 => x"38",
          5753 => x"a0",
          5754 => x"84",
          5755 => x"08",
          5756 => x"08",
          5757 => x"b1",
          5758 => x"33",
          5759 => x"54",
          5760 => x"33",
          5761 => x"e4",
          5762 => x"81",
          5763 => x"d4",
          5764 => x"33",
          5765 => x"63",
          5766 => x"78",
          5767 => x"db",
          5768 => x"a3",
          5769 => x"84",
          5770 => x"52",
          5771 => x"b8",
          5772 => x"bb",
          5773 => x"33",
          5774 => x"63",
          5775 => x"7d",
          5776 => x"2e",
          5777 => x"7a",
          5778 => x"e4",
          5779 => x"2e",
          5780 => x"d8",
          5781 => x"3d",
          5782 => x"bd",
          5783 => x"5b",
          5784 => x"1f",
          5785 => x"5f",
          5786 => x"56",
          5787 => x"80",
          5788 => x"56",
          5789 => x"ff",
          5790 => x"75",
          5791 => x"18",
          5792 => x"af",
          5793 => x"79",
          5794 => x"8a",
          5795 => x"70",
          5796 => x"08",
          5797 => x"7e",
          5798 => x"17",
          5799 => x"38",
          5800 => x"38",
          5801 => x"76",
          5802 => x"05",
          5803 => x"26",
          5804 => x"5e",
          5805 => x"81",
          5806 => x"78",
          5807 => x"0d",
          5808 => x"71",
          5809 => x"07",
          5810 => x"16",
          5811 => x"71",
          5812 => x"3d",
          5813 => x"ff",
          5814 => x"59",
          5815 => x"96",
          5816 => x"16",
          5817 => x"17",
          5818 => x"81",
          5819 => x"38",
          5820 => x"b4",
          5821 => x"b8",
          5822 => x"08",
          5823 => x"55",
          5824 => x"f6",
          5825 => x"17",
          5826 => x"33",
          5827 => x"fb",
          5828 => x"08",
          5829 => x"0b",
          5830 => x"83",
          5831 => x"43",
          5832 => x"09",
          5833 => x"39",
          5834 => x"59",
          5835 => x"5e",
          5836 => x"80",
          5837 => x"5a",
          5838 => x"34",
          5839 => x"39",
          5840 => x"b8",
          5841 => x"f7",
          5842 => x"56",
          5843 => x"54",
          5844 => x"53",
          5845 => x"22",
          5846 => x"2e",
          5847 => x"75",
          5848 => x"33",
          5849 => x"08",
          5850 => x"94",
          5851 => x"2e",
          5852 => x"70",
          5853 => x"2e",
          5854 => x"51",
          5855 => x"08",
          5856 => x"53",
          5857 => x"08",
          5858 => x"74",
          5859 => x"31",
          5860 => x"80",
          5861 => x"81",
          5862 => x"08",
          5863 => x"70",
          5864 => x"78",
          5865 => x"74",
          5866 => x"e4",
          5867 => x"2e",
          5868 => x"38",
          5869 => x"53",
          5870 => x"38",
          5871 => x"81",
          5872 => x"84",
          5873 => x"90",
          5874 => x"55",
          5875 => x"16",
          5876 => x"2e",
          5877 => x"94",
          5878 => x"74",
          5879 => x"90",
          5880 => x"90",
          5881 => x"78",
          5882 => x"78",
          5883 => x"80",
          5884 => x"0d",
          5885 => x"15",
          5886 => x"38",
          5887 => x"80",
          5888 => x"e4",
          5889 => x"16",
          5890 => x"80",
          5891 => x"12",
          5892 => x"78",
          5893 => x"74",
          5894 => x"89",
          5895 => x"2e",
          5896 => x"fe",
          5897 => x"89",
          5898 => x"fe",
          5899 => x"82",
          5900 => x"06",
          5901 => x"08",
          5902 => x"74",
          5903 => x"e4",
          5904 => x"2e",
          5905 => x"2e",
          5906 => x"88",
          5907 => x"dc",
          5908 => x"0b",
          5909 => x"04",
          5910 => x"75",
          5911 => x"3d",
          5912 => x"51",
          5913 => x"55",
          5914 => x"38",
          5915 => x"b8",
          5916 => x"76",
          5917 => x"97",
          5918 => x"b8",
          5919 => x"33",
          5920 => x"24",
          5921 => x"2a",
          5922 => x"80",
          5923 => x"33",
          5924 => x"7d",
          5925 => x"78",
          5926 => x"0c",
          5927 => x"23",
          5928 => x"3f",
          5929 => x"2e",
          5930 => x"38",
          5931 => x"55",
          5932 => x"17",
          5933 => x"71",
          5934 => x"0c",
          5935 => x"0d",
          5936 => x"9e",
          5937 => x"96",
          5938 => x"8e",
          5939 => x"57",
          5940 => x"52",
          5941 => x"0c",
          5942 => x"0d",
          5943 => x"c3",
          5944 => x"52",
          5945 => x"54",
          5946 => x"58",
          5947 => x"38",
          5948 => x"38",
          5949 => x"38",
          5950 => x"53",
          5951 => x"53",
          5952 => x"38",
          5953 => x"52",
          5954 => x"b8",
          5955 => x"84",
          5956 => x"a6",
          5957 => x"92",
          5958 => x"be",
          5959 => x"70",
          5960 => x"b8",
          5961 => x"84",
          5962 => x"75",
          5963 => x"e2",
          5964 => x"8e",
          5965 => x"70",
          5966 => x"b8",
          5967 => x"39",
          5968 => x"3f",
          5969 => x"0c",
          5970 => x"51",
          5971 => x"08",
          5972 => x"72",
          5973 => x"ed",
          5974 => x"3d",
          5975 => x"a5",
          5976 => x"b8",
          5977 => x"84",
          5978 => x"65",
          5979 => x"84",
          5980 => x"08",
          5981 => x"70",
          5982 => x"97",
          5983 => x"52",
          5984 => x"84",
          5985 => x"86",
          5986 => x"0d",
          5987 => x"5f",
          5988 => x"96",
          5989 => x"e4",
          5990 => x"38",
          5991 => x"08",
          5992 => x"59",
          5993 => x"7f",
          5994 => x"3d",
          5995 => x"33",
          5996 => x"38",
          5997 => x"08",
          5998 => x"7b",
          5999 => x"17",
          6000 => x"17",
          6001 => x"38",
          6002 => x"81",
          6003 => x"84",
          6004 => x"ff",
          6005 => x"7f",
          6006 => x"76",
          6007 => x"38",
          6008 => x"82",
          6009 => x"2b",
          6010 => x"88",
          6011 => x"fe",
          6012 => x"25",
          6013 => x"06",
          6014 => x"54",
          6015 => x"fe",
          6016 => x"18",
          6017 => x"77",
          6018 => x"0c",
          6019 => x"17",
          6020 => x"18",
          6021 => x"81",
          6022 => x"38",
          6023 => x"b4",
          6024 => x"b8",
          6025 => x"08",
          6026 => x"55",
          6027 => x"b0",
          6028 => x"18",
          6029 => x"33",
          6030 => x"fe",
          6031 => x"59",
          6032 => x"80",
          6033 => x"80",
          6034 => x"2e",
          6035 => x"30",
          6036 => x"25",
          6037 => x"5c",
          6038 => x"38",
          6039 => x"84",
          6040 => x"18",
          6041 => x"05",
          6042 => x"2b",
          6043 => x"82",
          6044 => x"5d",
          6045 => x"83",
          6046 => x"bf",
          6047 => x"0c",
          6048 => x"81",
          6049 => x"83",
          6050 => x"f7",
          6051 => x"80",
          6052 => x"80",
          6053 => x"80",
          6054 => x"18",
          6055 => x"da",
          6056 => x"dc",
          6057 => x"d4",
          6058 => x"81",
          6059 => x"2e",
          6060 => x"73",
          6061 => x"81",
          6062 => x"57",
          6063 => x"16",
          6064 => x"80",
          6065 => x"8c",
          6066 => x"78",
          6067 => x"38",
          6068 => x"84",
          6069 => x"78",
          6070 => x"73",
          6071 => x"84",
          6072 => x"08",
          6073 => x"e4",
          6074 => x"b8",
          6075 => x"80",
          6076 => x"81",
          6077 => x"38",
          6078 => x"08",
          6079 => x"af",
          6080 => x"16",
          6081 => x"34",
          6082 => x"38",
          6083 => x"f6",
          6084 => x"06",
          6085 => x"08",
          6086 => x"90",
          6087 => x"0b",
          6088 => x"17",
          6089 => x"3f",
          6090 => x"c2",
          6091 => x"81",
          6092 => x"58",
          6093 => x"27",
          6094 => x"98",
          6095 => x"81",
          6096 => x"a1",
          6097 => x"08",
          6098 => x"97",
          6099 => x"ff",
          6100 => x"55",
          6101 => x"73",
          6102 => x"84",
          6103 => x"08",
          6104 => x"e4",
          6105 => x"b8",
          6106 => x"80",
          6107 => x"89",
          6108 => x"38",
          6109 => x"08",
          6110 => x"38",
          6111 => x"33",
          6112 => x"78",
          6113 => x"80",
          6114 => x"fc",
          6115 => x"82",
          6116 => x"e4",
          6117 => x"90",
          6118 => x"84",
          6119 => x"54",
          6120 => x"33",
          6121 => x"e4",
          6122 => x"bb",
          6123 => x"3d",
          6124 => x"ff",
          6125 => x"56",
          6126 => x"38",
          6127 => x"0d",
          6128 => x"9b",
          6129 => x"3f",
          6130 => x"e4",
          6131 => x"33",
          6132 => x"86",
          6133 => x"5b",
          6134 => x"ee",
          6135 => x"87",
          6136 => x"3d",
          6137 => x"71",
          6138 => x"5c",
          6139 => x"38",
          6140 => x"80",
          6141 => x"18",
          6142 => x"5f",
          6143 => x"8f",
          6144 => x"3f",
          6145 => x"e4",
          6146 => x"08",
          6147 => x"84",
          6148 => x"08",
          6149 => x"0c",
          6150 => x"94",
          6151 => x"2b",
          6152 => x"98",
          6153 => x"88",
          6154 => x"38",
          6155 => x"5d",
          6156 => x"74",
          6157 => x"84",
          6158 => x"08",
          6159 => x"77",
          6160 => x"2e",
          6161 => x"7a",
          6162 => x"89",
          6163 => x"fd",
          6164 => x"7d",
          6165 => x"e4",
          6166 => x"0d",
          6167 => x"56",
          6168 => x"82",
          6169 => x"55",
          6170 => x"dd",
          6171 => x"52",
          6172 => x"3f",
          6173 => x"38",
          6174 => x"0c",
          6175 => x"08",
          6176 => x"18",
          6177 => x"ec",
          6178 => x"de",
          6179 => x"b8",
          6180 => x"75",
          6181 => x"38",
          6182 => x"b4",
          6183 => x"33",
          6184 => x"84",
          6185 => x"06",
          6186 => x"83",
          6187 => x"08",
          6188 => x"74",
          6189 => x"82",
          6190 => x"81",
          6191 => x"17",
          6192 => x"52",
          6193 => x"3f",
          6194 => x"79",
          6195 => x"78",
          6196 => x"e4",
          6197 => x"2e",
          6198 => x"81",
          6199 => x"08",
          6200 => x"74",
          6201 => x"84",
          6202 => x"08",
          6203 => x"58",
          6204 => x"16",
          6205 => x"07",
          6206 => x"77",
          6207 => x"fd",
          6208 => x"84",
          6209 => x"81",
          6210 => x"82",
          6211 => x"a0",
          6212 => x"b8",
          6213 => x"80",
          6214 => x"0c",
          6215 => x"52",
          6216 => x"bf",
          6217 => x"b8",
          6218 => x"b8",
          6219 => x"b8",
          6220 => x"cb",
          6221 => x"85",
          6222 => x"74",
          6223 => x"8f",
          6224 => x"3f",
          6225 => x"84",
          6226 => x"84",
          6227 => x"38",
          6228 => x"cb",
          6229 => x"b8",
          6230 => x"57",
          6231 => x"18",
          6232 => x"75",
          6233 => x"76",
          6234 => x"58",
          6235 => x"84",
          6236 => x"81",
          6237 => x"f4",
          6238 => x"77",
          6239 => x"77",
          6240 => x"51",
          6241 => x"08",
          6242 => x"39",
          6243 => x"b4",
          6244 => x"81",
          6245 => x"3f",
          6246 => x"38",
          6247 => x"b4",
          6248 => x"74",
          6249 => x"82",
          6250 => x"81",
          6251 => x"17",
          6252 => x"52",
          6253 => x"3f",
          6254 => x"08",
          6255 => x"38",
          6256 => x"38",
          6257 => x"3f",
          6258 => x"e4",
          6259 => x"b8",
          6260 => x"84",
          6261 => x"38",
          6262 => x"f9",
          6263 => x"f3",
          6264 => x"19",
          6265 => x"90",
          6266 => x"17",
          6267 => x"34",
          6268 => x"38",
          6269 => x"0d",
          6270 => x"ff",
          6271 => x"2e",
          6272 => x"0b",
          6273 => x"81",
          6274 => x"f4",
          6275 => x"34",
          6276 => x"34",
          6277 => x"75",
          6278 => x"d0",
          6279 => x"1a",
          6280 => x"59",
          6281 => x"88",
          6282 => x"75",
          6283 => x"38",
          6284 => x"b8",
          6285 => x"05",
          6286 => x"34",
          6287 => x"56",
          6288 => x"7e",
          6289 => x"57",
          6290 => x"2a",
          6291 => x"33",
          6292 => x"7d",
          6293 => x"51",
          6294 => x"08",
          6295 => x"38",
          6296 => x"17",
          6297 => x"34",
          6298 => x"0b",
          6299 => x"77",
          6300 => x"78",
          6301 => x"83",
          6302 => x"0b",
          6303 => x"83",
          6304 => x"3f",
          6305 => x"b8",
          6306 => x"90",
          6307 => x"74",
          6308 => x"34",
          6309 => x"7a",
          6310 => x"55",
          6311 => x"a0",
          6312 => x"58",
          6313 => x"58",
          6314 => x"5c",
          6315 => x"0b",
          6316 => x"83",
          6317 => x"3f",
          6318 => x"39",
          6319 => x"08",
          6320 => x"9b",
          6321 => x"70",
          6322 => x"81",
          6323 => x"2e",
          6324 => x"fe",
          6325 => x"ab",
          6326 => x"84",
          6327 => x"75",
          6328 => x"04",
          6329 => x"52",
          6330 => x"af",
          6331 => x"b8",
          6332 => x"05",
          6333 => x"7c",
          6334 => x"3d",
          6335 => x"05",
          6336 => x"34",
          6337 => x"3d",
          6338 => x"75",
          6339 => x"81",
          6340 => x"ef",
          6341 => x"ff",
          6342 => x"56",
          6343 => x"6a",
          6344 => x"88",
          6345 => x"0d",
          6346 => x"ff",
          6347 => x"91",
          6348 => x"d0",
          6349 => x"fa",
          6350 => x"70",
          6351 => x"7a",
          6352 => x"81",
          6353 => x"58",
          6354 => x"16",
          6355 => x"9f",
          6356 => x"e0",
          6357 => x"75",
          6358 => x"77",
          6359 => x"ff",
          6360 => x"70",
          6361 => x"58",
          6362 => x"1c",
          6363 => x"fd",
          6364 => x"ff",
          6365 => x"38",
          6366 => x"fe",
          6367 => x"a8",
          6368 => x"84",
          6369 => x"b8",
          6370 => x"81",
          6371 => x"8d",
          6372 => x"84",
          6373 => x"58",
          6374 => x"80",
          6375 => x"81",
          6376 => x"57",
          6377 => x"02",
          6378 => x"8b",
          6379 => x"40",
          6380 => x"57",
          6381 => x"0b",
          6382 => x"84",
          6383 => x"2e",
          6384 => x"2e",
          6385 => x"9a",
          6386 => x"33",
          6387 => x"82",
          6388 => x"fe",
          6389 => x"c7",
          6390 => x"b0",
          6391 => x"2e",
          6392 => x"b4",
          6393 => x"17",
          6394 => x"54",
          6395 => x"33",
          6396 => x"e4",
          6397 => x"81",
          6398 => x"7b",
          6399 => x"bf",
          6400 => x"2e",
          6401 => x"83",
          6402 => x"f2",
          6403 => x"80",
          6404 => x"83",
          6405 => x"90",
          6406 => x"7d",
          6407 => x"34",
          6408 => x"78",
          6409 => x"57",
          6410 => x"74",
          6411 => x"84",
          6412 => x"08",
          6413 => x"19",
          6414 => x"77",
          6415 => x"59",
          6416 => x"81",
          6417 => x"16",
          6418 => x"bd",
          6419 => x"85",
          6420 => x"17",
          6421 => x"19",
          6422 => x"83",
          6423 => x"a5",
          6424 => x"ae",
          6425 => x"b8",
          6426 => x"82",
          6427 => x"74",
          6428 => x"fe",
          6429 => x"84",
          6430 => x"82",
          6431 => x"0d",
          6432 => x"71",
          6433 => x"07",
          6434 => x"b8",
          6435 => x"84",
          6436 => x"38",
          6437 => x"0d",
          6438 => x"7b",
          6439 => x"94",
          6440 => x"7a",
          6441 => x"84",
          6442 => x"16",
          6443 => x"e4",
          6444 => x"27",
          6445 => x"7c",
          6446 => x"38",
          6447 => x"08",
          6448 => x"51",
          6449 => x"fa",
          6450 => x"b8",
          6451 => x"5b",
          6452 => x"b8",
          6453 => x"e4",
          6454 => x"a8",
          6455 => x"5d",
          6456 => x"8e",
          6457 => x"2e",
          6458 => x"54",
          6459 => x"53",
          6460 => x"e0",
          6461 => x"ec",
          6462 => x"02",
          6463 => x"57",
          6464 => x"97",
          6465 => x"b8",
          6466 => x"80",
          6467 => x"0c",
          6468 => x"52",
          6469 => x"d7",
          6470 => x"b8",
          6471 => x"05",
          6472 => x"73",
          6473 => x"09",
          6474 => x"06",
          6475 => x"17",
          6476 => x"34",
          6477 => x"b8",
          6478 => x"3d",
          6479 => x"82",
          6480 => x"3d",
          6481 => x"e4",
          6482 => x"2e",
          6483 => x"96",
          6484 => x"96",
          6485 => x"3f",
          6486 => x"e4",
          6487 => x"33",
          6488 => x"d2",
          6489 => x"22",
          6490 => x"76",
          6491 => x"74",
          6492 => x"77",
          6493 => x"73",
          6494 => x"83",
          6495 => x"3f",
          6496 => x"0c",
          6497 => x"6b",
          6498 => x"cc",
          6499 => x"c5",
          6500 => x"e4",
          6501 => x"07",
          6502 => x"2e",
          6503 => x"56",
          6504 => x"78",
          6505 => x"2e",
          6506 => x"5a",
          6507 => x"7c",
          6508 => x"b4",
          6509 => x"83",
          6510 => x"2e",
          6511 => x"54",
          6512 => x"33",
          6513 => x"e4",
          6514 => x"81",
          6515 => x"78",
          6516 => x"80",
          6517 => x"80",
          6518 => x"a7",
          6519 => x"33",
          6520 => x"88",
          6521 => x"07",
          6522 => x"0c",
          6523 => x"84",
          6524 => x"7c",
          6525 => x"70",
          6526 => x"b8",
          6527 => x"80",
          6528 => x"09",
          6529 => x"34",
          6530 => x"b4",
          6531 => x"81",
          6532 => x"3f",
          6533 => x"2e",
          6534 => x"b8",
          6535 => x"08",
          6536 => x"08",
          6537 => x"fe",
          6538 => x"82",
          6539 => x"77",
          6540 => x"05",
          6541 => x"fe",
          6542 => x"76",
          6543 => x"51",
          6544 => x"08",
          6545 => x"39",
          6546 => x"3f",
          6547 => x"e4",
          6548 => x"08",
          6549 => x"59",
          6550 => x"59",
          6551 => x"59",
          6552 => x"1c",
          6553 => x"2e",
          6554 => x"70",
          6555 => x"ea",
          6556 => x"ba",
          6557 => x"3d",
          6558 => x"ff",
          6559 => x"56",
          6560 => x"8f",
          6561 => x"76",
          6562 => x"55",
          6563 => x"70",
          6564 => x"58",
          6565 => x"a2",
          6566 => x"ff",
          6567 => x"f5",
          6568 => x"ff",
          6569 => x"95",
          6570 => x"08",
          6571 => x"08",
          6572 => x"2e",
          6573 => x"83",
          6574 => x"5b",
          6575 => x"38",
          6576 => x"81",
          6577 => x"57",
          6578 => x"74",
          6579 => x"75",
          6580 => x"38",
          6581 => x"79",
          6582 => x"77",
          6583 => x"74",
          6584 => x"1a",
          6585 => x"34",
          6586 => x"70",
          6587 => x"77",
          6588 => x"33",
          6589 => x"bc",
          6590 => x"b7",
          6591 => x"5c",
          6592 => x"38",
          6593 => x"45",
          6594 => x"52",
          6595 => x"e4",
          6596 => x"2e",
          6597 => x"e4",
          6598 => x"52",
          6599 => x"e4",
          6600 => x"fd",
          6601 => x"e4",
          6602 => x"f4",
          6603 => x"75",
          6604 => x"e4",
          6605 => x"c1",
          6606 => x"8b",
          6607 => x"81",
          6608 => x"58",
          6609 => x"7d",
          6610 => x"51",
          6611 => x"08",
          6612 => x"7a",
          6613 => x"9c",
          6614 => x"09",
          6615 => x"79",
          6616 => x"75",
          6617 => x"3f",
          6618 => x"e4",
          6619 => x"84",
          6620 => x"5c",
          6621 => x"b4",
          6622 => x"18",
          6623 => x"06",
          6624 => x"b8",
          6625 => x"d5",
          6626 => x"2e",
          6627 => x"b4",
          6628 => x"78",
          6629 => x"57",
          6630 => x"74",
          6631 => x"5c",
          6632 => x"1a",
          6633 => x"52",
          6634 => x"b8",
          6635 => x"80",
          6636 => x"84",
          6637 => x"fd",
          6638 => x"76",
          6639 => x"55",
          6640 => x"8b",
          6641 => x"55",
          6642 => x"70",
          6643 => x"74",
          6644 => x"81",
          6645 => x"58",
          6646 => x"fd",
          6647 => x"7d",
          6648 => x"51",
          6649 => x"08",
          6650 => x"df",
          6651 => x"7a",
          6652 => x"ec",
          6653 => x"09",
          6654 => x"e4",
          6655 => x"a8",
          6656 => x"08",
          6657 => x"74",
          6658 => x"08",
          6659 => x"52",
          6660 => x"b8",
          6661 => x"80",
          6662 => x"81",
          6663 => x"e7",
          6664 => x"18",
          6665 => x"52",
          6666 => x"3f",
          6667 => x"62",
          6668 => x"5e",
          6669 => x"9f",
          6670 => x"97",
          6671 => x"8f",
          6672 => x"59",
          6673 => x"80",
          6674 => x"91",
          6675 => x"79",
          6676 => x"08",
          6677 => x"81",
          6678 => x"2e",
          6679 => x"70",
          6680 => x"5c",
          6681 => x"7a",
          6682 => x"2a",
          6683 => x"08",
          6684 => x"78",
          6685 => x"26",
          6686 => x"5b",
          6687 => x"d8",
          6688 => x"9c",
          6689 => x"55",
          6690 => x"dc",
          6691 => x"81",
          6692 => x"c5",
          6693 => x"bb",
          6694 => x"c2",
          6695 => x"b8",
          6696 => x"0b",
          6697 => x"04",
          6698 => x"3f",
          6699 => x"73",
          6700 => x"56",
          6701 => x"8e",
          6702 => x"2e",
          6703 => x"2e",
          6704 => x"7e",
          6705 => x"e4",
          6706 => x"a3",
          6707 => x"59",
          6708 => x"12",
          6709 => x"38",
          6710 => x"0c",
          6711 => x"7b",
          6712 => x"05",
          6713 => x"26",
          6714 => x"16",
          6715 => x"7c",
          6716 => x"39",
          6717 => x"80",
          6718 => x"c5",
          6719 => x"1b",
          6720 => x"08",
          6721 => x"3d",
          6722 => x"33",
          6723 => x"08",
          6724 => x"85",
          6725 => x"33",
          6726 => x"2e",
          6727 => x"ba",
          6728 => x"33",
          6729 => x"75",
          6730 => x"08",
          6731 => x"80",
          6732 => x"11",
          6733 => x"5b",
          6734 => x"a9",
          6735 => x"06",
          6736 => x"7b",
          6737 => x"06",
          6738 => x"9f",
          6739 => x"51",
          6740 => x"08",
          6741 => x"2e",
          6742 => x"26",
          6743 => x"55",
          6744 => x"88",
          6745 => x"38",
          6746 => x"38",
          6747 => x"e7",
          6748 => x"89",
          6749 => x"47",
          6750 => x"65",
          6751 => x"5f",
          6752 => x"80",
          6753 => x"53",
          6754 => x"3f",
          6755 => x"95",
          6756 => x"83",
          6757 => x"59",
          6758 => x"2e",
          6759 => x"90",
          6760 => x"44",
          6761 => x"83",
          6762 => x"33",
          6763 => x"81",
          6764 => x"75",
          6765 => x"11",
          6766 => x"71",
          6767 => x"72",
          6768 => x"5c",
          6769 => x"a3",
          6770 => x"4f",
          6771 => x"80",
          6772 => x"57",
          6773 => x"61",
          6774 => x"63",
          6775 => x"06",
          6776 => x"81",
          6777 => x"6e",
          6778 => x"62",
          6779 => x"38",
          6780 => x"e6",
          6781 => x"9d",
          6782 => x"e6",
          6783 => x"22",
          6784 => x"38",
          6785 => x"78",
          6786 => x"e4",
          6787 => x"e4",
          6788 => x"0b",
          6789 => x"e4",
          6790 => x"05",
          6791 => x"2a",
          6792 => x"7d",
          6793 => x"70",
          6794 => x"44",
          6795 => x"1d",
          6796 => x"31",
          6797 => x"38",
          6798 => x"70",
          6799 => x"3f",
          6800 => x"2e",
          6801 => x"81",
          6802 => x"0b",
          6803 => x"38",
          6804 => x"74",
          6805 => x"5b",
          6806 => x"b8",
          6807 => x"f0",
          6808 => x"93",
          6809 => x"0d",
          6810 => x"d0",
          6811 => x"57",
          6812 => x"77",
          6813 => x"77",
          6814 => x"83",
          6815 => x"57",
          6816 => x"76",
          6817 => x"12",
          6818 => x"38",
          6819 => x"44",
          6820 => x"89",
          6821 => x"59",
          6822 => x"47",
          6823 => x"38",
          6824 => x"70",
          6825 => x"07",
          6826 => x"ce",
          6827 => x"83",
          6828 => x"f9",
          6829 => x"81",
          6830 => x"81",
          6831 => x"38",
          6832 => x"e4",
          6833 => x"5f",
          6834 => x"fe",
          6835 => x"fb",
          6836 => x"83",
          6837 => x"3d",
          6838 => x"06",
          6839 => x"f5",
          6840 => x"43",
          6841 => x"9f",
          6842 => x"77",
          6843 => x"f5",
          6844 => x"0c",
          6845 => x"04",
          6846 => x"38",
          6847 => x"81",
          6848 => x"38",
          6849 => x"70",
          6850 => x"74",
          6851 => x"59",
          6852 => x"33",
          6853 => x"15",
          6854 => x"45",
          6855 => x"34",
          6856 => x"ff",
          6857 => x"34",
          6858 => x"05",
          6859 => x"83",
          6860 => x"91",
          6861 => x"49",
          6862 => x"75",
          6863 => x"75",
          6864 => x"93",
          6865 => x"61",
          6866 => x"34",
          6867 => x"99",
          6868 => x"80",
          6869 => x"05",
          6870 => x"9d",
          6871 => x"61",
          6872 => x"b8",
          6873 => x"9f",
          6874 => x"38",
          6875 => x"a8",
          6876 => x"80",
          6877 => x"ff",
          6878 => x"34",
          6879 => x"05",
          6880 => x"a9",
          6881 => x"05",
          6882 => x"70",
          6883 => x"05",
          6884 => x"38",
          6885 => x"69",
          6886 => x"aa",
          6887 => x"52",
          6888 => x"57",
          6889 => x"60",
          6890 => x"38",
          6891 => x"81",
          6892 => x"f4",
          6893 => x"2e",
          6894 => x"57",
          6895 => x"76",
          6896 => x"55",
          6897 => x"76",
          6898 => x"05",
          6899 => x"64",
          6900 => x"26",
          6901 => x"53",
          6902 => x"3f",
          6903 => x"84",
          6904 => x"81",
          6905 => x"f4",
          6906 => x"5b",
          6907 => x"7f",
          6908 => x"62",
          6909 => x"55",
          6910 => x"74",
          6911 => x"fe",
          6912 => x"85",
          6913 => x"57",
          6914 => x"83",
          6915 => x"ff",
          6916 => x"82",
          6917 => x"c1",
          6918 => x"7d",
          6919 => x"59",
          6920 => x"ff",
          6921 => x"69",
          6922 => x"be",
          6923 => x"81",
          6924 => x"78",
          6925 => x"05",
          6926 => x"62",
          6927 => x"67",
          6928 => x"82",
          6929 => x"05",
          6930 => x"05",
          6931 => x"67",
          6932 => x"83",
          6933 => x"61",
          6934 => x"ca",
          6935 => x"61",
          6936 => x"58",
          6937 => x"98",
          6938 => x"34",
          6939 => x"51",
          6940 => x"b8",
          6941 => x"80",
          6942 => x"81",
          6943 => x"38",
          6944 => x"0c",
          6945 => x"04",
          6946 => x"64",
          6947 => x"ae",
          6948 => x"83",
          6949 => x"2e",
          6950 => x"83",
          6951 => x"70",
          6952 => x"86",
          6953 => x"52",
          6954 => x"b8",
          6955 => x"70",
          6956 => x"0b",
          6957 => x"05",
          6958 => x"27",
          6959 => x"39",
          6960 => x"26",
          6961 => x"77",
          6962 => x"8e",
          6963 => x"44",
          6964 => x"43",
          6965 => x"34",
          6966 => x"05",
          6967 => x"a2",
          6968 => x"61",
          6969 => x"61",
          6970 => x"c4",
          6971 => x"34",
          6972 => x"7c",
          6973 => x"5c",
          6974 => x"2a",
          6975 => x"98",
          6976 => x"82",
          6977 => x"05",
          6978 => x"61",
          6979 => x"34",
          6980 => x"b2",
          6981 => x"ff",
          6982 => x"61",
          6983 => x"c7",
          6984 => x"76",
          6985 => x"81",
          6986 => x"80",
          6987 => x"05",
          6988 => x"34",
          6989 => x"b8",
          6990 => x"79",
          6991 => x"84",
          6992 => x"90",
          6993 => x"b2",
          6994 => x"08",
          6995 => x"b4",
          6996 => x"b8",
          6997 => x"f0",
          6998 => x"ff",
          6999 => x"6a",
          7000 => x"34",
          7001 => x"85",
          7002 => x"ff",
          7003 => x"05",
          7004 => x"61",
          7005 => x"57",
          7006 => x"53",
          7007 => x"3f",
          7008 => x"70",
          7009 => x"76",
          7010 => x"70",
          7011 => x"d2",
          7012 => x"e1",
          7013 => x"c1",
          7014 => x"05",
          7015 => x"34",
          7016 => x"80",
          7017 => x"ff",
          7018 => x"34",
          7019 => x"e9",
          7020 => x"61",
          7021 => x"40",
          7022 => x"61",
          7023 => x"ed",
          7024 => x"34",
          7025 => x"d5",
          7026 => x"54",
          7027 => x"fe",
          7028 => x"53",
          7029 => x"3f",
          7030 => x"f4",
          7031 => x"7b",
          7032 => x"78",
          7033 => x"3d",
          7034 => x"79",
          7035 => x"2e",
          7036 => x"33",
          7037 => x"76",
          7038 => x"57",
          7039 => x"24",
          7040 => x"76",
          7041 => x"e4",
          7042 => x"0d",
          7043 => x"59",
          7044 => x"84",
          7045 => x"38",
          7046 => x"56",
          7047 => x"74",
          7048 => x"0c",
          7049 => x"0d",
          7050 => x"53",
          7051 => x"9e",
          7052 => x"70",
          7053 => x"1b",
          7054 => x"56",
          7055 => x"ff",
          7056 => x"0d",
          7057 => x"58",
          7058 => x"76",
          7059 => x"55",
          7060 => x"0c",
          7061 => x"56",
          7062 => x"77",
          7063 => x"34",
          7064 => x"38",
          7065 => x"18",
          7066 => x"38",
          7067 => x"54",
          7068 => x"9d",
          7069 => x"38",
          7070 => x"84",
          7071 => x"9f",
          7072 => x"c0",
          7073 => x"a2",
          7074 => x"72",
          7075 => x"56",
          7076 => x"51",
          7077 => x"84",
          7078 => x"fd",
          7079 => x"05",
          7080 => x"ff",
          7081 => x"06",
          7082 => x"3d",
          7083 => x"54",
          7084 => x"e9",
          7085 => x"e6",
          7086 => x"38",
          7087 => x"53",
          7088 => x"71",
          7089 => x"51",
          7090 => x"81",
          7091 => x"85",
          7092 => x"92",
          7093 => x"22",
          7094 => x"26",
          7095 => x"e4",
          7096 => x"b5",
          7097 => x"81",
          7098 => x"e4",
          7099 => x"0c",
          7100 => x"0d",
          7101 => x"80",
          7102 => x"83",
          7103 => x"26",
          7104 => x"56",
          7105 => x"73",
          7106 => x"70",
          7107 => x"22",
          7108 => x"ff",
          7109 => x"24",
          7110 => x"15",
          7111 => x"73",
          7112 => x"07",
          7113 => x"38",
          7114 => x"87",
          7115 => x"ff",
          7116 => x"71",
          7117 => x"73",
          7118 => x"ff",
          7119 => x"39",
          7120 => x"06",
          7121 => x"83",
          7122 => x"e6",
          7123 => x"51",
          7124 => x"ff",
          7125 => x"70",
          7126 => x"39",
          7127 => x"57",
          7128 => x"81",
          7129 => x"ff",
          7130 => x"75",
          7131 => x"52",
          7132 => x"00",
          7133 => x"ff",
          7134 => x"00",
          7135 => x"00",
          7136 => x"00",
          7137 => x"00",
          7138 => x"00",
          7139 => x"00",
          7140 => x"00",
          7141 => x"00",
          7142 => x"00",
          7143 => x"00",
          7144 => x"00",
          7145 => x"00",
          7146 => x"00",
          7147 => x"00",
          7148 => x"00",
          7149 => x"00",
          7150 => x"00",
          7151 => x"00",
          7152 => x"00",
          7153 => x"00",
          7154 => x"00",
          7155 => x"00",
          7156 => x"00",
          7157 => x"00",
          7158 => x"00",
          7159 => x"00",
          7160 => x"00",
          7161 => x"00",
          7162 => x"00",
          7163 => x"00",
          7164 => x"00",
          7165 => x"00",
          7166 => x"00",
          7167 => x"00",
          7168 => x"00",
          7169 => x"00",
          7170 => x"00",
          7171 => x"00",
          7172 => x"00",
          7173 => x"00",
          7174 => x"00",
          7175 => x"00",
          7176 => x"00",
          7177 => x"00",
          7178 => x"00",
          7179 => x"00",
          7180 => x"00",
          7181 => x"00",
          7182 => x"00",
          7183 => x"00",
          7184 => x"00",
          7185 => x"00",
          7186 => x"00",
          7187 => x"00",
          7188 => x"00",
          7189 => x"00",
          7190 => x"00",
          7191 => x"00",
          7192 => x"00",
          7193 => x"00",
          7194 => x"00",
          7195 => x"00",
          7196 => x"00",
          7197 => x"00",
          7198 => x"00",
          7199 => x"00",
          7200 => x"00",
          7201 => x"00",
          7202 => x"00",
          7203 => x"00",
          7204 => x"00",
          7205 => x"00",
          7206 => x"00",
          7207 => x"00",
          7208 => x"00",
          7209 => x"00",
          7210 => x"00",
          7211 => x"00",
          7212 => x"00",
          7213 => x"00",
          7214 => x"00",
          7215 => x"00",
          7216 => x"00",
          7217 => x"00",
          7218 => x"00",
          7219 => x"00",
          7220 => x"00",
          7221 => x"00",
          7222 => x"00",
          7223 => x"00",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"00",
          7230 => x"00",
          7231 => x"00",
          7232 => x"00",
          7233 => x"00",
          7234 => x"00",
          7235 => x"00",
          7236 => x"00",
          7237 => x"00",
          7238 => x"00",
          7239 => x"00",
          7240 => x"00",
          7241 => x"00",
          7242 => x"00",
          7243 => x"00",
          7244 => x"00",
          7245 => x"00",
          7246 => x"00",
          7247 => x"00",
          7248 => x"00",
          7249 => x"00",
          7250 => x"00",
          7251 => x"00",
          7252 => x"00",
          7253 => x"00",
          7254 => x"00",
          7255 => x"00",
          7256 => x"00",
          7257 => x"00",
          7258 => x"00",
          7259 => x"00",
          7260 => x"00",
          7261 => x"00",
          7262 => x"00",
          7263 => x"00",
          7264 => x"00",
          7265 => x"00",
          7266 => x"00",
          7267 => x"00",
          7268 => x"00",
          7269 => x"00",
          7270 => x"00",
          7271 => x"00",
          7272 => x"00",
          7273 => x"00",
          7274 => x"00",
          7275 => x"00",
          7276 => x"00",
          7277 => x"00",
          7278 => x"00",
          7279 => x"00",
          7280 => x"00",
          7281 => x"00",
          7282 => x"00",
          7283 => x"00",
          7284 => x"00",
          7285 => x"00",
          7286 => x"00",
          7287 => x"00",
          7288 => x"00",
          7289 => x"00",
          7290 => x"00",
          7291 => x"00",
          7292 => x"00",
          7293 => x"00",
          7294 => x"00",
          7295 => x"00",
          7296 => x"00",
          7297 => x"00",
          7298 => x"00",
          7299 => x"00",
          7300 => x"00",
          7301 => x"00",
          7302 => x"00",
          7303 => x"00",
          7304 => x"00",
          7305 => x"00",
          7306 => x"00",
          7307 => x"00",
          7308 => x"00",
          7309 => x"00",
          7310 => x"00",
          7311 => x"00",
          7312 => x"00",
          7313 => x"00",
          7314 => x"00",
          7315 => x"00",
          7316 => x"00",
          7317 => x"00",
          7318 => x"00",
          7319 => x"00",
          7320 => x"00",
          7321 => x"00",
          7322 => x"00",
          7323 => x"00",
          7324 => x"00",
          7325 => x"00",
          7326 => x"00",
          7327 => x"00",
          7328 => x"00",
          7329 => x"00",
          7330 => x"00",
          7331 => x"00",
          7332 => x"00",
          7333 => x"00",
          7334 => x"00",
          7335 => x"00",
          7336 => x"00",
          7337 => x"00",
          7338 => x"00",
          7339 => x"00",
          7340 => x"00",
          7341 => x"00",
          7342 => x"00",
          7343 => x"00",
          7344 => x"00",
          7345 => x"00",
          7346 => x"00",
          7347 => x"00",
          7348 => x"00",
          7349 => x"00",
          7350 => x"00",
          7351 => x"00",
          7352 => x"00",
          7353 => x"00",
          7354 => x"00",
          7355 => x"00",
          7356 => x"00",
          7357 => x"00",
          7358 => x"00",
          7359 => x"00",
          7360 => x"00",
          7361 => x"00",
          7362 => x"00",
          7363 => x"00",
          7364 => x"00",
          7365 => x"00",
          7366 => x"00",
          7367 => x"00",
          7368 => x"00",
          7369 => x"00",
          7370 => x"00",
          7371 => x"74",
          7372 => x"74",
          7373 => x"74",
          7374 => x"64",
          7375 => x"63",
          7376 => x"61",
          7377 => x"79",
          7378 => x"66",
          7379 => x"70",
          7380 => x"6d",
          7381 => x"68",
          7382 => x"68",
          7383 => x"63",
          7384 => x"6a",
          7385 => x"61",
          7386 => x"74",
          7387 => x"00",
          7388 => x"00",
          7389 => x"7a",
          7390 => x"69",
          7391 => x"69",
          7392 => x"00",
          7393 => x"55",
          7394 => x"65",
          7395 => x"50",
          7396 => x"72",
          7397 => x"72",
          7398 => x"54",
          7399 => x"20",
          7400 => x"6c",
          7401 => x"49",
          7402 => x"69",
          7403 => x"6f",
          7404 => x"46",
          7405 => x"6c",
          7406 => x"54",
          7407 => x"20",
          7408 => x"6f",
          7409 => x"6c",
          7410 => x"46",
          7411 => x"62",
          7412 => x"4e",
          7413 => x"74",
          7414 => x"6c",
          7415 => x"20",
          7416 => x"6e",
          7417 => x"44",
          7418 => x"20",
          7419 => x"2e",
          7420 => x"65",
          7421 => x"20",
          7422 => x"6c",
          7423 => x"53",
          7424 => x"69",
          7425 => x"65",
          7426 => x"46",
          7427 => x"64",
          7428 => x"6c",
          7429 => x"46",
          7430 => x"65",
          7431 => x"73",
          7432 => x"41",
          7433 => x"65",
          7434 => x"49",
          7435 => x"66",
          7436 => x"2e",
          7437 => x"61",
          7438 => x"64",
          7439 => x"69",
          7440 => x"64",
          7441 => x"20",
          7442 => x"64",
          7443 => x"72",
          7444 => x"6f",
          7445 => x"20",
          7446 => x"53",
          7447 => x"00",
          7448 => x"20",
          7449 => x"73",
          7450 => x"20",
          7451 => x"65",
          7452 => x"72",
          7453 => x"25",
          7454 => x"3a",
          7455 => x"00",
          7456 => x"7c",
          7457 => x"25",
          7458 => x"20",
          7459 => x"00",
          7460 => x"2a",
          7461 => x"30",
          7462 => x"32",
          7463 => x"66",
          7464 => x"2c",
          7465 => x"32",
          7466 => x"73",
          7467 => x"5a",
          7468 => x"72",
          7469 => x"6e",
          7470 => x"55",
          7471 => x"20",
          7472 => x"70",
          7473 => x"31",
          7474 => x"65",
          7475 => x"55",
          7476 => x"20",
          7477 => x"70",
          7478 => x"30",
          7479 => x"65",
          7480 => x"49",
          7481 => x"20",
          7482 => x"70",
          7483 => x"4c",
          7484 => x"65",
          7485 => x"50",
          7486 => x"72",
          7487 => x"54",
          7488 => x"74",
          7489 => x"53",
          7490 => x"75",
          7491 => x"2e",
          7492 => x"6c",
          7493 => x"65",
          7494 => x"61",
          7495 => x"2e",
          7496 => x"7a",
          7497 => x"68",
          7498 => x"65",
          7499 => x"69",
          7500 => x"20",
          7501 => x"20",
          7502 => x"73",
          7503 => x"6d",
          7504 => x"2e",
          7505 => x"25",
          7506 => x"30",
          7507 => x"63",
          7508 => x"00",
          7509 => x"62",
          7510 => x"25",
          7511 => x"00",
          7512 => x"20",
          7513 => x"6e",
          7514 => x"52",
          7515 => x"6e",
          7516 => x"63",
          7517 => x"2e",
          7518 => x"69",
          7519 => x"20",
          7520 => x"20",
          7521 => x"43",
          7522 => x"75",
          7523 => x"64",
          7524 => x"0a",
          7525 => x"75",
          7526 => x"64",
          7527 => x"6c",
          7528 => x"25",
          7529 => x"38",
          7530 => x"25",
          7531 => x"34",
          7532 => x"61",
          7533 => x"00",
          7534 => x"78",
          7535 => x"3e",
          7536 => x"30",
          7537 => x"43",
          7538 => x"2e",
          7539 => x"58",
          7540 => x"43",
          7541 => x"2e",
          7542 => x"44",
          7543 => x"6f",
          7544 => x"70",
          7545 => x"25",
          7546 => x"73",
          7547 => x"72",
          7548 => x"73",
          7549 => x"6e",
          7550 => x"63",
          7551 => x"6d",
          7552 => x"3f",
          7553 => x"64",
          7554 => x"25",
          7555 => x"25",
          7556 => x"43",
          7557 => x"61",
          7558 => x"3a",
          7559 => x"73",
          7560 => x"65",
          7561 => x"41",
          7562 => x"73",
          7563 => x"43",
          7564 => x"74",
          7565 => x"20",
          7566 => x"20",
          7567 => x"00",
          7568 => x"43",
          7569 => x"72",
          7570 => x"20",
          7571 => x"20",
          7572 => x"00",
          7573 => x"53",
          7574 => x"61",
          7575 => x"65",
          7576 => x"20",
          7577 => x"00",
          7578 => x"3a",
          7579 => x"5a",
          7580 => x"20",
          7581 => x"20",
          7582 => x"20",
          7583 => x"00",
          7584 => x"53",
          7585 => x"6c",
          7586 => x"71",
          7587 => x"20",
          7588 => x"34",
          7589 => x"20",
          7590 => x"62",
          7591 => x"41",
          7592 => x"20",
          7593 => x"64",
          7594 => x"7a",
          7595 => x"53",
          7596 => x"6f",
          7597 => x"20",
          7598 => x"20",
          7599 => x"34",
          7600 => x"20",
          7601 => x"20",
          7602 => x"20",
          7603 => x"4c",
          7604 => x"57",
          7605 => x"20",
          7606 => x"42",
          7607 => x"00",
          7608 => x"49",
          7609 => x"4c",
          7610 => x"65",
          7611 => x"29",
          7612 => x"54",
          7613 => x"20",
          7614 => x"73",
          7615 => x"29",
          7616 => x"53",
          7617 => x"20",
          7618 => x"65",
          7619 => x"29",
          7620 => x"52",
          7621 => x"20",
          7622 => x"25",
          7623 => x"20",
          7624 => x"20",
          7625 => x"30",
          7626 => x"29",
          7627 => x"49",
          7628 => x"4d",
          7629 => x"25",
          7630 => x"20",
          7631 => x"4d",
          7632 => x"30",
          7633 => x"29",
          7634 => x"57",
          7635 => x"20",
          7636 => x"25",
          7637 => x"20",
          7638 => x"6f",
          7639 => x"67",
          7640 => x"6f",
          7641 => x"00",
          7642 => x"6c",
          7643 => x"75",
          7644 => x"00",
          7645 => x"00",
          7646 => x"00",
          7647 => x"01",
          7648 => x"00",
          7649 => x"00",
          7650 => x"01",
          7651 => x"00",
          7652 => x"00",
          7653 => x"01",
          7654 => x"00",
          7655 => x"00",
          7656 => x"01",
          7657 => x"00",
          7658 => x"00",
          7659 => x"01",
          7660 => x"00",
          7661 => x"00",
          7662 => x"04",
          7663 => x"00",
          7664 => x"00",
          7665 => x"04",
          7666 => x"00",
          7667 => x"00",
          7668 => x"04",
          7669 => x"00",
          7670 => x"00",
          7671 => x"04",
          7672 => x"00",
          7673 => x"00",
          7674 => x"03",
          7675 => x"00",
          7676 => x"00",
          7677 => x"03",
          7678 => x"1b",
          7679 => x"1b",
          7680 => x"1b",
          7681 => x"1b",
          7682 => x"1b",
          7683 => x"1b",
          7684 => x"0e",
          7685 => x"0b",
          7686 => x"06",
          7687 => x"04",
          7688 => x"02",
          7689 => x"43",
          7690 => x"70",
          7691 => x"74",
          7692 => x"72",
          7693 => x"20",
          7694 => x"6e",
          7695 => x"6f",
          7696 => x"00",
          7697 => x"25",
          7698 => x"73",
          7699 => x"65",
          7700 => x"73",
          7701 => x"68",
          7702 => x"66",
          7703 => x"45",
          7704 => x"3e",
          7705 => x"1b",
          7706 => x"1b",
          7707 => x"1b",
          7708 => x"1b",
          7709 => x"1b",
          7710 => x"1b",
          7711 => x"1b",
          7712 => x"1b",
          7713 => x"1b",
          7714 => x"1b",
          7715 => x"1b",
          7716 => x"1b",
          7717 => x"1b",
          7718 => x"1b",
          7719 => x"1b",
          7720 => x"1b",
          7721 => x"00",
          7722 => x"00",
          7723 => x"2c",
          7724 => x"64",
          7725 => x"25",
          7726 => x"44",
          7727 => x"25",
          7728 => x"2c",
          7729 => x"25",
          7730 => x"3a",
          7731 => x"2c",
          7732 => x"64",
          7733 => x"52",
          7734 => x"75",
          7735 => x"55",
          7736 => x"25",
          7737 => x"44",
          7738 => x"25",
          7739 => x"48",
          7740 => x"00",
          7741 => x"65",
          7742 => x"6e",
          7743 => x"53",
          7744 => x"3e",
          7745 => x"2b",
          7746 => x"46",
          7747 => x"32",
          7748 => x"53",
          7749 => x"4e",
          7750 => x"20",
          7751 => x"20",
          7752 => x"41",
          7753 => x"41",
          7754 => x"00",
          7755 => x"00",
          7756 => x"01",
          7757 => x"14",
          7758 => x"80",
          7759 => x"45",
          7760 => x"90",
          7761 => x"59",
          7762 => x"41",
          7763 => x"a8",
          7764 => x"b0",
          7765 => x"b8",
          7766 => x"c0",
          7767 => x"c8",
          7768 => x"d0",
          7769 => x"d8",
          7770 => x"e0",
          7771 => x"e8",
          7772 => x"f0",
          7773 => x"f8",
          7774 => x"2b",
          7775 => x"5c",
          7776 => x"7f",
          7777 => x"00",
          7778 => x"00",
          7779 => x"00",
          7780 => x"00",
          7781 => x"00",
          7782 => x"00",
          7783 => x"00",
          7784 => x"00",
          7785 => x"00",
          7786 => x"00",
          7787 => x"00",
          7788 => x"20",
          7789 => x"00",
          7790 => x"00",
          7791 => x"00",
          7792 => x"00",
          7793 => x"25",
          7794 => x"25",
          7795 => x"25",
          7796 => x"25",
          7797 => x"25",
          7798 => x"25",
          7799 => x"25",
          7800 => x"25",
          7801 => x"25",
          7802 => x"25",
          7803 => x"25",
          7804 => x"25",
          7805 => x"03",
          7806 => x"00",
          7807 => x"03",
          7808 => x"03",
          7809 => x"22",
          7810 => x"00",
          7811 => x"00",
          7812 => x"25",
          7813 => x"00",
          7814 => x"00",
          7815 => x"01",
          7816 => x"01",
          7817 => x"01",
          7818 => x"01",
          7819 => x"01",
          7820 => x"01",
          7821 => x"01",
          7822 => x"01",
          7823 => x"01",
          7824 => x"01",
          7825 => x"01",
          7826 => x"01",
          7827 => x"01",
          7828 => x"01",
          7829 => x"01",
          7830 => x"01",
          7831 => x"01",
          7832 => x"01",
          7833 => x"01",
          7834 => x"01",
          7835 => x"01",
          7836 => x"01",
          7837 => x"01",
          7838 => x"01",
          7839 => x"00",
          7840 => x"01",
          7841 => x"02",
          7842 => x"02",
          7843 => x"02",
          7844 => x"01",
          7845 => x"01",
          7846 => x"02",
          7847 => x"02",
          7848 => x"01",
          7849 => x"02",
          7850 => x"01",
          7851 => x"02",
          7852 => x"02",
          7853 => x"02",
          7854 => x"02",
          7855 => x"02",
          7856 => x"01",
          7857 => x"02",
          7858 => x"01",
          7859 => x"02",
          7860 => x"02",
          7861 => x"00",
          7862 => x"03",
          7863 => x"03",
          7864 => x"03",
          7865 => x"03",
          7866 => x"03",
          7867 => x"01",
          7868 => x"03",
          7869 => x"03",
          7870 => x"03",
          7871 => x"07",
          7872 => x"01",
          7873 => x"00",
          7874 => x"05",
          7875 => x"1d",
          7876 => x"01",
          7877 => x"06",
          7878 => x"06",
          7879 => x"06",
          7880 => x"1f",
          7881 => x"1f",
          7882 => x"1f",
          7883 => x"1f",
          7884 => x"1f",
          7885 => x"1f",
          7886 => x"1f",
          7887 => x"1f",
          7888 => x"1f",
          7889 => x"1f",
          7890 => x"06",
          7891 => x"00",
          7892 => x"1f",
          7893 => x"21",
          7894 => x"21",
          7895 => x"04",
          7896 => x"01",
          7897 => x"01",
          7898 => x"03",
          7899 => x"00",
          7900 => x"00",
          7901 => x"00",
          7902 => x"00",
          7903 => x"00",
          7904 => x"00",
          7905 => x"00",
          7906 => x"00",
          7907 => x"00",
          7908 => x"00",
          7909 => x"00",
          7910 => x"00",
          7911 => x"00",
          7912 => x"00",
          7913 => x"00",
          7914 => x"00",
          7915 => x"00",
          7916 => x"00",
          7917 => x"00",
          7918 => x"00",
          7919 => x"00",
          7920 => x"00",
          7921 => x"00",
          7922 => x"00",
          7923 => x"00",
          7924 => x"00",
          7925 => x"00",
          7926 => x"00",
          7927 => x"00",
          7928 => x"00",
          7929 => x"00",
          7930 => x"00",
          7931 => x"00",
          7932 => x"00",
          7933 => x"00",
          7934 => x"00",
          7935 => x"00",
          7936 => x"00",
          7937 => x"00",
          7938 => x"00",
          7939 => x"00",
          7940 => x"00",
          7941 => x"00",
          7942 => x"00",
          7943 => x"00",
          7944 => x"00",
          7945 => x"00",
          7946 => x"00",
          7947 => x"00",
          7948 => x"00",
          7949 => x"00",
          7950 => x"00",
          7951 => x"00",
          7952 => x"00",
          7953 => x"00",
          7954 => x"00",
          7955 => x"00",
          7956 => x"00",
          7957 => x"00",
          7958 => x"00",
          7959 => x"00",
          7960 => x"01",
          7961 => x"00",
          7962 => x"00",
          7963 => x"05",
          7964 => x"00",
          7965 => x"01",
          7966 => x"01",
          7967 => x"00",
          7968 => x"00",
          7969 => x"00",
          7970 => x"00",
          7971 => x"00",
          7972 => x"00",
          7973 => x"00",
          7974 => x"00",
          7975 => x"00",
          7976 => x"00",
          7977 => x"00",
          7978 => x"00",
          7979 => x"01",
          7980 => x"01",
          7981 => x"02",
          7982 => x"1b",
          7983 => x"79",
          7984 => x"71",
          7985 => x"69",
          7986 => x"61",
          7987 => x"31",
          7988 => x"5c",
          7989 => x"f6",
          7990 => x"08",
          7991 => x"80",
          7992 => x"1b",
          7993 => x"59",
          7994 => x"51",
          7995 => x"49",
          7996 => x"41",
          7997 => x"31",
          7998 => x"5c",
          7999 => x"f6",
          8000 => x"08",
          8001 => x"80",
          8002 => x"1b",
          8003 => x"59",
          8004 => x"51",
          8005 => x"49",
          8006 => x"41",
          8007 => x"21",
          8008 => x"7c",
          8009 => x"f7",
          8010 => x"fb",
          8011 => x"85",
          8012 => x"1b",
          8013 => x"19",
          8014 => x"11",
          8015 => x"09",
          8016 => x"01",
          8017 => x"f0",
          8018 => x"f0",
          8019 => x"f0",
          8020 => x"f0",
          8021 => x"80",
          8022 => x"bf",
          8023 => x"35",
          8024 => x"7c",
          8025 => x"3d",
          8026 => x"46",
          8027 => x"3f",
          8028 => x"d3",
          8029 => x"c6",
          8030 => x"f0",
          8031 => x"80",
          8032 => x"00",
          8033 => x"00",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"00",
          8045 => x"00",
          8046 => x"00",
          8047 => x"00",
          8048 => x"00",
          8049 => x"00",
          8050 => x"00",
          8051 => x"00",
          8052 => x"00",
          8053 => x"00",
          8054 => x"00",
          8055 => x"00",
          8056 => x"00",
          8057 => x"00",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"00",
          8063 => x"00",
          8064 => x"00",
          8065 => x"00",
          8066 => x"00",
          8067 => x"00",
          8068 => x"00",
          8069 => x"00",
          8070 => x"00",
          8071 => x"00",
          8072 => x"00",
          8073 => x"00",
          8074 => x"00",
          8075 => x"00",
          8076 => x"00",
          8077 => x"00",
          8078 => x"00",
          8079 => x"00",
          8080 => x"00",
          8081 => x"00",
          8082 => x"00",
          8083 => x"00",
          8084 => x"00",
          8085 => x"00",
          8086 => x"00",
          8087 => x"00",
          8088 => x"00",
          8089 => x"00",
          8090 => x"00",
          8091 => x"00",
          8092 => x"00",
          8093 => x"00",
          8094 => x"00",
          8095 => x"00",
          8096 => x"00",
          8097 => x"00",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"00",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"00",
          8108 => x"00",
          8109 => x"00",
          8110 => x"00",
          8111 => x"00",
          8112 => x"00",
          8113 => x"00",
          8114 => x"00",
          8115 => x"00",
          8116 => x"00",
          8117 => x"00",
          8118 => x"00",
          8119 => x"00",
          8120 => x"00",
          8121 => x"00",
          8122 => x"00",
          8123 => x"00",
          8124 => x"00",
          8125 => x"00",
          8126 => x"00",
          8127 => x"00",
          8128 => x"00",
          8129 => x"00",
          8130 => x"00",
          8131 => x"00",
          8132 => x"00",
          8133 => x"00",
          8134 => x"00",
          8135 => x"00",
          8136 => x"00",
          8137 => x"00",
          8138 => x"00",
          8139 => x"00",
          8140 => x"00",
          8141 => x"00",
          8142 => x"00",
          8143 => x"00",
          8144 => x"00",
          8145 => x"00",
          8146 => x"00",
          8147 => x"00",
          8148 => x"00",
          8149 => x"00",
          8150 => x"00",
          8151 => x"00",
          8152 => x"00",
          8153 => x"00",
          8154 => x"00",
          8155 => x"00",
          8156 => x"00",
          8157 => x"00",
          8158 => x"00",
          8159 => x"00",
          8160 => x"00",
          8161 => x"00",
          8162 => x"00",
          8163 => x"00",
          8164 => x"00",
          8165 => x"00",
          8166 => x"00",
          8167 => x"00",
          8168 => x"00",
          8169 => x"00",
          8170 => x"00",
          8171 => x"00",
          8172 => x"00",
          8173 => x"00",
          8174 => x"00",
          8175 => x"00",
          8176 => x"00",
          8177 => x"00",
          8178 => x"00",
          8179 => x"00",
          8180 => x"00",
          8181 => x"00",
          8182 => x"00",
          8183 => x"00",
          8184 => x"00",
          8185 => x"00",
          8186 => x"00",
          8187 => x"00",
          8188 => x"00",
          8189 => x"00",
          8190 => x"00",
          8191 => x"00",
          8192 => x"00",
          8193 => x"00",
          8194 => x"00",
          8195 => x"00",
          8196 => x"00",
          8197 => x"00",
          8198 => x"00",
          8199 => x"00",
          8200 => x"00",
          8201 => x"00",
          8202 => x"00",
          8203 => x"00",
          8204 => x"00",
          8205 => x"00",
          8206 => x"00",
          8207 => x"00",
          8208 => x"00",
          8209 => x"00",
          8210 => x"00",
          8211 => x"00",
          8212 => x"00",
          8213 => x"00",
          8214 => x"00",
          8215 => x"00",
          8216 => x"00",
          8217 => x"00",
          8218 => x"00",
          8219 => x"00",
          8220 => x"00",
          8221 => x"00",
          8222 => x"00",
          8223 => x"00",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"00",
          8235 => x"00",
          8236 => x"00",
          8237 => x"00",
          8238 => x"00",
          8239 => x"00",
          8240 => x"00",
          8241 => x"00",
          8242 => x"00",
          8243 => x"00",
          8244 => x"00",
          8245 => x"00",
          8246 => x"00",
          8247 => x"00",
          8248 => x"00",
          8249 => x"00",
          8250 => x"00",
          8251 => x"00",
          8252 => x"00",
          8253 => x"00",
          8254 => x"00",
          8255 => x"00",
          8256 => x"00",
          8257 => x"00",
          8258 => x"00",
          8259 => x"00",
          8260 => x"00",
          8261 => x"00",
          8262 => x"00",
          8263 => x"00",
          8264 => x"00",
          8265 => x"00",
          8266 => x"00",
          8267 => x"00",
          8268 => x"00",
          8269 => x"00",
          8270 => x"00",
          8271 => x"00",
          8272 => x"00",
          8273 => x"00",
          8274 => x"00",
          8275 => x"00",
          8276 => x"00",
          8277 => x"00",
          8278 => x"00",
          8279 => x"00",
          8280 => x"00",
          8281 => x"00",
          8282 => x"00",
          8283 => x"00",
          8284 => x"00",
          8285 => x"00",
          8286 => x"00",
          8287 => x"00",
          8288 => x"00",
          8289 => x"00",
          8290 => x"00",
          8291 => x"00",
          8292 => x"00",
          8293 => x"00",
          8294 => x"00",
          8295 => x"00",
          8296 => x"00",
          8297 => x"00",
          8298 => x"00",
          8299 => x"00",
          8300 => x"00",
          8301 => x"00",
          8302 => x"00",
          8303 => x"00",
          8304 => x"00",
          8305 => x"00",
          8306 => x"00",
          8307 => x"00",
          8308 => x"00",
          8309 => x"00",
          8310 => x"00",
          8311 => x"00",
          8312 => x"00",
          8313 => x"00",
          8314 => x"00",
          8315 => x"00",
          8316 => x"00",
          8317 => x"00",
          8318 => x"00",
          8319 => x"00",
          8320 => x"00",
          8321 => x"00",
          8322 => x"00",
          8323 => x"00",
          8324 => x"00",
          8325 => x"00",
          8326 => x"00",
          8327 => x"00",
          8328 => x"00",
          8329 => x"00",
          8330 => x"00",
          8331 => x"00",
          8332 => x"00",
          8333 => x"00",
          8334 => x"00",
          8335 => x"00",
          8336 => x"00",
          8337 => x"00",
          8338 => x"00",
          8339 => x"00",
          8340 => x"00",
          8341 => x"00",
          8342 => x"00",
          8343 => x"00",
          8344 => x"00",
          8345 => x"00",
          8346 => x"00",
          8347 => x"00",
          8348 => x"00",
          8349 => x"00",
          8350 => x"00",
          8351 => x"00",
          8352 => x"00",
          8353 => x"00",
          8354 => x"00",
          8355 => x"00",
          8356 => x"00",
          8357 => x"00",
          8358 => x"00",
          8359 => x"00",
          8360 => x"00",
          8361 => x"00",
          8362 => x"00",
          8363 => x"00",
          8364 => x"00",
          8365 => x"00",
          8366 => x"00",
          8367 => x"00",
          8368 => x"00",
          8369 => x"00",
          8370 => x"00",
          8371 => x"00",
          8372 => x"00",
          8373 => x"00",
          8374 => x"00",
          8375 => x"00",
          8376 => x"00",
          8377 => x"00",
          8378 => x"00",
          8379 => x"00",
          8380 => x"00",
          8381 => x"00",
          8382 => x"00",
          8383 => x"00",
          8384 => x"00",
          8385 => x"00",
          8386 => x"00",
          8387 => x"00",
          8388 => x"00",
          8389 => x"00",
          8390 => x"00",
          8391 => x"00",
          8392 => x"00",
          8393 => x"00",
          8394 => x"00",
          8395 => x"00",
          8396 => x"00",
          8397 => x"00",
          8398 => x"00",
          8399 => x"00",
          8400 => x"00",
          8401 => x"00",
          8402 => x"00",
          8403 => x"00",
          8404 => x"00",
          8405 => x"00",
          8406 => x"00",
          8407 => x"00",
          8408 => x"00",
          8409 => x"00",
          8410 => x"00",
          8411 => x"00",
          8412 => x"00",
          8413 => x"00",
          8414 => x"00",
          8415 => x"00",
          8416 => x"00",
          8417 => x"00",
          8418 => x"00",
          8419 => x"00",
          8420 => x"00",
          8421 => x"00",
          8422 => x"00",
          8423 => x"00",
          8424 => x"00",
          8425 => x"00",
          8426 => x"00",
          8427 => x"00",
          8428 => x"00",
          8429 => x"00",
          8430 => x"00",
          8431 => x"00",
          8432 => x"00",
          8433 => x"00",
          8434 => x"00",
          8435 => x"00",
          8436 => x"00",
          8437 => x"00",
          8438 => x"00",
          8439 => x"00",
          8440 => x"00",
          8441 => x"00",
          8442 => x"00",
          8443 => x"00",
          8444 => x"00",
          8445 => x"00",
          8446 => x"00",
          8447 => x"00",
          8448 => x"00",
          8449 => x"00",
          8450 => x"00",
          8451 => x"00",
          8452 => x"00",
          8453 => x"00",
          8454 => x"00",
          8455 => x"00",
          8456 => x"00",
          8457 => x"00",
          8458 => x"00",
          8459 => x"00",
          8460 => x"00",
          8461 => x"00",
          8462 => x"00",
          8463 => x"00",
          8464 => x"00",
          8465 => x"00",
          8466 => x"00",
          8467 => x"00",
          8468 => x"00",
          8469 => x"00",
          8470 => x"00",
          8471 => x"00",
          8472 => x"00",
          8473 => x"00",
          8474 => x"00",
          8475 => x"00",
          8476 => x"00",
          8477 => x"00",
          8478 => x"00",
          8479 => x"00",
          8480 => x"00",
          8481 => x"00",
          8482 => x"00",
          8483 => x"00",
          8484 => x"00",
          8485 => x"00",
          8486 => x"00",
          8487 => x"00",
          8488 => x"00",
          8489 => x"00",
          8490 => x"00",
          8491 => x"00",
          8492 => x"00",
          8493 => x"00",
          8494 => x"00",
          8495 => x"00",
          8496 => x"00",
          8497 => x"00",
          8498 => x"00",
          8499 => x"00",
          8500 => x"00",
          8501 => x"00",
          8502 => x"00",
          8503 => x"00",
          8504 => x"00",
          8505 => x"00",
          8506 => x"00",
          8507 => x"00",
          8508 => x"00",
          8509 => x"00",
          8510 => x"00",
          8511 => x"00",
          8512 => x"00",
          8513 => x"00",
          8514 => x"00",
          8515 => x"00",
          8516 => x"00",
          8517 => x"00",
          8518 => x"00",
          8519 => x"00",
          8520 => x"00",
          8521 => x"00",
          8522 => x"00",
          8523 => x"00",
          8524 => x"00",
          8525 => x"00",
          8526 => x"00",
          8527 => x"00",
          8528 => x"00",
          8529 => x"00",
          8530 => x"00",
          8531 => x"00",
          8532 => x"00",
          8533 => x"00",
          8534 => x"00",
          8535 => x"00",
          8536 => x"00",
          8537 => x"00",
          8538 => x"00",
          8539 => x"00",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"00",
          8544 => x"00",
          8545 => x"00",
          8546 => x"00",
          8547 => x"00",
          8548 => x"00",
          8549 => x"00",
          8550 => x"00",
          8551 => x"00",
          8552 => x"00",
          8553 => x"00",
          8554 => x"00",
          8555 => x"00",
          8556 => x"00",
          8557 => x"00",
          8558 => x"00",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"00",
          8573 => x"00",
          8574 => x"00",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
          8818 => x"00",
          8819 => x"00",
          8820 => x"00",
          8821 => x"00",
          8822 => x"00",
          8823 => x"00",
          8824 => x"00",
          8825 => x"00",
          8826 => x"00",
          8827 => x"00",
          8828 => x"00",
          8829 => x"00",
          8830 => x"00",
          8831 => x"00",
          8832 => x"00",
          8833 => x"00",
          8834 => x"00",
          8835 => x"00",
          8836 => x"00",
          8837 => x"00",
          8838 => x"00",
          8839 => x"00",
          8840 => x"00",
          8841 => x"00",
          8842 => x"00",
          8843 => x"00",
          8844 => x"00",
          8845 => x"00",
          8846 => x"00",
          8847 => x"00",
          8848 => x"00",
          8849 => x"00",
          8850 => x"00",
          8851 => x"00",
          8852 => x"00",
          8853 => x"00",
          8854 => x"00",
          8855 => x"00",
          8856 => x"00",
          8857 => x"00",
          8858 => x"00",
          8859 => x"00",
          8860 => x"00",
          8861 => x"00",
          8862 => x"00",
          8863 => x"00",
          8864 => x"00",
          8865 => x"00",
          8866 => x"00",
          8867 => x"00",
          8868 => x"00",
          8869 => x"00",
          8870 => x"00",
          8871 => x"00",
          8872 => x"00",
          8873 => x"00",
          8874 => x"00",
          8875 => x"00",
          8876 => x"00",
          8877 => x"00",
          8878 => x"00",
          8879 => x"00",
          8880 => x"00",
          8881 => x"00",
          8882 => x"00",
          8883 => x"00",
          8884 => x"00",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"00",
          8923 => x"00",
          8924 => x"00",
          8925 => x"00",
          8926 => x"00",
          8927 => x"00",
          8928 => x"00",
          8929 => x"00",
          8930 => x"00",
          8931 => x"00",
          8932 => x"00",
          8933 => x"00",
          8934 => x"00",
          8935 => x"00",
          8936 => x"00",
          8937 => x"00",
          8938 => x"00",
          8939 => x"00",
          8940 => x"00",
          8941 => x"00",
          8942 => x"00",
          8943 => x"00",
          8944 => x"00",
          8945 => x"00",
          8946 => x"00",
          8947 => x"00",
          8948 => x"00",
          8949 => x"00",
          8950 => x"00",
          8951 => x"00",
          8952 => x"00",
          8953 => x"00",
          8954 => x"00",
          8955 => x"00",
          8956 => x"00",
          8957 => x"00",
          8958 => x"00",
          8959 => x"00",
          8960 => x"00",
          8961 => x"00",
          8962 => x"00",
          8963 => x"00",
          8964 => x"00",
          8965 => x"00",
          8966 => x"00",
          8967 => x"00",
          8968 => x"00",
          8969 => x"00",
          8970 => x"00",
          8971 => x"00",
          8972 => x"00",
          8973 => x"00",
          8974 => x"00",
          8975 => x"00",
          8976 => x"00",
          8977 => x"00",
          8978 => x"00",
          8979 => x"00",
          8980 => x"00",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"00",
          9020 => x"00",
          9021 => x"00",
          9022 => x"00",
          9023 => x"00",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"00",
          9028 => x"00",
          9029 => x"00",
          9030 => x"00",
          9031 => x"00",
          9032 => x"00",
          9033 => x"00",
          9034 => x"00",
          9035 => x"00",
          9036 => x"00",
          9037 => x"00",
          9038 => x"00",
          9039 => x"00",
          9040 => x"00",
          9041 => x"00",
          9042 => x"00",
          9043 => x"00",
          9044 => x"00",
          9045 => x"00",
          9046 => x"00",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"00",
          9052 => x"00",
          9053 => x"00",
          9054 => x"00",
          9055 => x"00",
          9056 => x"00",
          9057 => x"00",
          9058 => x"00",
          9059 => x"00",
          9060 => x"00",
          9061 => x"00",
          9062 => x"00",
          9063 => x"00",
          9064 => x"00",
          9065 => x"00",
          9066 => x"00",
          9067 => x"00",
          9068 => x"ce",
          9069 => x"fc",
          9070 => x"c4",
          9071 => x"eb",
          9072 => x"64",
          9073 => x"2f",
          9074 => x"24",
          9075 => x"51",
          9076 => x"04",
          9077 => x"0c",
          9078 => x"14",
          9079 => x"59",
          9080 => x"84",
          9081 => x"8c",
          9082 => x"94",
          9083 => x"80",
          9084 => x"00",
          9085 => x"00",
          9086 => x"00",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"00",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"00",
          9097 => x"00",
          9098 => x"00",
          9099 => x"00",
          9100 => x"00",
        others => X"00"
    );

    signal RAM0_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM1_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM2_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM3_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM4_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM5_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM6_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM7_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM0_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM1_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM2_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM3_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM4_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM5_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM6_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM7_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal lowDataA          :     std_logic_vector(WORD_32BIT_RANGE);   -- Low word in 64 bit output from RAM matrix.
    signal highDataA         :     std_logic_vector(WORD_32BIT_RANGE);   -- High word in 64 bit output from RAM matrix.
    signal lowDataB          :     std_logic_vector(WORD_32BIT_RANGE);   -- Low word in 64 bit output from RAM matrix.
    signal highDataB         :     std_logic_vector(WORD_32BIT_RANGE);   -- High word in 64 bit output from RAM matrix.

begin

    -- Correctly assign the Little Endian value to the correct array, byte writes the data is in '7 downto 0', h-word writes
    -- the data is in '15 downto 0', word writes the data is in '31 downto 0'. Long words (64bits) are treated as two words for Endianness,
    -- and not as one continuous long word, this is because the ZPU is 32bit even when accessing a 64bit chunk.
    --
    RAM0_DATA <= memAWrite(7 downto 0)   when memAAddr(2) = '0'
                 else (others => '0');
    RAM1_DATA <= memAWrite(15 downto 8)  when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(15 downto 8)  when memAAddr(2) = '0' and (memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM4_DATA <= memAWrite(7 downto 0)   when memAAddr(2) = '1'
                 else (others => '0');
    RAM5_DATA <= memAWrite(15 downto 8)  when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM6_DATA <= memAWrite(23 downto 16) when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(7 downto 0);
    RAM7_DATA <= memAWrite(31 downto 24) when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(15 downto 8)  when memAAddr(2) = '1' and (memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "011") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "01"))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "010") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "01"))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "001") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "00"))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "000") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "00"))
                 else '0';
    RAM4_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "111") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "11"))
                 else '0';
    RAM5_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "110") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "11"))
                 else '0';
    RAM6_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "101") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "10"))
                 else '0';
    RAM7_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "100") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "10"))
                 else '0';

    memARead  <= lowDataA  when memAAddr(2) = '0'
                 else
                 highDataA;
    memBRead  <= lowDataB & highDataB;

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM0_DATA;
            else
                lowDataA(7 downto 0)    <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM1_DATA;
            else
                lowDataA(15 downto 8)   <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM2_DATA;
            else
                lowDataA(23 downto 16)  <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM3_DATA;
            else
                lowDataA(31 downto 24)  <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 4 - Port A - bits 39 to 32 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM4_WREN = '1' then
                RAM4(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM4_DATA;
            else
                highDataA(7 downto 0)   <= RAM4(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 5 - Port A - bits 47 to 40 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM5_WREN = '1' then
                RAM5(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM5_DATA;
            else
                highDataA(15 downto 8)  <= RAM5(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 6 - Port A - bits 56 to 48
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM6_WREN = '1' then
                RAM6(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM6_DATA;
            else
                highDataA(23 downto 16) <= RAM6(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 7 - Port A - bits 63 to 57 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM7_WREN = '1' then
                RAM7(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM7_DATA;
            else
                highDataA(31 downto 24) <= RAM7(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;


    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(7 downto 0);
                lowDataB(7 downto 0)    <= memBWrite(7 downto 0);
            else
                lowDataB(7 downto 0)    <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(15 downto 8);
                lowDataB(15 downto 8)    <= memBWrite(15 downto 8);
            else
                lowDataB(15 downto 8)    <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(23 downto 16);
                lowDataB(23 downto 16)  <= memBWrite(23 downto 16);
            else
                lowDataB(23 downto 16)  <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(31 downto 24);
                lowDataB(31 downto 24)  <= memBWrite(31 downto 24);
            else
                lowDataB(31 downto 24)  <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 4 - Port B - bits 39 downto 32
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM4(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(39 downto 32);
                highDataB(7 downto 0)   <= memBWrite(39 downto 32);
            else
                highDataB(7 downto 0)   <= RAM4(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 5 - Port B - bits 47 downto 40
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM5(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(47 downto 40);
                highDataB(15 downto 8)  <= memBWrite(47 downto 40);
            else
                highDataB(15 downto 8)  <= RAM5(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 6 - Port B - bits 55 downto 48
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM6(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(55 downto 48);
                highDataB(23 downto 16)  <= memBWrite(55 downto 48);
            else
                highDataB(23 downto 16)  <= RAM6(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 7 - Port B - bits 63 downto 56 
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM7(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(63 downto 56);
                highDataB(31 downto 24)  <= memBWrite(63 downto 56);
            else
                highDataB(31 downto 24)  <= RAM7(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

end arch;
