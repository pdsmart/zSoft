-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b83ff",
             1 => x"f80d0b0b",
             2 => x"0b93b704",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b93",
            73 => x"9b040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b92fe",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b8299",
           162 => x"a0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"93830400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b80cf",
           171 => x"942d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b80d1",
           179 => x"802d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"95040b0b",
           269 => x"0b8ca404",
           270 => x"0b0b0b8c",
           271 => x"b3040b0b",
           272 => x"0b8cc204",
           273 => x"0b0b0b8c",
           274 => x"d1040b0b",
           275 => x"0b8ce004",
           276 => x"0b0b0b8c",
           277 => x"ef040b0b",
           278 => x"0b8cfe04",
           279 => x"0b0b0b8d",
           280 => x"8d040b0b",
           281 => x"0b8d9c04",
           282 => x"0b0b0b8d",
           283 => x"ab040b0b",
           284 => x"0b8dbb04",
           285 => x"0b0b0b8d",
           286 => x"cb040b0b",
           287 => x"0b8ddb04",
           288 => x"0b0b0b8d",
           289 => x"eb040b0b",
           290 => x"0b8dfb04",
           291 => x"0b0b0b8e",
           292 => x"8b040b0b",
           293 => x"0b8e9b04",
           294 => x"0b0b0b8e",
           295 => x"ab040b0b",
           296 => x"0b8ebb04",
           297 => x"0b0b0b8e",
           298 => x"cb040b0b",
           299 => x"0b8edb04",
           300 => x"0b0b0b8e",
           301 => x"eb040b0b",
           302 => x"0b8efb04",
           303 => x"0b0b0b8f",
           304 => x"8b040b0b",
           305 => x"0b8f9b04",
           306 => x"0b0b0b8f",
           307 => x"ab040b0b",
           308 => x"0b8fbb04",
           309 => x"0b0b0b8f",
           310 => x"cb040b0b",
           311 => x"0b8fdb04",
           312 => x"0b0b0b8f",
           313 => x"eb040b0b",
           314 => x"0b8ffb04",
           315 => x"0b0b0b90",
           316 => x"8b040b0b",
           317 => x"0b909b04",
           318 => x"0b0b0b90",
           319 => x"ab040b0b",
           320 => x"0b90bb04",
           321 => x"0b0b0b90",
           322 => x"cb040b0b",
           323 => x"0b90db04",
           324 => x"0b0b0b90",
           325 => x"eb040b0b",
           326 => x"0b90fb04",
           327 => x"0b0b0b91",
           328 => x"8b040b0b",
           329 => x"0b919b04",
           330 => x"0b0b0b91",
           331 => x"ab040b0b",
           332 => x"0b91bb04",
           333 => x"0b0b0b91",
           334 => x"cb040b0b",
           335 => x"0b91db04",
           336 => x"0b0b0b91",
           337 => x"eb040b0b",
           338 => x"0b91fb04",
           339 => x"0b0b0b92",
           340 => x"8b040b0b",
           341 => x"0b929b04",
           342 => x"0b0b0b92",
           343 => x"ab040b0b",
           344 => x"0b92bb04",
           345 => x"0b0b0b92",
           346 => x"cb04ffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0482bba4",
           386 => x"0c80f8f5",
           387 => x"2d82bba4",
           388 => x"0882e090",
           389 => x"0482bba4",
           390 => x"0cbed22d",
           391 => x"82bba408",
           392 => x"82e09004",
           393 => x"82bba40c",
           394 => x"bb832d82",
           395 => x"bba40882",
           396 => x"e0900482",
           397 => x"bba40cb4",
           398 => x"fc2d82bb",
           399 => x"a40882e0",
           400 => x"900482bb",
           401 => x"a40c94ab",
           402 => x"2d82bba4",
           403 => x"0882e090",
           404 => x"0482bba4",
           405 => x"0cbce22d",
           406 => x"82bba408",
           407 => x"82e09004",
           408 => x"82bba40c",
           409 => x"b5b22d82",
           410 => x"bba40882",
           411 => x"e0900482",
           412 => x"bba40caf",
           413 => x"ab2d82bb",
           414 => x"a40882e0",
           415 => x"900482bb",
           416 => x"a40c93d6",
           417 => x"2d82bba4",
           418 => x"0882e090",
           419 => x"0482bba4",
           420 => x"0c96be2d",
           421 => x"82bba408",
           422 => x"82e09004",
           423 => x"82bba40c",
           424 => x"97cb2d82",
           425 => x"bba40882",
           426 => x"e0900482",
           427 => x"bba40c80",
           428 => x"fc9f2d82",
           429 => x"bba40882",
           430 => x"e0900482",
           431 => x"bba40c80",
           432 => x"fcfd2d82",
           433 => x"bba40882",
           434 => x"e0900482",
           435 => x"bba40c80",
           436 => x"f4b92d82",
           437 => x"bba40882",
           438 => x"e0900482",
           439 => x"bba40c80",
           440 => x"f6b12d82",
           441 => x"bba40882",
           442 => x"e0900482",
           443 => x"bba40c80",
           444 => x"f7e42d82",
           445 => x"bba40882",
           446 => x"e0900482",
           447 => x"bba40c81",
           448 => x"dc842d82",
           449 => x"bba40882",
           450 => x"e0900482",
           451 => x"bba40c81",
           452 => x"e8f52d82",
           453 => x"bba40882",
           454 => x"e0900482",
           455 => x"bba40c81",
           456 => x"e0e92d82",
           457 => x"bba40882",
           458 => x"e0900482",
           459 => x"bba40c81",
           460 => x"e3e62d82",
           461 => x"bba40882",
           462 => x"e0900482",
           463 => x"bba40c81",
           464 => x"ee842d82",
           465 => x"bba40882",
           466 => x"e0900482",
           467 => x"bba40c81",
           468 => x"f6e42d82",
           469 => x"bba40882",
           470 => x"e0900482",
           471 => x"bba40c81",
           472 => x"e7d72d82",
           473 => x"bba40882",
           474 => x"e0900482",
           475 => x"bba40c81",
           476 => x"f1a32d82",
           477 => x"bba40882",
           478 => x"e0900482",
           479 => x"bba40c81",
           480 => x"f2c22d82",
           481 => x"bba40882",
           482 => x"e0900482",
           483 => x"bba40c81",
           484 => x"f2e12d82",
           485 => x"bba40882",
           486 => x"e0900482",
           487 => x"bba40c81",
           488 => x"facb2d82",
           489 => x"bba40882",
           490 => x"e0900482",
           491 => x"bba40c81",
           492 => x"f8b12d82",
           493 => x"bba40882",
           494 => x"e0900482",
           495 => x"bba40c81",
           496 => x"fd9f2d82",
           497 => x"bba40882",
           498 => x"e0900482",
           499 => x"bba40c81",
           500 => x"f3e52d82",
           501 => x"bba40882",
           502 => x"e0900482",
           503 => x"bba40c82",
           504 => x"809f2d82",
           505 => x"bba40882",
           506 => x"e0900482",
           507 => x"bba40c82",
           508 => x"81a02d82",
           509 => x"bba40882",
           510 => x"e0900482",
           511 => x"bba40c81",
           512 => x"e9d52d82",
           513 => x"bba40882",
           514 => x"e0900482",
           515 => x"bba40c81",
           516 => x"e9ae2d82",
           517 => x"bba40882",
           518 => x"e0900482",
           519 => x"bba40c81",
           520 => x"ead92d82",
           521 => x"bba40882",
           522 => x"e0900482",
           523 => x"bba40c81",
           524 => x"f4bc2d82",
           525 => x"bba40882",
           526 => x"e0900482",
           527 => x"bba40c82",
           528 => x"82912d82",
           529 => x"bba40882",
           530 => x"e0900482",
           531 => x"bba40c82",
           532 => x"849b2d82",
           533 => x"bba40882",
           534 => x"e0900482",
           535 => x"bba40c82",
           536 => x"87dd2d82",
           537 => x"bba40882",
           538 => x"e0900482",
           539 => x"bba40c81",
           540 => x"dba32d82",
           541 => x"bba40882",
           542 => x"e0900482",
           543 => x"bba40c82",
           544 => x"8ac92d82",
           545 => x"bba40882",
           546 => x"e0900482",
           547 => x"bba40c82",
           548 => x"98fe2d82",
           549 => x"bba40882",
           550 => x"e0900482",
           551 => x"bba40c82",
           552 => x"96ea2d82",
           553 => x"bba40882",
           554 => x"e0900482",
           555 => x"bba40c81",
           556 => x"acde2d82",
           557 => x"bba40882",
           558 => x"e0900482",
           559 => x"bba40c81",
           560 => x"aec82d82",
           561 => x"bba40882",
           562 => x"e0900482",
           563 => x"bba40c81",
           564 => x"b0ac2d82",
           565 => x"bba40882",
           566 => x"e0900482",
           567 => x"bba40c80",
           568 => x"f4e22d82",
           569 => x"bba40882",
           570 => x"e0900482",
           571 => x"bba40c80",
           572 => x"f6862d82",
           573 => x"bba40882",
           574 => x"e0900482",
           575 => x"bba40c80",
           576 => x"f9ea2d82",
           577 => x"bba40882",
           578 => x"e0900482",
           579 => x"bba40c80",
           580 => x"d6962d82",
           581 => x"bba40882",
           582 => x"e0900482",
           583 => x"bba40c81",
           584 => x"a6f22d82",
           585 => x"bba40882",
           586 => x"e0900482",
           587 => x"bba40c81",
           588 => x"a79a2d82",
           589 => x"bba40882",
           590 => x"e0900482",
           591 => x"bba40c81",
           592 => x"ab922d82",
           593 => x"bba40882",
           594 => x"e0900482",
           595 => x"bba40c81",
           596 => x"a3dc2d82",
           597 => x"bba40882",
           598 => x"e090043c",
           599 => x"04000010",
           600 => x"10101010",
           601 => x"10101010",
           602 => x"10101010",
           603 => x"10101010",
           604 => x"10101010",
           605 => x"10101010",
           606 => x"10101010",
           607 => x"10105351",
           608 => x"04000073",
           609 => x"81ff0673",
           610 => x"83060981",
           611 => x"05830510",
           612 => x"10102b07",
           613 => x"72fc060c",
           614 => x"51510472",
           615 => x"72807281",
           616 => x"06ff0509",
           617 => x"72060571",
           618 => x"1052720a",
           619 => x"100a5372",
           620 => x"ed385151",
           621 => x"53510482",
           622 => x"bb987082",
           623 => x"d2f4278e",
           624 => x"38807170",
           625 => x"8405530c",
           626 => x"0b0b0b93",
           627 => x"ba048c81",
           628 => x"5180f2fe",
           629 => x"040082bb",
           630 => x"a4080282",
           631 => x"bba40cfb",
           632 => x"3d0d82bb",
           633 => x"a4088c05",
           634 => x"7082bba4",
           635 => x"08fc050c",
           636 => x"82bba408",
           637 => x"fc050854",
           638 => x"82bba408",
           639 => x"88050853",
           640 => x"82d2ec08",
           641 => x"5254849a",
           642 => x"3f82bb98",
           643 => x"087082bb",
           644 => x"a408f805",
           645 => x"0c82bba4",
           646 => x"08f80508",
           647 => x"7082bb98",
           648 => x"0c515487",
           649 => x"3d0d82bb",
           650 => x"a40c0482",
           651 => x"bba40802",
           652 => x"82bba40c",
           653 => x"fb3d0d82",
           654 => x"bba40890",
           655 => x"05088511",
           656 => x"33708132",
           657 => x"70810651",
           658 => x"51515271",
           659 => x"8f38800b",
           660 => x"82bba408",
           661 => x"8c050825",
           662 => x"83388d39",
           663 => x"800b82bb",
           664 => x"a408f405",
           665 => x"0c81c439",
           666 => x"82bba408",
           667 => x"8c0508ff",
           668 => x"0582bba4",
           669 => x"088c050c",
           670 => x"800b82bb",
           671 => x"a408f805",
           672 => x"0c82bba4",
           673 => x"08880508",
           674 => x"82bba408",
           675 => x"fc050c82",
           676 => x"bba408f8",
           677 => x"05088a2e",
           678 => x"80f63880",
           679 => x"0b82bba4",
           680 => x"088c0508",
           681 => x"2580e938",
           682 => x"82bba408",
           683 => x"90050851",
           684 => x"abb23f82",
           685 => x"bb980870",
           686 => x"82bba408",
           687 => x"f8050c52",
           688 => x"82bba408",
           689 => x"f80508ff",
           690 => x"2e098106",
           691 => x"8d38800b",
           692 => x"82bba408",
           693 => x"f4050c80",
           694 => x"d23982bb",
           695 => x"a408fc05",
           696 => x"0882bba4",
           697 => x"08f80508",
           698 => x"53537173",
           699 => x"3482bba4",
           700 => x"088c0508",
           701 => x"ff0582bb",
           702 => x"a4088c05",
           703 => x"0c82bba4",
           704 => x"08fc0508",
           705 => x"810582bb",
           706 => x"a408fc05",
           707 => x"0cff8039",
           708 => x"82bba408",
           709 => x"fc050852",
           710 => x"80723482",
           711 => x"bba40888",
           712 => x"05087082",
           713 => x"bba408f4",
           714 => x"050c5282",
           715 => x"bba408f4",
           716 => x"050882bb",
           717 => x"980c873d",
           718 => x"0d82bba4",
           719 => x"0c0482bb",
           720 => x"a4080282",
           721 => x"bba40cf4",
           722 => x"3d0d860b",
           723 => x"82bba408",
           724 => x"e5053482",
           725 => x"bba40888",
           726 => x"050882bb",
           727 => x"a408e005",
           728 => x"0cfe0a0b",
           729 => x"82bba408",
           730 => x"e8050c82",
           731 => x"bba40890",
           732 => x"057082bb",
           733 => x"a408fc05",
           734 => x"0c82bba4",
           735 => x"08fc0508",
           736 => x"5482bba4",
           737 => x"088c0508",
           738 => x"5382bba4",
           739 => x"08e00570",
           740 => x"53515481",
           741 => x"8d3f82bb",
           742 => x"98087082",
           743 => x"bba408dc",
           744 => x"050c82bb",
           745 => x"a408ec05",
           746 => x"0882bba4",
           747 => x"08880508",
           748 => x"05515480",
           749 => x"743482bb",
           750 => x"a408dc05",
           751 => x"087082bb",
           752 => x"980c548e",
           753 => x"3d0d82bb",
           754 => x"a40c0482",
           755 => x"bba40802",
           756 => x"82bba40c",
           757 => x"fb3d0d82",
           758 => x"bba40890",
           759 => x"057082bb",
           760 => x"a408fc05",
           761 => x"0c82bba4",
           762 => x"08fc0508",
           763 => x"5482bba4",
           764 => x"088c0508",
           765 => x"5382bba4",
           766 => x"08880508",
           767 => x"5254a33f",
           768 => x"82bb9808",
           769 => x"7082bba4",
           770 => x"08f8050c",
           771 => x"82bba408",
           772 => x"f8050870",
           773 => x"82bb980c",
           774 => x"5154873d",
           775 => x"0d82bba4",
           776 => x"0c0482bb",
           777 => x"a4080282",
           778 => x"bba40ced",
           779 => x"3d0d800b",
           780 => x"82bba408",
           781 => x"e4052382",
           782 => x"bba40888",
           783 => x"05085380",
           784 => x"0b8c140c",
           785 => x"82bba408",
           786 => x"88050885",
           787 => x"11337081",
           788 => x"2a708132",
           789 => x"70810651",
           790 => x"51515153",
           791 => x"72802e8d",
           792 => x"38ff0b82",
           793 => x"bba408e0",
           794 => x"050c96ac",
           795 => x"3982bba4",
           796 => x"088c0508",
           797 => x"53723353",
           798 => x"7282bba4",
           799 => x"08f80534",
           800 => x"7281ff06",
           801 => x"5372802e",
           802 => x"95fa3882",
           803 => x"bba4088c",
           804 => x"05088105",
           805 => x"82bba408",
           806 => x"8c050c82",
           807 => x"bba408e4",
           808 => x"05227081",
           809 => x"06515372",
           810 => x"802e958b",
           811 => x"3882bba4",
           812 => x"08f80533",
           813 => x"53af7327",
           814 => x"81fc3882",
           815 => x"bba408f8",
           816 => x"05335372",
           817 => x"b92681ee",
           818 => x"3882bba4",
           819 => x"08f80533",
           820 => x"5372b02e",
           821 => x"09810680",
           822 => x"c53882bb",
           823 => x"a408e805",
           824 => x"3370982b",
           825 => x"70982c51",
           826 => x"515372b2",
           827 => x"3882bba4",
           828 => x"08e40522",
           829 => x"70832a70",
           830 => x"81327081",
           831 => x"06515151",
           832 => x"5372802e",
           833 => x"993882bb",
           834 => x"a408e405",
           835 => x"22708280",
           836 => x"07515372",
           837 => x"82bba408",
           838 => x"e40523fe",
           839 => x"d03982bb",
           840 => x"a408e805",
           841 => x"3370982b",
           842 => x"70982c70",
           843 => x"70832b72",
           844 => x"11731151",
           845 => x"51515351",
           846 => x"55537282",
           847 => x"bba408e8",
           848 => x"053482bb",
           849 => x"a408e805",
           850 => x"335482bb",
           851 => x"a408f805",
           852 => x"337015d0",
           853 => x"11515153",
           854 => x"7282bba4",
           855 => x"08e80534",
           856 => x"82bba408",
           857 => x"e8053370",
           858 => x"982b7098",
           859 => x"2c515153",
           860 => x"7280258b",
           861 => x"3880ff0b",
           862 => x"82bba408",
           863 => x"e8053482",
           864 => x"bba408e4",
           865 => x"05227083",
           866 => x"2a708106",
           867 => x"51515372",
           868 => x"fddb3882",
           869 => x"bba408e8",
           870 => x"05337088",
           871 => x"2b70902b",
           872 => x"70902c70",
           873 => x"882c5151",
           874 => x"51515372",
           875 => x"82bba408",
           876 => x"ec0523fd",
           877 => x"b83982bb",
           878 => x"a408e405",
           879 => x"2270832a",
           880 => x"70810651",
           881 => x"51537280",
           882 => x"2e9d3882",
           883 => x"bba408e8",
           884 => x"05337098",
           885 => x"2b70982c",
           886 => x"51515372",
           887 => x"8a38810b",
           888 => x"82bba408",
           889 => x"e8053482",
           890 => x"bba408f8",
           891 => x"0533e011",
           892 => x"82bba408",
           893 => x"c4050c53",
           894 => x"82bba408",
           895 => x"c4050880",
           896 => x"d8269294",
           897 => x"3882bba4",
           898 => x"08c40508",
           899 => x"70822b82",
           900 => x"9aec1170",
           901 => x"08515151",
           902 => x"53720482",
           903 => x"bba408e4",
           904 => x"05227090",
           905 => x"07515372",
           906 => x"82bba408",
           907 => x"e4052382",
           908 => x"bba408e4",
           909 => x"052270a0",
           910 => x"07515372",
           911 => x"82bba408",
           912 => x"e40523fc",
           913 => x"a83982bb",
           914 => x"a408e405",
           915 => x"22708180",
           916 => x"07515372",
           917 => x"82bba408",
           918 => x"e40523fc",
           919 => x"903982bb",
           920 => x"a408e405",
           921 => x"227080c0",
           922 => x"07515372",
           923 => x"82bba408",
           924 => x"e40523fb",
           925 => x"f83982bb",
           926 => x"a408e405",
           927 => x"22708807",
           928 => x"51537282",
           929 => x"bba408e4",
           930 => x"0523800b",
           931 => x"82bba408",
           932 => x"e80534fb",
           933 => x"d83982bb",
           934 => x"a408e405",
           935 => x"22708407",
           936 => x"51537282",
           937 => x"bba408e4",
           938 => x"0523fbc1",
           939 => x"39bf0b82",
           940 => x"bba408fc",
           941 => x"053482bb",
           942 => x"a408ec05",
           943 => x"22ff1151",
           944 => x"537282bb",
           945 => x"a408ec05",
           946 => x"2380e30b",
           947 => x"82bba408",
           948 => x"f805348d",
           949 => x"a83982bb",
           950 => x"a4089005",
           951 => x"0882bba4",
           952 => x"08900508",
           953 => x"840582bb",
           954 => x"a4089005",
           955 => x"0c700851",
           956 => x"537282bb",
           957 => x"a408fc05",
           958 => x"3482bba4",
           959 => x"08ec0522",
           960 => x"ff115153",
           961 => x"7282bba4",
           962 => x"08ec0523",
           963 => x"8cef3982",
           964 => x"bba40890",
           965 => x"050882bb",
           966 => x"a4089005",
           967 => x"08840582",
           968 => x"bba40890",
           969 => x"050c7008",
           970 => x"82bba408",
           971 => x"fc050c82",
           972 => x"bba408e4",
           973 => x"05227083",
           974 => x"2a708106",
           975 => x"51515153",
           976 => x"72802eab",
           977 => x"3882bba4",
           978 => x"08e80533",
           979 => x"70982b53",
           980 => x"72982c53",
           981 => x"82bba408",
           982 => x"fc050852",
           983 => x"53adfa3f",
           984 => x"82bb9808",
           985 => x"537282bb",
           986 => x"a408f405",
           987 => x"23993982",
           988 => x"bba408fc",
           989 => x"050851a8",
           990 => x"ac3f82bb",
           991 => x"98085372",
           992 => x"82bba408",
           993 => x"f4052382",
           994 => x"bba408ec",
           995 => x"05225382",
           996 => x"bba408f4",
           997 => x"05227371",
           998 => x"31545472",
           999 => x"82bba408",
          1000 => x"ec05238b",
          1001 => x"d83982bb",
          1002 => x"a4089005",
          1003 => x"0882bba4",
          1004 => x"08900508",
          1005 => x"840582bb",
          1006 => x"a4089005",
          1007 => x"0c700882",
          1008 => x"bba408fc",
          1009 => x"050c82bb",
          1010 => x"a408e405",
          1011 => x"2270832a",
          1012 => x"70810651",
          1013 => x"51515372",
          1014 => x"802eab38",
          1015 => x"82bba408",
          1016 => x"e8053370",
          1017 => x"982b5372",
          1018 => x"982c5382",
          1019 => x"bba408fc",
          1020 => x"05085253",
          1021 => x"ace33f82",
          1022 => x"bb980853",
          1023 => x"7282bba4",
          1024 => x"08f40523",
          1025 => x"993982bb",
          1026 => x"a408fc05",
          1027 => x"0851a795",
          1028 => x"3f82bb98",
          1029 => x"08537282",
          1030 => x"bba408f4",
          1031 => x"052382bb",
          1032 => x"a408ec05",
          1033 => x"225382bb",
          1034 => x"a408f405",
          1035 => x"22737131",
          1036 => x"54547282",
          1037 => x"bba408ec",
          1038 => x"05238ac1",
          1039 => x"3982bba4",
          1040 => x"08e40522",
          1041 => x"70822a70",
          1042 => x"81065151",
          1043 => x"5372802e",
          1044 => x"a43882bb",
          1045 => x"a4089005",
          1046 => x"0882bba4",
          1047 => x"08900508",
          1048 => x"840582bb",
          1049 => x"a4089005",
          1050 => x"0c700882",
          1051 => x"bba408dc",
          1052 => x"050c53a2",
          1053 => x"3982bba4",
          1054 => x"08900508",
          1055 => x"82bba408",
          1056 => x"90050884",
          1057 => x"0582bba4",
          1058 => x"0890050c",
          1059 => x"700882bb",
          1060 => x"a408dc05",
          1061 => x"0c5382bb",
          1062 => x"a408dc05",
          1063 => x"0882bba4",
          1064 => x"08fc050c",
          1065 => x"82bba408",
          1066 => x"fc050880",
          1067 => x"25a43882",
          1068 => x"bba408e4",
          1069 => x"05227082",
          1070 => x"07515372",
          1071 => x"82bba408",
          1072 => x"e4052382",
          1073 => x"bba408fc",
          1074 => x"05083082",
          1075 => x"bba408fc",
          1076 => x"050c82bb",
          1077 => x"a408e405",
          1078 => x"2270ffbf",
          1079 => x"06515372",
          1080 => x"82bba408",
          1081 => x"e4052381",
          1082 => x"af39880b",
          1083 => x"82bba408",
          1084 => x"f40523a9",
          1085 => x"3982bba4",
          1086 => x"08e40522",
          1087 => x"7080c007",
          1088 => x"51537282",
          1089 => x"bba408e4",
          1090 => x"052380f8",
          1091 => x"0b82bba4",
          1092 => x"08f80534",
          1093 => x"900b82bb",
          1094 => x"a408f405",
          1095 => x"2382bba4",
          1096 => x"08e40522",
          1097 => x"70822a70",
          1098 => x"81065151",
          1099 => x"5372802e",
          1100 => x"a43882bb",
          1101 => x"a4089005",
          1102 => x"0882bba4",
          1103 => x"08900508",
          1104 => x"840582bb",
          1105 => x"a4089005",
          1106 => x"0c700882",
          1107 => x"bba408d8",
          1108 => x"050c53a2",
          1109 => x"3982bba4",
          1110 => x"08900508",
          1111 => x"82bba408",
          1112 => x"90050884",
          1113 => x"0582bba4",
          1114 => x"0890050c",
          1115 => x"700882bb",
          1116 => x"a408d805",
          1117 => x"0c5382bb",
          1118 => x"a408d805",
          1119 => x"0882bba4",
          1120 => x"08fc050c",
          1121 => x"82bba408",
          1122 => x"e4052270",
          1123 => x"cf065153",
          1124 => x"7282bba4",
          1125 => x"08e40523",
          1126 => x"82bba80b",
          1127 => x"82bba408",
          1128 => x"f0050c82",
          1129 => x"bba408f0",
          1130 => x"050882bb",
          1131 => x"a408f405",
          1132 => x"2282bba4",
          1133 => x"08fc0508",
          1134 => x"71557054",
          1135 => x"565455af",
          1136 => x"953f82bb",
          1137 => x"98085372",
          1138 => x"753482bb",
          1139 => x"a408f005",
          1140 => x"0882bba4",
          1141 => x"08d4050c",
          1142 => x"82bba408",
          1143 => x"f0050870",
          1144 => x"33515389",
          1145 => x"7327a438",
          1146 => x"82bba408",
          1147 => x"f0050853",
          1148 => x"72335482",
          1149 => x"bba408f8",
          1150 => x"05337015",
          1151 => x"df115151",
          1152 => x"537282bb",
          1153 => x"a408d005",
          1154 => x"34973982",
          1155 => x"bba408f0",
          1156 => x"05085372",
          1157 => x"33b01151",
          1158 => x"537282bb",
          1159 => x"a408d005",
          1160 => x"3482bba4",
          1161 => x"08d40508",
          1162 => x"5382bba4",
          1163 => x"08d00533",
          1164 => x"733482bb",
          1165 => x"a408f005",
          1166 => x"08810582",
          1167 => x"bba408f0",
          1168 => x"050c82bb",
          1169 => x"a408f405",
          1170 => x"22705382",
          1171 => x"bba408fc",
          1172 => x"05085253",
          1173 => x"adcd3f82",
          1174 => x"bb980870",
          1175 => x"82bba408",
          1176 => x"fc050c53",
          1177 => x"82bba408",
          1178 => x"fc050880",
          1179 => x"2e8438fe",
          1180 => x"b23982bb",
          1181 => x"a408f005",
          1182 => x"0882bba8",
          1183 => x"54557254",
          1184 => x"74707531",
          1185 => x"51537282",
          1186 => x"bba408fc",
          1187 => x"053482bb",
          1188 => x"a408e405",
          1189 => x"2270b206",
          1190 => x"51537280",
          1191 => x"2e943882",
          1192 => x"bba408ec",
          1193 => x"0522ff11",
          1194 => x"51537282",
          1195 => x"bba408ec",
          1196 => x"052382bb",
          1197 => x"a408e405",
          1198 => x"2270862a",
          1199 => x"70810651",
          1200 => x"51537280",
          1201 => x"2e80e738",
          1202 => x"82bba408",
          1203 => x"ec052270",
          1204 => x"902b82bb",
          1205 => x"a408cc05",
          1206 => x"0c82bba4",
          1207 => x"08cc0508",
          1208 => x"902c82bb",
          1209 => x"a408cc05",
          1210 => x"0c82bba4",
          1211 => x"08f40522",
          1212 => x"51537290",
          1213 => x"2e098106",
          1214 => x"953882bb",
          1215 => x"a408cc05",
          1216 => x"08fe0553",
          1217 => x"7282bba4",
          1218 => x"08c80523",
          1219 => x"933982bb",
          1220 => x"a408cc05",
          1221 => x"08ff0553",
          1222 => x"7282bba4",
          1223 => x"08c80523",
          1224 => x"82bba408",
          1225 => x"c8052282",
          1226 => x"bba408ec",
          1227 => x"052382bb",
          1228 => x"a408e405",
          1229 => x"2270832a",
          1230 => x"70810651",
          1231 => x"51537280",
          1232 => x"2e80d038",
          1233 => x"82bba408",
          1234 => x"e8053370",
          1235 => x"982b7098",
          1236 => x"2c82bba4",
          1237 => x"08fc0533",
          1238 => x"57515153",
          1239 => x"72742497",
          1240 => x"3882bba4",
          1241 => x"08e40522",
          1242 => x"70f70651",
          1243 => x"537282bb",
          1244 => x"a408e405",
          1245 => x"239d3982",
          1246 => x"bba408e8",
          1247 => x"05335382",
          1248 => x"bba408fc",
          1249 => x"05337371",
          1250 => x"31545472",
          1251 => x"82bba408",
          1252 => x"e8053482",
          1253 => x"bba408e4",
          1254 => x"05227083",
          1255 => x"2a708106",
          1256 => x"51515372",
          1257 => x"802eb138",
          1258 => x"82bba408",
          1259 => x"e8053370",
          1260 => x"882b7090",
          1261 => x"2b70902c",
          1262 => x"70882c51",
          1263 => x"51515153",
          1264 => x"725482bb",
          1265 => x"a408ec05",
          1266 => x"22707531",
          1267 => x"51537282",
          1268 => x"bba408ec",
          1269 => x"0523af39",
          1270 => x"82bba408",
          1271 => x"fc053370",
          1272 => x"882b7090",
          1273 => x"2b70902c",
          1274 => x"70882c51",
          1275 => x"51515153",
          1276 => x"725482bb",
          1277 => x"a408ec05",
          1278 => x"22707531",
          1279 => x"51537282",
          1280 => x"bba408ec",
          1281 => x"052382bb",
          1282 => x"a408e405",
          1283 => x"22708380",
          1284 => x"06515372",
          1285 => x"b03882bb",
          1286 => x"a408ec05",
          1287 => x"22ff1154",
          1288 => x"547282bb",
          1289 => x"a408ec05",
          1290 => x"2373902b",
          1291 => x"70902c51",
          1292 => x"53807325",
          1293 => x"903882bb",
          1294 => x"a4088805",
          1295 => x"0852a051",
          1296 => x"96903fd2",
          1297 => x"3982bba4",
          1298 => x"08e40522",
          1299 => x"70812a70",
          1300 => x"81065151",
          1301 => x"5372802e",
          1302 => x"913882bb",
          1303 => x"a4088805",
          1304 => x"0852ad51",
          1305 => x"95ec3f80",
          1306 => x"c73982bb",
          1307 => x"a408e405",
          1308 => x"2270842a",
          1309 => x"70810651",
          1310 => x"51537280",
          1311 => x"2e903882",
          1312 => x"bba40888",
          1313 => x"050852ab",
          1314 => x"5195c73f",
          1315 => x"a33982bb",
          1316 => x"a408e405",
          1317 => x"2270852a",
          1318 => x"70810651",
          1319 => x"51537280",
          1320 => x"2e8e3882",
          1321 => x"bba40888",
          1322 => x"050852a0",
          1323 => x"5195a33f",
          1324 => x"82bba408",
          1325 => x"e4052270",
          1326 => x"862a7081",
          1327 => x"06515153",
          1328 => x"72802eb1",
          1329 => x"3882bba4",
          1330 => x"08880508",
          1331 => x"52b05195",
          1332 => x"813f82bb",
          1333 => x"a408f405",
          1334 => x"22537290",
          1335 => x"2e098106",
          1336 => x"943882bb",
          1337 => x"a4088805",
          1338 => x"085282bb",
          1339 => x"a408f805",
          1340 => x"335194de",
          1341 => x"3f82bba4",
          1342 => x"08e40522",
          1343 => x"70882a70",
          1344 => x"81065151",
          1345 => x"5372802e",
          1346 => x"b03882bb",
          1347 => x"a408ec05",
          1348 => x"22ff1154",
          1349 => x"547282bb",
          1350 => x"a408ec05",
          1351 => x"2373902b",
          1352 => x"70902c51",
          1353 => x"53807325",
          1354 => x"903882bb",
          1355 => x"a4088805",
          1356 => x"0852b051",
          1357 => x"949c3fd2",
          1358 => x"3982bba4",
          1359 => x"08e40522",
          1360 => x"70832a70",
          1361 => x"81065151",
          1362 => x"5372802e",
          1363 => x"b03882bb",
          1364 => x"a408e805",
          1365 => x"33ff1154",
          1366 => x"547282bb",
          1367 => x"a408e805",
          1368 => x"3473982b",
          1369 => x"70982c51",
          1370 => x"53807325",
          1371 => x"903882bb",
          1372 => x"a4088805",
          1373 => x"0852b051",
          1374 => x"93d83fd2",
          1375 => x"3982bba4",
          1376 => x"08e40522",
          1377 => x"70872a70",
          1378 => x"81065151",
          1379 => x"5372b038",
          1380 => x"82bba408",
          1381 => x"ec0522ff",
          1382 => x"11545472",
          1383 => x"82bba408",
          1384 => x"ec052373",
          1385 => x"902b7090",
          1386 => x"2c515380",
          1387 => x"73259038",
          1388 => x"82bba408",
          1389 => x"88050852",
          1390 => x"a0519396",
          1391 => x"3fd23982",
          1392 => x"bba408f8",
          1393 => x"05335372",
          1394 => x"80e32e09",
          1395 => x"81069738",
          1396 => x"82bba408",
          1397 => x"88050852",
          1398 => x"82bba408",
          1399 => x"fc053351",
          1400 => x"92f03f81",
          1401 => x"ee3982bb",
          1402 => x"a408f805",
          1403 => x"33537280",
          1404 => x"f32e0981",
          1405 => x"0680cb38",
          1406 => x"82bba408",
          1407 => x"f40522ff",
          1408 => x"11515372",
          1409 => x"82bba408",
          1410 => x"f4052372",
          1411 => x"83ffff06",
          1412 => x"537283ff",
          1413 => x"ff2e81bb",
          1414 => x"3882bba4",
          1415 => x"08880508",
          1416 => x"5282bba4",
          1417 => x"08fc0508",
          1418 => x"70335282",
          1419 => x"bba408fc",
          1420 => x"05088105",
          1421 => x"82bba408",
          1422 => x"fc050c53",
          1423 => x"92943fff",
          1424 => x"b73982bb",
          1425 => x"a408f805",
          1426 => x"33537280",
          1427 => x"d32e0981",
          1428 => x"0680cb38",
          1429 => x"82bba408",
          1430 => x"f40522ff",
          1431 => x"11515372",
          1432 => x"82bba408",
          1433 => x"f4052372",
          1434 => x"83ffff06",
          1435 => x"537283ff",
          1436 => x"ff2e80df",
          1437 => x"3882bba4",
          1438 => x"08880508",
          1439 => x"5282bba4",
          1440 => x"08fc0508",
          1441 => x"70335253",
          1442 => x"91c83f82",
          1443 => x"bba408fc",
          1444 => x"05088105",
          1445 => x"82bba408",
          1446 => x"fc050cff",
          1447 => x"b73982bb",
          1448 => x"a408f005",
          1449 => x"0882bba8",
          1450 => x"2ea93882",
          1451 => x"bba40888",
          1452 => x"05085282",
          1453 => x"bba408f0",
          1454 => x"0508ff05",
          1455 => x"82bba408",
          1456 => x"f0050c82",
          1457 => x"bba408f0",
          1458 => x"05087033",
          1459 => x"52539182",
          1460 => x"3fcc3982",
          1461 => x"bba408e4",
          1462 => x"05227087",
          1463 => x"2a708106",
          1464 => x"51515372",
          1465 => x"802e80c3",
          1466 => x"3882bba4",
          1467 => x"08ec0522",
          1468 => x"ff115454",
          1469 => x"7282bba4",
          1470 => x"08ec0523",
          1471 => x"73902b70",
          1472 => x"902c5153",
          1473 => x"807325a3",
          1474 => x"3882bba4",
          1475 => x"08880508",
          1476 => x"52a05190",
          1477 => x"bd3fd239",
          1478 => x"82bba408",
          1479 => x"88050852",
          1480 => x"82bba408",
          1481 => x"f8053351",
          1482 => x"90a83f80",
          1483 => x"0b82bba4",
          1484 => x"08e40523",
          1485 => x"eab73982",
          1486 => x"bba408f8",
          1487 => x"05335372",
          1488 => x"a52e0981",
          1489 => x"06a83881",
          1490 => x"0b82bba4",
          1491 => x"08e40523",
          1492 => x"800b82bb",
          1493 => x"a408ec05",
          1494 => x"23800b82",
          1495 => x"bba408e8",
          1496 => x"05348a0b",
          1497 => x"82bba408",
          1498 => x"f40523ea",
          1499 => x"803982bb",
          1500 => x"a4088805",
          1501 => x"085282bb",
          1502 => x"a408f805",
          1503 => x"33518fd2",
          1504 => x"3fe9ea39",
          1505 => x"82bba408",
          1506 => x"8805088c",
          1507 => x"11087082",
          1508 => x"bba408e0",
          1509 => x"050c5153",
          1510 => x"82bba408",
          1511 => x"e0050882",
          1512 => x"bb980c95",
          1513 => x"3d0d82bb",
          1514 => x"a40c0482",
          1515 => x"bba40802",
          1516 => x"82bba40c",
          1517 => x"f73d0d80",
          1518 => x"0b82bba4",
          1519 => x"08f00534",
          1520 => x"82bba408",
          1521 => x"8c050853",
          1522 => x"80730c82",
          1523 => x"bba40888",
          1524 => x"05087008",
          1525 => x"51537233",
          1526 => x"537282bb",
          1527 => x"a408f805",
          1528 => x"347281ff",
          1529 => x"065372a0",
          1530 => x"2e098106",
          1531 => x"913882bb",
          1532 => x"a4088805",
          1533 => x"08700881",
          1534 => x"05710c53",
          1535 => x"ce3982bb",
          1536 => x"a408f805",
          1537 => x"335372ad",
          1538 => x"2e098106",
          1539 => x"a438810b",
          1540 => x"82bba408",
          1541 => x"f0053482",
          1542 => x"bba40888",
          1543 => x"05087008",
          1544 => x"8105710c",
          1545 => x"70085153",
          1546 => x"723382bb",
          1547 => x"a408f805",
          1548 => x"3482bba4",
          1549 => x"08f80533",
          1550 => x"5372b02e",
          1551 => x"09810681",
          1552 => x"dc3882bb",
          1553 => x"a4088805",
          1554 => x"08700881",
          1555 => x"05710c70",
          1556 => x"08515372",
          1557 => x"3382bba4",
          1558 => x"08f80534",
          1559 => x"82bba408",
          1560 => x"f8053382",
          1561 => x"bba408e8",
          1562 => x"050c82bb",
          1563 => x"a408e805",
          1564 => x"0880e22e",
          1565 => x"b63882bb",
          1566 => x"a408e805",
          1567 => x"0880f82e",
          1568 => x"843880cd",
          1569 => x"39900b82",
          1570 => x"bba408f4",
          1571 => x"053482bb",
          1572 => x"a4088805",
          1573 => x"08700881",
          1574 => x"05710c70",
          1575 => x"08515372",
          1576 => x"3382bba4",
          1577 => x"08f80534",
          1578 => x"81a43982",
          1579 => x"0b82bba4",
          1580 => x"08f40534",
          1581 => x"82bba408",
          1582 => x"88050870",
          1583 => x"08810571",
          1584 => x"0c700851",
          1585 => x"53723382",
          1586 => x"bba408f8",
          1587 => x"053480fe",
          1588 => x"3982bba4",
          1589 => x"08f80533",
          1590 => x"5372a026",
          1591 => x"8d38810b",
          1592 => x"82bba408",
          1593 => x"ec050c83",
          1594 => x"803982bb",
          1595 => x"a408f805",
          1596 => x"3353af73",
          1597 => x"27903882",
          1598 => x"bba408f8",
          1599 => x"05335372",
          1600 => x"b9268338",
          1601 => x"8d39800b",
          1602 => x"82bba408",
          1603 => x"ec050c82",
          1604 => x"d839880b",
          1605 => x"82bba408",
          1606 => x"f40534b2",
          1607 => x"3982bba4",
          1608 => x"08f80533",
          1609 => x"53af7327",
          1610 => x"903882bb",
          1611 => x"a408f805",
          1612 => x"335372b9",
          1613 => x"2683388d",
          1614 => x"39800b82",
          1615 => x"bba408ec",
          1616 => x"050c82a5",
          1617 => x"398a0b82",
          1618 => x"bba408f4",
          1619 => x"0534800b",
          1620 => x"82bba408",
          1621 => x"fc050c82",
          1622 => x"bba408f8",
          1623 => x"053353a0",
          1624 => x"732781cf",
          1625 => x"3882bba4",
          1626 => x"08f80533",
          1627 => x"5380e073",
          1628 => x"27943882",
          1629 => x"bba408f8",
          1630 => x"0533e011",
          1631 => x"51537282",
          1632 => x"bba408f8",
          1633 => x"053482bb",
          1634 => x"a408f805",
          1635 => x"33d01151",
          1636 => x"537282bb",
          1637 => x"a408f805",
          1638 => x"3482bba4",
          1639 => x"08f80533",
          1640 => x"53907327",
          1641 => x"ad3882bb",
          1642 => x"a408f805",
          1643 => x"33f91151",
          1644 => x"537282bb",
          1645 => x"a408f805",
          1646 => x"3482bba4",
          1647 => x"08f80533",
          1648 => x"53728926",
          1649 => x"8d38800b",
          1650 => x"82bba408",
          1651 => x"ec050c81",
          1652 => x"983982bb",
          1653 => x"a408f805",
          1654 => x"3382bba4",
          1655 => x"08f40533",
          1656 => x"54547274",
          1657 => x"268d3880",
          1658 => x"0b82bba4",
          1659 => x"08ec050c",
          1660 => x"80f73982",
          1661 => x"bba408f4",
          1662 => x"05337082",
          1663 => x"bba408fc",
          1664 => x"05082982",
          1665 => x"bba408f8",
          1666 => x"05337012",
          1667 => x"82bba408",
          1668 => x"fc050c82",
          1669 => x"bba40888",
          1670 => x"05087008",
          1671 => x"8105710c",
          1672 => x"70085151",
          1673 => x"52555372",
          1674 => x"3382bba4",
          1675 => x"08f80534",
          1676 => x"fea53982",
          1677 => x"bba408f0",
          1678 => x"05335372",
          1679 => x"802e9038",
          1680 => x"82bba408",
          1681 => x"fc050830",
          1682 => x"82bba408",
          1683 => x"fc050c82",
          1684 => x"bba4088c",
          1685 => x"050882bb",
          1686 => x"a408fc05",
          1687 => x"08710c53",
          1688 => x"810b82bb",
          1689 => x"a408ec05",
          1690 => x"0c82bba4",
          1691 => x"08ec0508",
          1692 => x"82bb980c",
          1693 => x"8b3d0d82",
          1694 => x"bba40c04",
          1695 => x"82bba408",
          1696 => x"0282bba4",
          1697 => x"0cfd3d0d",
          1698 => x"82d2e808",
          1699 => x"5382bba4",
          1700 => x"088c0508",
          1701 => x"5282bba4",
          1702 => x"08880508",
          1703 => x"51df8c3f",
          1704 => x"82bb9808",
          1705 => x"7082bb98",
          1706 => x"0c54853d",
          1707 => x"0d82bba4",
          1708 => x"0c0482bb",
          1709 => x"a4080282",
          1710 => x"bba40cf7",
          1711 => x"3d0d800b",
          1712 => x"82bba408",
          1713 => x"f0053482",
          1714 => x"bba4088c",
          1715 => x"05085380",
          1716 => x"730c82bb",
          1717 => x"a4088805",
          1718 => x"08700851",
          1719 => x"53723353",
          1720 => x"7282bba4",
          1721 => x"08f80534",
          1722 => x"7281ff06",
          1723 => x"5372a02e",
          1724 => x"09810691",
          1725 => x"3882bba4",
          1726 => x"08880508",
          1727 => x"70088105",
          1728 => x"710c53ce",
          1729 => x"3982bba4",
          1730 => x"08f80533",
          1731 => x"5372ad2e",
          1732 => x"098106a4",
          1733 => x"38810b82",
          1734 => x"bba408f0",
          1735 => x"053482bb",
          1736 => x"a4088805",
          1737 => x"08700881",
          1738 => x"05710c70",
          1739 => x"08515372",
          1740 => x"3382bba4",
          1741 => x"08f80534",
          1742 => x"82bba408",
          1743 => x"f8053353",
          1744 => x"72b02e09",
          1745 => x"810681dc",
          1746 => x"3882bba4",
          1747 => x"08880508",
          1748 => x"70088105",
          1749 => x"710c7008",
          1750 => x"51537233",
          1751 => x"82bba408",
          1752 => x"f8053482",
          1753 => x"bba408f8",
          1754 => x"053382bb",
          1755 => x"a408e805",
          1756 => x"0c82bba4",
          1757 => x"08e80508",
          1758 => x"80e22eb6",
          1759 => x"3882bba4",
          1760 => x"08e80508",
          1761 => x"80f82e84",
          1762 => x"3880cd39",
          1763 => x"900b82bb",
          1764 => x"a408f405",
          1765 => x"3482bba4",
          1766 => x"08880508",
          1767 => x"70088105",
          1768 => x"710c7008",
          1769 => x"51537233",
          1770 => x"82bba408",
          1771 => x"f8053481",
          1772 => x"a439820b",
          1773 => x"82bba408",
          1774 => x"f4053482",
          1775 => x"bba40888",
          1776 => x"05087008",
          1777 => x"8105710c",
          1778 => x"70085153",
          1779 => x"723382bb",
          1780 => x"a408f805",
          1781 => x"3480fe39",
          1782 => x"82bba408",
          1783 => x"f8053353",
          1784 => x"72a0268d",
          1785 => x"38810b82",
          1786 => x"bba408ec",
          1787 => x"050c8380",
          1788 => x"3982bba4",
          1789 => x"08f80533",
          1790 => x"53af7327",
          1791 => x"903882bb",
          1792 => x"a408f805",
          1793 => x"335372b9",
          1794 => x"2683388d",
          1795 => x"39800b82",
          1796 => x"bba408ec",
          1797 => x"050c82d8",
          1798 => x"39880b82",
          1799 => x"bba408f4",
          1800 => x"0534b239",
          1801 => x"82bba408",
          1802 => x"f8053353",
          1803 => x"af732790",
          1804 => x"3882bba4",
          1805 => x"08f80533",
          1806 => x"5372b926",
          1807 => x"83388d39",
          1808 => x"800b82bb",
          1809 => x"a408ec05",
          1810 => x"0c82a539",
          1811 => x"8a0b82bb",
          1812 => x"a408f405",
          1813 => x"34800b82",
          1814 => x"bba408fc",
          1815 => x"050c82bb",
          1816 => x"a408f805",
          1817 => x"3353a073",
          1818 => x"2781cf38",
          1819 => x"82bba408",
          1820 => x"f8053353",
          1821 => x"80e07327",
          1822 => x"943882bb",
          1823 => x"a408f805",
          1824 => x"33e01151",
          1825 => x"537282bb",
          1826 => x"a408f805",
          1827 => x"3482bba4",
          1828 => x"08f80533",
          1829 => x"d0115153",
          1830 => x"7282bba4",
          1831 => x"08f80534",
          1832 => x"82bba408",
          1833 => x"f8053353",
          1834 => x"907327ad",
          1835 => x"3882bba4",
          1836 => x"08f80533",
          1837 => x"f9115153",
          1838 => x"7282bba4",
          1839 => x"08f80534",
          1840 => x"82bba408",
          1841 => x"f8053353",
          1842 => x"7289268d",
          1843 => x"38800b82",
          1844 => x"bba408ec",
          1845 => x"050c8198",
          1846 => x"3982bba4",
          1847 => x"08f80533",
          1848 => x"82bba408",
          1849 => x"f4053354",
          1850 => x"54727426",
          1851 => x"8d38800b",
          1852 => x"82bba408",
          1853 => x"ec050c80",
          1854 => x"f73982bb",
          1855 => x"a408f405",
          1856 => x"337082bb",
          1857 => x"a408fc05",
          1858 => x"082982bb",
          1859 => x"a408f805",
          1860 => x"33701282",
          1861 => x"bba408fc",
          1862 => x"050c82bb",
          1863 => x"a4088805",
          1864 => x"08700881",
          1865 => x"05710c70",
          1866 => x"08515152",
          1867 => x"55537233",
          1868 => x"82bba408",
          1869 => x"f80534fe",
          1870 => x"a53982bb",
          1871 => x"a408f005",
          1872 => x"33537280",
          1873 => x"2e903882",
          1874 => x"bba408fc",
          1875 => x"05083082",
          1876 => x"bba408fc",
          1877 => x"050c82bb",
          1878 => x"a4088c05",
          1879 => x"0882bba4",
          1880 => x"08fc0508",
          1881 => x"710c5381",
          1882 => x"0b82bba4",
          1883 => x"08ec050c",
          1884 => x"82bba408",
          1885 => x"ec050882",
          1886 => x"bb980c8b",
          1887 => x"3d0d82bb",
          1888 => x"a40c0482",
          1889 => x"bba40802",
          1890 => x"82bba40c",
          1891 => x"fb3d0d80",
          1892 => x"0b82bba4",
          1893 => x"08f8050c",
          1894 => x"82d2ec08",
          1895 => x"85113370",
          1896 => x"812a7081",
          1897 => x"32708106",
          1898 => x"51515151",
          1899 => x"5372802e",
          1900 => x"8d38ff0b",
          1901 => x"82bba408",
          1902 => x"f4050c81",
          1903 => x"923982bb",
          1904 => x"a4088805",
          1905 => x"08537233",
          1906 => x"82bba408",
          1907 => x"88050881",
          1908 => x"0582bba4",
          1909 => x"0888050c",
          1910 => x"537282bb",
          1911 => x"a408fc05",
          1912 => x"347281ff",
          1913 => x"06537280",
          1914 => x"2eb03882",
          1915 => x"d2ec0882",
          1916 => x"d2ec0853",
          1917 => x"82bba408",
          1918 => x"fc053352",
          1919 => x"90110851",
          1920 => x"53722d82",
          1921 => x"bb980853",
          1922 => x"72802eff",
          1923 => x"b138ff0b",
          1924 => x"82bba408",
          1925 => x"f8050cff",
          1926 => x"a53982d2",
          1927 => x"ec0882d2",
          1928 => x"ec085353",
          1929 => x"8a519013",
          1930 => x"0853722d",
          1931 => x"82bb9808",
          1932 => x"5372802e",
          1933 => x"8a38ff0b",
          1934 => x"82bba408",
          1935 => x"f8050c82",
          1936 => x"bba408f8",
          1937 => x"05087082",
          1938 => x"bba408f4",
          1939 => x"050c5382",
          1940 => x"bba408f4",
          1941 => x"050882bb",
          1942 => x"980c873d",
          1943 => x"0d82bba4",
          1944 => x"0c0482bb",
          1945 => x"a4080282",
          1946 => x"bba40cfb",
          1947 => x"3d0d800b",
          1948 => x"82bba408",
          1949 => x"f8050c82",
          1950 => x"bba4088c",
          1951 => x"05088511",
          1952 => x"3370812a",
          1953 => x"70813270",
          1954 => x"81065151",
          1955 => x"51515372",
          1956 => x"802e8d38",
          1957 => x"ff0b82bb",
          1958 => x"a408f405",
          1959 => x"0c80f339",
          1960 => x"82bba408",
          1961 => x"88050853",
          1962 => x"723382bb",
          1963 => x"a4088805",
          1964 => x"08810582",
          1965 => x"bba40888",
          1966 => x"050c5372",
          1967 => x"82bba408",
          1968 => x"fc053472",
          1969 => x"81ff0653",
          1970 => x"72802eb6",
          1971 => x"3882bba4",
          1972 => x"088c0508",
          1973 => x"82bba408",
          1974 => x"8c050853",
          1975 => x"82bba408",
          1976 => x"fc053352",
          1977 => x"90110851",
          1978 => x"53722d82",
          1979 => x"bb980853",
          1980 => x"72802eff",
          1981 => x"ab38ff0b",
          1982 => x"82bba408",
          1983 => x"f8050cff",
          1984 => x"9f3982bb",
          1985 => x"a408f805",
          1986 => x"087082bb",
          1987 => x"a408f405",
          1988 => x"0c5382bb",
          1989 => x"a408f405",
          1990 => x"0882bb98",
          1991 => x"0c873d0d",
          1992 => x"82bba40c",
          1993 => x"0482bba4",
          1994 => x"080282bb",
          1995 => x"a40cfe3d",
          1996 => x"0d82d2ec",
          1997 => x"085282bb",
          1998 => x"a4088805",
          1999 => x"0851933f",
          2000 => x"82bb9808",
          2001 => x"7082bb98",
          2002 => x"0c53843d",
          2003 => x"0d82bba4",
          2004 => x"0c0482bb",
          2005 => x"a4080282",
          2006 => x"bba40cfb",
          2007 => x"3d0d82bb",
          2008 => x"a4088c05",
          2009 => x"08851133",
          2010 => x"70812a70",
          2011 => x"81327081",
          2012 => x"06515151",
          2013 => x"51537280",
          2014 => x"2e8d38ff",
          2015 => x"0b82bba4",
          2016 => x"08fc050c",
          2017 => x"81cb3982",
          2018 => x"bba4088c",
          2019 => x"05088511",
          2020 => x"3370822a",
          2021 => x"70810651",
          2022 => x"51515372",
          2023 => x"802e80db",
          2024 => x"3882bba4",
          2025 => x"088c0508",
          2026 => x"82bba408",
          2027 => x"8c050854",
          2028 => x"548c1408",
          2029 => x"88140825",
          2030 => x"9f3882bb",
          2031 => x"a4088c05",
          2032 => x"08700870",
          2033 => x"82bba408",
          2034 => x"88050852",
          2035 => x"57545472",
          2036 => x"75347308",
          2037 => x"8105740c",
          2038 => x"82bba408",
          2039 => x"8c05088c",
          2040 => x"11088105",
          2041 => x"8c120c82",
          2042 => x"bba40888",
          2043 => x"05087082",
          2044 => x"bba408fc",
          2045 => x"050c5153",
          2046 => x"80d73982",
          2047 => x"bba4088c",
          2048 => x"050882bb",
          2049 => x"a4088c05",
          2050 => x"085382bb",
          2051 => x"a4088805",
          2052 => x"087081ff",
          2053 => x"06539012",
          2054 => x"08515454",
          2055 => x"722d82bb",
          2056 => x"98085372",
          2057 => x"a33882bb",
          2058 => x"a4088c05",
          2059 => x"088c1108",
          2060 => x"81058c12",
          2061 => x"0c82bba4",
          2062 => x"08880508",
          2063 => x"7082bba4",
          2064 => x"08fc050c",
          2065 => x"51538a39",
          2066 => x"ff0b82bb",
          2067 => x"a408fc05",
          2068 => x"0c82bba4",
          2069 => x"08fc0508",
          2070 => x"82bb980c",
          2071 => x"873d0d82",
          2072 => x"bba40c04",
          2073 => x"82bba408",
          2074 => x"0282bba4",
          2075 => x"0cf93d0d",
          2076 => x"82bba408",
          2077 => x"88050885",
          2078 => x"11337081",
          2079 => x"32708106",
          2080 => x"51515152",
          2081 => x"71802e8d",
          2082 => x"38ff0b82",
          2083 => x"bba408f8",
          2084 => x"050c8394",
          2085 => x"3982bba4",
          2086 => x"08880508",
          2087 => x"85113370",
          2088 => x"862a7081",
          2089 => x"06515151",
          2090 => x"5271802e",
          2091 => x"80c53882",
          2092 => x"bba40888",
          2093 => x"050882bb",
          2094 => x"a4088805",
          2095 => x"08535385",
          2096 => x"123370ff",
          2097 => x"bf065152",
          2098 => x"71851434",
          2099 => x"82bba408",
          2100 => x"8805088c",
          2101 => x"11088105",
          2102 => x"8c120c82",
          2103 => x"bba40888",
          2104 => x"05088411",
          2105 => x"337082bb",
          2106 => x"a408f805",
          2107 => x"0c515152",
          2108 => x"82b63982",
          2109 => x"bba40888",
          2110 => x"05088511",
          2111 => x"3370822a",
          2112 => x"70810651",
          2113 => x"51515271",
          2114 => x"802e80d7",
          2115 => x"3882bba4",
          2116 => x"08880508",
          2117 => x"70087033",
          2118 => x"82bba408",
          2119 => x"fc050c51",
          2120 => x"5282bba4",
          2121 => x"08fc0508",
          2122 => x"a93882bb",
          2123 => x"a4088805",
          2124 => x"0882bba4",
          2125 => x"08880508",
          2126 => x"53538512",
          2127 => x"3370a007",
          2128 => x"51527185",
          2129 => x"1434ff0b",
          2130 => x"82bba408",
          2131 => x"f8050c81",
          2132 => x"d73982bb",
          2133 => x"a4088805",
          2134 => x"08700881",
          2135 => x"05710c52",
          2136 => x"81a13982",
          2137 => x"bba40888",
          2138 => x"050882bb",
          2139 => x"a4088805",
          2140 => x"08529411",
          2141 => x"08515271",
          2142 => x"2d82bb98",
          2143 => x"087082bb",
          2144 => x"a408fc05",
          2145 => x"0c5282bb",
          2146 => x"a408fc05",
          2147 => x"08802580",
          2148 => x"f23882bb",
          2149 => x"a4088805",
          2150 => x"0882bba4",
          2151 => x"08f4050c",
          2152 => x"82bba408",
          2153 => x"88050885",
          2154 => x"113382bb",
          2155 => x"a408f005",
          2156 => x"0c5282bb",
          2157 => x"a408fc05",
          2158 => x"08ff2e09",
          2159 => x"81069538",
          2160 => x"82bba408",
          2161 => x"f0050890",
          2162 => x"07527182",
          2163 => x"bba408ec",
          2164 => x"05349339",
          2165 => x"82bba408",
          2166 => x"f00508a0",
          2167 => x"07527182",
          2168 => x"bba408ec",
          2169 => x"053482bb",
          2170 => x"a408f405",
          2171 => x"085282bb",
          2172 => x"a408ec05",
          2173 => x"33851334",
          2174 => x"ff0b82bb",
          2175 => x"a408f805",
          2176 => x"0ca63982",
          2177 => x"bba40888",
          2178 => x"05088c11",
          2179 => x"0881058c",
          2180 => x"120c82bb",
          2181 => x"a408fc05",
          2182 => x"087081ff",
          2183 => x"067082bb",
          2184 => x"a408f805",
          2185 => x"0c515152",
          2186 => x"82bba408",
          2187 => x"f8050882",
          2188 => x"bb980c89",
          2189 => x"3d0d82bb",
          2190 => x"a40c0482",
          2191 => x"bba40802",
          2192 => x"82bba40c",
          2193 => x"fd3d0d82",
          2194 => x"bba40888",
          2195 => x"050882bb",
          2196 => x"a408fc05",
          2197 => x"0c82bba4",
          2198 => x"088c0508",
          2199 => x"82bba408",
          2200 => x"f8050c82",
          2201 => x"bba40890",
          2202 => x"0508802e",
          2203 => x"82a23882",
          2204 => x"bba408f8",
          2205 => x"050882bb",
          2206 => x"a408fc05",
          2207 => x"082681ac",
          2208 => x"3882bba4",
          2209 => x"08f80508",
          2210 => x"82bba408",
          2211 => x"90050805",
          2212 => x"5182bba4",
          2213 => x"08fc0508",
          2214 => x"71278190",
          2215 => x"3882bba4",
          2216 => x"08fc0508",
          2217 => x"82bba408",
          2218 => x"90050805",
          2219 => x"82bba408",
          2220 => x"fc050c82",
          2221 => x"bba408f8",
          2222 => x"050882bb",
          2223 => x"a4089005",
          2224 => x"080582bb",
          2225 => x"a408f805",
          2226 => x"0c82bba4",
          2227 => x"08900508",
          2228 => x"810582bb",
          2229 => x"a4089005",
          2230 => x"0c82bba4",
          2231 => x"08900508",
          2232 => x"ff0582bb",
          2233 => x"a4089005",
          2234 => x"0c82bba4",
          2235 => x"08900508",
          2236 => x"802e819c",
          2237 => x"3882bba4",
          2238 => x"08fc0508",
          2239 => x"ff0582bb",
          2240 => x"a408fc05",
          2241 => x"0c82bba4",
          2242 => x"08f80508",
          2243 => x"ff0582bb",
          2244 => x"a408f805",
          2245 => x"0c82bba4",
          2246 => x"08fc0508",
          2247 => x"82bba408",
          2248 => x"f8050853",
          2249 => x"51713371",
          2250 => x"34ffae39",
          2251 => x"82bba408",
          2252 => x"90050881",
          2253 => x"0582bba4",
          2254 => x"0890050c",
          2255 => x"82bba408",
          2256 => x"900508ff",
          2257 => x"0582bba4",
          2258 => x"0890050c",
          2259 => x"82bba408",
          2260 => x"90050880",
          2261 => x"2eba3882",
          2262 => x"bba408f8",
          2263 => x"05085170",
          2264 => x"3382bba4",
          2265 => x"08f80508",
          2266 => x"810582bb",
          2267 => x"a408f805",
          2268 => x"0c82bba4",
          2269 => x"08fc0508",
          2270 => x"52527171",
          2271 => x"3482bba4",
          2272 => x"08fc0508",
          2273 => x"810582bb",
          2274 => x"a408fc05",
          2275 => x"0cffad39",
          2276 => x"82bba408",
          2277 => x"88050870",
          2278 => x"82bb980c",
          2279 => x"51853d0d",
          2280 => x"82bba40c",
          2281 => x"0482bba4",
          2282 => x"080282bb",
          2283 => x"a40cfe3d",
          2284 => x"0d82bba4",
          2285 => x"08880508",
          2286 => x"82bba408",
          2287 => x"fc050c82",
          2288 => x"bba408fc",
          2289 => x"05085271",
          2290 => x"3382bba4",
          2291 => x"08fc0508",
          2292 => x"810582bb",
          2293 => x"a408fc05",
          2294 => x"0c7081ff",
          2295 => x"06515170",
          2296 => x"802e8338",
          2297 => x"da3982bb",
          2298 => x"a408fc05",
          2299 => x"08ff0582",
          2300 => x"bba408fc",
          2301 => x"050c82bb",
          2302 => x"a408fc05",
          2303 => x"0882bba4",
          2304 => x"08880508",
          2305 => x"317082bb",
          2306 => x"980c5184",
          2307 => x"3d0d82bb",
          2308 => x"a40c0482",
          2309 => x"bba40802",
          2310 => x"82bba40c",
          2311 => x"fe3d0d82",
          2312 => x"bba40888",
          2313 => x"050882bb",
          2314 => x"a408fc05",
          2315 => x"0c82bba4",
          2316 => x"088c0508",
          2317 => x"52713382",
          2318 => x"bba4088c",
          2319 => x"05088105",
          2320 => x"82bba408",
          2321 => x"8c050c82",
          2322 => x"bba408fc",
          2323 => x"05085351",
          2324 => x"70723482",
          2325 => x"bba408fc",
          2326 => x"05088105",
          2327 => x"82bba408",
          2328 => x"fc050c70",
          2329 => x"81ff0651",
          2330 => x"70802e84",
          2331 => x"38ffbe39",
          2332 => x"82bba408",
          2333 => x"88050870",
          2334 => x"82bb980c",
          2335 => x"51843d0d",
          2336 => x"82bba40c",
          2337 => x"0482bba4",
          2338 => x"080282bb",
          2339 => x"a40cfd3d",
          2340 => x"0d82bba4",
          2341 => x"08880508",
          2342 => x"82bba408",
          2343 => x"fc050c82",
          2344 => x"bba4088c",
          2345 => x"050882bb",
          2346 => x"a408f805",
          2347 => x"0c82bba4",
          2348 => x"08900508",
          2349 => x"802e80e5",
          2350 => x"3882bba4",
          2351 => x"08900508",
          2352 => x"810582bb",
          2353 => x"a4089005",
          2354 => x"0c82bba4",
          2355 => x"08900508",
          2356 => x"ff0582bb",
          2357 => x"a4089005",
          2358 => x"0c82bba4",
          2359 => x"08900508",
          2360 => x"802eba38",
          2361 => x"82bba408",
          2362 => x"f8050851",
          2363 => x"703382bb",
          2364 => x"a408f805",
          2365 => x"08810582",
          2366 => x"bba408f8",
          2367 => x"050c82bb",
          2368 => x"a408fc05",
          2369 => x"08525271",
          2370 => x"713482bb",
          2371 => x"a408fc05",
          2372 => x"08810582",
          2373 => x"bba408fc",
          2374 => x"050cffad",
          2375 => x"3982bba4",
          2376 => x"08880508",
          2377 => x"7082bb98",
          2378 => x"0c51853d",
          2379 => x"0d82bba4",
          2380 => x"0c0482bb",
          2381 => x"a4080282",
          2382 => x"bba40cfd",
          2383 => x"3d0d82bb",
          2384 => x"a4089005",
          2385 => x"08802e81",
          2386 => x"f43882bb",
          2387 => x"a4088c05",
          2388 => x"08527133",
          2389 => x"82bba408",
          2390 => x"8c050881",
          2391 => x"0582bba4",
          2392 => x"088c050c",
          2393 => x"82bba408",
          2394 => x"88050870",
          2395 => x"337281ff",
          2396 => x"06535454",
          2397 => x"5171712e",
          2398 => x"843880ce",
          2399 => x"3982bba4",
          2400 => x"08880508",
          2401 => x"52713382",
          2402 => x"bba40888",
          2403 => x"05088105",
          2404 => x"82bba408",
          2405 => x"88050c70",
          2406 => x"81ff0651",
          2407 => x"51708d38",
          2408 => x"800b82bb",
          2409 => x"a408fc05",
          2410 => x"0c819b39",
          2411 => x"82bba408",
          2412 => x"900508ff",
          2413 => x"0582bba4",
          2414 => x"0890050c",
          2415 => x"82bba408",
          2416 => x"90050880",
          2417 => x"2e8438ff",
          2418 => x"813982bb",
          2419 => x"a4089005",
          2420 => x"08802e80",
          2421 => x"e83882bb",
          2422 => x"a4088805",
          2423 => x"08703352",
          2424 => x"53708d38",
          2425 => x"ff0b82bb",
          2426 => x"a408fc05",
          2427 => x"0c80d739",
          2428 => x"82bba408",
          2429 => x"8c0508ff",
          2430 => x"0582bba4",
          2431 => x"088c050c",
          2432 => x"82bba408",
          2433 => x"8c050870",
          2434 => x"33525270",
          2435 => x"8c38810b",
          2436 => x"82bba408",
          2437 => x"fc050cae",
          2438 => x"3982bba4",
          2439 => x"08880508",
          2440 => x"703382bb",
          2441 => x"a4088c05",
          2442 => x"08703372",
          2443 => x"71317082",
          2444 => x"bba408fc",
          2445 => x"050c5355",
          2446 => x"5252538a",
          2447 => x"39800b82",
          2448 => x"bba408fc",
          2449 => x"050c82bb",
          2450 => x"a408fc05",
          2451 => x"0882bb98",
          2452 => x"0c853d0d",
          2453 => x"82bba40c",
          2454 => x"0482bba4",
          2455 => x"080282bb",
          2456 => x"a40cfd3d",
          2457 => x"0d82bba4",
          2458 => x"08880508",
          2459 => x"82bba408",
          2460 => x"f8050c82",
          2461 => x"bba4088c",
          2462 => x"05088d38",
          2463 => x"800b82bb",
          2464 => x"a408fc05",
          2465 => x"0c80ec39",
          2466 => x"82bba408",
          2467 => x"f8050852",
          2468 => x"713382bb",
          2469 => x"a408f805",
          2470 => x"08810582",
          2471 => x"bba408f8",
          2472 => x"050c7081",
          2473 => x"ff065151",
          2474 => x"70802e9f",
          2475 => x"3882bba4",
          2476 => x"088c0508",
          2477 => x"ff0582bb",
          2478 => x"a4088c05",
          2479 => x"0c82bba4",
          2480 => x"088c0508",
          2481 => x"ff2e8438",
          2482 => x"ffbe3982",
          2483 => x"bba408f8",
          2484 => x"0508ff05",
          2485 => x"82bba408",
          2486 => x"f8050c82",
          2487 => x"bba408f8",
          2488 => x"050882bb",
          2489 => x"a4088805",
          2490 => x"08317082",
          2491 => x"bba408fc",
          2492 => x"050c5182",
          2493 => x"bba408fc",
          2494 => x"050882bb",
          2495 => x"980c853d",
          2496 => x"0d82bba4",
          2497 => x"0c0482bb",
          2498 => x"a4080282",
          2499 => x"bba40cfe",
          2500 => x"3d0d82bb",
          2501 => x"a4088805",
          2502 => x"0882bba4",
          2503 => x"08fc050c",
          2504 => x"82bba408",
          2505 => x"90050880",
          2506 => x"2e80d438",
          2507 => x"82bba408",
          2508 => x"90050881",
          2509 => x"0582bba4",
          2510 => x"0890050c",
          2511 => x"82bba408",
          2512 => x"900508ff",
          2513 => x"0582bba4",
          2514 => x"0890050c",
          2515 => x"82bba408",
          2516 => x"90050880",
          2517 => x"2ea93882",
          2518 => x"bba4088c",
          2519 => x"05085170",
          2520 => x"82bba408",
          2521 => x"fc050852",
          2522 => x"52717134",
          2523 => x"82bba408",
          2524 => x"fc050881",
          2525 => x"0582bba4",
          2526 => x"08fc050c",
          2527 => x"ffbe3982",
          2528 => x"bba40888",
          2529 => x"05087082",
          2530 => x"bb980c51",
          2531 => x"843d0d82",
          2532 => x"bba40c04",
          2533 => x"82bba408",
          2534 => x"0282bba4",
          2535 => x"0cf93d0d",
          2536 => x"800b82bb",
          2537 => x"a408fc05",
          2538 => x"0c82bba4",
          2539 => x"08880508",
          2540 => x"8025b938",
          2541 => x"82bba408",
          2542 => x"88050830",
          2543 => x"82bba408",
          2544 => x"88050c80",
          2545 => x"0b82bba4",
          2546 => x"08f4050c",
          2547 => x"82bba408",
          2548 => x"fc05088a",
          2549 => x"38810b82",
          2550 => x"bba408f4",
          2551 => x"050c82bb",
          2552 => x"a408f405",
          2553 => x"0882bba4",
          2554 => x"08fc050c",
          2555 => x"82bba408",
          2556 => x"8c050880",
          2557 => x"25b93882",
          2558 => x"bba4088c",
          2559 => x"05083082",
          2560 => x"bba4088c",
          2561 => x"050c800b",
          2562 => x"82bba408",
          2563 => x"f0050c82",
          2564 => x"bba408fc",
          2565 => x"05088a38",
          2566 => x"810b82bb",
          2567 => x"a408f005",
          2568 => x"0c82bba4",
          2569 => x"08f00508",
          2570 => x"82bba408",
          2571 => x"fc050c80",
          2572 => x"5382bba4",
          2573 => x"088c0508",
          2574 => x"5282bba4",
          2575 => x"08880508",
          2576 => x"5182c53f",
          2577 => x"82bb9808",
          2578 => x"7082bba4",
          2579 => x"08f8050c",
          2580 => x"5482bba4",
          2581 => x"08fc0508",
          2582 => x"802e9038",
          2583 => x"82bba408",
          2584 => x"f8050830",
          2585 => x"82bba408",
          2586 => x"f8050c82",
          2587 => x"bba408f8",
          2588 => x"05087082",
          2589 => x"bb980c54",
          2590 => x"893d0d82",
          2591 => x"bba40c04",
          2592 => x"82bba408",
          2593 => x"0282bba4",
          2594 => x"0cfb3d0d",
          2595 => x"800b82bb",
          2596 => x"a408fc05",
          2597 => x"0c82bba4",
          2598 => x"08880508",
          2599 => x"80259938",
          2600 => x"82bba408",
          2601 => x"88050830",
          2602 => x"82bba408",
          2603 => x"88050c81",
          2604 => x"0b82bba4",
          2605 => x"08fc050c",
          2606 => x"82bba408",
          2607 => x"8c050880",
          2608 => x"25903882",
          2609 => x"bba4088c",
          2610 => x"05083082",
          2611 => x"bba4088c",
          2612 => x"050c8153",
          2613 => x"82bba408",
          2614 => x"8c050852",
          2615 => x"82bba408",
          2616 => x"88050851",
          2617 => x"81a23f82",
          2618 => x"bb980870",
          2619 => x"82bba408",
          2620 => x"f8050c54",
          2621 => x"82bba408",
          2622 => x"fc050880",
          2623 => x"2e903882",
          2624 => x"bba408f8",
          2625 => x"05083082",
          2626 => x"bba408f8",
          2627 => x"050c82bb",
          2628 => x"a408f805",
          2629 => x"087082bb",
          2630 => x"980c5487",
          2631 => x"3d0d82bb",
          2632 => x"a40c0482",
          2633 => x"bba40802",
          2634 => x"82bba40c",
          2635 => x"fd3d0d80",
          2636 => x"5382bba4",
          2637 => x"088c0508",
          2638 => x"5282bba4",
          2639 => x"08880508",
          2640 => x"5180c53f",
          2641 => x"82bb9808",
          2642 => x"7082bb98",
          2643 => x"0c54853d",
          2644 => x"0d82bba4",
          2645 => x"0c0482bb",
          2646 => x"a4080282",
          2647 => x"bba40cfd",
          2648 => x"3d0d8153",
          2649 => x"82bba408",
          2650 => x"8c050852",
          2651 => x"82bba408",
          2652 => x"88050851",
          2653 => x"933f82bb",
          2654 => x"98087082",
          2655 => x"bb980c54",
          2656 => x"853d0d82",
          2657 => x"bba40c04",
          2658 => x"82bba408",
          2659 => x"0282bba4",
          2660 => x"0cfd3d0d",
          2661 => x"810b82bb",
          2662 => x"a408fc05",
          2663 => x"0c800b82",
          2664 => x"bba408f8",
          2665 => x"050c82bb",
          2666 => x"a4088c05",
          2667 => x"0882bba4",
          2668 => x"08880508",
          2669 => x"27b93882",
          2670 => x"bba408fc",
          2671 => x"0508802e",
          2672 => x"ae38800b",
          2673 => x"82bba408",
          2674 => x"8c050824",
          2675 => x"a23882bb",
          2676 => x"a4088c05",
          2677 => x"081082bb",
          2678 => x"a4088c05",
          2679 => x"0c82bba4",
          2680 => x"08fc0508",
          2681 => x"1082bba4",
          2682 => x"08fc050c",
          2683 => x"ffb83982",
          2684 => x"bba408fc",
          2685 => x"0508802e",
          2686 => x"80e13882",
          2687 => x"bba4088c",
          2688 => x"050882bb",
          2689 => x"a4088805",
          2690 => x"0826ad38",
          2691 => x"82bba408",
          2692 => x"88050882",
          2693 => x"bba4088c",
          2694 => x"05083182",
          2695 => x"bba40888",
          2696 => x"050c82bb",
          2697 => x"a408f805",
          2698 => x"0882bba4",
          2699 => x"08fc0508",
          2700 => x"0782bba4",
          2701 => x"08f8050c",
          2702 => x"82bba408",
          2703 => x"fc050881",
          2704 => x"2a82bba4",
          2705 => x"08fc050c",
          2706 => x"82bba408",
          2707 => x"8c050881",
          2708 => x"2a82bba4",
          2709 => x"088c050c",
          2710 => x"ff953982",
          2711 => x"bba40890",
          2712 => x"0508802e",
          2713 => x"933882bb",
          2714 => x"a4088805",
          2715 => x"087082bb",
          2716 => x"a408f405",
          2717 => x"0c519139",
          2718 => x"82bba408",
          2719 => x"f8050870",
          2720 => x"82bba408",
          2721 => x"f4050c51",
          2722 => x"82bba408",
          2723 => x"f4050882",
          2724 => x"bb980c85",
          2725 => x"3d0d82bb",
          2726 => x"a40c04f9",
          2727 => x"3d0d7970",
          2728 => x"08705656",
          2729 => x"5874802e",
          2730 => x"80e33895",
          2731 => x"39750851",
          2732 => x"f1f33f82",
          2733 => x"bb980815",
          2734 => x"780c8516",
          2735 => x"335480cd",
          2736 => x"39743354",
          2737 => x"73a02e09",
          2738 => x"81068638",
          2739 => x"811555f1",
          2740 => x"39805776",
          2741 => x"902982b6",
          2742 => x"98057008",
          2743 => x"5256f1c5",
          2744 => x"3f82bb98",
          2745 => x"08537452",
          2746 => x"750851f4",
          2747 => x"c53f82bb",
          2748 => x"98088b38",
          2749 => x"84163354",
          2750 => x"73812eff",
          2751 => x"b0388117",
          2752 => x"7081ff06",
          2753 => x"58549977",
          2754 => x"27c938ff",
          2755 => x"547382bb",
          2756 => x"980c893d",
          2757 => x"0d04ff3d",
          2758 => x"0d735271",
          2759 => x"9326818e",
          2760 => x"38718429",
          2761 => x"8299b005",
          2762 => x"52710804",
          2763 => x"829efc51",
          2764 => x"81803982",
          2765 => x"9f885180",
          2766 => x"f939829f",
          2767 => x"9c5180f2",
          2768 => x"39829fb0",
          2769 => x"5180eb39",
          2770 => x"829fc051",
          2771 => x"80e43982",
          2772 => x"9fd05180",
          2773 => x"dd39829f",
          2774 => x"e45180d6",
          2775 => x"39829ff4",
          2776 => x"5180cf39",
          2777 => x"82a08c51",
          2778 => x"80c83982",
          2779 => x"a0a45180",
          2780 => x"c13982a0",
          2781 => x"bc51bb39",
          2782 => x"82a0d851",
          2783 => x"b53982a0",
          2784 => x"ec51af39",
          2785 => x"82a19851",
          2786 => x"a93982a1",
          2787 => x"ac51a339",
          2788 => x"82a1cc51",
          2789 => x"9d3982a1",
          2790 => x"e0519739",
          2791 => x"82a1f851",
          2792 => x"913982a2",
          2793 => x"90518b39",
          2794 => x"82a2a851",
          2795 => x"853982a2",
          2796 => x"b451e3cf",
          2797 => x"3f833d0d",
          2798 => x"04fb3d0d",
          2799 => x"77795656",
          2800 => x"7487e726",
          2801 => x"8a387452",
          2802 => x"7587e829",
          2803 => x"51903987",
          2804 => x"e8527451",
          2805 => x"facd3f82",
          2806 => x"bb980852",
          2807 => x"7551fac3",
          2808 => x"3f82bb98",
          2809 => x"08547953",
          2810 => x"755282a2",
          2811 => x"c451ffbb",
          2812 => x"e53f873d",
          2813 => x"0d04ec3d",
          2814 => x"0d660284",
          2815 => x"0580e305",
          2816 => x"335b5780",
          2817 => x"68783070",
          2818 => x"7a077325",
          2819 => x"51575959",
          2820 => x"78567787",
          2821 => x"ff268338",
          2822 => x"81567476",
          2823 => x"077081ff",
          2824 => x"06515593",
          2825 => x"56748182",
          2826 => x"38815376",
          2827 => x"528c3d70",
          2828 => x"52568183",
          2829 => x"cf3f82bb",
          2830 => x"98085782",
          2831 => x"bb9808b9",
          2832 => x"3882bb98",
          2833 => x"0887c098",
          2834 => x"880c82bb",
          2835 => x"98085996",
          2836 => x"3dd40554",
          2837 => x"84805377",
          2838 => x"52755181",
          2839 => x"888b3f82",
          2840 => x"bb980857",
          2841 => x"82bb9808",
          2842 => x"90387a55",
          2843 => x"74802e89",
          2844 => x"38741975",
          2845 => x"195959d7",
          2846 => x"39963dd8",
          2847 => x"0551818f",
          2848 => x"f43f7630",
          2849 => x"70780780",
          2850 => x"257b3070",
          2851 => x"9f2a7206",
          2852 => x"51575156",
          2853 => x"74802e90",
          2854 => x"3882a2e8",
          2855 => x"5387c098",
          2856 => x"88085278",
          2857 => x"51fe923f",
          2858 => x"76567582",
          2859 => x"bb980c96",
          2860 => x"3d0d04f8",
          2861 => x"3d0d7c02",
          2862 => x"8405b705",
          2863 => x"335859ff",
          2864 => x"5880537b",
          2865 => x"527a51fe",
          2866 => x"ad3f82bb",
          2867 => x"9808a638",
          2868 => x"76802e88",
          2869 => x"3876812e",
          2870 => x"9a389a39",
          2871 => x"62566155",
          2872 => x"605482bb",
          2873 => x"98537f52",
          2874 => x"7e51782d",
          2875 => x"82bb9808",
          2876 => x"58833978",
          2877 => x"047782bb",
          2878 => x"980c8a3d",
          2879 => x"0d04f33d",
          2880 => x"0d7f6163",
          2881 => x"028c0580",
          2882 => x"cf053373",
          2883 => x"73156841",
          2884 => x"5f5c5c5e",
          2885 => x"5e5e7a52",
          2886 => x"82a2f051",
          2887 => x"ffb9b73f",
          2888 => x"82a2f851",
          2889 => x"e0dd3f80",
          2890 => x"55747927",
          2891 => x"80fd387b",
          2892 => x"902e8938",
          2893 => x"7ba02ea6",
          2894 => x"3880c439",
          2895 => x"74185372",
          2896 => x"7a278e38",
          2897 => x"72225282",
          2898 => x"a2fc51ff",
          2899 => x"b9883f88",
          2900 => x"3982a388",
          2901 => x"51e0ac3f",
          2902 => x"82155580",
          2903 => x"c1397418",
          2904 => x"53727a27",
          2905 => x"8e387208",
          2906 => x"5282a2f0",
          2907 => x"51ffb8e6",
          2908 => x"3f883982",
          2909 => x"a38451e0",
          2910 => x"8a3f8415",
          2911 => x"55a03974",
          2912 => x"1853727a",
          2913 => x"278e3872",
          2914 => x"335282a3",
          2915 => x"9051ffb8",
          2916 => x"c53f8839",
          2917 => x"82a39851",
          2918 => x"dfe93f81",
          2919 => x"155582d2",
          2920 => x"ec0852a0",
          2921 => x"51e3ab3f",
          2922 => x"feff3982",
          2923 => x"a39c51df",
          2924 => x"d23f8055",
          2925 => x"74792780",
          2926 => x"c6387418",
          2927 => x"70335553",
          2928 => x"8056727a",
          2929 => x"27833881",
          2930 => x"5680539f",
          2931 => x"74278338",
          2932 => x"81537573",
          2933 => x"067081ff",
          2934 => x"06515372",
          2935 => x"802e9038",
          2936 => x"7380fe26",
          2937 => x"8a3882d2",
          2938 => x"ec085273",
          2939 => x"51883982",
          2940 => x"d2ec0852",
          2941 => x"a051e2da",
          2942 => x"3f811555",
          2943 => x"ffb63982",
          2944 => x"a3a051de",
          2945 => x"fe3f7818",
          2946 => x"791c5c58",
          2947 => x"a0ef3f82",
          2948 => x"bb980898",
          2949 => x"2b70982c",
          2950 => x"515776a0",
          2951 => x"2e098106",
          2952 => x"aa38a0d9",
          2953 => x"3f82bb98",
          2954 => x"08982b70",
          2955 => x"982c70a0",
          2956 => x"32703072",
          2957 => x"9b327030",
          2958 => x"70720773",
          2959 => x"75070651",
          2960 => x"58585957",
          2961 => x"51578073",
          2962 => x"24d83876",
          2963 => x"9b2e0981",
          2964 => x"06853880",
          2965 => x"538c397c",
          2966 => x"1e537278",
          2967 => x"26fdb738",
          2968 => x"ff537282",
          2969 => x"bb980c8f",
          2970 => x"3d0d04fc",
          2971 => x"3d0d029b",
          2972 => x"053382a3",
          2973 => x"a45382a3",
          2974 => x"ac5255ff",
          2975 => x"b6d83f82",
          2976 => x"b9f02251",
          2977 => x"a9ca3f82",
          2978 => x"a3b85482",
          2979 => x"a3c45382",
          2980 => x"b9f13352",
          2981 => x"82a3cc51",
          2982 => x"ffb6bb3f",
          2983 => x"74802e84",
          2984 => x"38a4fc3f",
          2985 => x"863d0d04",
          2986 => x"fe3d0d87",
          2987 => x"c0968008",
          2988 => x"53aaa73f",
          2989 => x"81519cb2",
          2990 => x"3f82a3e8",
          2991 => x"519dc73f",
          2992 => x"80519ca6",
          2993 => x"3f72812a",
          2994 => x"70810651",
          2995 => x"5271802e",
          2996 => x"92388151",
          2997 => x"9c943f82",
          2998 => x"a484519d",
          2999 => x"a93f8051",
          3000 => x"9c883f72",
          3001 => x"822a7081",
          3002 => x"06515271",
          3003 => x"802e9238",
          3004 => x"81519bf6",
          3005 => x"3f82a498",
          3006 => x"519d8b3f",
          3007 => x"80519bea",
          3008 => x"3f72832a",
          3009 => x"70810651",
          3010 => x"5271802e",
          3011 => x"92388151",
          3012 => x"9bd83f82",
          3013 => x"a4a8519c",
          3014 => x"ed3f8051",
          3015 => x"9bcc3f72",
          3016 => x"842a7081",
          3017 => x"06515271",
          3018 => x"802e9238",
          3019 => x"81519bba",
          3020 => x"3f82a4bc",
          3021 => x"519ccf3f",
          3022 => x"80519bae",
          3023 => x"3f72852a",
          3024 => x"70810651",
          3025 => x"5271802e",
          3026 => x"92388151",
          3027 => x"9b9c3f82",
          3028 => x"a4d0519c",
          3029 => x"b13f8051",
          3030 => x"9b903f72",
          3031 => x"862a7081",
          3032 => x"06515271",
          3033 => x"802e9238",
          3034 => x"81519afe",
          3035 => x"3f82a4e4",
          3036 => x"519c933f",
          3037 => x"80519af2",
          3038 => x"3f72872a",
          3039 => x"70810651",
          3040 => x"5271802e",
          3041 => x"92388151",
          3042 => x"9ae03f82",
          3043 => x"a4f8519b",
          3044 => x"f53f8051",
          3045 => x"9ad43f72",
          3046 => x"882a7081",
          3047 => x"06515271",
          3048 => x"802e9238",
          3049 => x"81519ac2",
          3050 => x"3f82a58c",
          3051 => x"519bd73f",
          3052 => x"80519ab6",
          3053 => x"3fa8ab3f",
          3054 => x"843d0d04",
          3055 => x"fb3d0d77",
          3056 => x"028405a3",
          3057 => x"05337055",
          3058 => x"56568052",
          3059 => x"7551eeb6",
          3060 => x"3f0b0b82",
          3061 => x"b6943354",
          3062 => x"73a93881",
          3063 => x"5382a5cc",
          3064 => x"5282d298",
          3065 => x"5180fc9c",
          3066 => x"3f82bb98",
          3067 => x"08307082",
          3068 => x"bb980807",
          3069 => x"80258271",
          3070 => x"31515154",
          3071 => x"730b0b82",
          3072 => x"b694340b",
          3073 => x"0b82b694",
          3074 => x"33547381",
          3075 => x"2e098106",
          3076 => x"af3882d2",
          3077 => x"98537452",
          3078 => x"755181b6",
          3079 => x"cd3f82bb",
          3080 => x"9808802e",
          3081 => x"8b3882bb",
          3082 => x"980851da",
          3083 => x"d63f9139",
          3084 => x"82d29851",
          3085 => x"8188be3f",
          3086 => x"820b0b0b",
          3087 => x"82b69434",
          3088 => x"0b0b82b6",
          3089 => x"94335473",
          3090 => x"822e0981",
          3091 => x"068c3882",
          3092 => x"a5dc5374",
          3093 => x"527551ae",
          3094 => x"953f800b",
          3095 => x"82bb980c",
          3096 => x"873d0d04",
          3097 => x"cd3d0d80",
          3098 => x"707182d2",
          3099 => x"940c405e",
          3100 => x"81527d51",
          3101 => x"80cae83f",
          3102 => x"82bb9808",
          3103 => x"81ff065a",
          3104 => x"797e2e09",
          3105 => x"8106a338",
          3106 => x"973d5a83",
          3107 => x"5382a5e8",
          3108 => x"527951e7",
          3109 => x"f03f7d53",
          3110 => x"795282bc",
          3111 => x"c45180fa",
          3112 => x"823f82bb",
          3113 => x"98087e2e",
          3114 => x"883882a5",
          3115 => x"ec5191c8",
          3116 => x"39817040",
          3117 => x"5e82a6a4",
          3118 => x"51d9c83f",
          3119 => x"973d7047",
          3120 => x"5b80f852",
          3121 => x"7a51fdf4",
          3122 => x"3fb53dff",
          3123 => x"840551f3",
          3124 => x"ca3f82bb",
          3125 => x"9808902b",
          3126 => x"70902c51",
          3127 => x"5a7980c1",
          3128 => x"2e89d438",
          3129 => x"7980c124",
          3130 => x"80d93879",
          3131 => x"ab2e83b9",
          3132 => x"3879ab24",
          3133 => x"a4387982",
          3134 => x"2e81b338",
          3135 => x"7982248a",
          3136 => x"3879802e",
          3137 => x"ffaf388e",
          3138 => x"ed397984",
          3139 => x"2e828338",
          3140 => x"79942e82",
          3141 => x"ad388ede",
          3142 => x"3979bd2e",
          3143 => x"84ff3879",
          3144 => x"bd249038",
          3145 => x"79b02e83",
          3146 => x"a63879bc",
          3147 => x"2e848838",
          3148 => x"8ec43979",
          3149 => x"bf2e85c6",
          3150 => x"387980c0",
          3151 => x"2e86bd38",
          3152 => x"8eb43979",
          3153 => x"80d52e8d",
          3154 => x"90387980",
          3155 => x"d524b038",
          3156 => x"7980d02e",
          3157 => x"8cc93879",
          3158 => x"80d02492",
          3159 => x"387980c2",
          3160 => x"2e89f638",
          3161 => x"7980c32e",
          3162 => x"8b9b388e",
          3163 => x"89397980",
          3164 => x"d12e8cba",
          3165 => x"387980d4",
          3166 => x"2e8cc238",
          3167 => x"8df83979",
          3168 => x"81822e8d",
          3169 => x"d1387981",
          3170 => x"82249238",
          3171 => x"7980f82e",
          3172 => x"8ce33879",
          3173 => x"80f92e8d",
          3174 => x"80388dda",
          3175 => x"39798183",
          3176 => x"2e8dc138",
          3177 => x"7981852e",
          3178 => x"8dc6388d",
          3179 => x"c939b53d",
          3180 => x"ff801153",
          3181 => x"ff840551",
          3182 => x"d1f83f82",
          3183 => x"bb980888",
          3184 => x"3882a6a8",
          3185 => x"518fb139",
          3186 => x"b53dfefc",
          3187 => x"1153ff84",
          3188 => x"0551d1de",
          3189 => x"3f82bb98",
          3190 => x"08802e88",
          3191 => x"38816425",
          3192 => x"83388044",
          3193 => x"0280cf05",
          3194 => x"33520280",
          3195 => x"d3053351",
          3196 => x"80c7ec3f",
          3197 => x"82bb9808",
          3198 => x"81ff065a",
          3199 => x"798d3882",
          3200 => x"a6b851d6",
          3201 => x"fe3f815f",
          3202 => x"fdab3982",
          3203 => x"a6c8518e",
          3204 => x"e739b53d",
          3205 => x"ff801153",
          3206 => x"ff840551",
          3207 => x"d1943f82",
          3208 => x"bb980880",
          3209 => x"2efd8e38",
          3210 => x"80538052",
          3211 => x"0280d305",
          3212 => x"335180cb",
          3213 => x"f73f82bb",
          3214 => x"98085282",
          3215 => x"a6e0518c",
          3216 => x"8e39b53d",
          3217 => x"ff801153",
          3218 => x"ff840551",
          3219 => x"d0e43f82",
          3220 => x"bb980880",
          3221 => x"2e873864",
          3222 => x"8926fcd9",
          3223 => x"38b53dfe",
          3224 => x"fc1153ff",
          3225 => x"840551d0",
          3226 => x"c93f82bb",
          3227 => x"98088638",
          3228 => x"82bb9808",
          3229 => x"44645382",
          3230 => x"a6e8527a",
          3231 => x"51ffb1be",
          3232 => x"3f0280cf",
          3233 => x"0533537a",
          3234 => x"526484b4",
          3235 => x"2982bcc4",
          3236 => x"055180f6",
          3237 => x"8e3f82bb",
          3238 => x"98088190",
          3239 => x"3882a6b8",
          3240 => x"51d5e03f",
          3241 => x"815efc8d",
          3242 => x"39b53dff",
          3243 => x"8405518f",
          3244 => x"b13f82bb",
          3245 => x"9808b63d",
          3246 => x"ff840552",
          3247 => x"5c90c73f",
          3248 => x"815382bb",
          3249 => x"9808527b",
          3250 => x"51f2ab3f",
          3251 => x"80d539b5",
          3252 => x"3dff8405",
          3253 => x"518f8b3f",
          3254 => x"82bb9808",
          3255 => x"b63dff84",
          3256 => x"05525c90",
          3257 => x"a13f82bb",
          3258 => x"9808b63d",
          3259 => x"ff840552",
          3260 => x"5b90933f",
          3261 => x"82bb9808",
          3262 => x"b63dff84",
          3263 => x"05525a90",
          3264 => x"853f82d2",
          3265 => x"e85982b9",
          3266 => x"bc5882bb",
          3267 => x"c8578056",
          3268 => x"805582bb",
          3269 => x"980881ff",
          3270 => x"06547953",
          3271 => x"7a527b51",
          3272 => x"f3913f82",
          3273 => x"bb980880",
          3274 => x"2efb8a38",
          3275 => x"82bb9808",
          3276 => x"51efe33f",
          3277 => x"faff39b5",
          3278 => x"3dff8011",
          3279 => x"53ff8405",
          3280 => x"51ceef3f",
          3281 => x"82bb9808",
          3282 => x"802efae9",
          3283 => x"38b53dfe",
          3284 => x"fc1153ff",
          3285 => x"840551ce",
          3286 => x"d93f82bb",
          3287 => x"9808802e",
          3288 => x"fad338b5",
          3289 => x"3dfef811",
          3290 => x"53ff8405",
          3291 => x"51cec33f",
          3292 => x"82bb9808",
          3293 => x"863882bb",
          3294 => x"98084382",
          3295 => x"a6ec51d4",
          3296 => x"823f6464",
          3297 => x"5d5b7a7c",
          3298 => x"2781ea38",
          3299 => x"625a797b",
          3300 => x"7084055d",
          3301 => x"0c7b7b26",
          3302 => x"f53881d9",
          3303 => x"39b53dff",
          3304 => x"801153ff",
          3305 => x"840551ce",
          3306 => x"893f82bb",
          3307 => x"9808802e",
          3308 => x"fa8338b5",
          3309 => x"3dfefc11",
          3310 => x"53ff8405",
          3311 => x"51cdf33f",
          3312 => x"82bb9808",
          3313 => x"802ef9ed",
          3314 => x"38b53dfe",
          3315 => x"f81153ff",
          3316 => x"840551cd",
          3317 => x"dd3f82bb",
          3318 => x"9808802e",
          3319 => x"f9d73882",
          3320 => x"a6fc51d3",
          3321 => x"9e3f645b",
          3322 => x"7a642781",
          3323 => x"8838625a",
          3324 => x"7a708105",
          3325 => x"5c337a34",
          3326 => x"62810543",
          3327 => x"eb39b53d",
          3328 => x"ff801153",
          3329 => x"ff840551",
          3330 => x"cda83f82",
          3331 => x"bb980880",
          3332 => x"2ef9a238",
          3333 => x"b53dfefc",
          3334 => x"1153ff84",
          3335 => x"0551cd92",
          3336 => x"3f82bb98",
          3337 => x"08802ef9",
          3338 => x"8c38b53d",
          3339 => x"fef81153",
          3340 => x"ff840551",
          3341 => x"ccfc3f82",
          3342 => x"bb980880",
          3343 => x"2ef8f638",
          3344 => x"82a78851",
          3345 => x"d2bd3f64",
          3346 => x"5b7a6427",
          3347 => x"a8386270",
          3348 => x"337c335f",
          3349 => x"5b5c797d",
          3350 => x"2e923879",
          3351 => x"557b547a",
          3352 => x"33537a52",
          3353 => x"82a79851",
          3354 => x"ffaaeb3f",
          3355 => x"811b6381",
          3356 => x"05445bd5",
          3357 => x"3982a7b0",
          3358 => x"5189fd39",
          3359 => x"b53dff80",
          3360 => x"1153ff84",
          3361 => x"0551ccaa",
          3362 => x"3f82bb98",
          3363 => x"0880df38",
          3364 => x"82ba8433",
          3365 => x"5a79802e",
          3366 => x"893882b9",
          3367 => x"bc084580",
          3368 => x"cd3982ba",
          3369 => x"85335a79",
          3370 => x"802e8838",
          3371 => x"82b9c408",
          3372 => x"45bc3982",
          3373 => x"ba86335a",
          3374 => x"79802e88",
          3375 => x"3882b9cc",
          3376 => x"0845ab39",
          3377 => x"82ba8733",
          3378 => x"5a79802e",
          3379 => x"883882b9",
          3380 => x"d408459a",
          3381 => x"3982ba82",
          3382 => x"335a7980",
          3383 => x"2e883882",
          3384 => x"b9dc0845",
          3385 => x"893982b9",
          3386 => x"ec08fc80",
          3387 => x"0545b53d",
          3388 => x"fefc1153",
          3389 => x"ff840551",
          3390 => x"cbb83f82",
          3391 => x"bb980880",
          3392 => x"de3882ba",
          3393 => x"84335a79",
          3394 => x"802e8938",
          3395 => x"82b9c008",
          3396 => x"4480cc39",
          3397 => x"82ba8533",
          3398 => x"5a79802e",
          3399 => x"883882b9",
          3400 => x"c80844bb",
          3401 => x"3982ba86",
          3402 => x"335a7980",
          3403 => x"2e883882",
          3404 => x"b9d00844",
          3405 => x"aa3982ba",
          3406 => x"87335a79",
          3407 => x"802e8838",
          3408 => x"82b9d808",
          3409 => x"44993982",
          3410 => x"ba82335a",
          3411 => x"79802e88",
          3412 => x"3882b9e0",
          3413 => x"08448839",
          3414 => x"82b9ec08",
          3415 => x"880544b5",
          3416 => x"3dfef811",
          3417 => x"53ff8405",
          3418 => x"51cac73f",
          3419 => x"82bb9808",
          3420 => x"802ea738",
          3421 => x"80635d5d",
          3422 => x"7b882e83",
          3423 => x"38815d7b",
          3424 => x"90327030",
          3425 => x"7072079f",
          3426 => x"2a706006",
          3427 => x"51515b5b",
          3428 => x"79802e88",
          3429 => x"387ba02e",
          3430 => x"83388843",
          3431 => x"82a7b451",
          3432 => x"cfe13fa0",
          3433 => x"55645462",
          3434 => x"53635264",
          3435 => x"51eecf3f",
          3436 => x"82a7c451",
          3437 => x"87c239b5",
          3438 => x"3dff8011",
          3439 => x"53ff8405",
          3440 => x"51c9ef3f",
          3441 => x"82bb9808",
          3442 => x"802ef5e9",
          3443 => x"38b53dfe",
          3444 => x"fc1153ff",
          3445 => x"840551c9",
          3446 => x"d93f82bb",
          3447 => x"9808802e",
          3448 => x"a438645a",
          3449 => x"0280cf05",
          3450 => x"337a3464",
          3451 => x"810545b5",
          3452 => x"3dfefc11",
          3453 => x"53ff8405",
          3454 => x"51c9b73f",
          3455 => x"82bb9808",
          3456 => x"e138f5b1",
          3457 => x"39647033",
          3458 => x"545282a7",
          3459 => x"d051ffa7",
          3460 => x"c53f80f8",
          3461 => x"527a51c8",
          3462 => x"e33f7a46",
          3463 => x"7a335a79",
          3464 => x"ae2ef591",
          3465 => x"389f7a27",
          3466 => x"9f38b53d",
          3467 => x"fefc1153",
          3468 => x"ff840551",
          3469 => x"c8fc3f82",
          3470 => x"bb980880",
          3471 => x"2e913864",
          3472 => x"5a0280cf",
          3473 => x"05337a34",
          3474 => x"64810545",
          3475 => x"ffb73982",
          3476 => x"a7dc51ce",
          3477 => x"ae3fffad",
          3478 => x"39b53dfe",
          3479 => x"f41153ff",
          3480 => x"840551c2",
          3481 => x"c63f82bb",
          3482 => x"9808802e",
          3483 => x"f4c738b5",
          3484 => x"3dfef011",
          3485 => x"53ff8405",
          3486 => x"51c2b03f",
          3487 => x"82bb9808",
          3488 => x"802ea638",
          3489 => x"615a0280",
          3490 => x"c205227a",
          3491 => x"7082055c",
          3492 => x"237942b5",
          3493 => x"3dfef011",
          3494 => x"53ff8405",
          3495 => x"51c28c3f",
          3496 => x"82bb9808",
          3497 => x"df38f48d",
          3498 => x"39617022",
          3499 => x"545282a7",
          3500 => x"e451ffa6",
          3501 => x"a13f80f8",
          3502 => x"527a51c7",
          3503 => x"bf3f7a46",
          3504 => x"7a335a79",
          3505 => x"ae2ef3ed",
          3506 => x"38799f26",
          3507 => x"87386182",
          3508 => x"0542d639",
          3509 => x"b53dfef0",
          3510 => x"1153ff84",
          3511 => x"0551c1cb",
          3512 => x"3f82bb98",
          3513 => x"08802e93",
          3514 => x"38615a02",
          3515 => x"80c20522",
          3516 => x"7a708205",
          3517 => x"5c237942",
          3518 => x"ffaf3982",
          3519 => x"a7dc51cd",
          3520 => x"823fffa5",
          3521 => x"39b53dfe",
          3522 => x"f41153ff",
          3523 => x"840551c1",
          3524 => x"9a3f82bb",
          3525 => x"9808802e",
          3526 => x"f39b38b5",
          3527 => x"3dfef011",
          3528 => x"53ff8405",
          3529 => x"51c1843f",
          3530 => x"82bb9808",
          3531 => x"802ea038",
          3532 => x"6161710c",
          3533 => x"5a618405",
          3534 => x"42b53dfe",
          3535 => x"f01153ff",
          3536 => x"840551c0",
          3537 => x"e63f82bb",
          3538 => x"9808e538",
          3539 => x"f2e73961",
          3540 => x"70085452",
          3541 => x"82a7f051",
          3542 => x"ffa4fb3f",
          3543 => x"80f8527a",
          3544 => x"51c6993f",
          3545 => x"7a467a33",
          3546 => x"5a79ae2e",
          3547 => x"f2c7389f",
          3548 => x"7a279b38",
          3549 => x"b53dfef0",
          3550 => x"1153ff84",
          3551 => x"0551c0ab",
          3552 => x"3f82bb98",
          3553 => x"08802e8d",
          3554 => x"38616171",
          3555 => x"0c5a6184",
          3556 => x"0542ffbb",
          3557 => x"3982a7dc",
          3558 => x"51cbe83f",
          3559 => x"ffb13982",
          3560 => x"a7fc51cb",
          3561 => x"de3f8251",
          3562 => x"988b3ff2",
          3563 => x"883982a8",
          3564 => x"9451cbcf",
          3565 => x"3fa25197",
          3566 => x"e03ff1f9",
          3567 => x"3982a8ac",
          3568 => x"51cbc03f",
          3569 => x"8480810b",
          3570 => x"87c09484",
          3571 => x"0c848081",
          3572 => x"0b87c094",
          3573 => x"940cf1dd",
          3574 => x"3982a8c0",
          3575 => x"51cba43f",
          3576 => x"8c80830b",
          3577 => x"87c09484",
          3578 => x"0c8c8083",
          3579 => x"0b87c094",
          3580 => x"940cf1c1",
          3581 => x"39b53dff",
          3582 => x"801153ff",
          3583 => x"840551c5",
          3584 => x"b13f82bb",
          3585 => x"9808802e",
          3586 => x"f1ab3864",
          3587 => x"5282a8d4",
          3588 => x"51ffa3c2",
          3589 => x"3f645a79",
          3590 => x"04b53dff",
          3591 => x"801153ff",
          3592 => x"840551c5",
          3593 => x"8d3f82bb",
          3594 => x"9808802e",
          3595 => x"f1873864",
          3596 => x"5282a8f0",
          3597 => x"51ffa39e",
          3598 => x"3f645a79",
          3599 => x"2d82bb98",
          3600 => x"08802ef0",
          3601 => x"f03882bb",
          3602 => x"98085282",
          3603 => x"a98c51ff",
          3604 => x"a3843ff0",
          3605 => x"e03982a9",
          3606 => x"a851caa7",
          3607 => x"3fffa2d7",
          3608 => x"3ff0d239",
          3609 => x"82a9c451",
          3610 => x"ca993f80",
          3611 => x"5affa839",
          3612 => x"91ad3ff0",
          3613 => x"c0397a46",
          3614 => x"7a335a79",
          3615 => x"802ef0b5",
          3616 => x"387e7e06",
          3617 => x"5a79802e",
          3618 => x"81d638b5",
          3619 => x"3dff8405",
          3620 => x"5183cf3f",
          3621 => x"82bb9808",
          3622 => x"5c815d7c",
          3623 => x"822eb238",
          3624 => x"7c822489",
          3625 => x"387c812e",
          3626 => x"8c3880cd",
          3627 => x"397c832e",
          3628 => x"b03880c5",
          3629 => x"3982a9d8",
          3630 => x"567b5582",
          3631 => x"a9dc5480",
          3632 => x"5382a9e0",
          3633 => x"52b53dff",
          3634 => x"b00551ff",
          3635 => x"a4f03fbb",
          3636 => x"3982aa80",
          3637 => x"52b53dff",
          3638 => x"b00551ff",
          3639 => x"a4e03fab",
          3640 => x"397b5582",
          3641 => x"a9dc5480",
          3642 => x"5382a9f0",
          3643 => x"52b53dff",
          3644 => x"b00551ff",
          3645 => x"a4c83f93",
          3646 => x"397b5480",
          3647 => x"5382a9fc",
          3648 => x"52b53dff",
          3649 => x"b00551ff",
          3650 => x"a4b43f82",
          3651 => x"d2e85982",
          3652 => x"b9bc5882",
          3653 => x"bbc85780",
          3654 => x"56655580",
          3655 => x"5482e080",
          3656 => x"5382e080",
          3657 => x"52b53dff",
          3658 => x"b00551e7",
          3659 => x"863f82bb",
          3660 => x"980882bb",
          3661 => x"98080970",
          3662 => x"30707207",
          3663 => x"8025515c",
          3664 => x"5c40805b",
          3665 => x"7c832683",
          3666 => x"38815b79",
          3667 => x"7b065a79",
          3668 => x"802e8d38",
          3669 => x"811d7081",
          3670 => x"ff065e5a",
          3671 => x"7cfebc38",
          3672 => x"7e81327e",
          3673 => x"8132075a",
          3674 => x"798a387f",
          3675 => x"ff2e0981",
          3676 => x"06eec238",
          3677 => x"82aa8451",
          3678 => x"c8893fee",
          3679 => x"b839f53d",
          3680 => x"0d800b82",
          3681 => x"bbc83487",
          3682 => x"c0948c70",
          3683 => x"08545587",
          3684 => x"84805272",
          3685 => x"51df8c3f",
          3686 => x"82bb9808",
          3687 => x"902b7508",
          3688 => x"55538784",
          3689 => x"80527351",
          3690 => x"def93f72",
          3691 => x"82bb9808",
          3692 => x"07750c87",
          3693 => x"c0949c70",
          3694 => x"08545587",
          3695 => x"84805272",
          3696 => x"51dee03f",
          3697 => x"82bb9808",
          3698 => x"902b7508",
          3699 => x"55538784",
          3700 => x"80527351",
          3701 => x"decd3f72",
          3702 => x"82bb9808",
          3703 => x"07750c8c",
          3704 => x"80830b87",
          3705 => x"c094840c",
          3706 => x"8c80830b",
          3707 => x"87c09494",
          3708 => x"0c80fa82",
          3709 => x"5a80fcee",
          3710 => x"5b830284",
          3711 => x"05990534",
          3712 => x"805c82d2",
          3713 => x"e80b873d",
          3714 => x"7088130c",
          3715 => x"70720c82",
          3716 => x"d2ec0c54",
          3717 => x"89bd3f93",
          3718 => x"c13f82aa",
          3719 => x"9451c6e3",
          3720 => x"3f82aaa0",
          3721 => x"51c6dc3f",
          3722 => x"80dda851",
          3723 => x"92e63f81",
          3724 => x"51e8b83f",
          3725 => x"ecae3f80",
          3726 => x"04fe3d0d",
          3727 => x"80528353",
          3728 => x"71882b52",
          3729 => x"87d93f82",
          3730 => x"bb980881",
          3731 => x"ff067207",
          3732 => x"ff145452",
          3733 => x"728025e8",
          3734 => x"387182bb",
          3735 => x"980c843d",
          3736 => x"0d04fc3d",
          3737 => x"0d767008",
          3738 => x"54558073",
          3739 => x"52547274",
          3740 => x"2e818a38",
          3741 => x"72335170",
          3742 => x"a02e0981",
          3743 => x"06863881",
          3744 => x"1353f139",
          3745 => x"72335170",
          3746 => x"a22e0981",
          3747 => x"06863881",
          3748 => x"13538154",
          3749 => x"72527381",
          3750 => x"2e098106",
          3751 => x"9f388439",
          3752 => x"81125280",
          3753 => x"72335254",
          3754 => x"70a22e83",
          3755 => x"38815470",
          3756 => x"802e9d38",
          3757 => x"73ea3898",
          3758 => x"39811252",
          3759 => x"80723352",
          3760 => x"5470a02e",
          3761 => x"83388154",
          3762 => x"70802e84",
          3763 => x"3873ea38",
          3764 => x"80723352",
          3765 => x"5470a02e",
          3766 => x"09810683",
          3767 => x"38815470",
          3768 => x"a2327030",
          3769 => x"70802576",
          3770 => x"07515151",
          3771 => x"70802e88",
          3772 => x"38807270",
          3773 => x"81055434",
          3774 => x"71750c72",
          3775 => x"517082bb",
          3776 => x"980c863d",
          3777 => x"0d04fc3d",
          3778 => x"0d765372",
          3779 => x"08802e92",
          3780 => x"38863dfc",
          3781 => x"05527251",
          3782 => x"ffb9903f",
          3783 => x"82bb9808",
          3784 => x"85388053",
          3785 => x"83397453",
          3786 => x"7282bb98",
          3787 => x"0c863d0d",
          3788 => x"04fc3d0d",
          3789 => x"76821133",
          3790 => x"ff055253",
          3791 => x"8152708b",
          3792 => x"26819838",
          3793 => x"831333ff",
          3794 => x"05518252",
          3795 => x"709e2681",
          3796 => x"8a388413",
          3797 => x"33518352",
          3798 => x"70972680",
          3799 => x"fe388513",
          3800 => x"33518452",
          3801 => x"70bb2680",
          3802 => x"f2388613",
          3803 => x"33518552",
          3804 => x"70bb2680",
          3805 => x"e6388813",
          3806 => x"22558652",
          3807 => x"7487e726",
          3808 => x"80d9388a",
          3809 => x"13225487",
          3810 => x"527387e7",
          3811 => x"2680cc38",
          3812 => x"810b87c0",
          3813 => x"989c0c72",
          3814 => x"2287c098",
          3815 => x"bc0c8213",
          3816 => x"3387c098",
          3817 => x"b80c8313",
          3818 => x"3387c098",
          3819 => x"b40c8413",
          3820 => x"3387c098",
          3821 => x"b00c8513",
          3822 => x"3387c098",
          3823 => x"ac0c8613",
          3824 => x"3387c098",
          3825 => x"a80c7487",
          3826 => x"c098a40c",
          3827 => x"7387c098",
          3828 => x"a00c800b",
          3829 => x"87c0989c",
          3830 => x"0c805271",
          3831 => x"82bb980c",
          3832 => x"863d0d04",
          3833 => x"f33d0d7f",
          3834 => x"5b87c098",
          3835 => x"9c5d817d",
          3836 => x"0c87c098",
          3837 => x"bc085e7d",
          3838 => x"7b2387c0",
          3839 => x"98b8085a",
          3840 => x"79821c34",
          3841 => x"87c098b4",
          3842 => x"085a7983",
          3843 => x"1c3487c0",
          3844 => x"98b0085a",
          3845 => x"79841c34",
          3846 => x"87c098ac",
          3847 => x"085a7985",
          3848 => x"1c3487c0",
          3849 => x"98a8085a",
          3850 => x"79861c34",
          3851 => x"87c098a4",
          3852 => x"085c7b88",
          3853 => x"1c2387c0",
          3854 => x"98a0085a",
          3855 => x"798a1c23",
          3856 => x"807d0c79",
          3857 => x"83ffff06",
          3858 => x"597b83ff",
          3859 => x"ff065886",
          3860 => x"1b335785",
          3861 => x"1b335684",
          3862 => x"1b335583",
          3863 => x"1b335482",
          3864 => x"1b33537d",
          3865 => x"83ffff06",
          3866 => x"5282aab8",
          3867 => x"51ff9ae6",
          3868 => x"3f8f3d0d",
          3869 => x"04fb3d0d",
          3870 => x"029f0533",
          3871 => x"82b9b833",
          3872 => x"7081ff06",
          3873 => x"58555587",
          3874 => x"c0948451",
          3875 => x"75802e86",
          3876 => x"3887c094",
          3877 => x"94517008",
          3878 => x"70962a70",
          3879 => x"81065354",
          3880 => x"5270802e",
          3881 => x"8c387191",
          3882 => x"2a708106",
          3883 => x"515170d7",
          3884 => x"38728132",
          3885 => x"70810651",
          3886 => x"5170802e",
          3887 => x"8d387193",
          3888 => x"2a708106",
          3889 => x"515170ff",
          3890 => x"be387381",
          3891 => x"ff065187",
          3892 => x"c0948052",
          3893 => x"70802e86",
          3894 => x"3887c094",
          3895 => x"90527472",
          3896 => x"0c7482bb",
          3897 => x"980c873d",
          3898 => x"0d04ff3d",
          3899 => x"0d028f05",
          3900 => x"33703070",
          3901 => x"9f2a5152",
          3902 => x"527082b9",
          3903 => x"b834833d",
          3904 => x"0d04f93d",
          3905 => x"0d02a705",
          3906 => x"3358778a",
          3907 => x"2e098106",
          3908 => x"87387a52",
          3909 => x"8d51eb3f",
          3910 => x"82b9b833",
          3911 => x"7081ff06",
          3912 => x"585687c0",
          3913 => x"94845376",
          3914 => x"802e8638",
          3915 => x"87c09494",
          3916 => x"53720870",
          3917 => x"962a7081",
          3918 => x"06555654",
          3919 => x"72802e8c",
          3920 => x"3873912a",
          3921 => x"70810651",
          3922 => x"5372d738",
          3923 => x"74813270",
          3924 => x"81065153",
          3925 => x"72802e8d",
          3926 => x"3873932a",
          3927 => x"70810651",
          3928 => x"5372ffbe",
          3929 => x"387581ff",
          3930 => x"065387c0",
          3931 => x"94805472",
          3932 => x"802e8638",
          3933 => x"87c09490",
          3934 => x"5477740c",
          3935 => x"800b82bb",
          3936 => x"980c893d",
          3937 => x"0d04f93d",
          3938 => x"0d795480",
          3939 => x"74337081",
          3940 => x"ff065353",
          3941 => x"5770772e",
          3942 => x"80fc3871",
          3943 => x"81ff0681",
          3944 => x"1582b9b8",
          3945 => x"337081ff",
          3946 => x"06595755",
          3947 => x"5887c094",
          3948 => x"84517580",
          3949 => x"2e863887",
          3950 => x"c0949451",
          3951 => x"70087096",
          3952 => x"2a708106",
          3953 => x"53545270",
          3954 => x"802e8c38",
          3955 => x"71912a70",
          3956 => x"81065151",
          3957 => x"70d73872",
          3958 => x"81327081",
          3959 => x"06515170",
          3960 => x"802e8d38",
          3961 => x"71932a70",
          3962 => x"81065151",
          3963 => x"70ffbe38",
          3964 => x"7481ff06",
          3965 => x"5187c094",
          3966 => x"80527080",
          3967 => x"2e863887",
          3968 => x"c0949052",
          3969 => x"77720c81",
          3970 => x"17743370",
          3971 => x"81ff0653",
          3972 => x"535770ff",
          3973 => x"86387682",
          3974 => x"bb980c89",
          3975 => x"3d0d04fe",
          3976 => x"3d0d82b9",
          3977 => x"b8337081",
          3978 => x"ff065452",
          3979 => x"87c09484",
          3980 => x"5172802e",
          3981 => x"863887c0",
          3982 => x"94945170",
          3983 => x"0870822a",
          3984 => x"70810651",
          3985 => x"51517080",
          3986 => x"2ee23871",
          3987 => x"81ff0651",
          3988 => x"87c09480",
          3989 => x"5270802e",
          3990 => x"863887c0",
          3991 => x"94905271",
          3992 => x"087081ff",
          3993 => x"0682bb98",
          3994 => x"0c51843d",
          3995 => x"0d04ffaf",
          3996 => x"3f82bb98",
          3997 => x"0881ff06",
          3998 => x"82bb980c",
          3999 => x"04fe3d0d",
          4000 => x"82b9b833",
          4001 => x"7081ff06",
          4002 => x"525387c0",
          4003 => x"94845270",
          4004 => x"802e8638",
          4005 => x"87c09494",
          4006 => x"52710870",
          4007 => x"822a7081",
          4008 => x"06515151",
          4009 => x"ff527080",
          4010 => x"2ea03872",
          4011 => x"81ff0651",
          4012 => x"87c09480",
          4013 => x"5270802e",
          4014 => x"863887c0",
          4015 => x"94905271",
          4016 => x"0870982b",
          4017 => x"70982c51",
          4018 => x"53517182",
          4019 => x"bb980c84",
          4020 => x"3d0d04ff",
          4021 => x"3d0d87c0",
          4022 => x"9e800870",
          4023 => x"9c2a8a06",
          4024 => x"51517080",
          4025 => x"2e84b438",
          4026 => x"87c09ea4",
          4027 => x"0882b9bc",
          4028 => x"0c87c09e",
          4029 => x"a80882b9",
          4030 => x"c00c87c0",
          4031 => x"9e940882",
          4032 => x"b9c40c87",
          4033 => x"c09e9808",
          4034 => x"82b9c80c",
          4035 => x"87c09e9c",
          4036 => x"0882b9cc",
          4037 => x"0c87c09e",
          4038 => x"a00882b9",
          4039 => x"d00c87c0",
          4040 => x"9eac0882",
          4041 => x"b9d40c87",
          4042 => x"c09eb008",
          4043 => x"82b9d80c",
          4044 => x"87c09eb4",
          4045 => x"0882b9dc",
          4046 => x"0c87c09e",
          4047 => x"b80882b9",
          4048 => x"e00c87c0",
          4049 => x"9ebc0882",
          4050 => x"b9e40c87",
          4051 => x"c09ec008",
          4052 => x"82b9e80c",
          4053 => x"87c09ec4",
          4054 => x"0882b9ec",
          4055 => x"0c87c09e",
          4056 => x"80085170",
          4057 => x"82b9f023",
          4058 => x"87c09e84",
          4059 => x"0882b9f4",
          4060 => x"0c87c09e",
          4061 => x"880882b9",
          4062 => x"f80c87c0",
          4063 => x"9e8c0882",
          4064 => x"b9fc0c81",
          4065 => x"0b82ba80",
          4066 => x"34800b87",
          4067 => x"c09e9008",
          4068 => x"7084800a",
          4069 => x"06515252",
          4070 => x"70802e83",
          4071 => x"38815271",
          4072 => x"82ba8134",
          4073 => x"800b87c0",
          4074 => x"9e900870",
          4075 => x"88800a06",
          4076 => x"51525270",
          4077 => x"802e8338",
          4078 => x"81527182",
          4079 => x"ba823480",
          4080 => x"0b87c09e",
          4081 => x"90087090",
          4082 => x"800a0651",
          4083 => x"52527080",
          4084 => x"2e833881",
          4085 => x"527182ba",
          4086 => x"8334800b",
          4087 => x"87c09e90",
          4088 => x"08708880",
          4089 => x"80065152",
          4090 => x"5270802e",
          4091 => x"83388152",
          4092 => x"7182ba84",
          4093 => x"34800b87",
          4094 => x"c09e9008",
          4095 => x"70a08080",
          4096 => x"06515252",
          4097 => x"70802e83",
          4098 => x"38815271",
          4099 => x"82ba8534",
          4100 => x"800b87c0",
          4101 => x"9e900870",
          4102 => x"90808006",
          4103 => x"51525270",
          4104 => x"802e8338",
          4105 => x"81527182",
          4106 => x"ba863480",
          4107 => x"0b87c09e",
          4108 => x"90087084",
          4109 => x"80800651",
          4110 => x"52527080",
          4111 => x"2e833881",
          4112 => x"527182ba",
          4113 => x"8734800b",
          4114 => x"87c09e90",
          4115 => x"08708280",
          4116 => x"80065152",
          4117 => x"5270802e",
          4118 => x"83388152",
          4119 => x"7182ba88",
          4120 => x"34800b87",
          4121 => x"c09e9008",
          4122 => x"70818080",
          4123 => x"06515252",
          4124 => x"70802e83",
          4125 => x"38815271",
          4126 => x"82ba8934",
          4127 => x"800b87c0",
          4128 => x"9e900870",
          4129 => x"80c08006",
          4130 => x"51525270",
          4131 => x"802e8338",
          4132 => x"81527182",
          4133 => x"ba8a3480",
          4134 => x"0b87c09e",
          4135 => x"900870a0",
          4136 => x"80065152",
          4137 => x"5270802e",
          4138 => x"83388152",
          4139 => x"7182ba8b",
          4140 => x"3487c09e",
          4141 => x"90087098",
          4142 => x"8006708a",
          4143 => x"2a515151",
          4144 => x"7082ba8c",
          4145 => x"34800b87",
          4146 => x"c09e9008",
          4147 => x"70848006",
          4148 => x"51525270",
          4149 => x"802e8338",
          4150 => x"81527182",
          4151 => x"ba8d3487",
          4152 => x"c09e9008",
          4153 => x"7083f006",
          4154 => x"70842a51",
          4155 => x"51517082",
          4156 => x"ba8e3480",
          4157 => x"0b87c09e",
          4158 => x"90087088",
          4159 => x"06515252",
          4160 => x"70802e83",
          4161 => x"38815271",
          4162 => x"82ba8f34",
          4163 => x"87c09e90",
          4164 => x"08708706",
          4165 => x"51517082",
          4166 => x"ba903483",
          4167 => x"3d0d04fb",
          4168 => x"3d0d82aa",
          4169 => x"d051ffb8",
          4170 => x"da3f82ba",
          4171 => x"80335473",
          4172 => x"802e8938",
          4173 => x"82aae451",
          4174 => x"ffb8c83f",
          4175 => x"82aaf851",
          4176 => x"ffb8c03f",
          4177 => x"82ba8233",
          4178 => x"5473802e",
          4179 => x"943882b9",
          4180 => x"dc0882b9",
          4181 => x"e0081154",
          4182 => x"5282ab90",
          4183 => x"51ff90f6",
          4184 => x"3f82ba87",
          4185 => x"33547380",
          4186 => x"2e943882",
          4187 => x"b9d40882",
          4188 => x"b9d80811",
          4189 => x"545282ab",
          4190 => x"ac51ff90",
          4191 => x"d93f82ba",
          4192 => x"84335473",
          4193 => x"802e9438",
          4194 => x"82b9bc08",
          4195 => x"82b9c008",
          4196 => x"11545282",
          4197 => x"abc851ff",
          4198 => x"90bc3f82",
          4199 => x"ba853354",
          4200 => x"73802e94",
          4201 => x"3882b9c4",
          4202 => x"0882b9c8",
          4203 => x"08115452",
          4204 => x"82abe451",
          4205 => x"ff909f3f",
          4206 => x"82ba8633",
          4207 => x"5473802e",
          4208 => x"943882b9",
          4209 => x"cc0882b9",
          4210 => x"d0081154",
          4211 => x"5282ac80",
          4212 => x"51ff9082",
          4213 => x"3f82ba8b",
          4214 => x"33547380",
          4215 => x"2e8e3882",
          4216 => x"ba8c3352",
          4217 => x"82ac9c51",
          4218 => x"ff8feb3f",
          4219 => x"82ba8f33",
          4220 => x"5473802e",
          4221 => x"8e3882ba",
          4222 => x"90335282",
          4223 => x"acbc51ff",
          4224 => x"8fd43f82",
          4225 => x"ba8d3354",
          4226 => x"73802e8e",
          4227 => x"3882ba8e",
          4228 => x"335282ac",
          4229 => x"dc51ff8f",
          4230 => x"bd3f82ba",
          4231 => x"81335473",
          4232 => x"802e8938",
          4233 => x"82acfc51",
          4234 => x"ffb6d83f",
          4235 => x"82ba8333",
          4236 => x"5473802e",
          4237 => x"893882ad",
          4238 => x"9051ffb6",
          4239 => x"c63f82ba",
          4240 => x"88335473",
          4241 => x"802e8938",
          4242 => x"82ad9c51",
          4243 => x"ffb6b43f",
          4244 => x"82ba8933",
          4245 => x"5473802e",
          4246 => x"893882ad",
          4247 => x"a851ffb6",
          4248 => x"a23f82ba",
          4249 => x"8a335473",
          4250 => x"802e8938",
          4251 => x"82adb451",
          4252 => x"ffb6903f",
          4253 => x"82adc051",
          4254 => x"ffb6883f",
          4255 => x"82b9e408",
          4256 => x"5282adcc",
          4257 => x"51ff8ece",
          4258 => x"3f82b9e8",
          4259 => x"085282ad",
          4260 => x"f451ff8e",
          4261 => x"c13f82b9",
          4262 => x"ec085282",
          4263 => x"ae9c51ff",
          4264 => x"8eb43f82",
          4265 => x"aec451ff",
          4266 => x"b5d93f82",
          4267 => x"b9f02252",
          4268 => x"82aecc51",
          4269 => x"ff8e9f3f",
          4270 => x"82b9f408",
          4271 => x"56bd84c0",
          4272 => x"527551cc",
          4273 => x"de3f82bb",
          4274 => x"9808bd84",
          4275 => x"c0297671",
          4276 => x"31545482",
          4277 => x"bb980852",
          4278 => x"82aef451",
          4279 => x"ff8df73f",
          4280 => x"82ba8733",
          4281 => x"5473802e",
          4282 => x"a93882b9",
          4283 => x"f80856bd",
          4284 => x"84c05275",
          4285 => x"51ccac3f",
          4286 => x"82bb9808",
          4287 => x"bd84c029",
          4288 => x"76713154",
          4289 => x"5482bb98",
          4290 => x"085282af",
          4291 => x"a051ff8d",
          4292 => x"c53f82ba",
          4293 => x"82335473",
          4294 => x"802ea938",
          4295 => x"82b9fc08",
          4296 => x"56bd84c0",
          4297 => x"527551cb",
          4298 => x"fa3f82bb",
          4299 => x"9808bd84",
          4300 => x"c0297671",
          4301 => x"31545482",
          4302 => x"bb980852",
          4303 => x"82afcc51",
          4304 => x"ff8d933f",
          4305 => x"82a7b051",
          4306 => x"ffb4b83f",
          4307 => x"873d0d04",
          4308 => x"fe3d0d02",
          4309 => x"920533ff",
          4310 => x"05527184",
          4311 => x"26aa3871",
          4312 => x"8429829a",
          4313 => x"80055271",
          4314 => x"080482af",
          4315 => x"f8519d39",
          4316 => x"82b08051",
          4317 => x"973982b0",
          4318 => x"88519139",
          4319 => x"82b09051",
          4320 => x"8b3982b0",
          4321 => x"94518539",
          4322 => x"82b09c51",
          4323 => x"ffb3f43f",
          4324 => x"843d0d04",
          4325 => x"7188800c",
          4326 => x"04ff3d0d",
          4327 => x"87c09684",
          4328 => x"70085252",
          4329 => x"80720c70",
          4330 => x"74077082",
          4331 => x"ba940c72",
          4332 => x"0c833d0d",
          4333 => x"04ff3d0d",
          4334 => x"87c09684",
          4335 => x"700882ba",
          4336 => x"940c5280",
          4337 => x"720c7309",
          4338 => x"7082ba94",
          4339 => x"08067082",
          4340 => x"ba940c73",
          4341 => x"0c51833d",
          4342 => x"0d04800b",
          4343 => x"87c09684",
          4344 => x"0c0482ba",
          4345 => x"940887c0",
          4346 => x"96840c04",
          4347 => x"fd3d0d76",
          4348 => x"982b7098",
          4349 => x"2c79982b",
          4350 => x"70982c72",
          4351 => x"10137082",
          4352 => x"2b515351",
          4353 => x"54515180",
          4354 => x"0b82b0a8",
          4355 => x"12335553",
          4356 => x"7174259c",
          4357 => x"3882b0a4",
          4358 => x"11081202",
          4359 => x"84059705",
          4360 => x"33713352",
          4361 => x"52527072",
          4362 => x"2e098106",
          4363 => x"83388153",
          4364 => x"7282bb98",
          4365 => x"0c853d0d",
          4366 => x"04fc3d0d",
          4367 => x"78028405",
          4368 => x"9f053371",
          4369 => x"33545553",
          4370 => x"71802ea2",
          4371 => x"388851ff",
          4372 => x"b5d33fa0",
          4373 => x"51ffb5cd",
          4374 => x"3f8851ff",
          4375 => x"b5c73f72",
          4376 => x"33ff0552",
          4377 => x"71733471",
          4378 => x"81ff0652",
          4379 => x"db397651",
          4380 => x"ffb2903f",
          4381 => x"73733486",
          4382 => x"3d0d04f6",
          4383 => x"3d0d7c02",
          4384 => x"8405b705",
          4385 => x"33028805",
          4386 => x"bb053382",
          4387 => x"baf03370",
          4388 => x"842982ba",
          4389 => x"98057008",
          4390 => x"5159595a",
          4391 => x"58597480",
          4392 => x"2e863874",
          4393 => x"519ab53f",
          4394 => x"82baf033",
          4395 => x"70842982",
          4396 => x"ba980581",
          4397 => x"19705458",
          4398 => x"565a9db6",
          4399 => x"3f82bb98",
          4400 => x"08750c82",
          4401 => x"baf03370",
          4402 => x"842982ba",
          4403 => x"98057008",
          4404 => x"51565a74",
          4405 => x"802ea738",
          4406 => x"75537852",
          4407 => x"7451ffbf",
          4408 => x"a43f82ba",
          4409 => x"f0338105",
          4410 => x"557482ba",
          4411 => x"f0347481",
          4412 => x"ff065593",
          4413 => x"75278738",
          4414 => x"800b82ba",
          4415 => x"f0347780",
          4416 => x"2eb63882",
          4417 => x"baec0856",
          4418 => x"75802eac",
          4419 => x"3882bae8",
          4420 => x"335574a4",
          4421 => x"388c3dfc",
          4422 => x"05547653",
          4423 => x"78527551",
          4424 => x"80d9c33f",
          4425 => x"82baec08",
          4426 => x"528a5181",
          4427 => x"8ed03f82",
          4428 => x"baec0851",
          4429 => x"80dda03f",
          4430 => x"8c3d0d04",
          4431 => x"fd3d0d82",
          4432 => x"ba985393",
          4433 => x"54720852",
          4434 => x"71802e89",
          4435 => x"38715199",
          4436 => x"8b3f8073",
          4437 => x"0cff1484",
          4438 => x"14545473",
          4439 => x"8025e638",
          4440 => x"800b82ba",
          4441 => x"f03482ba",
          4442 => x"ec085271",
          4443 => x"802e9538",
          4444 => x"715180de",
          4445 => x"803f82ba",
          4446 => x"ec085198",
          4447 => x"df3f800b",
          4448 => x"82baec0c",
          4449 => x"853d0d04",
          4450 => x"dc3d0d81",
          4451 => x"57805282",
          4452 => x"baec0851",
          4453 => x"80e2ed3f",
          4454 => x"82bb9808",
          4455 => x"80d33882",
          4456 => x"baec0853",
          4457 => x"80f85288",
          4458 => x"3d705256",
          4459 => x"818bbb3f",
          4460 => x"82bb9808",
          4461 => x"802eba38",
          4462 => x"7551ffbb",
          4463 => x"e83f82bb",
          4464 => x"98085580",
          4465 => x"0b82bb98",
          4466 => x"08259d38",
          4467 => x"82bb9808",
          4468 => x"ff057017",
          4469 => x"55558074",
          4470 => x"34755376",
          4471 => x"52811782",
          4472 => x"b3985257",
          4473 => x"ff87ef3f",
          4474 => x"74ff2e09",
          4475 => x"8106ffaf",
          4476 => x"38a63d0d",
          4477 => x"04d93d0d",
          4478 => x"aa3d08ad",
          4479 => x"3d085a5a",
          4480 => x"81705858",
          4481 => x"805282ba",
          4482 => x"ec085180",
          4483 => x"e1f63f82",
          4484 => x"bb980881",
          4485 => x"9538ff0b",
          4486 => x"82baec08",
          4487 => x"545580f8",
          4488 => x"528b3d70",
          4489 => x"5256818a",
          4490 => x"c13f82bb",
          4491 => x"9808802e",
          4492 => x"a5387551",
          4493 => x"ffbaee3f",
          4494 => x"82bb9808",
          4495 => x"81185855",
          4496 => x"800b82bb",
          4497 => x"9808258e",
          4498 => x"3882bb98",
          4499 => x"08ff0570",
          4500 => x"17555580",
          4501 => x"74347409",
          4502 => x"70307072",
          4503 => x"079f2a51",
          4504 => x"55557877",
          4505 => x"2e853873",
          4506 => x"ffac3882",
          4507 => x"baec088c",
          4508 => x"11085351",
          4509 => x"80e18d3f",
          4510 => x"82bb9808",
          4511 => x"802e8938",
          4512 => x"82b3a451",
          4513 => x"ffadfc3f",
          4514 => x"78772e09",
          4515 => x"81069b38",
          4516 => x"75527951",
          4517 => x"ffbafc3f",
          4518 => x"7951ffba",
          4519 => x"883fab3d",
          4520 => x"085482bb",
          4521 => x"98087434",
          4522 => x"80587782",
          4523 => x"bb980ca9",
          4524 => x"3d0d04f6",
          4525 => x"3d0d7c7e",
          4526 => x"715c7172",
          4527 => x"3357595a",
          4528 => x"5873a02e",
          4529 => x"098106a2",
          4530 => x"38783378",
          4531 => x"05567776",
          4532 => x"27983881",
          4533 => x"17705b70",
          4534 => x"71335658",
          4535 => x"5573a02e",
          4536 => x"09810686",
          4537 => x"38757526",
          4538 => x"ea388054",
          4539 => x"73882982",
          4540 => x"baf40570",
          4541 => x"085255ff",
          4542 => x"b9ab3f82",
          4543 => x"bb980853",
          4544 => x"79527408",
          4545 => x"51ffbcaa",
          4546 => x"3f82bb98",
          4547 => x"0880c638",
          4548 => x"84153355",
          4549 => x"74812e88",
          4550 => x"3874822e",
          4551 => x"8838b639",
          4552 => x"fce63fad",
          4553 => x"39811a5a",
          4554 => x"8c3dfc11",
          4555 => x"53f80551",
          4556 => x"ffa6ff3f",
          4557 => x"82bb9808",
          4558 => x"802e9a38",
          4559 => x"ff1b5378",
          4560 => x"527751fd",
          4561 => x"b03f82bb",
          4562 => x"980881ff",
          4563 => x"06557485",
          4564 => x"38745491",
          4565 => x"39811470",
          4566 => x"81ff0651",
          4567 => x"54827427",
          4568 => x"ff8a3880",
          4569 => x"547382bb",
          4570 => x"980c8c3d",
          4571 => x"0d04d33d",
          4572 => x"0db03d08",
          4573 => x"b23d08b4",
          4574 => x"3d08595f",
          4575 => x"5a800baf",
          4576 => x"3d3482ba",
          4577 => x"f03382ba",
          4578 => x"ec08555b",
          4579 => x"7381cb38",
          4580 => x"7382bae8",
          4581 => x"33555573",
          4582 => x"83388155",
          4583 => x"76802e81",
          4584 => x"bc388170",
          4585 => x"76065556",
          4586 => x"73802e81",
          4587 => x"ad38a851",
          4588 => x"97c03f82",
          4589 => x"bb980882",
          4590 => x"baec0c82",
          4591 => x"bb980880",
          4592 => x"2e819238",
          4593 => x"93537652",
          4594 => x"82bb9808",
          4595 => x"5180ccb4",
          4596 => x"3f82bb98",
          4597 => x"08802e8c",
          4598 => x"3882b3d0",
          4599 => x"51ffaba3",
          4600 => x"3f80f739",
          4601 => x"82bb9808",
          4602 => x"5b82baec",
          4603 => x"085380f8",
          4604 => x"52903d70",
          4605 => x"52548186",
          4606 => x"f13f82bb",
          4607 => x"98085682",
          4608 => x"bb980874",
          4609 => x"2e098106",
          4610 => x"80d03882",
          4611 => x"bb980851",
          4612 => x"ffb7923f",
          4613 => x"82bb9808",
          4614 => x"55800b82",
          4615 => x"bb980825",
          4616 => x"a93882bb",
          4617 => x"9808ff05",
          4618 => x"70175555",
          4619 => x"80743480",
          4620 => x"537481ff",
          4621 => x"06527551",
          4622 => x"f8c13f81",
          4623 => x"1b7081ff",
          4624 => x"065c5493",
          4625 => x"7b278338",
          4626 => x"805b74ff",
          4627 => x"2e098106",
          4628 => x"ff973886",
          4629 => x"397582ba",
          4630 => x"e834768c",
          4631 => x"3882baec",
          4632 => x"08802e84",
          4633 => x"38f9d53f",
          4634 => x"8f3d5dec",
          4635 => x"903f82bb",
          4636 => x"9808982b",
          4637 => x"70982c51",
          4638 => x"5978ff2e",
          4639 => x"ee387881",
          4640 => x"ff0682d2",
          4641 => x"c4337098",
          4642 => x"2b70982c",
          4643 => x"82d2c033",
          4644 => x"70982b70",
          4645 => x"972c7198",
          4646 => x"2c057084",
          4647 => x"2982b0a4",
          4648 => x"05700815",
          4649 => x"70335151",
          4650 => x"51515959",
          4651 => x"51595d58",
          4652 => x"81567378",
          4653 => x"2e80e938",
          4654 => x"777427b4",
          4655 => x"38748180",
          4656 => x"0a2981ff",
          4657 => x"0a057098",
          4658 => x"2c515580",
          4659 => x"752480ce",
          4660 => x"38765374",
          4661 => x"527751f6",
          4662 => x"933f82bb",
          4663 => x"980881ff",
          4664 => x"06547380",
          4665 => x"2ed73874",
          4666 => x"82d2c034",
          4667 => x"8156b139",
          4668 => x"7481800a",
          4669 => x"2981800a",
          4670 => x"0570982c",
          4671 => x"7081ff06",
          4672 => x"56515573",
          4673 => x"95269738",
          4674 => x"76537452",
          4675 => x"7751f5dc",
          4676 => x"3f82bb98",
          4677 => x"0881ff06",
          4678 => x"5473cc38",
          4679 => x"d3398056",
          4680 => x"75802e80",
          4681 => x"ca38811c",
          4682 => x"557482d2",
          4683 => x"c4347498",
          4684 => x"2b70982c",
          4685 => x"82d2c033",
          4686 => x"70982b70",
          4687 => x"982c7010",
          4688 => x"1170822b",
          4689 => x"82b0a811",
          4690 => x"335e5151",
          4691 => x"51575851",
          4692 => x"5574772e",
          4693 => x"098106fe",
          4694 => x"923882b0",
          4695 => x"ac14087d",
          4696 => x"0c800b82",
          4697 => x"d2c43480",
          4698 => x"0b82d2c0",
          4699 => x"34923975",
          4700 => x"82d2c434",
          4701 => x"7582d2c0",
          4702 => x"3478af3d",
          4703 => x"34757d0c",
          4704 => x"7e547395",
          4705 => x"26fde138",
          4706 => x"73842982",
          4707 => x"9a940554",
          4708 => x"73080482",
          4709 => x"d2cc3354",
          4710 => x"737e2efd",
          4711 => x"cb3882d2",
          4712 => x"c8335573",
          4713 => x"7527ab38",
          4714 => x"74982b70",
          4715 => x"982c5155",
          4716 => x"7375249e",
          4717 => x"38741a54",
          4718 => x"73338115",
          4719 => x"34748180",
          4720 => x"0a2981ff",
          4721 => x"0a057098",
          4722 => x"2c82d2cc",
          4723 => x"33565155",
          4724 => x"df3982d2",
          4725 => x"cc338111",
          4726 => x"56547482",
          4727 => x"d2cc3473",
          4728 => x"1a54ae3d",
          4729 => x"33743482",
          4730 => x"d2c83354",
          4731 => x"737e2589",
          4732 => x"38811454",
          4733 => x"7382d2c8",
          4734 => x"3482d2cc",
          4735 => x"33708180",
          4736 => x"0a2981ff",
          4737 => x"0a057098",
          4738 => x"2c82d2c8",
          4739 => x"335a5156",
          4740 => x"56747725",
          4741 => x"a338741a",
          4742 => x"70335254",
          4743 => x"ffaa863f",
          4744 => x"7481800a",
          4745 => x"2981800a",
          4746 => x"0570982c",
          4747 => x"82d2c833",
          4748 => x"56515573",
          4749 => x"7524df38",
          4750 => x"82d2cc33",
          4751 => x"70982b70",
          4752 => x"982c82d2",
          4753 => x"c8335a51",
          4754 => x"56567477",
          4755 => x"25fc9938",
          4756 => x"8851ffa9",
          4757 => x"d03f7481",
          4758 => x"800a2981",
          4759 => x"800a0570",
          4760 => x"982c82d2",
          4761 => x"c8335651",
          4762 => x"55737524",
          4763 => x"e338fbf8",
          4764 => x"39837a34",
          4765 => x"800b811b",
          4766 => x"3482d2cc",
          4767 => x"53805282",
          4768 => x"a98851f3",
          4769 => x"b43f81e4",
          4770 => x"3982d2cc",
          4771 => x"337081ff",
          4772 => x"06555573",
          4773 => x"802efbd0",
          4774 => x"3882d2c8",
          4775 => x"33ff0554",
          4776 => x"7382d2c8",
          4777 => x"34ff1554",
          4778 => x"7382d2cc",
          4779 => x"348851ff",
          4780 => x"a8f33f82",
          4781 => x"d2cc3370",
          4782 => x"982b7098",
          4783 => x"2c82d2c8",
          4784 => x"33575156",
          4785 => x"57747425",
          4786 => x"a838741a",
          4787 => x"54811433",
          4788 => x"74347333",
          4789 => x"51ffa8cd",
          4790 => x"3f748180",
          4791 => x"0a298180",
          4792 => x"0a057098",
          4793 => x"2c82d2c8",
          4794 => x"33585155",
          4795 => x"757524da",
          4796 => x"38a051ff",
          4797 => x"a8af3f82",
          4798 => x"d2cc3370",
          4799 => x"982b7098",
          4800 => x"2c82d2c8",
          4801 => x"33575156",
          4802 => x"57747424",
          4803 => x"fada3888",
          4804 => x"51ffa891",
          4805 => x"3f748180",
          4806 => x"0a298180",
          4807 => x"0a057098",
          4808 => x"2c82d2c8",
          4809 => x"33585155",
          4810 => x"757525e3",
          4811 => x"38fab939",
          4812 => x"82d2c833",
          4813 => x"7a055480",
          4814 => x"74348a51",
          4815 => x"ffa7e63f",
          4816 => x"82d2c852",
          4817 => x"7951f6eb",
          4818 => x"3f82bb98",
          4819 => x"0881ff06",
          4820 => x"54739638",
          4821 => x"82d2c833",
          4822 => x"5473802e",
          4823 => x"8f388153",
          4824 => x"73527951",
          4825 => x"f2953f84",
          4826 => x"39807a34",
          4827 => x"800b82d2",
          4828 => x"cc34800b",
          4829 => x"82d2c834",
          4830 => x"7982bb98",
          4831 => x"0caf3d0d",
          4832 => x"0482d2cc",
          4833 => x"33547380",
          4834 => x"2ef9dd38",
          4835 => x"8851ffa7",
          4836 => x"943f82d2",
          4837 => x"cc33ff05",
          4838 => x"547382d2",
          4839 => x"cc347381",
          4840 => x"ff0654e2",
          4841 => x"3982d2cc",
          4842 => x"3382d2c8",
          4843 => x"33555573",
          4844 => x"752ef9b4",
          4845 => x"38ff1454",
          4846 => x"7382d2c8",
          4847 => x"3474982b",
          4848 => x"70982c75",
          4849 => x"81ff0656",
          4850 => x"51557474",
          4851 => x"25a83874",
          4852 => x"1a548114",
          4853 => x"33743473",
          4854 => x"3351ffa6",
          4855 => x"c83f7481",
          4856 => x"800a2981",
          4857 => x"800a0570",
          4858 => x"982c82d2",
          4859 => x"c8335851",
          4860 => x"55757524",
          4861 => x"da38a051",
          4862 => x"ffa6aa3f",
          4863 => x"82d2cc33",
          4864 => x"70982b70",
          4865 => x"982c82d2",
          4866 => x"c8335751",
          4867 => x"56577474",
          4868 => x"24f8d538",
          4869 => x"8851ffa6",
          4870 => x"8c3f7481",
          4871 => x"800a2981",
          4872 => x"800a0570",
          4873 => x"982c82d2",
          4874 => x"c8335851",
          4875 => x"55757525",
          4876 => x"e338f8b4",
          4877 => x"3982d2cc",
          4878 => x"337081ff",
          4879 => x"0682d2c8",
          4880 => x"33595654",
          4881 => x"747727f8",
          4882 => x"9f388114",
          4883 => x"547382d2",
          4884 => x"cc34741a",
          4885 => x"70335254",
          4886 => x"ffa5ca3f",
          4887 => x"82d2cc33",
          4888 => x"7081ff06",
          4889 => x"82d2c833",
          4890 => x"58565475",
          4891 => x"7526db38",
          4892 => x"f7f63982",
          4893 => x"d2cc5380",
          4894 => x"5282a988",
          4895 => x"51efba3f",
          4896 => x"800b82d2",
          4897 => x"cc34800b",
          4898 => x"82d2c834",
          4899 => x"f7da397a",
          4900 => x"b03882ba",
          4901 => x"e4085574",
          4902 => x"802ea638",
          4903 => x"7451ffae",
          4904 => x"843f82bb",
          4905 => x"980882d2",
          4906 => x"c83482bb",
          4907 => x"980881ff",
          4908 => x"06810553",
          4909 => x"74527951",
          4910 => x"ffafca3f",
          4911 => x"935b81c0",
          4912 => x"397a8429",
          4913 => x"82ba9805",
          4914 => x"fc110856",
          4915 => x"5474802e",
          4916 => x"a7387451",
          4917 => x"ffadce3f",
          4918 => x"82bb9808",
          4919 => x"82d2c834",
          4920 => x"82bb9808",
          4921 => x"81ff0681",
          4922 => x"05537452",
          4923 => x"7951ffaf",
          4924 => x"943fff1b",
          4925 => x"5480fa39",
          4926 => x"73085574",
          4927 => x"802ef6e8",
          4928 => x"387451ff",
          4929 => x"ad9f3f99",
          4930 => x"397a932e",
          4931 => x"098106ae",
          4932 => x"3882ba98",
          4933 => x"08557480",
          4934 => x"2ea43874",
          4935 => x"51ffad85",
          4936 => x"3f82bb98",
          4937 => x"0882d2c8",
          4938 => x"3482bb98",
          4939 => x"0881ff06",
          4940 => x"81055374",
          4941 => x"527951ff",
          4942 => x"aecb3f80",
          4943 => x"c3397a84",
          4944 => x"2982ba9c",
          4945 => x"05700856",
          4946 => x"5474802e",
          4947 => x"ab387451",
          4948 => x"ffacd23f",
          4949 => x"82bb9808",
          4950 => x"82d2c834",
          4951 => x"82bb9808",
          4952 => x"81ff0681",
          4953 => x"05537452",
          4954 => x"7951ffae",
          4955 => x"983f811b",
          4956 => x"547381ff",
          4957 => x"065b8939",
          4958 => x"7482d2c8",
          4959 => x"34747a34",
          4960 => x"82d2cc53",
          4961 => x"82d2c833",
          4962 => x"527951ed",
          4963 => x"ac3ff5d8",
          4964 => x"3982d2cc",
          4965 => x"337081ff",
          4966 => x"0682d2c8",
          4967 => x"33595654",
          4968 => x"747727f5",
          4969 => x"c3388114",
          4970 => x"547382d2",
          4971 => x"cc34741a",
          4972 => x"70335254",
          4973 => x"ffa2ee3f",
          4974 => x"f5ae3982",
          4975 => x"d2cc3354",
          4976 => x"73802ef5",
          4977 => x"a3388851",
          4978 => x"ffa2da3f",
          4979 => x"82d2cc33",
          4980 => x"ff055473",
          4981 => x"82d2cc34",
          4982 => x"f58e39f9",
          4983 => x"3d0d83c0",
          4984 => x"800b82bb",
          4985 => x"900c8480",
          4986 => x"0b82bb8c",
          4987 => x"23a08053",
          4988 => x"805283c0",
          4989 => x"8051ffb2",
          4990 => x"8d3f82bb",
          4991 => x"90085480",
          4992 => x"58777434",
          4993 => x"81577681",
          4994 => x"153482bb",
          4995 => x"90085477",
          4996 => x"84153476",
          4997 => x"85153482",
          4998 => x"bb900854",
          4999 => x"77861534",
          5000 => x"76871534",
          5001 => x"82bb9008",
          5002 => x"82bb8c22",
          5003 => x"ff05fe80",
          5004 => x"80077083",
          5005 => x"ffff0670",
          5006 => x"882a5851",
          5007 => x"55567488",
          5008 => x"17347389",
          5009 => x"173482bb",
          5010 => x"8c227088",
          5011 => x"2982bb90",
          5012 => x"0805f811",
          5013 => x"51555577",
          5014 => x"82153476",
          5015 => x"83153489",
          5016 => x"3d0d04ff",
          5017 => x"3d0d7352",
          5018 => x"81518472",
          5019 => x"278f38fb",
          5020 => x"12832a82",
          5021 => x"117083ff",
          5022 => x"ff065151",
          5023 => x"517082bb",
          5024 => x"980c833d",
          5025 => x"0d04f93d",
          5026 => x"0d02a605",
          5027 => x"22028405",
          5028 => x"aa052271",
          5029 => x"0582bb90",
          5030 => x"0871832b",
          5031 => x"71117483",
          5032 => x"2b731170",
          5033 => x"33811233",
          5034 => x"71882b07",
          5035 => x"02a405ae",
          5036 => x"05227181",
          5037 => x"ffff0607",
          5038 => x"70882a53",
          5039 => x"51525954",
          5040 => x"5b5b5753",
          5041 => x"54557177",
          5042 => x"34708118",
          5043 => x"3482bb90",
          5044 => x"08147588",
          5045 => x"2a525470",
          5046 => x"82153474",
          5047 => x"83153482",
          5048 => x"bb900870",
          5049 => x"17703381",
          5050 => x"12337188",
          5051 => x"2b077083",
          5052 => x"2b8ffff8",
          5053 => x"06515256",
          5054 => x"52710573",
          5055 => x"83ffff06",
          5056 => x"70882a54",
          5057 => x"54517182",
          5058 => x"12347281",
          5059 => x"ff065372",
          5060 => x"83123482",
          5061 => x"bb900816",
          5062 => x"56717634",
          5063 => x"72811734",
          5064 => x"893d0d04",
          5065 => x"fb3d0d82",
          5066 => x"bb900802",
          5067 => x"84059e05",
          5068 => x"2270832b",
          5069 => x"72118611",
          5070 => x"33871233",
          5071 => x"718b2b71",
          5072 => x"832b0758",
          5073 => x"5b595255",
          5074 => x"52720584",
          5075 => x"12338513",
          5076 => x"3371882b",
          5077 => x"0770882a",
          5078 => x"54565652",
          5079 => x"70841334",
          5080 => x"73851334",
          5081 => x"82bb9008",
          5082 => x"70148411",
          5083 => x"33851233",
          5084 => x"718b2b71",
          5085 => x"832b0756",
          5086 => x"59575272",
          5087 => x"05861233",
          5088 => x"87133371",
          5089 => x"882b0770",
          5090 => x"882a5456",
          5091 => x"56527086",
          5092 => x"13347387",
          5093 => x"133482bb",
          5094 => x"90081370",
          5095 => x"33811233",
          5096 => x"71882b07",
          5097 => x"7081ffff",
          5098 => x"0670882a",
          5099 => x"53515353",
          5100 => x"53717334",
          5101 => x"70811434",
          5102 => x"873d0d04",
          5103 => x"fa3d0d02",
          5104 => x"a2052282",
          5105 => x"bb900871",
          5106 => x"832b7111",
          5107 => x"70338112",
          5108 => x"3371882b",
          5109 => x"07708829",
          5110 => x"15703381",
          5111 => x"12337198",
          5112 => x"2b71902b",
          5113 => x"07535f53",
          5114 => x"55525a56",
          5115 => x"57535471",
          5116 => x"802580f6",
          5117 => x"387251fe",
          5118 => x"ab3f82bb",
          5119 => x"90087016",
          5120 => x"70338112",
          5121 => x"33718b2b",
          5122 => x"71832b07",
          5123 => x"74117033",
          5124 => x"81123371",
          5125 => x"882b0770",
          5126 => x"832b8fff",
          5127 => x"f8065152",
          5128 => x"5451535a",
          5129 => x"58537205",
          5130 => x"74882a54",
          5131 => x"52728213",
          5132 => x"34738313",
          5133 => x"3482bb90",
          5134 => x"08701670",
          5135 => x"33811233",
          5136 => x"718b2b71",
          5137 => x"832b0756",
          5138 => x"59575572",
          5139 => x"05703381",
          5140 => x"12337188",
          5141 => x"2b077081",
          5142 => x"ffff0670",
          5143 => x"882a5751",
          5144 => x"52585272",
          5145 => x"74347181",
          5146 => x"1534883d",
          5147 => x"0d04fb3d",
          5148 => x"0d82bb90",
          5149 => x"08028405",
          5150 => x"9e052270",
          5151 => x"832b7211",
          5152 => x"82113383",
          5153 => x"1233718b",
          5154 => x"2b71832b",
          5155 => x"07595b59",
          5156 => x"52565273",
          5157 => x"05713381",
          5158 => x"13337188",
          5159 => x"2b07028c",
          5160 => x"05a20522",
          5161 => x"71077088",
          5162 => x"2a535153",
          5163 => x"53537173",
          5164 => x"34708114",
          5165 => x"3482bb90",
          5166 => x"08701570",
          5167 => x"33811233",
          5168 => x"718b2b71",
          5169 => x"832b0756",
          5170 => x"59575272",
          5171 => x"05821233",
          5172 => x"83133371",
          5173 => x"882b0770",
          5174 => x"882a5455",
          5175 => x"56527082",
          5176 => x"13347283",
          5177 => x"133482bb",
          5178 => x"90081482",
          5179 => x"11338312",
          5180 => x"3371882b",
          5181 => x"0782bb98",
          5182 => x"0c525487",
          5183 => x"3d0d04f7",
          5184 => x"3d0d7b82",
          5185 => x"bb900831",
          5186 => x"832a7083",
          5187 => x"ffff0670",
          5188 => x"535753fd",
          5189 => x"a73f82bb",
          5190 => x"90087683",
          5191 => x"2b711182",
          5192 => x"11338312",
          5193 => x"33718b2b",
          5194 => x"71832b07",
          5195 => x"75117033",
          5196 => x"81123371",
          5197 => x"982b7190",
          5198 => x"2b075342",
          5199 => x"4051535b",
          5200 => x"58555954",
          5201 => x"7280258d",
          5202 => x"38828080",
          5203 => x"527551fe",
          5204 => x"9d3f8184",
          5205 => x"39841433",
          5206 => x"85153371",
          5207 => x"8b2b7183",
          5208 => x"2b077611",
          5209 => x"79882a53",
          5210 => x"51555855",
          5211 => x"76861434",
          5212 => x"7581ff06",
          5213 => x"56758714",
          5214 => x"3482bb90",
          5215 => x"08701984",
          5216 => x"12338513",
          5217 => x"3371882b",
          5218 => x"0770882a",
          5219 => x"54575b56",
          5220 => x"53728416",
          5221 => x"34738516",
          5222 => x"3482bb90",
          5223 => x"08185380",
          5224 => x"0b861434",
          5225 => x"800b8714",
          5226 => x"3482bb90",
          5227 => x"08537684",
          5228 => x"14347585",
          5229 => x"143482bb",
          5230 => x"90081870",
          5231 => x"33811233",
          5232 => x"71882b07",
          5233 => x"70828080",
          5234 => x"0770882a",
          5235 => x"53515556",
          5236 => x"54747434",
          5237 => x"72811534",
          5238 => x"8b3d0d04",
          5239 => x"ff3d0d73",
          5240 => x"5282bb90",
          5241 => x"088438f7",
          5242 => x"f23f7180",
          5243 => x"2e863871",
          5244 => x"51fe8c3f",
          5245 => x"833d0d04",
          5246 => x"f53d0d80",
          5247 => x"7e5258f8",
          5248 => x"e23f82bb",
          5249 => x"980883ff",
          5250 => x"ff0682bb",
          5251 => x"90088411",
          5252 => x"33851233",
          5253 => x"71882b07",
          5254 => x"705f5956",
          5255 => x"585a81ff",
          5256 => x"ff597578",
          5257 => x"2e80cb38",
          5258 => x"75882917",
          5259 => x"70338112",
          5260 => x"3371882b",
          5261 => x"077081ff",
          5262 => x"ff067931",
          5263 => x"7083ffff",
          5264 => x"06707f27",
          5265 => x"52535156",
          5266 => x"59557779",
          5267 => x"278a3873",
          5268 => x"802e8538",
          5269 => x"75785a5b",
          5270 => x"84153385",
          5271 => x"16337188",
          5272 => x"2b075754",
          5273 => x"75c23878",
          5274 => x"81ffff2e",
          5275 => x"85387a79",
          5276 => x"59568076",
          5277 => x"832b82bb",
          5278 => x"90081170",
          5279 => x"33811233",
          5280 => x"71882b07",
          5281 => x"7081ffff",
          5282 => x"0651525a",
          5283 => x"565c5573",
          5284 => x"752e8338",
          5285 => x"81558054",
          5286 => x"79782681",
          5287 => x"cc387454",
          5288 => x"74802e81",
          5289 => x"c438777a",
          5290 => x"2e098106",
          5291 => x"89387551",
          5292 => x"f8f23f81",
          5293 => x"ac398280",
          5294 => x"80537952",
          5295 => x"7551f7c6",
          5296 => x"3f82bb90",
          5297 => x"08701c86",
          5298 => x"11338712",
          5299 => x"33718b2b",
          5300 => x"71832b07",
          5301 => x"535a5e55",
          5302 => x"74057a17",
          5303 => x"7083ffff",
          5304 => x"0670882a",
          5305 => x"5c595654",
          5306 => x"78841534",
          5307 => x"7681ff06",
          5308 => x"57768515",
          5309 => x"3482bb90",
          5310 => x"0875832b",
          5311 => x"7111721e",
          5312 => x"86113387",
          5313 => x"12337188",
          5314 => x"2b077088",
          5315 => x"2a535b5e",
          5316 => x"535a5654",
          5317 => x"73861934",
          5318 => x"75871934",
          5319 => x"82bb9008",
          5320 => x"701c8411",
          5321 => x"33851233",
          5322 => x"718b2b71",
          5323 => x"832b0753",
          5324 => x"5d5a5574",
          5325 => x"05547886",
          5326 => x"15347687",
          5327 => x"153482bb",
          5328 => x"90087016",
          5329 => x"711d8411",
          5330 => x"33851233",
          5331 => x"71882b07",
          5332 => x"70882a53",
          5333 => x"5a5f5256",
          5334 => x"54738416",
          5335 => x"34758516",
          5336 => x"3482bb90",
          5337 => x"081b8405",
          5338 => x"547382bb",
          5339 => x"980c8d3d",
          5340 => x"0d04fe3d",
          5341 => x"0d745282",
          5342 => x"bb900884",
          5343 => x"38f4dc3f",
          5344 => x"71537180",
          5345 => x"2e8b3871",
          5346 => x"51fced3f",
          5347 => x"82bb9808",
          5348 => x"537282bb",
          5349 => x"980c843d",
          5350 => x"0d04ee3d",
          5351 => x"0d646640",
          5352 => x"5c807042",
          5353 => x"4082bb90",
          5354 => x"08602e09",
          5355 => x"81068438",
          5356 => x"f4a93f7b",
          5357 => x"8e387e51",
          5358 => x"ffb83f82",
          5359 => x"bb980854",
          5360 => x"83c7397e",
          5361 => x"8b387b51",
          5362 => x"fc923f7e",
          5363 => x"5483ba39",
          5364 => x"7e51f58f",
          5365 => x"3f82bb98",
          5366 => x"0883ffff",
          5367 => x"0682bb90",
          5368 => x"087d7131",
          5369 => x"832a7083",
          5370 => x"ffff0670",
          5371 => x"832b7311",
          5372 => x"70338112",
          5373 => x"3371882b",
          5374 => x"07707531",
          5375 => x"7083ffff",
          5376 => x"06708829",
          5377 => x"fc057388",
          5378 => x"291a7033",
          5379 => x"81123371",
          5380 => x"882b0770",
          5381 => x"902b5344",
          5382 => x"4e534841",
          5383 => x"525c545b",
          5384 => x"415c565b",
          5385 => x"5b738025",
          5386 => x"8f387681",
          5387 => x"ffff0675",
          5388 => x"317083ff",
          5389 => x"ff064254",
          5390 => x"82163383",
          5391 => x"17337188",
          5392 => x"2b077088",
          5393 => x"291c7033",
          5394 => x"81123371",
          5395 => x"982b7190",
          5396 => x"2b075347",
          5397 => x"45525654",
          5398 => x"7380258b",
          5399 => x"38787531",
          5400 => x"7083ffff",
          5401 => x"06415477",
          5402 => x"7b2781fe",
          5403 => x"38601854",
          5404 => x"737b2e09",
          5405 => x"81068f38",
          5406 => x"7851f6c0",
          5407 => x"3f7a83ff",
          5408 => x"ff065881",
          5409 => x"e5397f8e",
          5410 => x"387a7424",
          5411 => x"89387851",
          5412 => x"f6aa3f81",
          5413 => x"a5397f18",
          5414 => x"557a7524",
          5415 => x"80c83879",
          5416 => x"1d821133",
          5417 => x"83123371",
          5418 => x"882b0753",
          5419 => x"5754f4f4",
          5420 => x"3f805278",
          5421 => x"51f7b73f",
          5422 => x"82bb9808",
          5423 => x"83ffff06",
          5424 => x"7e547c53",
          5425 => x"70832b82",
          5426 => x"bb900811",
          5427 => x"84055355",
          5428 => x"59ff9ae7",
          5429 => x"3f82bb90",
          5430 => x"08148405",
          5431 => x"7583ffff",
          5432 => x"06595c81",
          5433 => x"85396015",
          5434 => x"547a7424",
          5435 => x"80d43878",
          5436 => x"51f5c93f",
          5437 => x"82bb9008",
          5438 => x"1d821133",
          5439 => x"83123371",
          5440 => x"882b0753",
          5441 => x"4354f49c",
          5442 => x"3f805278",
          5443 => x"51f6df3f",
          5444 => x"82bb9808",
          5445 => x"83ffff06",
          5446 => x"7e547c53",
          5447 => x"70832b82",
          5448 => x"bb900811",
          5449 => x"84055355",
          5450 => x"59ff9a8f",
          5451 => x"3f82bb90",
          5452 => x"08148405",
          5453 => x"60620519",
          5454 => x"555c7383",
          5455 => x"ffff0658",
          5456 => x"a9397b7f",
          5457 => x"5254f9b0",
          5458 => x"3f82bb98",
          5459 => x"085c82bb",
          5460 => x"9808802e",
          5461 => x"93387d53",
          5462 => x"735282bb",
          5463 => x"980851ff",
          5464 => x"9ea33f73",
          5465 => x"51f7983f",
          5466 => x"7a587a78",
          5467 => x"27993880",
          5468 => x"537a5278",
          5469 => x"51f28f3f",
          5470 => x"7a19832b",
          5471 => x"82bb9008",
          5472 => x"05840551",
          5473 => x"f6f93f7b",
          5474 => x"547382bb",
          5475 => x"980c943d",
          5476 => x"0d04fc3d",
          5477 => x"0d777729",
          5478 => x"705254fb",
          5479 => x"d53f82bb",
          5480 => x"98085582",
          5481 => x"bb980880",
          5482 => x"2e8e3873",
          5483 => x"53805282",
          5484 => x"bb980851",
          5485 => x"ffa2cf3f",
          5486 => x"7482bb98",
          5487 => x"0c863d0d",
          5488 => x"04ff3d0d",
          5489 => x"028f0533",
          5490 => x"51815270",
          5491 => x"72268738",
          5492 => x"82bb9411",
          5493 => x"33527182",
          5494 => x"bb980c83",
          5495 => x"3d0d04fc",
          5496 => x"3d0d029b",
          5497 => x"05330284",
          5498 => x"059f0533",
          5499 => x"56538351",
          5500 => x"72812680",
          5501 => x"e0387284",
          5502 => x"2b87c092",
          5503 => x"8c115351",
          5504 => x"88547480",
          5505 => x"2e843881",
          5506 => x"88547372",
          5507 => x"0c87c092",
          5508 => x"8c115181",
          5509 => x"710c850b",
          5510 => x"87c0988c",
          5511 => x"0c705271",
          5512 => x"08708206",
          5513 => x"51517080",
          5514 => x"2e8a3887",
          5515 => x"c0988c08",
          5516 => x"5170ec38",
          5517 => x"7108fc80",
          5518 => x"80065271",
          5519 => x"923887c0",
          5520 => x"988c0851",
          5521 => x"70802e87",
          5522 => x"387182bb",
          5523 => x"94143482",
          5524 => x"bb941333",
          5525 => x"517082bb",
          5526 => x"980c863d",
          5527 => x"0d04f33d",
          5528 => x"0d606264",
          5529 => x"028c05bf",
          5530 => x"05335740",
          5531 => x"585b8374",
          5532 => x"525afecd",
          5533 => x"3f82bb98",
          5534 => x"0881067a",
          5535 => x"54527181",
          5536 => x"be387172",
          5537 => x"75842b87",
          5538 => x"c0928011",
          5539 => x"87c0928c",
          5540 => x"1287c092",
          5541 => x"8413415a",
          5542 => x"40575a58",
          5543 => x"850b87c0",
          5544 => x"988c0c76",
          5545 => x"7d0c8476",
          5546 => x"0c750870",
          5547 => x"852a7081",
          5548 => x"06515354",
          5549 => x"71802e8e",
          5550 => x"387b0852",
          5551 => x"717b7081",
          5552 => x"055d3481",
          5553 => x"19598074",
          5554 => x"a2065353",
          5555 => x"71732e83",
          5556 => x"38815378",
          5557 => x"83ff268f",
          5558 => x"3872802e",
          5559 => x"8a3887c0",
          5560 => x"988c0852",
          5561 => x"71c33887",
          5562 => x"c0988c08",
          5563 => x"5271802e",
          5564 => x"87387884",
          5565 => x"802e9938",
          5566 => x"81760c87",
          5567 => x"c0928c15",
          5568 => x"53720870",
          5569 => x"82065152",
          5570 => x"71f738ff",
          5571 => x"1a5a8d39",
          5572 => x"84801781",
          5573 => x"197081ff",
          5574 => x"065a5357",
          5575 => x"79802e90",
          5576 => x"3873fc80",
          5577 => x"80065271",
          5578 => x"87387d78",
          5579 => x"26feed38",
          5580 => x"73fc8080",
          5581 => x"06527180",
          5582 => x"2e833881",
          5583 => x"52715372",
          5584 => x"82bb980c",
          5585 => x"8f3d0d04",
          5586 => x"f33d0d60",
          5587 => x"6264028c",
          5588 => x"05bf0533",
          5589 => x"5740585b",
          5590 => x"83598074",
          5591 => x"5258fce1",
          5592 => x"3f82bb98",
          5593 => x"08810679",
          5594 => x"54527178",
          5595 => x"2e098106",
          5596 => x"81b13877",
          5597 => x"74842b87",
          5598 => x"c0928011",
          5599 => x"87c0928c",
          5600 => x"1287c092",
          5601 => x"84134059",
          5602 => x"5f565a85",
          5603 => x"0b87c098",
          5604 => x"8c0c767d",
          5605 => x"0c82760c",
          5606 => x"80587508",
          5607 => x"70842a70",
          5608 => x"81065153",
          5609 => x"5471802e",
          5610 => x"8c387a70",
          5611 => x"81055c33",
          5612 => x"7c0c8118",
          5613 => x"5873812a",
          5614 => x"70810651",
          5615 => x"5271802e",
          5616 => x"8a3887c0",
          5617 => x"988c0852",
          5618 => x"71d03887",
          5619 => x"c0988c08",
          5620 => x"5271802e",
          5621 => x"87387784",
          5622 => x"802e9938",
          5623 => x"81760c87",
          5624 => x"c0928c15",
          5625 => x"53720870",
          5626 => x"82065152",
          5627 => x"71f738ff",
          5628 => x"19598d39",
          5629 => x"811a7081",
          5630 => x"ff068480",
          5631 => x"19595b52",
          5632 => x"78802e90",
          5633 => x"3873fc80",
          5634 => x"80065271",
          5635 => x"87387d7a",
          5636 => x"26fef838",
          5637 => x"73fc8080",
          5638 => x"06527180",
          5639 => x"2e833881",
          5640 => x"52715372",
          5641 => x"82bb980c",
          5642 => x"8f3d0d04",
          5643 => x"fa3d0d7a",
          5644 => x"028405a3",
          5645 => x"05330288",
          5646 => x"05a70533",
          5647 => x"71545456",
          5648 => x"57fafe3f",
          5649 => x"82bb9808",
          5650 => x"81065383",
          5651 => x"547280fe",
          5652 => x"38850b87",
          5653 => x"c0988c0c",
          5654 => x"81567176",
          5655 => x"2e80dc38",
          5656 => x"71762493",
          5657 => x"3874842b",
          5658 => x"87c0928c",
          5659 => x"11545471",
          5660 => x"802e8d38",
          5661 => x"80d43971",
          5662 => x"832e80c6",
          5663 => x"3880cb39",
          5664 => x"72087081",
          5665 => x"2a708106",
          5666 => x"51515271",
          5667 => x"802e8a38",
          5668 => x"87c0988c",
          5669 => x"085271e8",
          5670 => x"3887c098",
          5671 => x"8c085271",
          5672 => x"96388173",
          5673 => x"0c87c092",
          5674 => x"8c145372",
          5675 => x"08708206",
          5676 => x"515271f7",
          5677 => x"38963980",
          5678 => x"56923988",
          5679 => x"800a770c",
          5680 => x"85398180",
          5681 => x"770c7256",
          5682 => x"83398456",
          5683 => x"75547382",
          5684 => x"bb980c88",
          5685 => x"3d0d04fe",
          5686 => x"3d0d7481",
          5687 => x"11337133",
          5688 => x"71882b07",
          5689 => x"82bb980c",
          5690 => x"5351843d",
          5691 => x"0d04fd3d",
          5692 => x"0d758311",
          5693 => x"33821233",
          5694 => x"71902b71",
          5695 => x"882b0781",
          5696 => x"14337072",
          5697 => x"07882b75",
          5698 => x"33710782",
          5699 => x"bb980c52",
          5700 => x"53545654",
          5701 => x"52853d0d",
          5702 => x"04ff3d0d",
          5703 => x"73028405",
          5704 => x"92052252",
          5705 => x"52707270",
          5706 => x"81055434",
          5707 => x"70882a51",
          5708 => x"70723483",
          5709 => x"3d0d04ff",
          5710 => x"3d0d7375",
          5711 => x"52527072",
          5712 => x"70810554",
          5713 => x"3470882a",
          5714 => x"51707270",
          5715 => x"81055434",
          5716 => x"70882a51",
          5717 => x"70727081",
          5718 => x"05543470",
          5719 => x"882a5170",
          5720 => x"7234833d",
          5721 => x"0d04fe3d",
          5722 => x"0d767577",
          5723 => x"54545170",
          5724 => x"802e9238",
          5725 => x"71708105",
          5726 => x"53337370",
          5727 => x"81055534",
          5728 => x"ff1151eb",
          5729 => x"39843d0d",
          5730 => x"04fe3d0d",
          5731 => x"75777654",
          5732 => x"52537272",
          5733 => x"70810554",
          5734 => x"34ff1151",
          5735 => x"70f43884",
          5736 => x"3d0d04fc",
          5737 => x"3d0d7877",
          5738 => x"79565653",
          5739 => x"74708105",
          5740 => x"56337470",
          5741 => x"81055633",
          5742 => x"717131ff",
          5743 => x"16565252",
          5744 => x"5272802e",
          5745 => x"86387180",
          5746 => x"2ee23871",
          5747 => x"82bb980c",
          5748 => x"863d0d04",
          5749 => x"fe3d0d74",
          5750 => x"76545189",
          5751 => x"3971732e",
          5752 => x"8a388111",
          5753 => x"51703352",
          5754 => x"71f33870",
          5755 => x"3382bb98",
          5756 => x"0c843d0d",
          5757 => x"04800b82",
          5758 => x"bb980c04",
          5759 => x"800b82bb",
          5760 => x"980c04f7",
          5761 => x"3d0d7b56",
          5762 => x"800b8317",
          5763 => x"33565a74",
          5764 => x"7a2e80d6",
          5765 => x"388154b0",
          5766 => x"160853b4",
          5767 => x"16705381",
          5768 => x"17335259",
          5769 => x"faa23f82",
          5770 => x"bb98087a",
          5771 => x"2e098106",
          5772 => x"b73882bb",
          5773 => x"98088317",
          5774 => x"34b01608",
          5775 => x"70a41808",
          5776 => x"319c1808",
          5777 => x"59565874",
          5778 => x"77279f38",
          5779 => x"82163355",
          5780 => x"74822e09",
          5781 => x"81069338",
          5782 => x"81547618",
          5783 => x"53785281",
          5784 => x"163351f9",
          5785 => x"e33f8339",
          5786 => x"815a7982",
          5787 => x"bb980c8b",
          5788 => x"3d0d04fa",
          5789 => x"3d0d787a",
          5790 => x"56568057",
          5791 => x"74b01708",
          5792 => x"2eaf3875",
          5793 => x"51fefc3f",
          5794 => x"82bb9808",
          5795 => x"5782bb98",
          5796 => x"089f3881",
          5797 => x"547453b4",
          5798 => x"16528116",
          5799 => x"3351f7be",
          5800 => x"3f82bb98",
          5801 => x"08802e85",
          5802 => x"38ff5581",
          5803 => x"5774b017",
          5804 => x"0c7682bb",
          5805 => x"980c883d",
          5806 => x"0d04f83d",
          5807 => x"0d7a7052",
          5808 => x"57fec03f",
          5809 => x"82bb9808",
          5810 => x"5882bb98",
          5811 => x"08819138",
          5812 => x"76335574",
          5813 => x"832e0981",
          5814 => x"0680f038",
          5815 => x"84173359",
          5816 => x"78812e09",
          5817 => x"810680e3",
          5818 => x"38848053",
          5819 => x"82bb9808",
          5820 => x"52b41770",
          5821 => x"5256fd91",
          5822 => x"3f82d4d5",
          5823 => x"5284b217",
          5824 => x"51fc963f",
          5825 => x"848b85a4",
          5826 => x"d2527551",
          5827 => x"fca93f86",
          5828 => x"8a85e4f2",
          5829 => x"52849817",
          5830 => x"51fc9c3f",
          5831 => x"90170852",
          5832 => x"849c1751",
          5833 => x"fc913f8c",
          5834 => x"17085284",
          5835 => x"a01751fc",
          5836 => x"863fa017",
          5837 => x"08810570",
          5838 => x"b0190c79",
          5839 => x"55537552",
          5840 => x"81173351",
          5841 => x"f8823f77",
          5842 => x"84183480",
          5843 => x"53805281",
          5844 => x"173351f9",
          5845 => x"d73f82bb",
          5846 => x"9808802e",
          5847 => x"83388158",
          5848 => x"7782bb98",
          5849 => x"0c8a3d0d",
          5850 => x"04fb3d0d",
          5851 => x"77fe1a98",
          5852 => x"1208fe05",
          5853 => x"55565480",
          5854 => x"56747327",
          5855 => x"8d388a14",
          5856 => x"22757129",
          5857 => x"ac160805",
          5858 => x"57537582",
          5859 => x"bb980c87",
          5860 => x"3d0d04f9",
          5861 => x"3d0d7a7a",
          5862 => x"70085654",
          5863 => x"57817727",
          5864 => x"81df3876",
          5865 => x"98150827",
          5866 => x"81d738ff",
          5867 => x"74335458",
          5868 => x"72822e80",
          5869 => x"f5387282",
          5870 => x"24893872",
          5871 => x"812e8d38",
          5872 => x"81bf3972",
          5873 => x"832e818e",
          5874 => x"3881b639",
          5875 => x"76812a17",
          5876 => x"70892aa4",
          5877 => x"16080553",
          5878 => x"745255fd",
          5879 => x"963f82bb",
          5880 => x"9808819f",
          5881 => x"387483ff",
          5882 => x"0614b411",
          5883 => x"33811770",
          5884 => x"892aa418",
          5885 => x"08055576",
          5886 => x"54575753",
          5887 => x"fcf53f82",
          5888 => x"bb980880",
          5889 => x"fe387483",
          5890 => x"ff0614b4",
          5891 => x"11337088",
          5892 => x"2b780779",
          5893 => x"81067184",
          5894 => x"2a5c5258",
          5895 => x"51537280",
          5896 => x"e238759f",
          5897 => x"ff065880",
          5898 => x"da397688",
          5899 => x"2aa41508",
          5900 => x"05527351",
          5901 => x"fcbd3f82",
          5902 => x"bb980880",
          5903 => x"c6387610",
          5904 => x"83fe0674",
          5905 => x"05b40551",
          5906 => x"f98d3f82",
          5907 => x"bb980883",
          5908 => x"ffff0658",
          5909 => x"ae397687",
          5910 => x"2aa41508",
          5911 => x"05527351",
          5912 => x"fc913f82",
          5913 => x"bb98089b",
          5914 => x"3876822b",
          5915 => x"83fc0674",
          5916 => x"05b40551",
          5917 => x"f8f83f82",
          5918 => x"bb9808f0",
          5919 => x"0a065883",
          5920 => x"39815877",
          5921 => x"82bb980c",
          5922 => x"893d0d04",
          5923 => x"f83d0d7a",
          5924 => x"7c7e5a58",
          5925 => x"56825981",
          5926 => x"7727829e",
          5927 => x"38769817",
          5928 => x"08278296",
          5929 => x"38753353",
          5930 => x"72792e81",
          5931 => x"9d387279",
          5932 => x"24893872",
          5933 => x"812e8d38",
          5934 => x"82803972",
          5935 => x"832e81b8",
          5936 => x"3881f739",
          5937 => x"76812a17",
          5938 => x"70892aa4",
          5939 => x"18080553",
          5940 => x"765255fb",
          5941 => x"9e3f82bb",
          5942 => x"98085982",
          5943 => x"bb980881",
          5944 => x"d9387483",
          5945 => x"ff0616b4",
          5946 => x"05811678",
          5947 => x"81065956",
          5948 => x"54775376",
          5949 => x"802e8f38",
          5950 => x"77842b9f",
          5951 => x"f0067433",
          5952 => x"8f067107",
          5953 => x"51537274",
          5954 => x"34810b83",
          5955 => x"17347489",
          5956 => x"2aa41708",
          5957 => x"05527551",
          5958 => x"fad93f82",
          5959 => x"bb980859",
          5960 => x"82bb9808",
          5961 => x"81943874",
          5962 => x"83ff0616",
          5963 => x"b4057884",
          5964 => x"2a545476",
          5965 => x"8f387788",
          5966 => x"2a743381",
          5967 => x"f006718f",
          5968 => x"06075153",
          5969 => x"72743480",
          5970 => x"ec397688",
          5971 => x"2aa41708",
          5972 => x"05527551",
          5973 => x"fa9d3f82",
          5974 => x"bb980859",
          5975 => x"82bb9808",
          5976 => x"80d83877",
          5977 => x"83ffff06",
          5978 => x"52761083",
          5979 => x"fe067605",
          5980 => x"b40551f7",
          5981 => x"a43fbe39",
          5982 => x"76872aa4",
          5983 => x"17080552",
          5984 => x"7551f9ef",
          5985 => x"3f82bb98",
          5986 => x"085982bb",
          5987 => x"9808ab38",
          5988 => x"77f00a06",
          5989 => x"77822b83",
          5990 => x"fc067018",
          5991 => x"b4057054",
          5992 => x"515454f6",
          5993 => x"c93f82bb",
          5994 => x"98088f0a",
          5995 => x"06740752",
          5996 => x"7251f783",
          5997 => x"3f810b83",
          5998 => x"17347882",
          5999 => x"bb980c8a",
          6000 => x"3d0d04f8",
          6001 => x"3d0d7a7c",
          6002 => x"7e720859",
          6003 => x"56565981",
          6004 => x"7527a438",
          6005 => x"74981708",
          6006 => x"279d3873",
          6007 => x"802eaa38",
          6008 => x"ff537352",
          6009 => x"7551fda4",
          6010 => x"3f82bb98",
          6011 => x"085482bb",
          6012 => x"980880f2",
          6013 => x"38933982",
          6014 => x"5480eb39",
          6015 => x"815480e6",
          6016 => x"3982bb98",
          6017 => x"085480de",
          6018 => x"39745278",
          6019 => x"51fb843f",
          6020 => x"82bb9808",
          6021 => x"5882bb98",
          6022 => x"08802e80",
          6023 => x"c73882bb",
          6024 => x"9808812e",
          6025 => x"d23882bb",
          6026 => x"9808ff2e",
          6027 => x"cf388053",
          6028 => x"74527551",
          6029 => x"fcd63f82",
          6030 => x"bb9808c5",
          6031 => x"38981608",
          6032 => x"fe119018",
          6033 => x"08575557",
          6034 => x"74742790",
          6035 => x"38811590",
          6036 => x"170c8416",
          6037 => x"33810754",
          6038 => x"73841734",
          6039 => x"77557678",
          6040 => x"26ffa638",
          6041 => x"80547382",
          6042 => x"bb980c8a",
          6043 => x"3d0d04f6",
          6044 => x"3d0d7c7e",
          6045 => x"7108595b",
          6046 => x"5b799538",
          6047 => x"8c170858",
          6048 => x"77802e88",
          6049 => x"38981708",
          6050 => x"7826b238",
          6051 => x"8158ae39",
          6052 => x"79527a51",
          6053 => x"f9fd3f81",
          6054 => x"557482bb",
          6055 => x"98082782",
          6056 => x"e03882bb",
          6057 => x"98085582",
          6058 => x"bb9808ff",
          6059 => x"2e82d238",
          6060 => x"98170882",
          6061 => x"bb980826",
          6062 => x"82c73879",
          6063 => x"58901708",
          6064 => x"70565473",
          6065 => x"802e82b9",
          6066 => x"38777a2e",
          6067 => x"09810680",
          6068 => x"e238811a",
          6069 => x"56981708",
          6070 => x"76268338",
          6071 => x"82567552",
          6072 => x"7a51f9af",
          6073 => x"3f805982",
          6074 => x"bb980881",
          6075 => x"2e098106",
          6076 => x"863882bb",
          6077 => x"98085982",
          6078 => x"bb980809",
          6079 => x"70307072",
          6080 => x"07802570",
          6081 => x"7c0782bb",
          6082 => x"98085451",
          6083 => x"51555573",
          6084 => x"81ef3882",
          6085 => x"bb980880",
          6086 => x"2e95388c",
          6087 => x"17085481",
          6088 => x"74279038",
          6089 => x"73981808",
          6090 => x"27893873",
          6091 => x"58853975",
          6092 => x"80db3877",
          6093 => x"56811656",
          6094 => x"98170876",
          6095 => x"26893882",
          6096 => x"56757826",
          6097 => x"81ac3875",
          6098 => x"527a51f8",
          6099 => x"c63f82bb",
          6100 => x"9808802e",
          6101 => x"b8388059",
          6102 => x"82bb9808",
          6103 => x"812e0981",
          6104 => x"06863882",
          6105 => x"bb980859",
          6106 => x"82bb9808",
          6107 => x"09703070",
          6108 => x"72078025",
          6109 => x"707c0751",
          6110 => x"51555573",
          6111 => x"80f83875",
          6112 => x"782e0981",
          6113 => x"06ffae38",
          6114 => x"735580f5",
          6115 => x"39ff5375",
          6116 => x"527651f9",
          6117 => x"f73f82bb",
          6118 => x"980882bb",
          6119 => x"98083070",
          6120 => x"82bb9808",
          6121 => x"07802551",
          6122 => x"55557980",
          6123 => x"2e943873",
          6124 => x"802e8f38",
          6125 => x"75537952",
          6126 => x"7651f9d0",
          6127 => x"3f82bb98",
          6128 => x"085574a5",
          6129 => x"38758c18",
          6130 => x"0c981708",
          6131 => x"fe059018",
          6132 => x"08565474",
          6133 => x"74268638",
          6134 => x"ff159018",
          6135 => x"0c841733",
          6136 => x"81075473",
          6137 => x"84183497",
          6138 => x"39ff5674",
          6139 => x"812e9038",
          6140 => x"8c398055",
          6141 => x"8c3982bb",
          6142 => x"98085585",
          6143 => x"39815675",
          6144 => x"557482bb",
          6145 => x"980c8c3d",
          6146 => x"0d04f83d",
          6147 => x"0d7a7052",
          6148 => x"55f3f03f",
          6149 => x"82bb9808",
          6150 => x"58815682",
          6151 => x"bb980880",
          6152 => x"d8387b52",
          6153 => x"7451f6c1",
          6154 => x"3f82bb98",
          6155 => x"0882bb98",
          6156 => x"08b0170c",
          6157 => x"59848053",
          6158 => x"7752b415",
          6159 => x"705257f2",
          6160 => x"c83f7756",
          6161 => x"84398116",
          6162 => x"568a1522",
          6163 => x"58757827",
          6164 => x"97388154",
          6165 => x"75195376",
          6166 => x"52811533",
          6167 => x"51ede93f",
          6168 => x"82bb9808",
          6169 => x"802edf38",
          6170 => x"8a152276",
          6171 => x"32703070",
          6172 => x"7207709f",
          6173 => x"2a535156",
          6174 => x"567582bb",
          6175 => x"980c8a3d",
          6176 => x"0d04f83d",
          6177 => x"0d7a7c71",
          6178 => x"08585657",
          6179 => x"74f0800a",
          6180 => x"2680f138",
          6181 => x"749f0653",
          6182 => x"7280e938",
          6183 => x"7490180c",
          6184 => x"88170854",
          6185 => x"73aa3875",
          6186 => x"33538273",
          6187 => x"278838a8",
          6188 => x"16085473",
          6189 => x"9b387485",
          6190 => x"2a53820b",
          6191 => x"8817225a",
          6192 => x"58727927",
          6193 => x"80fe38a8",
          6194 => x"16089818",
          6195 => x"0c80cd39",
          6196 => x"8a162270",
          6197 => x"892b5458",
          6198 => x"727526b2",
          6199 => x"38735276",
          6200 => x"51f5b03f",
          6201 => x"82bb9808",
          6202 => x"5482bb98",
          6203 => x"08ff2ebd",
          6204 => x"38810b82",
          6205 => x"bb980827",
          6206 => x"8b389816",
          6207 => x"0882bb98",
          6208 => x"08268538",
          6209 => x"8258bd39",
          6210 => x"74733155",
          6211 => x"cb397352",
          6212 => x"7551f4d5",
          6213 => x"3f82bb98",
          6214 => x"0898180c",
          6215 => x"7394180c",
          6216 => x"98170853",
          6217 => x"82587280",
          6218 => x"2e9a3885",
          6219 => x"39815894",
          6220 => x"3974892a",
          6221 => x"1398180c",
          6222 => x"7483ff06",
          6223 => x"16b4059c",
          6224 => x"180c8058",
          6225 => x"7782bb98",
          6226 => x"0c8a3d0d",
          6227 => x"04f83d0d",
          6228 => x"7a700890",
          6229 => x"1208a005",
          6230 => x"595754f0",
          6231 => x"800a7727",
          6232 => x"8638800b",
          6233 => x"98150c98",
          6234 => x"14085384",
          6235 => x"5572802e",
          6236 => x"81cb3876",
          6237 => x"83ff0658",
          6238 => x"7781b538",
          6239 => x"81139815",
          6240 => x"0c941408",
          6241 => x"55749238",
          6242 => x"76852a88",
          6243 => x"17225653",
          6244 => x"74732681",
          6245 => x"9b3880c0",
          6246 => x"398a1622",
          6247 => x"ff057789",
          6248 => x"2a065372",
          6249 => x"818a3874",
          6250 => x"527351f3",
          6251 => x"e63f82bb",
          6252 => x"98085382",
          6253 => x"55810b82",
          6254 => x"bb980827",
          6255 => x"80ff3881",
          6256 => x"5582bb98",
          6257 => x"08ff2e80",
          6258 => x"f4389816",
          6259 => x"0882bb98",
          6260 => x"082680ca",
          6261 => x"387b8a38",
          6262 => x"7798150c",
          6263 => x"845580dd",
          6264 => x"39941408",
          6265 => x"527351f9",
          6266 => x"863f82bb",
          6267 => x"98085387",
          6268 => x"5582bb98",
          6269 => x"08802e80",
          6270 => x"c4388255",
          6271 => x"82bb9808",
          6272 => x"812eba38",
          6273 => x"815582bb",
          6274 => x"9808ff2e",
          6275 => x"b03882bb",
          6276 => x"98085275",
          6277 => x"51fbf33f",
          6278 => x"82bb9808",
          6279 => x"a0387294",
          6280 => x"150c7252",
          6281 => x"7551f2c1",
          6282 => x"3f82bb98",
          6283 => x"0898150c",
          6284 => x"7690150c",
          6285 => x"7716b405",
          6286 => x"9c150c80",
          6287 => x"557482bb",
          6288 => x"980c8a3d",
          6289 => x"0d04f73d",
          6290 => x"0d7b7d71",
          6291 => x"085b5b57",
          6292 => x"80527651",
          6293 => x"fcac3f82",
          6294 => x"bb980854",
          6295 => x"82bb9808",
          6296 => x"80ec3882",
          6297 => x"bb980856",
          6298 => x"98170852",
          6299 => x"7851f083",
          6300 => x"3f82bb98",
          6301 => x"085482bb",
          6302 => x"980880d2",
          6303 => x"3882bb98",
          6304 => x"089c1808",
          6305 => x"70335154",
          6306 => x"587281e5",
          6307 => x"2e098106",
          6308 => x"83388158",
          6309 => x"82bb9808",
          6310 => x"55728338",
          6311 => x"81557775",
          6312 => x"07537280",
          6313 => x"2e8e3881",
          6314 => x"1656757a",
          6315 => x"2e098106",
          6316 => x"8838a539",
          6317 => x"82bb9808",
          6318 => x"56815276",
          6319 => x"51fd8e3f",
          6320 => x"82bb9808",
          6321 => x"5482bb98",
          6322 => x"08802eff",
          6323 => x"9b387384",
          6324 => x"2e098106",
          6325 => x"83388754",
          6326 => x"7382bb98",
          6327 => x"0c8b3d0d",
          6328 => x"04fd3d0d",
          6329 => x"769a1152",
          6330 => x"54ebec3f",
          6331 => x"82bb9808",
          6332 => x"83ffff06",
          6333 => x"76703351",
          6334 => x"53537183",
          6335 => x"2e098106",
          6336 => x"90389414",
          6337 => x"51ebd03f",
          6338 => x"82bb9808",
          6339 => x"902b7307",
          6340 => x"537282bb",
          6341 => x"980c853d",
          6342 => x"0d04fc3d",
          6343 => x"0d777970",
          6344 => x"83ffff06",
          6345 => x"549a1253",
          6346 => x"5555ebed",
          6347 => x"3f767033",
          6348 => x"51537283",
          6349 => x"2e098106",
          6350 => x"8b387390",
          6351 => x"2a529415",
          6352 => x"51ebd63f",
          6353 => x"863d0d04",
          6354 => x"f73d0d7b",
          6355 => x"7d5b5584",
          6356 => x"75085a58",
          6357 => x"98150880",
          6358 => x"2e818a38",
          6359 => x"98150852",
          6360 => x"7851ee8f",
          6361 => x"3f82bb98",
          6362 => x"085882bb",
          6363 => x"980880f5",
          6364 => x"389c1508",
          6365 => x"70335553",
          6366 => x"73863884",
          6367 => x"5880e639",
          6368 => x"8b133370",
          6369 => x"bf067081",
          6370 => x"ff065851",
          6371 => x"53728616",
          6372 => x"3482bb98",
          6373 => x"08537381",
          6374 => x"e52e8338",
          6375 => x"815373ae",
          6376 => x"2ea93881",
          6377 => x"70740654",
          6378 => x"5772802e",
          6379 => x"9e38758f",
          6380 => x"2e993882",
          6381 => x"bb980876",
          6382 => x"df065454",
          6383 => x"72882e09",
          6384 => x"81068338",
          6385 => x"7654737a",
          6386 => x"2ea03880",
          6387 => x"527451fa",
          6388 => x"fc3f82bb",
          6389 => x"98085882",
          6390 => x"bb980889",
          6391 => x"38981508",
          6392 => x"fefa3886",
          6393 => x"39800b98",
          6394 => x"160c7782",
          6395 => x"bb980c8b",
          6396 => x"3d0d04fb",
          6397 => x"3d0d7770",
          6398 => x"08575481",
          6399 => x"527351fc",
          6400 => x"c53f82bb",
          6401 => x"98085582",
          6402 => x"bb9808b4",
          6403 => x"38981408",
          6404 => x"527551ec",
          6405 => x"de3f82bb",
          6406 => x"98085582",
          6407 => x"bb9808a0",
          6408 => x"38a05382",
          6409 => x"bb980852",
          6410 => x"9c140851",
          6411 => x"eadb3f8b",
          6412 => x"53a01452",
          6413 => x"9c140851",
          6414 => x"eaac3f81",
          6415 => x"0b831734",
          6416 => x"7482bb98",
          6417 => x"0c873d0d",
          6418 => x"04fd3d0d",
          6419 => x"75700898",
          6420 => x"12085470",
          6421 => x"535553ec",
          6422 => x"9a3f82bb",
          6423 => x"98088d38",
          6424 => x"9c130853",
          6425 => x"e5733481",
          6426 => x"0b831534",
          6427 => x"853d0d04",
          6428 => x"fa3d0d78",
          6429 => x"7a575780",
          6430 => x"0b891734",
          6431 => x"98170880",
          6432 => x"2e818238",
          6433 => x"80708918",
          6434 => x"5555559c",
          6435 => x"17081470",
          6436 => x"33811656",
          6437 => x"515271a0",
          6438 => x"2ea83871",
          6439 => x"852e0981",
          6440 => x"06843881",
          6441 => x"e5527389",
          6442 => x"2e098106",
          6443 => x"8b38ae73",
          6444 => x"70810555",
          6445 => x"34811555",
          6446 => x"71737081",
          6447 => x"05553481",
          6448 => x"15558a74",
          6449 => x"27c53875",
          6450 => x"15880552",
          6451 => x"800b8113",
          6452 => x"349c1708",
          6453 => x"528b1233",
          6454 => x"8817349c",
          6455 => x"17089c11",
          6456 => x"5252e88a",
          6457 => x"3f82bb98",
          6458 => x"08760c96",
          6459 => x"1251e7e7",
          6460 => x"3f82bb98",
          6461 => x"08861723",
          6462 => x"981251e7",
          6463 => x"da3f82bb",
          6464 => x"98088417",
          6465 => x"23883d0d",
          6466 => x"04f33d0d",
          6467 => x"7f70085e",
          6468 => x"5b806170",
          6469 => x"33515555",
          6470 => x"73af2e83",
          6471 => x"38815573",
          6472 => x"80dc2e91",
          6473 => x"3874802e",
          6474 => x"8c38941d",
          6475 => x"08881c0c",
          6476 => x"aa398115",
          6477 => x"41806170",
          6478 => x"33565656",
          6479 => x"73af2e09",
          6480 => x"81068338",
          6481 => x"81567380",
          6482 => x"dc327030",
          6483 => x"70802578",
          6484 => x"07515154",
          6485 => x"73dc3873",
          6486 => x"881c0c60",
          6487 => x"70335154",
          6488 => x"739f2696",
          6489 => x"38ff800b",
          6490 => x"ab1c3480",
          6491 => x"527a51f6",
          6492 => x"913f82bb",
          6493 => x"98085585",
          6494 => x"9839913d",
          6495 => x"61a01d5c",
          6496 => x"5a5e8b53",
          6497 => x"a0527951",
          6498 => x"e7ff3f80",
          6499 => x"70595788",
          6500 => x"7933555c",
          6501 => x"73ae2e09",
          6502 => x"810680d4",
          6503 => x"38781870",
          6504 => x"33811a71",
          6505 => x"ae327030",
          6506 => x"709f2a73",
          6507 => x"82260751",
          6508 => x"51535a57",
          6509 => x"54738c38",
          6510 => x"79175475",
          6511 => x"74348117",
          6512 => x"57db3975",
          6513 => x"af327030",
          6514 => x"709f2a51",
          6515 => x"51547580",
          6516 => x"dc2e8c38",
          6517 => x"73802e87",
          6518 => x"3875a026",
          6519 => x"82bd3877",
          6520 => x"197e0ca4",
          6521 => x"54a07627",
          6522 => x"82bd38a0",
          6523 => x"5482b839",
          6524 => x"78187033",
          6525 => x"811a5a57",
          6526 => x"54a07627",
          6527 => x"81fc3875",
          6528 => x"af327030",
          6529 => x"7780dc32",
          6530 => x"70307280",
          6531 => x"25718025",
          6532 => x"07515156",
          6533 => x"51557380",
          6534 => x"2eac3884",
          6535 => x"39811858",
          6536 => x"80781a70",
          6537 => x"33515555",
          6538 => x"73af2e09",
          6539 => x"81068338",
          6540 => x"81557380",
          6541 => x"dc327030",
          6542 => x"70802577",
          6543 => x"07515154",
          6544 => x"73db3881",
          6545 => x"b53975ae",
          6546 => x"2e098106",
          6547 => x"83388154",
          6548 => x"767c2774",
          6549 => x"07547380",
          6550 => x"2ea2387b",
          6551 => x"8b327030",
          6552 => x"77ae3270",
          6553 => x"30728025",
          6554 => x"719f2a07",
          6555 => x"53515651",
          6556 => x"557481a7",
          6557 => x"3888578b",
          6558 => x"5cfef539",
          6559 => x"75982b54",
          6560 => x"7380258c",
          6561 => x"387580ff",
          6562 => x"0682b4e0",
          6563 => x"11335754",
          6564 => x"7551e6e1",
          6565 => x"3f82bb98",
          6566 => x"08802eb2",
          6567 => x"38781870",
          6568 => x"33811a71",
          6569 => x"545a5654",
          6570 => x"e6d23f82",
          6571 => x"bb980880",
          6572 => x"2e80e838",
          6573 => x"ff1c5476",
          6574 => x"742780df",
          6575 => x"38791754",
          6576 => x"75743481",
          6577 => x"177a1155",
          6578 => x"57747434",
          6579 => x"a7397552",
          6580 => x"82b48051",
          6581 => x"e5fe3f82",
          6582 => x"bb9808bf",
          6583 => x"38ff9f16",
          6584 => x"54739926",
          6585 => x"8938e016",
          6586 => x"7081ff06",
          6587 => x"57547917",
          6588 => x"54757434",
          6589 => x"811757fd",
          6590 => x"f7397719",
          6591 => x"7e0c7680",
          6592 => x"2e993879",
          6593 => x"33547381",
          6594 => x"e52e0981",
          6595 => x"06843885",
          6596 => x"7a348454",
          6597 => x"a076278f",
          6598 => x"388b3986",
          6599 => x"5581f239",
          6600 => x"845680f3",
          6601 => x"39805473",
          6602 => x"8b1b3480",
          6603 => x"7b085852",
          6604 => x"7a51f2ce",
          6605 => x"3f82bb98",
          6606 => x"085682bb",
          6607 => x"980880d7",
          6608 => x"38981b08",
          6609 => x"527651e6",
          6610 => x"aa3f82bb",
          6611 => x"98085682",
          6612 => x"bb980880",
          6613 => x"c2389c1b",
          6614 => x"08703355",
          6615 => x"5573802e",
          6616 => x"ffbe388b",
          6617 => x"1533bf06",
          6618 => x"5473861c",
          6619 => x"348b1533",
          6620 => x"70832a70",
          6621 => x"81065155",
          6622 => x"58739238",
          6623 => x"8b537952",
          6624 => x"7451e49f",
          6625 => x"3f82bb98",
          6626 => x"08802e8b",
          6627 => x"3875527a",
          6628 => x"51f3ba3f",
          6629 => x"ff9f3975",
          6630 => x"ab1c3357",
          6631 => x"5574802e",
          6632 => x"bb387484",
          6633 => x"2e098106",
          6634 => x"80e73875",
          6635 => x"852a7081",
          6636 => x"0677822a",
          6637 => x"58515473",
          6638 => x"802e9638",
          6639 => x"75810654",
          6640 => x"73802efb",
          6641 => x"b538ff80",
          6642 => x"0bab1c34",
          6643 => x"805580c1",
          6644 => x"39758106",
          6645 => x"5473ba38",
          6646 => x"8555b639",
          6647 => x"75822a70",
          6648 => x"81065154",
          6649 => x"73ab3886",
          6650 => x"1b337084",
          6651 => x"2a708106",
          6652 => x"51555573",
          6653 => x"802ee138",
          6654 => x"901b0883",
          6655 => x"ff061db4",
          6656 => x"05527c51",
          6657 => x"f5db3f82",
          6658 => x"bb980888",
          6659 => x"1c0cfaea",
          6660 => x"397482bb",
          6661 => x"980c8f3d",
          6662 => x"0d04f63d",
          6663 => x"0d7c5bff",
          6664 => x"7b087071",
          6665 => x"7355595c",
          6666 => x"55597380",
          6667 => x"2e81c638",
          6668 => x"75708105",
          6669 => x"573370a0",
          6670 => x"26525271",
          6671 => x"ba2e8d38",
          6672 => x"70ee3871",
          6673 => x"ba2e0981",
          6674 => x"0681a538",
          6675 => x"7333d011",
          6676 => x"7081ff06",
          6677 => x"51525370",
          6678 => x"89269138",
          6679 => x"82147381",
          6680 => x"ff06d005",
          6681 => x"56527176",
          6682 => x"2e80f738",
          6683 => x"800b82b4",
          6684 => x"d0595577",
          6685 => x"087a5557",
          6686 => x"76708105",
          6687 => x"58337470",
          6688 => x"81055633",
          6689 => x"ff9f1253",
          6690 => x"53537099",
          6691 => x"268938e0",
          6692 => x"137081ff",
          6693 => x"065451ff",
          6694 => x"9f125170",
          6695 => x"99268938",
          6696 => x"e0127081",
          6697 => x"ff065351",
          6698 => x"7230709f",
          6699 => x"2a515172",
          6700 => x"722e0981",
          6701 => x"06853870",
          6702 => x"ffbe3872",
          6703 => x"30747732",
          6704 => x"70307072",
          6705 => x"079f2a73",
          6706 => x"9f2a0753",
          6707 => x"54545170",
          6708 => x"802e8f38",
          6709 => x"81158419",
          6710 => x"59558375",
          6711 => x"25ff9438",
          6712 => x"8b397483",
          6713 => x"24863874",
          6714 => x"767c0c59",
          6715 => x"78518639",
          6716 => x"82d2e433",
          6717 => x"517082bb",
          6718 => x"980c8c3d",
          6719 => x"0d04fa3d",
          6720 => x"0d785680",
          6721 => x"0b831734",
          6722 => x"ff0bb017",
          6723 => x"0c795275",
          6724 => x"51e2e03f",
          6725 => x"845582bb",
          6726 => x"98088180",
          6727 => x"3884b216",
          6728 => x"51dfb43f",
          6729 => x"82bb9808",
          6730 => x"83ffff06",
          6731 => x"54835573",
          6732 => x"82d4d52e",
          6733 => x"09810680",
          6734 => x"e338800b",
          6735 => x"b4173356",
          6736 => x"577481e9",
          6737 => x"2e098106",
          6738 => x"83388157",
          6739 => x"7481eb32",
          6740 => x"70307080",
          6741 => x"25790751",
          6742 => x"5154738a",
          6743 => x"387481e8",
          6744 => x"2e098106",
          6745 => x"b5388353",
          6746 => x"82b49052",
          6747 => x"80ea1651",
          6748 => x"e0b13f82",
          6749 => x"bb980855",
          6750 => x"82bb9808",
          6751 => x"802e9d38",
          6752 => x"855382b4",
          6753 => x"94528186",
          6754 => x"1651e097",
          6755 => x"3f82bb98",
          6756 => x"085582bb",
          6757 => x"9808802e",
          6758 => x"83388255",
          6759 => x"7482bb98",
          6760 => x"0c883d0d",
          6761 => x"04f23d0d",
          6762 => x"61028405",
          6763 => x"80cb0533",
          6764 => x"58558075",
          6765 => x"0c6051fc",
          6766 => x"e13f82bb",
          6767 => x"9808588b",
          6768 => x"56800b82",
          6769 => x"bb980824",
          6770 => x"86fc3882",
          6771 => x"bb980884",
          6772 => x"2982d2d0",
          6773 => x"05700855",
          6774 => x"538c5673",
          6775 => x"802e86e6",
          6776 => x"3873750c",
          6777 => x"7681fe06",
          6778 => x"74335457",
          6779 => x"72802eae",
          6780 => x"38811433",
          6781 => x"51d7ca3f",
          6782 => x"82bb9808",
          6783 => x"81ff0670",
          6784 => x"81065455",
          6785 => x"72983876",
          6786 => x"802e86b8",
          6787 => x"3874822a",
          6788 => x"70810651",
          6789 => x"538a5672",
          6790 => x"86ac3886",
          6791 => x"a7398074",
          6792 => x"34778115",
          6793 => x"34815281",
          6794 => x"143351d7",
          6795 => x"b23f82bb",
          6796 => x"980881ff",
          6797 => x"06708106",
          6798 => x"54558356",
          6799 => x"72868738",
          6800 => x"76802e8f",
          6801 => x"3874822a",
          6802 => x"70810651",
          6803 => x"538a5672",
          6804 => x"85f43880",
          6805 => x"70537452",
          6806 => x"5bfda33f",
          6807 => x"82bb9808",
          6808 => x"81ff0657",
          6809 => x"76822e09",
          6810 => x"810680e2",
          6811 => x"388c3d74",
          6812 => x"56588356",
          6813 => x"83f61533",
          6814 => x"70585372",
          6815 => x"802e8d38",
          6816 => x"83fa1551",
          6817 => x"dce83f82",
          6818 => x"bb980857",
          6819 => x"76787084",
          6820 => x"055a0cff",
          6821 => x"16901656",
          6822 => x"56758025",
          6823 => x"d738800b",
          6824 => x"8d3d5456",
          6825 => x"72708405",
          6826 => x"54085b83",
          6827 => x"577a802e",
          6828 => x"95387a52",
          6829 => x"7351fcc6",
          6830 => x"3f82bb98",
          6831 => x"0881ff06",
          6832 => x"57817727",
          6833 => x"89388116",
          6834 => x"56837627",
          6835 => x"d7388156",
          6836 => x"76842e84",
          6837 => x"f1388d56",
          6838 => x"76812684",
          6839 => x"e938bf14",
          6840 => x"51dbf43f",
          6841 => x"82bb9808",
          6842 => x"83ffff06",
          6843 => x"53728480",
          6844 => x"2e098106",
          6845 => x"84d03880",
          6846 => x"ca1451db",
          6847 => x"da3f82bb",
          6848 => x"980883ff",
          6849 => x"ff065877",
          6850 => x"8d3880d8",
          6851 => x"1451dbde",
          6852 => x"3f82bb98",
          6853 => x"0858779c",
          6854 => x"150c80c4",
          6855 => x"14338215",
          6856 => x"3480c414",
          6857 => x"33ff1170",
          6858 => x"81ff0651",
          6859 => x"54558d56",
          6860 => x"72812684",
          6861 => x"91387481",
          6862 => x"ff067871",
          6863 => x"2980c116",
          6864 => x"33525953",
          6865 => x"728a1523",
          6866 => x"72802e8b",
          6867 => x"38ff1373",
          6868 => x"06537280",
          6869 => x"2e86388d",
          6870 => x"5683eb39",
          6871 => x"80c51451",
          6872 => x"daf53f82",
          6873 => x"bb980853",
          6874 => x"82bb9808",
          6875 => x"88152372",
          6876 => x"8f06578d",
          6877 => x"567683ce",
          6878 => x"3880c714",
          6879 => x"51dad83f",
          6880 => x"82bb9808",
          6881 => x"83ffff06",
          6882 => x"55748d38",
          6883 => x"80d41451",
          6884 => x"dadc3f82",
          6885 => x"bb980855",
          6886 => x"80c21451",
          6887 => x"dab93f82",
          6888 => x"bb980883",
          6889 => x"ffff0653",
          6890 => x"8d567280",
          6891 => x"2e839738",
          6892 => x"88142278",
          6893 => x"1471842a",
          6894 => x"055a5a78",
          6895 => x"75268386",
          6896 => x"388a1422",
          6897 => x"52747931",
          6898 => x"51fefad7",
          6899 => x"3f82bb98",
          6900 => x"085582bb",
          6901 => x"9808802e",
          6902 => x"82ec3882",
          6903 => x"bb980880",
          6904 => x"fffffff5",
          6905 => x"26833883",
          6906 => x"577483ff",
          6907 => x"f5268338",
          6908 => x"8257749f",
          6909 => x"f5268538",
          6910 => x"81578939",
          6911 => x"8d567680",
          6912 => x"2e82c338",
          6913 => x"82157098",
          6914 => x"160c7ba0",
          6915 => x"160c731c",
          6916 => x"70a4170c",
          6917 => x"7a1dac17",
          6918 => x"0c545576",
          6919 => x"832e0981",
          6920 => x"06af3880",
          6921 => x"de1451d9",
          6922 => x"ae3f82bb",
          6923 => x"980883ff",
          6924 => x"ff06538d",
          6925 => x"5672828e",
          6926 => x"3879828a",
          6927 => x"3880e014",
          6928 => x"51d9ab3f",
          6929 => x"82bb9808",
          6930 => x"a8150c74",
          6931 => x"822b53a2",
          6932 => x"398d5679",
          6933 => x"802e81ee",
          6934 => x"387713a8",
          6935 => x"150c7415",
          6936 => x"5376822e",
          6937 => x"8d387410",
          6938 => x"1570812a",
          6939 => x"76810605",
          6940 => x"515383ff",
          6941 => x"13892a53",
          6942 => x"8d56729c",
          6943 => x"15082681",
          6944 => x"c538ff0b",
          6945 => x"90150cff",
          6946 => x"0b8c150c",
          6947 => x"ff800b84",
          6948 => x"15347683",
          6949 => x"2e098106",
          6950 => x"81923880",
          6951 => x"e41451d8",
          6952 => x"b63f82bb",
          6953 => x"980883ff",
          6954 => x"ff065372",
          6955 => x"812e0981",
          6956 => x"0680f938",
          6957 => x"811b5273",
          6958 => x"51dbb83f",
          6959 => x"82bb9808",
          6960 => x"80ea3882",
          6961 => x"bb980884",
          6962 => x"153484b2",
          6963 => x"1451d887",
          6964 => x"3f82bb98",
          6965 => x"0883ffff",
          6966 => x"06537282",
          6967 => x"d4d52e09",
          6968 => x"810680c8",
          6969 => x"38b41451",
          6970 => x"d8843f82",
          6971 => x"bb980884",
          6972 => x"8b85a4d2",
          6973 => x"2e098106",
          6974 => x"b3388498",
          6975 => x"1451d7ee",
          6976 => x"3f82bb98",
          6977 => x"08868a85",
          6978 => x"e4f22e09",
          6979 => x"81069d38",
          6980 => x"849c1451",
          6981 => x"d7d83f82",
          6982 => x"bb980890",
          6983 => x"150c84a0",
          6984 => x"1451d7ca",
          6985 => x"3f82bb98",
          6986 => x"088c150c",
          6987 => x"76743482",
          6988 => x"d2e02281",
          6989 => x"05537282",
          6990 => x"d2e02372",
          6991 => x"86152380",
          6992 => x"0b94150c",
          6993 => x"80567582",
          6994 => x"bb980c90",
          6995 => x"3d0d04fb",
          6996 => x"3d0d7754",
          6997 => x"89557380",
          6998 => x"2eb93873",
          6999 => x"08537280",
          7000 => x"2eb13872",
          7001 => x"33527180",
          7002 => x"2ea93886",
          7003 => x"13228415",
          7004 => x"22575271",
          7005 => x"762e0981",
          7006 => x"06993881",
          7007 => x"133351d0",
          7008 => x"c03f82bb",
          7009 => x"98088106",
          7010 => x"52718838",
          7011 => x"71740854",
          7012 => x"55833980",
          7013 => x"53787371",
          7014 => x"0c527482",
          7015 => x"bb980c87",
          7016 => x"3d0d04fa",
          7017 => x"3d0d02ab",
          7018 => x"05337a58",
          7019 => x"893dfc05",
          7020 => x"5256f4e6",
          7021 => x"3f8b5480",
          7022 => x"0b82bb98",
          7023 => x"0824bc38",
          7024 => x"82bb9808",
          7025 => x"842982d2",
          7026 => x"d0057008",
          7027 => x"55557380",
          7028 => x"2e843880",
          7029 => x"74347854",
          7030 => x"73802e84",
          7031 => x"38807434",
          7032 => x"78750c75",
          7033 => x"5475802e",
          7034 => x"92388053",
          7035 => x"893d7053",
          7036 => x"840551f7",
          7037 => x"b03f82bb",
          7038 => x"98085473",
          7039 => x"82bb980c",
          7040 => x"883d0d04",
          7041 => x"eb3d0d67",
          7042 => x"02840580",
          7043 => x"e7053359",
          7044 => x"59895478",
          7045 => x"802e84c8",
          7046 => x"3877bf06",
          7047 => x"7054983d",
          7048 => x"d0055399",
          7049 => x"3d840552",
          7050 => x"58f6fa3f",
          7051 => x"82bb9808",
          7052 => x"5582bb98",
          7053 => x"0884a438",
          7054 => x"7a5c6852",
          7055 => x"8c3d7052",
          7056 => x"56edc63f",
          7057 => x"82bb9808",
          7058 => x"5582bb98",
          7059 => x"08923802",
          7060 => x"80d70533",
          7061 => x"70982b55",
          7062 => x"57738025",
          7063 => x"83388655",
          7064 => x"779c0654",
          7065 => x"73802e81",
          7066 => x"ab387480",
          7067 => x"2e953874",
          7068 => x"842e0981",
          7069 => x"06aa3875",
          7070 => x"51eaf83f",
          7071 => x"82bb9808",
          7072 => x"559e3902",
          7073 => x"b2053391",
          7074 => x"06547381",
          7075 => x"b8387782",
          7076 => x"2a708106",
          7077 => x"51547380",
          7078 => x"2e8e3888",
          7079 => x"5583bc39",
          7080 => x"77880758",
          7081 => x"7483b438",
          7082 => x"77832a70",
          7083 => x"81065154",
          7084 => x"73802e81",
          7085 => x"af386252",
          7086 => x"7a51e8a5",
          7087 => x"3f82bb98",
          7088 => x"08568288",
          7089 => x"b20a5262",
          7090 => x"8e0551d4",
          7091 => x"ea3f6254",
          7092 => x"a00b8b15",
          7093 => x"34805362",
          7094 => x"527a51e8",
          7095 => x"bd3f8052",
          7096 => x"629c0551",
          7097 => x"d4d13f7a",
          7098 => x"54810b83",
          7099 => x"15347580",
          7100 => x"2e80f138",
          7101 => x"7ab01108",
          7102 => x"51548053",
          7103 => x"7552973d",
          7104 => x"d40551dd",
          7105 => x"be3f82bb",
          7106 => x"98085582",
          7107 => x"bb980882",
          7108 => x"ca38b739",
          7109 => x"7482c438",
          7110 => x"02b20533",
          7111 => x"70842a70",
          7112 => x"81065155",
          7113 => x"5673802e",
          7114 => x"86388455",
          7115 => x"82ad3977",
          7116 => x"812a7081",
          7117 => x"06515473",
          7118 => x"802ea938",
          7119 => x"75810654",
          7120 => x"73802ea0",
          7121 => x"38875582",
          7122 => x"92397352",
          7123 => x"7a51d6a3",
          7124 => x"3f82bb98",
          7125 => x"087bff18",
          7126 => x"8c120c55",
          7127 => x"5582bb98",
          7128 => x"0881f838",
          7129 => x"77832a70",
          7130 => x"81065154",
          7131 => x"73802e86",
          7132 => x"387780c0",
          7133 => x"07587ab0",
          7134 => x"1108a01b",
          7135 => x"0c63a41b",
          7136 => x"0c635370",
          7137 => x"5257e6d9",
          7138 => x"3f82bb98",
          7139 => x"0882bb98",
          7140 => x"08881b0c",
          7141 => x"639c0552",
          7142 => x"5ad2d33f",
          7143 => x"82bb9808",
          7144 => x"82bb9808",
          7145 => x"8c1b0c77",
          7146 => x"7a0c5686",
          7147 => x"1722841a",
          7148 => x"2377901a",
          7149 => x"34800b91",
          7150 => x"1a34800b",
          7151 => x"9c1a0c80",
          7152 => x"0b941a0c",
          7153 => x"77852a70",
          7154 => x"81065154",
          7155 => x"73802e81",
          7156 => x"8d3882bb",
          7157 => x"9808802e",
          7158 => x"81843882",
          7159 => x"bb980894",
          7160 => x"1a0c8a17",
          7161 => x"2270892b",
          7162 => x"7b525957",
          7163 => x"a8397652",
          7164 => x"7851d79f",
          7165 => x"3f82bb98",
          7166 => x"085782bb",
          7167 => x"98088126",
          7168 => x"83388255",
          7169 => x"82bb9808",
          7170 => x"ff2e0981",
          7171 => x"06833879",
          7172 => x"55757831",
          7173 => x"56743070",
          7174 => x"76078025",
          7175 => x"51547776",
          7176 => x"278a3881",
          7177 => x"70750655",
          7178 => x"5a73c338",
          7179 => x"76981a0c",
          7180 => x"74a93875",
          7181 => x"83ff0654",
          7182 => x"73802ea2",
          7183 => x"3876527a",
          7184 => x"51d6a63f",
          7185 => x"82bb9808",
          7186 => x"85388255",
          7187 => x"8e397589",
          7188 => x"2a82bb98",
          7189 => x"08059c1a",
          7190 => x"0c843980",
          7191 => x"790c7454",
          7192 => x"7382bb98",
          7193 => x"0c973d0d",
          7194 => x"04f23d0d",
          7195 => x"60636564",
          7196 => x"40405d59",
          7197 => x"807e0c90",
          7198 => x"3dfc0552",
          7199 => x"7851f9cf",
          7200 => x"3f82bb98",
          7201 => x"085582bb",
          7202 => x"98088a38",
          7203 => x"91193355",
          7204 => x"74802e86",
          7205 => x"38745682",
          7206 => x"c4399019",
          7207 => x"33810655",
          7208 => x"87567480",
          7209 => x"2e82b638",
          7210 => x"9539820b",
          7211 => x"911a3482",
          7212 => x"5682aa39",
          7213 => x"810b911a",
          7214 => x"34815682",
          7215 => x"a0398c19",
          7216 => x"08941a08",
          7217 => x"3155747c",
          7218 => x"27833874",
          7219 => x"5c7b802e",
          7220 => x"82893894",
          7221 => x"19087083",
          7222 => x"ff065656",
          7223 => x"7481b238",
          7224 => x"7e8a1122",
          7225 => x"ff057789",
          7226 => x"2a065b55",
          7227 => x"79a83875",
          7228 => x"87388819",
          7229 => x"08558f39",
          7230 => x"98190852",
          7231 => x"7851d593",
          7232 => x"3f82bb98",
          7233 => x"08558175",
          7234 => x"27ff9f38",
          7235 => x"74ff2eff",
          7236 => x"a3387498",
          7237 => x"1a0c9819",
          7238 => x"08527e51",
          7239 => x"d4cb3f82",
          7240 => x"bb980880",
          7241 => x"2eff8338",
          7242 => x"82bb9808",
          7243 => x"1a7c892a",
          7244 => x"59577780",
          7245 => x"2e80d638",
          7246 => x"771a7f8a",
          7247 => x"1122585c",
          7248 => x"55757527",
          7249 => x"8538757a",
          7250 => x"31587754",
          7251 => x"76537c52",
          7252 => x"811b3351",
          7253 => x"ca883f82",
          7254 => x"bb9808fe",
          7255 => x"d7387e83",
          7256 => x"11335656",
          7257 => x"74802e9f",
          7258 => x"38b01608",
          7259 => x"77315574",
          7260 => x"78279438",
          7261 => x"848053b4",
          7262 => x"1652b016",
          7263 => x"08773189",
          7264 => x"2b7d0551",
          7265 => x"cfe03f77",
          7266 => x"892b56b9",
          7267 => x"39769c1a",
          7268 => x"0c941908",
          7269 => x"83ff0684",
          7270 => x"80713157",
          7271 => x"557b7627",
          7272 => x"83387b56",
          7273 => x"9c190852",
          7274 => x"7e51d1c7",
          7275 => x"3f82bb98",
          7276 => x"08fe8138",
          7277 => x"75539419",
          7278 => x"0883ff06",
          7279 => x"1fb40552",
          7280 => x"7c51cfa2",
          7281 => x"3f7b7631",
          7282 => x"7e08177f",
          7283 => x"0c761e94",
          7284 => x"1b081894",
          7285 => x"1c0c5e5c",
          7286 => x"fdf33980",
          7287 => x"567582bb",
          7288 => x"980c903d",
          7289 => x"0d04f23d",
          7290 => x"0d606365",
          7291 => x"6440405d",
          7292 => x"58807e0c",
          7293 => x"903dfc05",
          7294 => x"527751f6",
          7295 => x"d23f82bb",
          7296 => x"98085582",
          7297 => x"bb98088a",
          7298 => x"38911833",
          7299 => x"5574802e",
          7300 => x"86387456",
          7301 => x"83b83990",
          7302 => x"18337081",
          7303 => x"2a708106",
          7304 => x"51565687",
          7305 => x"5674802e",
          7306 => x"83a43895",
          7307 => x"39820b91",
          7308 => x"19348256",
          7309 => x"83983981",
          7310 => x"0b911934",
          7311 => x"8156838e",
          7312 => x"39941808",
          7313 => x"7c115656",
          7314 => x"74762784",
          7315 => x"3875095c",
          7316 => x"7b802e82",
          7317 => x"ec389418",
          7318 => x"087083ff",
          7319 => x"06565674",
          7320 => x"81fd387e",
          7321 => x"8a1122ff",
          7322 => x"0577892a",
          7323 => x"065c557a",
          7324 => x"bf38758c",
          7325 => x"38881808",
          7326 => x"55749c38",
          7327 => x"7a528539",
          7328 => x"98180852",
          7329 => x"7751d7e7",
          7330 => x"3f82bb98",
          7331 => x"085582bb",
          7332 => x"9808802e",
          7333 => x"82ab3874",
          7334 => x"812eff91",
          7335 => x"3874ff2e",
          7336 => x"ff953874",
          7337 => x"98190c88",
          7338 => x"18088538",
          7339 => x"7488190c",
          7340 => x"7e55b015",
          7341 => x"089c1908",
          7342 => x"2e098106",
          7343 => x"8d387451",
          7344 => x"cec13f82",
          7345 => x"bb9808fe",
          7346 => x"ee389818",
          7347 => x"08527e51",
          7348 => x"d1973f82",
          7349 => x"bb980880",
          7350 => x"2efed238",
          7351 => x"82bb9808",
          7352 => x"1b7c892a",
          7353 => x"5a577880",
          7354 => x"2e80d538",
          7355 => x"781b7f8a",
          7356 => x"1122585b",
          7357 => x"55757527",
          7358 => x"8538757b",
          7359 => x"31597854",
          7360 => x"76537c52",
          7361 => x"811a3351",
          7362 => x"c8be3f82",
          7363 => x"bb9808fe",
          7364 => x"a6387eb0",
          7365 => x"11087831",
          7366 => x"56567479",
          7367 => x"279b3884",
          7368 => x"8053b016",
          7369 => x"08773189",
          7370 => x"2b7d0552",
          7371 => x"b41651cc",
          7372 => x"b53f7e55",
          7373 => x"800b8316",
          7374 => x"3478892b",
          7375 => x"5680db39",
          7376 => x"8c180894",
          7377 => x"19082693",
          7378 => x"387e51cd",
          7379 => x"b63f82bb",
          7380 => x"9808fde3",
          7381 => x"387e77b0",
          7382 => x"120c5576",
          7383 => x"9c190c94",
          7384 => x"180883ff",
          7385 => x"06848071",
          7386 => x"3157557b",
          7387 => x"76278338",
          7388 => x"7b569c18",
          7389 => x"08527e51",
          7390 => x"cdf93f82",
          7391 => x"bb9808fd",
          7392 => x"b6387553",
          7393 => x"7c529418",
          7394 => x"0883ff06",
          7395 => x"1fb40551",
          7396 => x"cbd43f7e",
          7397 => x"55810b83",
          7398 => x"16347b76",
          7399 => x"317e0817",
          7400 => x"7f0c761e",
          7401 => x"941a0818",
          7402 => x"70941c0c",
          7403 => x"8c1b0858",
          7404 => x"585e5c74",
          7405 => x"76278338",
          7406 => x"7555748c",
          7407 => x"190cfd90",
          7408 => x"39901833",
          7409 => x"80c00755",
          7410 => x"74901934",
          7411 => x"80567582",
          7412 => x"bb980c90",
          7413 => x"3d0d04f8",
          7414 => x"3d0d7a8b",
          7415 => x"3dfc0553",
          7416 => x"705256f2",
          7417 => x"ea3f82bb",
          7418 => x"98085782",
          7419 => x"bb980880",
          7420 => x"fb389016",
          7421 => x"3370862a",
          7422 => x"70810651",
          7423 => x"55557380",
          7424 => x"2e80e938",
          7425 => x"a0160852",
          7426 => x"7851cce7",
          7427 => x"3f82bb98",
          7428 => x"085782bb",
          7429 => x"980880d4",
          7430 => x"38a41608",
          7431 => x"8b1133a0",
          7432 => x"07555573",
          7433 => x"8b163488",
          7434 => x"16085374",
          7435 => x"52750851",
          7436 => x"dde83f8c",
          7437 => x"1608529c",
          7438 => x"1551c9fb",
          7439 => x"3f8288b2",
          7440 => x"0a529615",
          7441 => x"51c9f03f",
          7442 => x"76529215",
          7443 => x"51c9ca3f",
          7444 => x"7854810b",
          7445 => x"83153478",
          7446 => x"51ccdf3f",
          7447 => x"82bb9808",
          7448 => x"90173381",
          7449 => x"bf065557",
          7450 => x"73901734",
          7451 => x"7682bb98",
          7452 => x"0c8a3d0d",
          7453 => x"04fc3d0d",
          7454 => x"76705254",
          7455 => x"fed93f82",
          7456 => x"bb980853",
          7457 => x"82bb9808",
          7458 => x"9c38863d",
          7459 => x"fc055273",
          7460 => x"51f1bc3f",
          7461 => x"82bb9808",
          7462 => x"5382bb98",
          7463 => x"08873882",
          7464 => x"bb980874",
          7465 => x"0c7282bb",
          7466 => x"980c863d",
          7467 => x"0d04ff3d",
          7468 => x"0d843d51",
          7469 => x"e6e43f8b",
          7470 => x"52800b82",
          7471 => x"bb980824",
          7472 => x"8b3882bb",
          7473 => x"980882d2",
          7474 => x"e4348052",
          7475 => x"7182bb98",
          7476 => x"0c833d0d",
          7477 => x"04ef3d0d",
          7478 => x"8053933d",
          7479 => x"d0055294",
          7480 => x"3d51e9c1",
          7481 => x"3f82bb98",
          7482 => x"085582bb",
          7483 => x"980880e0",
          7484 => x"38765863",
          7485 => x"52933dd4",
          7486 => x"0551e08d",
          7487 => x"3f82bb98",
          7488 => x"085582bb",
          7489 => x"9808bc38",
          7490 => x"0280c705",
          7491 => x"3370982b",
          7492 => x"55567380",
          7493 => x"25893876",
          7494 => x"7a94120c",
          7495 => x"54b23902",
          7496 => x"a2053370",
          7497 => x"842a7081",
          7498 => x"06515556",
          7499 => x"73802e9e",
          7500 => x"38767f53",
          7501 => x"705254db",
          7502 => x"a83f82bb",
          7503 => x"98089415",
          7504 => x"0c8e3982",
          7505 => x"bb980884",
          7506 => x"2e098106",
          7507 => x"83388555",
          7508 => x"7482bb98",
          7509 => x"0c933d0d",
          7510 => x"04e43d0d",
          7511 => x"6f6f5b5b",
          7512 => x"807a3480",
          7513 => x"539e3dff",
          7514 => x"b805529f",
          7515 => x"3d51e8b5",
          7516 => x"3f82bb98",
          7517 => x"085782bb",
          7518 => x"980882fc",
          7519 => x"387b437a",
          7520 => x"7c941108",
          7521 => x"47555864",
          7522 => x"5473802e",
          7523 => x"81ed38a0",
          7524 => x"52933d70",
          7525 => x"5255d5ea",
          7526 => x"3f82bb98",
          7527 => x"085782bb",
          7528 => x"980882d4",
          7529 => x"3868527b",
          7530 => x"51c9c83f",
          7531 => x"82bb9808",
          7532 => x"5782bb98",
          7533 => x"0882c138",
          7534 => x"69527b51",
          7535 => x"daa33f82",
          7536 => x"bb980845",
          7537 => x"76527451",
          7538 => x"d5b83f82",
          7539 => x"bb980857",
          7540 => x"82bb9808",
          7541 => x"82a23880",
          7542 => x"527451da",
          7543 => x"eb3f82bb",
          7544 => x"98085782",
          7545 => x"bb9808a4",
          7546 => x"3869527b",
          7547 => x"51d9f23f",
          7548 => x"7382bb98",
          7549 => x"082ea638",
          7550 => x"76527451",
          7551 => x"d6cf3f82",
          7552 => x"bb980857",
          7553 => x"82bb9808",
          7554 => x"802ecc38",
          7555 => x"76842e09",
          7556 => x"81068638",
          7557 => x"825781e0",
          7558 => x"397681dc",
          7559 => x"389e3dff",
          7560 => x"bc055274",
          7561 => x"51dcc93f",
          7562 => x"76903d78",
          7563 => x"11811133",
          7564 => x"51565a56",
          7565 => x"73802e91",
          7566 => x"3802b905",
          7567 => x"55811681",
          7568 => x"16703356",
          7569 => x"565673f5",
          7570 => x"38811654",
          7571 => x"73782681",
          7572 => x"90387580",
          7573 => x"2e993878",
          7574 => x"16810555",
          7575 => x"ff186f11",
          7576 => x"ff18ff18",
          7577 => x"58585558",
          7578 => x"74337434",
          7579 => x"75ee38ff",
          7580 => x"186f1155",
          7581 => x"58af7434",
          7582 => x"fe8d3977",
          7583 => x"7b2e0981",
          7584 => x"068a38ff",
          7585 => x"186f1155",
          7586 => x"58af7434",
          7587 => x"800b82d2",
          7588 => x"e4337084",
          7589 => x"2982b4d0",
          7590 => x"05700870",
          7591 => x"33525c56",
          7592 => x"56567376",
          7593 => x"2e8d3881",
          7594 => x"16701a70",
          7595 => x"33515556",
          7596 => x"73f53882",
          7597 => x"16547378",
          7598 => x"26a73880",
          7599 => x"55747627",
          7600 => x"91387419",
          7601 => x"5473337a",
          7602 => x"7081055c",
          7603 => x"34811555",
          7604 => x"ec39ba7a",
          7605 => x"7081055c",
          7606 => x"3474ff2e",
          7607 => x"09810685",
          7608 => x"38915794",
          7609 => x"396e1881",
          7610 => x"19595473",
          7611 => x"337a7081",
          7612 => x"055c347a",
          7613 => x"7826ee38",
          7614 => x"807a3476",
          7615 => x"82bb980c",
          7616 => x"9e3d0d04",
          7617 => x"f73d0d7b",
          7618 => x"7d8d3dfc",
          7619 => x"05547153",
          7620 => x"5755ecbb",
          7621 => x"3f82bb98",
          7622 => x"085382bb",
          7623 => x"980882fa",
          7624 => x"38911533",
          7625 => x"537282f2",
          7626 => x"388c1508",
          7627 => x"54737627",
          7628 => x"92389015",
          7629 => x"3370812a",
          7630 => x"70810651",
          7631 => x"54577283",
          7632 => x"38735694",
          7633 => x"15085480",
          7634 => x"7094170c",
          7635 => x"5875782e",
          7636 => x"82973879",
          7637 => x"8a112270",
          7638 => x"892b5951",
          7639 => x"5373782e",
          7640 => x"b7387652",
          7641 => x"ff1651fe",
          7642 => x"e3b93f82",
          7643 => x"bb9808ff",
          7644 => x"15785470",
          7645 => x"535553fe",
          7646 => x"e3a93f82",
          7647 => x"bb980873",
          7648 => x"26963876",
          7649 => x"30707506",
          7650 => x"7094180c",
          7651 => x"77713198",
          7652 => x"18085758",
          7653 => x"5153b139",
          7654 => x"88150854",
          7655 => x"73a63873",
          7656 => x"527451cd",
          7657 => x"ca3f82bb",
          7658 => x"98085482",
          7659 => x"bb980881",
          7660 => x"2e819a38",
          7661 => x"82bb9808",
          7662 => x"ff2e819b",
          7663 => x"3882bb98",
          7664 => x"0888160c",
          7665 => x"7398160c",
          7666 => x"73802e81",
          7667 => x"9c387676",
          7668 => x"2780dc38",
          7669 => x"75773194",
          7670 => x"16081894",
          7671 => x"170c9016",
          7672 => x"3370812a",
          7673 => x"70810651",
          7674 => x"555a5672",
          7675 => x"802e9a38",
          7676 => x"73527451",
          7677 => x"ccf93f82",
          7678 => x"bb980854",
          7679 => x"82bb9808",
          7680 => x"943882bb",
          7681 => x"980856a7",
          7682 => x"39735274",
          7683 => x"51c7843f",
          7684 => x"82bb9808",
          7685 => x"5473ff2e",
          7686 => x"be388174",
          7687 => x"27af3879",
          7688 => x"53739814",
          7689 => x"0827a638",
          7690 => x"7398160c",
          7691 => x"ffa03994",
          7692 => x"15081694",
          7693 => x"160c7583",
          7694 => x"ff065372",
          7695 => x"802eaa38",
          7696 => x"73527951",
          7697 => x"c6a33f82",
          7698 => x"bb980894",
          7699 => x"38820b91",
          7700 => x"16348253",
          7701 => x"80c43981",
          7702 => x"0b911634",
          7703 => x"8153bb39",
          7704 => x"75892a82",
          7705 => x"bb980805",
          7706 => x"58941508",
          7707 => x"548c1508",
          7708 => x"74279038",
          7709 => x"738c160c",
          7710 => x"90153380",
          7711 => x"c0075372",
          7712 => x"90163473",
          7713 => x"83ff0653",
          7714 => x"72802e8c",
          7715 => x"38779c16",
          7716 => x"082e8538",
          7717 => x"779c160c",
          7718 => x"80537282",
          7719 => x"bb980c8b",
          7720 => x"3d0d04f9",
          7721 => x"3d0d7956",
          7722 => x"89547580",
          7723 => x"2e818a38",
          7724 => x"8053893d",
          7725 => x"fc05528a",
          7726 => x"3d840551",
          7727 => x"e1e73f82",
          7728 => x"bb980855",
          7729 => x"82bb9808",
          7730 => x"80ea3877",
          7731 => x"760c7a52",
          7732 => x"7551d8b5",
          7733 => x"3f82bb98",
          7734 => x"085582bb",
          7735 => x"980880c3",
          7736 => x"38ab1633",
          7737 => x"70982b55",
          7738 => x"57807424",
          7739 => x"a2388616",
          7740 => x"3370842a",
          7741 => x"70810651",
          7742 => x"55577380",
          7743 => x"2ead389c",
          7744 => x"16085277",
          7745 => x"51d3da3f",
          7746 => x"82bb9808",
          7747 => x"88170c77",
          7748 => x"54861422",
          7749 => x"84172374",
          7750 => x"527551ce",
          7751 => x"e53f82bb",
          7752 => x"98085574",
          7753 => x"842e0981",
          7754 => x"06853885",
          7755 => x"55863974",
          7756 => x"802e8438",
          7757 => x"80760c74",
          7758 => x"547382bb",
          7759 => x"980c893d",
          7760 => x"0d04fc3d",
          7761 => x"0d76873d",
          7762 => x"fc055370",
          7763 => x"5253e7ff",
          7764 => x"3f82bb98",
          7765 => x"08873882",
          7766 => x"bb980873",
          7767 => x"0c863d0d",
          7768 => x"04fb3d0d",
          7769 => x"7779893d",
          7770 => x"fc055471",
          7771 => x"535654e7",
          7772 => x"de3f82bb",
          7773 => x"98085382",
          7774 => x"bb980880",
          7775 => x"df387493",
          7776 => x"3882bb98",
          7777 => x"08527351",
          7778 => x"cdf83f82",
          7779 => x"bb980853",
          7780 => x"80ca3982",
          7781 => x"bb980852",
          7782 => x"7351d3ac",
          7783 => x"3f82bb98",
          7784 => x"085382bb",
          7785 => x"9808842e",
          7786 => x"09810685",
          7787 => x"38805387",
          7788 => x"3982bb98",
          7789 => x"08a63874",
          7790 => x"527351d5",
          7791 => x"b33f7252",
          7792 => x"7351cf89",
          7793 => x"3f82bb98",
          7794 => x"08843270",
          7795 => x"30707207",
          7796 => x"9f2c7082",
          7797 => x"bb980806",
          7798 => x"51515454",
          7799 => x"7282bb98",
          7800 => x"0c873d0d",
          7801 => x"04ee3d0d",
          7802 => x"65578053",
          7803 => x"893d7053",
          7804 => x"963d5256",
          7805 => x"dfaf3f82",
          7806 => x"bb980855",
          7807 => x"82bb9808",
          7808 => x"b2386452",
          7809 => x"7551d681",
          7810 => x"3f82bb98",
          7811 => x"085582bb",
          7812 => x"9808a038",
          7813 => x"0280cb05",
          7814 => x"3370982b",
          7815 => x"55587380",
          7816 => x"25853886",
          7817 => x"558d3976",
          7818 => x"802e8838",
          7819 => x"76527551",
          7820 => x"d4be3f74",
          7821 => x"82bb980c",
          7822 => x"943d0d04",
          7823 => x"f03d0d63",
          7824 => x"65555c80",
          7825 => x"53923dec",
          7826 => x"0552933d",
          7827 => x"51ded63f",
          7828 => x"82bb9808",
          7829 => x"5b82bb98",
          7830 => x"08828038",
          7831 => x"7c740c73",
          7832 => x"08981108",
          7833 => x"fe119013",
          7834 => x"08595658",
          7835 => x"55757426",
          7836 => x"9138757c",
          7837 => x"0c81e439",
          7838 => x"815b81cc",
          7839 => x"39825b81",
          7840 => x"c73982bb",
          7841 => x"98087533",
          7842 => x"55597381",
          7843 => x"2e098106",
          7844 => x"bf388275",
          7845 => x"5f577652",
          7846 => x"923df005",
          7847 => x"51c1f43f",
          7848 => x"82bb9808",
          7849 => x"ff2ed138",
          7850 => x"82bb9808",
          7851 => x"812ece38",
          7852 => x"82bb9808",
          7853 => x"307082bb",
          7854 => x"98080780",
          7855 => x"257a0581",
          7856 => x"197f5359",
          7857 => x"5a549814",
          7858 => x"087726ca",
          7859 => x"3880f939",
          7860 => x"a4150882",
          7861 => x"bb980857",
          7862 => x"58759838",
          7863 => x"77528118",
          7864 => x"7d5258ff",
          7865 => x"bf8d3f82",
          7866 => x"bb98085b",
          7867 => x"82bb9808",
          7868 => x"80d6387c",
          7869 => x"70337712",
          7870 => x"ff1a5d52",
          7871 => x"56547482",
          7872 => x"2e098106",
          7873 => x"9e38b414",
          7874 => x"51ffbbcb",
          7875 => x"3f82bb98",
          7876 => x"0883ffff",
          7877 => x"06703070",
          7878 => x"80251b82",
          7879 => x"19595b51",
          7880 => x"549b39b4",
          7881 => x"1451ffbb",
          7882 => x"c53f82bb",
          7883 => x"9808f00a",
          7884 => x"06703070",
          7885 => x"80251b84",
          7886 => x"19595b51",
          7887 => x"547583ff",
          7888 => x"067a5856",
          7889 => x"79ff9238",
          7890 => x"787c0c7c",
          7891 => x"7990120c",
          7892 => x"84113381",
          7893 => x"07565474",
          7894 => x"8415347a",
          7895 => x"82bb980c",
          7896 => x"923d0d04",
          7897 => x"f93d0d79",
          7898 => x"8a3dfc05",
          7899 => x"53705257",
          7900 => x"e3dd3f82",
          7901 => x"bb980856",
          7902 => x"82bb9808",
          7903 => x"81a83891",
          7904 => x"17335675",
          7905 => x"81a03890",
          7906 => x"17337081",
          7907 => x"2a708106",
          7908 => x"51555587",
          7909 => x"5573802e",
          7910 => x"818e3894",
          7911 => x"17085473",
          7912 => x"8c180827",
          7913 => x"81803873",
          7914 => x"9b3882bb",
          7915 => x"98085388",
          7916 => x"17085276",
          7917 => x"51c48c3f",
          7918 => x"82bb9808",
          7919 => x"7488190c",
          7920 => x"5680c939",
          7921 => x"98170852",
          7922 => x"7651ffbf",
          7923 => x"c63f82bb",
          7924 => x"9808ff2e",
          7925 => x"09810683",
          7926 => x"38815682",
          7927 => x"bb980881",
          7928 => x"2e098106",
          7929 => x"85388256",
          7930 => x"a33975a0",
          7931 => x"38775482",
          7932 => x"bb980898",
          7933 => x"15082794",
          7934 => x"38981708",
          7935 => x"5382bb98",
          7936 => x"08527651",
          7937 => x"c3bd3f82",
          7938 => x"bb980856",
          7939 => x"9417088c",
          7940 => x"180c9017",
          7941 => x"3380c007",
          7942 => x"54739018",
          7943 => x"3475802e",
          7944 => x"85387591",
          7945 => x"18347555",
          7946 => x"7482bb98",
          7947 => x"0c893d0d",
          7948 => x"04e23d0d",
          7949 => x"8253a03d",
          7950 => x"ffa40552",
          7951 => x"a13d51da",
          7952 => x"e43f82bb",
          7953 => x"98085582",
          7954 => x"bb980881",
          7955 => x"f5387845",
          7956 => x"a13d0852",
          7957 => x"953d7052",
          7958 => x"58d1ae3f",
          7959 => x"82bb9808",
          7960 => x"5582bb98",
          7961 => x"0881db38",
          7962 => x"0280fb05",
          7963 => x"3370852a",
          7964 => x"70810651",
          7965 => x"55568655",
          7966 => x"7381c738",
          7967 => x"75982b54",
          7968 => x"80742481",
          7969 => x"bd380280",
          7970 => x"d6053370",
          7971 => x"81065854",
          7972 => x"87557681",
          7973 => x"ad386b52",
          7974 => x"7851ccc5",
          7975 => x"3f82bb98",
          7976 => x"0874842a",
          7977 => x"70810651",
          7978 => x"55567380",
          7979 => x"2e80d438",
          7980 => x"785482bb",
          7981 => x"98089415",
          7982 => x"082e8186",
          7983 => x"38735a82",
          7984 => x"bb98085c",
          7985 => x"76528a3d",
          7986 => x"705254c7",
          7987 => x"b53f82bb",
          7988 => x"98085582",
          7989 => x"bb980880",
          7990 => x"e93882bb",
          7991 => x"98085273",
          7992 => x"51cce53f",
          7993 => x"82bb9808",
          7994 => x"5582bb98",
          7995 => x"08863887",
          7996 => x"5580cf39",
          7997 => x"82bb9808",
          7998 => x"842e8838",
          7999 => x"82bb9808",
          8000 => x"80c03877",
          8001 => x"51cec23f",
          8002 => x"82bb9808",
          8003 => x"82bb9808",
          8004 => x"307082bb",
          8005 => x"98080780",
          8006 => x"25515555",
          8007 => x"75802e94",
          8008 => x"3873802e",
          8009 => x"8f388053",
          8010 => x"75527751",
          8011 => x"c1953f82",
          8012 => x"bb980855",
          8013 => x"748c3878",
          8014 => x"51ffbafe",
          8015 => x"3f82bb98",
          8016 => x"08557482",
          8017 => x"bb980ca0",
          8018 => x"3d0d04e9",
          8019 => x"3d0d8253",
          8020 => x"993dc005",
          8021 => x"529a3d51",
          8022 => x"d8cb3f82",
          8023 => x"bb980854",
          8024 => x"82bb9808",
          8025 => x"82b03878",
          8026 => x"5e69528e",
          8027 => x"3d705258",
          8028 => x"cf973f82",
          8029 => x"bb980854",
          8030 => x"82bb9808",
          8031 => x"86388854",
          8032 => x"82943982",
          8033 => x"bb980884",
          8034 => x"2e098106",
          8035 => x"82883802",
          8036 => x"80df0533",
          8037 => x"70852a81",
          8038 => x"06515586",
          8039 => x"547481f6",
          8040 => x"38785a74",
          8041 => x"528a3d70",
          8042 => x"5257c1c3",
          8043 => x"3f82bb98",
          8044 => x"08755556",
          8045 => x"82bb9808",
          8046 => x"83388754",
          8047 => x"82bb9808",
          8048 => x"812e0981",
          8049 => x"06833882",
          8050 => x"5482bb98",
          8051 => x"08ff2e09",
          8052 => x"81068638",
          8053 => x"815481b4",
          8054 => x"397381b0",
          8055 => x"3882bb98",
          8056 => x"08527851",
          8057 => x"c4a43f82",
          8058 => x"bb980854",
          8059 => x"82bb9808",
          8060 => x"819a388b",
          8061 => x"53a052b4",
          8062 => x"1951ffb7",
          8063 => x"8c3f7854",
          8064 => x"ae0bb415",
          8065 => x"34785490",
          8066 => x"0bbf1534",
          8067 => x"8288b20a",
          8068 => x"5280ca19",
          8069 => x"51ffb69f",
          8070 => x"3f755378",
          8071 => x"b4115351",
          8072 => x"c9f83fa0",
          8073 => x"5378b411",
          8074 => x"5380d405",
          8075 => x"51ffb6b6",
          8076 => x"3f7854ae",
          8077 => x"0b80d515",
          8078 => x"347f5378",
          8079 => x"80d41153",
          8080 => x"51c9d73f",
          8081 => x"7854810b",
          8082 => x"83153477",
          8083 => x"51cba43f",
          8084 => x"82bb9808",
          8085 => x"5482bb98",
          8086 => x"08b23882",
          8087 => x"88b20a52",
          8088 => x"64960551",
          8089 => x"ffb5d03f",
          8090 => x"75536452",
          8091 => x"7851c9aa",
          8092 => x"3f645490",
          8093 => x"0b8b1534",
          8094 => x"7854810b",
          8095 => x"83153478",
          8096 => x"51ffb8b6",
          8097 => x"3f82bb98",
          8098 => x"08548b39",
          8099 => x"80537552",
          8100 => x"7651ffbe",
          8101 => x"ae3f7382",
          8102 => x"bb980c99",
          8103 => x"3d0d04da",
          8104 => x"3d0da93d",
          8105 => x"840551d2",
          8106 => x"f13f8253",
          8107 => x"a83dff84",
          8108 => x"0552a93d",
          8109 => x"51d5ee3f",
          8110 => x"82bb9808",
          8111 => x"5582bb98",
          8112 => x"0882d338",
          8113 => x"784da93d",
          8114 => x"08529d3d",
          8115 => x"705258cc",
          8116 => x"b83f82bb",
          8117 => x"98085582",
          8118 => x"bb980882",
          8119 => x"b9380281",
          8120 => x"9b053381",
          8121 => x"a0065486",
          8122 => x"557382aa",
          8123 => x"38a053a4",
          8124 => x"3d0852a8",
          8125 => x"3dff8805",
          8126 => x"51ffb4ea",
          8127 => x"3fac5377",
          8128 => x"52923d70",
          8129 => x"5254ffb4",
          8130 => x"dd3faa3d",
          8131 => x"08527351",
          8132 => x"cbf73f82",
          8133 => x"bb980855",
          8134 => x"82bb9808",
          8135 => x"9538636f",
          8136 => x"2e098106",
          8137 => x"883865a2",
          8138 => x"3d082e92",
          8139 => x"38885581",
          8140 => x"e53982bb",
          8141 => x"9808842e",
          8142 => x"09810681",
          8143 => x"b8387351",
          8144 => x"c9b13f82",
          8145 => x"bb980855",
          8146 => x"82bb9808",
          8147 => x"81c83868",
          8148 => x"569353a8",
          8149 => x"3dff9505",
          8150 => x"528d1651",
          8151 => x"ffb4873f",
          8152 => x"02af0533",
          8153 => x"8b17348b",
          8154 => x"16337084",
          8155 => x"2a708106",
          8156 => x"51555573",
          8157 => x"893874a0",
          8158 => x"0754738b",
          8159 => x"17347854",
          8160 => x"810b8315",
          8161 => x"348b1633",
          8162 => x"70842a70",
          8163 => x"81065155",
          8164 => x"5573802e",
          8165 => x"80e5386e",
          8166 => x"642e80df",
          8167 => x"38755278",
          8168 => x"51c6be3f",
          8169 => x"82bb9808",
          8170 => x"527851ff",
          8171 => x"b7bb3f82",
          8172 => x"5582bb98",
          8173 => x"08802e80",
          8174 => x"dd3882bb",
          8175 => x"98085278",
          8176 => x"51ffb5af",
          8177 => x"3f82bb98",
          8178 => x"087980d4",
          8179 => x"11585855",
          8180 => x"82bb9808",
          8181 => x"80c03881",
          8182 => x"16335473",
          8183 => x"ae2e0981",
          8184 => x"06993863",
          8185 => x"53755276",
          8186 => x"51c6af3f",
          8187 => x"7854810b",
          8188 => x"83153487",
          8189 => x"3982bb98",
          8190 => x"089c3877",
          8191 => x"51c8ca3f",
          8192 => x"82bb9808",
          8193 => x"5582bb98",
          8194 => x"088c3878",
          8195 => x"51ffb5aa",
          8196 => x"3f82bb98",
          8197 => x"08557482",
          8198 => x"bb980ca8",
          8199 => x"3d0d04ed",
          8200 => x"3d0d0280",
          8201 => x"db053302",
          8202 => x"840580df",
          8203 => x"05335757",
          8204 => x"8253953d",
          8205 => x"d0055296",
          8206 => x"3d51d2e9",
          8207 => x"3f82bb98",
          8208 => x"085582bb",
          8209 => x"980880cf",
          8210 => x"38785a65",
          8211 => x"52953dd4",
          8212 => x"0551c9b5",
          8213 => x"3f82bb98",
          8214 => x"085582bb",
          8215 => x"9808b838",
          8216 => x"0280cf05",
          8217 => x"3381a006",
          8218 => x"54865573",
          8219 => x"aa3875a7",
          8220 => x"06617109",
          8221 => x"8b123371",
          8222 => x"067a7406",
          8223 => x"07515755",
          8224 => x"56748b15",
          8225 => x"34785481",
          8226 => x"0b831534",
          8227 => x"7851ffb4",
          8228 => x"a93f82bb",
          8229 => x"98085574",
          8230 => x"82bb980c",
          8231 => x"953d0d04",
          8232 => x"ef3d0d64",
          8233 => x"56825393",
          8234 => x"3dd00552",
          8235 => x"943d51d1",
          8236 => x"f43f82bb",
          8237 => x"98085582",
          8238 => x"bb980880",
          8239 => x"cb387658",
          8240 => x"6352933d",
          8241 => x"d40551c8",
          8242 => x"c03f82bb",
          8243 => x"98085582",
          8244 => x"bb9808b4",
          8245 => x"380280c7",
          8246 => x"053381a0",
          8247 => x"06548655",
          8248 => x"73a63884",
          8249 => x"16228617",
          8250 => x"2271902b",
          8251 => x"07535496",
          8252 => x"1f51ffb0",
          8253 => x"c23f7654",
          8254 => x"810b8315",
          8255 => x"347651ff",
          8256 => x"b3b83f82",
          8257 => x"bb980855",
          8258 => x"7482bb98",
          8259 => x"0c933d0d",
          8260 => x"04ea3d0d",
          8261 => x"696b5c5a",
          8262 => x"8053983d",
          8263 => x"d0055299",
          8264 => x"3d51d181",
          8265 => x"3f82bb98",
          8266 => x"0882bb98",
          8267 => x"08307082",
          8268 => x"bb980807",
          8269 => x"80255155",
          8270 => x"5779802e",
          8271 => x"81853881",
          8272 => x"70750655",
          8273 => x"5573802e",
          8274 => x"80f9387b",
          8275 => x"5d805f80",
          8276 => x"528d3d70",
          8277 => x"5254ffbe",
          8278 => x"a93f82bb",
          8279 => x"98085782",
          8280 => x"bb980880",
          8281 => x"d1387452",
          8282 => x"7351c3dc",
          8283 => x"3f82bb98",
          8284 => x"085782bb",
          8285 => x"9808bf38",
          8286 => x"82bb9808",
          8287 => x"82bb9808",
          8288 => x"655b5956",
          8289 => x"78188119",
          8290 => x"7b185659",
          8291 => x"55743374",
          8292 => x"34811656",
          8293 => x"8a7827ec",
          8294 => x"388b5675",
          8295 => x"1a548074",
          8296 => x"3475802e",
          8297 => x"9e38ff16",
          8298 => x"701b7033",
          8299 => x"51555673",
          8300 => x"a02ee838",
          8301 => x"8e397684",
          8302 => x"2e098106",
          8303 => x"8638807a",
          8304 => x"34805776",
          8305 => x"30707807",
          8306 => x"80255154",
          8307 => x"7a802e80",
          8308 => x"c1387380",
          8309 => x"2ebc387b",
          8310 => x"a0110853",
          8311 => x"51ffb193",
          8312 => x"3f82bb98",
          8313 => x"085782bb",
          8314 => x"9808a738",
          8315 => x"7b703355",
          8316 => x"5580c356",
          8317 => x"73832e8b",
          8318 => x"3880e456",
          8319 => x"73842e83",
          8320 => x"38a75675",
          8321 => x"15b40551",
          8322 => x"ffade33f",
          8323 => x"82bb9808",
          8324 => x"7b0c7682",
          8325 => x"bb980c98",
          8326 => x"3d0d04e6",
          8327 => x"3d0d8253",
          8328 => x"9c3dffb8",
          8329 => x"05529d3d",
          8330 => x"51cefa3f",
          8331 => x"82bb9808",
          8332 => x"82bb9808",
          8333 => x"565482bb",
          8334 => x"98088398",
          8335 => x"388b53a0",
          8336 => x"528b3d70",
          8337 => x"5259ffae",
          8338 => x"c03f736d",
          8339 => x"70337081",
          8340 => x"ff065257",
          8341 => x"55579f74",
          8342 => x"2781bc38",
          8343 => x"78587481",
          8344 => x"ff066d81",
          8345 => x"054e7052",
          8346 => x"55ffaf89",
          8347 => x"3f82bb98",
          8348 => x"08802ea5",
          8349 => x"386c7033",
          8350 => x"70535754",
          8351 => x"ffaefd3f",
          8352 => x"82bb9808",
          8353 => x"802e8d38",
          8354 => x"74882b76",
          8355 => x"076d8105",
          8356 => x"4e558639",
          8357 => x"82bb9808",
          8358 => x"55ff9f15",
          8359 => x"7083ffff",
          8360 => x"06515473",
          8361 => x"99268a38",
          8362 => x"e0157083",
          8363 => x"ffff0656",
          8364 => x"5480ff75",
          8365 => x"27873882",
          8366 => x"b3e01533",
          8367 => x"5574802e",
          8368 => x"a3387452",
          8369 => x"82b5e051",
          8370 => x"ffae893f",
          8371 => x"82bb9808",
          8372 => x"933881ff",
          8373 => x"75278838",
          8374 => x"76892688",
          8375 => x"388b398a",
          8376 => x"77278638",
          8377 => x"865581ec",
          8378 => x"3981ff75",
          8379 => x"278f3874",
          8380 => x"882a5473",
          8381 => x"78708105",
          8382 => x"5a348117",
          8383 => x"57747870",
          8384 => x"81055a34",
          8385 => x"81176d70",
          8386 => x"337081ff",
          8387 => x"06525755",
          8388 => x"57739f26",
          8389 => x"fec8388b",
          8390 => x"3d335486",
          8391 => x"557381e5",
          8392 => x"2e81b138",
          8393 => x"76802e99",
          8394 => x"3802a705",
          8395 => x"55761570",
          8396 => x"33515473",
          8397 => x"a02e0981",
          8398 => x"068738ff",
          8399 => x"175776ed",
          8400 => x"38794180",
          8401 => x"43805291",
          8402 => x"3d705255",
          8403 => x"ffbab33f",
          8404 => x"82bb9808",
          8405 => x"5482bb98",
          8406 => x"0880f738",
          8407 => x"81527451",
          8408 => x"ffbfe53f",
          8409 => x"82bb9808",
          8410 => x"5482bb98",
          8411 => x"088d3876",
          8412 => x"80c43867",
          8413 => x"54e57434",
          8414 => x"80c63982",
          8415 => x"bb980884",
          8416 => x"2e098106",
          8417 => x"80cc3880",
          8418 => x"5476742e",
          8419 => x"80c43881",
          8420 => x"527451ff",
          8421 => x"bdb03f82",
          8422 => x"bb980854",
          8423 => x"82bb9808",
          8424 => x"b138a053",
          8425 => x"82bb9808",
          8426 => x"526751ff",
          8427 => x"abdb3f67",
          8428 => x"54880b8b",
          8429 => x"15348b53",
          8430 => x"78526751",
          8431 => x"ffaba73f",
          8432 => x"7954810b",
          8433 => x"83153479",
          8434 => x"51ffadee",
          8435 => x"3f82bb98",
          8436 => x"08547355",
          8437 => x"7482bb98",
          8438 => x"0c9c3d0d",
          8439 => x"04f23d0d",
          8440 => x"60620288",
          8441 => x"0580cb05",
          8442 => x"33933dfc",
          8443 => x"05557254",
          8444 => x"405e5ad2",
          8445 => x"da3f82bb",
          8446 => x"98085882",
          8447 => x"bb980882",
          8448 => x"bd38911a",
          8449 => x"33587782",
          8450 => x"b5387c80",
          8451 => x"2e97388c",
          8452 => x"1a085978",
          8453 => x"9038901a",
          8454 => x"3370812a",
          8455 => x"70810651",
          8456 => x"55557390",
          8457 => x"38875482",
          8458 => x"97398258",
          8459 => x"82903981",
          8460 => x"58828b39",
          8461 => x"7e8a1122",
          8462 => x"70892b70",
          8463 => x"557f5456",
          8464 => x"5656fec9",
          8465 => x"de3fff14",
          8466 => x"7d067030",
          8467 => x"7072079f",
          8468 => x"2a82bb98",
          8469 => x"08058c19",
          8470 => x"087c405a",
          8471 => x"5d555581",
          8472 => x"77278838",
          8473 => x"98160877",
          8474 => x"26833882",
          8475 => x"57767756",
          8476 => x"59805674",
          8477 => x"527951ff",
          8478 => x"ae993f81",
          8479 => x"157f5555",
          8480 => x"98140875",
          8481 => x"26833882",
          8482 => x"5582bb98",
          8483 => x"08812eff",
          8484 => x"993882bb",
          8485 => x"9808ff2e",
          8486 => x"ff953882",
          8487 => x"bb98088e",
          8488 => x"38811656",
          8489 => x"757b2e09",
          8490 => x"81068738",
          8491 => x"93397459",
          8492 => x"80567477",
          8493 => x"2e098106",
          8494 => x"ffb93887",
          8495 => x"5880ff39",
          8496 => x"7d802eba",
          8497 => x"38787b55",
          8498 => x"557a802e",
          8499 => x"b4388115",
          8500 => x"5673812e",
          8501 => x"09810683",
          8502 => x"38ff5675",
          8503 => x"5374527e",
          8504 => x"51ffafa8",
          8505 => x"3f82bb98",
          8506 => x"085882bb",
          8507 => x"980880ce",
          8508 => x"38748116",
          8509 => x"ff165656",
          8510 => x"5c73d338",
          8511 => x"8439ff19",
          8512 => x"5c7e7c8c",
          8513 => x"120c557d",
          8514 => x"802eb338",
          8515 => x"78881b0c",
          8516 => x"7c8c1b0c",
          8517 => x"901a3380",
          8518 => x"c0075473",
          8519 => x"901b3498",
          8520 => x"1508fe05",
          8521 => x"90160857",
          8522 => x"54757426",
          8523 => x"9138757b",
          8524 => x"3190160c",
          8525 => x"84153381",
          8526 => x"07547384",
          8527 => x"16347754",
          8528 => x"7382bb98",
          8529 => x"0c903d0d",
          8530 => x"04e93d0d",
          8531 => x"6b6d0288",
          8532 => x"0580eb05",
          8533 => x"339d3d54",
          8534 => x"5a5c59c5",
          8535 => x"bd3f8b56",
          8536 => x"800b82bb",
          8537 => x"9808248b",
          8538 => x"f83882bb",
          8539 => x"98088429",
          8540 => x"82d2d005",
          8541 => x"70085155",
          8542 => x"74802e84",
          8543 => x"38807534",
          8544 => x"82bb9808",
          8545 => x"81ff065f",
          8546 => x"81527e51",
          8547 => x"ffa0d03f",
          8548 => x"82bb9808",
          8549 => x"81ff0670",
          8550 => x"81065657",
          8551 => x"8356748b",
          8552 => x"c0387682",
          8553 => x"2a708106",
          8554 => x"51558a56",
          8555 => x"748bb238",
          8556 => x"993dfc05",
          8557 => x"5383527e",
          8558 => x"51ffa4f0",
          8559 => x"3f82bb98",
          8560 => x"08993867",
          8561 => x"5574802e",
          8562 => x"92387482",
          8563 => x"8080268b",
          8564 => x"38ff1575",
          8565 => x"06557480",
          8566 => x"2e833881",
          8567 => x"4878802e",
          8568 => x"87388480",
          8569 => x"79269238",
          8570 => x"7881800a",
          8571 => x"268b38ff",
          8572 => x"19790655",
          8573 => x"74802e86",
          8574 => x"3893568a",
          8575 => x"e4397889",
          8576 => x"2a6e892a",
          8577 => x"70892b77",
          8578 => x"59484359",
          8579 => x"7a833881",
          8580 => x"56613070",
          8581 => x"80257707",
          8582 => x"51559156",
          8583 => x"748ac238",
          8584 => x"993df805",
          8585 => x"5381527e",
          8586 => x"51ffa480",
          8587 => x"3f815682",
          8588 => x"bb98088a",
          8589 => x"ac387783",
          8590 => x"2a707706",
          8591 => x"82bb9808",
          8592 => x"43564574",
          8593 => x"8338bf41",
          8594 => x"66558e56",
          8595 => x"6075268a",
          8596 => x"90387461",
          8597 => x"31704855",
          8598 => x"80ff7527",
          8599 => x"8a833893",
          8600 => x"56788180",
          8601 => x"2689fa38",
          8602 => x"77812a70",
          8603 => x"81065643",
          8604 => x"74802e95",
          8605 => x"38778706",
          8606 => x"5574822e",
          8607 => x"838d3877",
          8608 => x"81065574",
          8609 => x"802e8383",
          8610 => x"38778106",
          8611 => x"55935682",
          8612 => x"5e74802e",
          8613 => x"89cb3878",
          8614 => x"5a7d832e",
          8615 => x"09810680",
          8616 => x"e13878ae",
          8617 => x"3866912a",
          8618 => x"57810b82",
          8619 => x"b6842256",
          8620 => x"5a74802e",
          8621 => x"9d387477",
          8622 => x"26983882",
          8623 => x"b6845679",
          8624 => x"10821770",
          8625 => x"2257575a",
          8626 => x"74802e86",
          8627 => x"38767527",
          8628 => x"ee387952",
          8629 => x"6651fec4",
          8630 => x"ca3f82bb",
          8631 => x"98088429",
          8632 => x"84870570",
          8633 => x"892a5e55",
          8634 => x"a05c800b",
          8635 => x"82bb9808",
          8636 => x"fc808a05",
          8637 => x"5644fdff",
          8638 => x"f00a7527",
          8639 => x"80ec3888",
          8640 => x"d33978ae",
          8641 => x"38668c2a",
          8642 => x"57810b82",
          8643 => x"b5f42256",
          8644 => x"5a74802e",
          8645 => x"9d387477",
          8646 => x"26983882",
          8647 => x"b5f45679",
          8648 => x"10821770",
          8649 => x"2257575a",
          8650 => x"74802e86",
          8651 => x"38767527",
          8652 => x"ee387952",
          8653 => x"6651fec3",
          8654 => x"ea3f82bb",
          8655 => x"98081084",
          8656 => x"055782bb",
          8657 => x"98089ff5",
          8658 => x"26963881",
          8659 => x"0b82bb98",
          8660 => x"081082bb",
          8661 => x"98080571",
          8662 => x"11722a83",
          8663 => x"0559565e",
          8664 => x"83ff1789",
          8665 => x"2a5d815c",
          8666 => x"a044601c",
          8667 => x"7d116505",
          8668 => x"697012ff",
          8669 => x"05713070",
          8670 => x"72067431",
          8671 => x"5c525957",
          8672 => x"59407d83",
          8673 => x"2e098106",
          8674 => x"8938761c",
          8675 => x"6018415c",
          8676 => x"8439761d",
          8677 => x"5d799029",
          8678 => x"18706231",
          8679 => x"68585155",
          8680 => x"74762687",
          8681 => x"af38757c",
          8682 => x"317d317a",
          8683 => x"53706531",
          8684 => x"5255fec2",
          8685 => x"ee3f82bb",
          8686 => x"9808587d",
          8687 => x"832e0981",
          8688 => x"069b3882",
          8689 => x"bb980883",
          8690 => x"fff52680",
          8691 => x"dd387887",
          8692 => x"83387981",
          8693 => x"2a5978fd",
          8694 => x"be3886f8",
          8695 => x"397d822e",
          8696 => x"09810680",
          8697 => x"c53883ff",
          8698 => x"f50b82bb",
          8699 => x"980827a0",
          8700 => x"38788f38",
          8701 => x"791a5574",
          8702 => x"80c02686",
          8703 => x"387459fd",
          8704 => x"96396281",
          8705 => x"06557480",
          8706 => x"2e8f3883",
          8707 => x"5efd8839",
          8708 => x"82bb9808",
          8709 => x"9ff52692",
          8710 => x"387886b8",
          8711 => x"38791a59",
          8712 => x"81807927",
          8713 => x"fcf13886",
          8714 => x"ab398055",
          8715 => x"7d812e09",
          8716 => x"81068338",
          8717 => x"7d559ff5",
          8718 => x"78278b38",
          8719 => x"74810655",
          8720 => x"8e567486",
          8721 => x"9c388480",
          8722 => x"5380527a",
          8723 => x"51ffa2b9",
          8724 => x"3f8b5382",
          8725 => x"b49c527a",
          8726 => x"51ffa28a",
          8727 => x"3f848052",
          8728 => x"8b1b51ff",
          8729 => x"a1b33f79",
          8730 => x"8d1c347b",
          8731 => x"83ffff06",
          8732 => x"528e1b51",
          8733 => x"ffa1a23f",
          8734 => x"810b901c",
          8735 => x"347d8332",
          8736 => x"70307096",
          8737 => x"2a848006",
          8738 => x"54515591",
          8739 => x"1b51ffa1",
          8740 => x"883f6655",
          8741 => x"7483ffff",
          8742 => x"26903874",
          8743 => x"83ffff06",
          8744 => x"52931b51",
          8745 => x"ffa0f23f",
          8746 => x"8a397452",
          8747 => x"a01b51ff",
          8748 => x"a1853ff8",
          8749 => x"0b951c34",
          8750 => x"bf52981b",
          8751 => x"51ffa0d9",
          8752 => x"3f81ff52",
          8753 => x"9a1b51ff",
          8754 => x"a0cf3f60",
          8755 => x"529c1b51",
          8756 => x"ffa0e43f",
          8757 => x"7d832e09",
          8758 => x"810680cb",
          8759 => x"388288b2",
          8760 => x"0a5280c3",
          8761 => x"1b51ffa0",
          8762 => x"ce3f7c52",
          8763 => x"a41b51ff",
          8764 => x"a0c53f82",
          8765 => x"52ac1b51",
          8766 => x"ffa0bc3f",
          8767 => x"8152b01b",
          8768 => x"51ffa095",
          8769 => x"3f8652b2",
          8770 => x"1b51ffa0",
          8771 => x"8c3fff80",
          8772 => x"0b80c01c",
          8773 => x"34a90b80",
          8774 => x"c21c3493",
          8775 => x"5382b4a8",
          8776 => x"5280c71b",
          8777 => x"51ae3982",
          8778 => x"88b20a52",
          8779 => x"a71b51ff",
          8780 => x"a0853f7c",
          8781 => x"83ffff06",
          8782 => x"52961b51",
          8783 => x"ff9fda3f",
          8784 => x"ff800ba4",
          8785 => x"1c34a90b",
          8786 => x"a61c3493",
          8787 => x"5382b4bc",
          8788 => x"52ab1b51",
          8789 => x"ffa08f3f",
          8790 => x"82d4d552",
          8791 => x"83fe1b70",
          8792 => x"5259ff9f",
          8793 => x"b43f8154",
          8794 => x"60537a52",
          8795 => x"7e51ff9b",
          8796 => x"d73f8156",
          8797 => x"82bb9808",
          8798 => x"83e7387d",
          8799 => x"832e0981",
          8800 => x"0680ee38",
          8801 => x"75546086",
          8802 => x"05537a52",
          8803 => x"7e51ff9b",
          8804 => x"b73f8480",
          8805 => x"5380527a",
          8806 => x"51ff9fed",
          8807 => x"3f848b85",
          8808 => x"a4d2527a",
          8809 => x"51ff9f8f",
          8810 => x"3f868a85",
          8811 => x"e4f25283",
          8812 => x"e41b51ff",
          8813 => x"9f813fff",
          8814 => x"185283e8",
          8815 => x"1b51ff9e",
          8816 => x"f63f8252",
          8817 => x"83ec1b51",
          8818 => x"ff9eec3f",
          8819 => x"82d4d552",
          8820 => x"7851ff9e",
          8821 => x"c43f7554",
          8822 => x"60870553",
          8823 => x"7a527e51",
          8824 => x"ff9ae53f",
          8825 => x"75546016",
          8826 => x"537a527e",
          8827 => x"51ff9ad8",
          8828 => x"3f655380",
          8829 => x"527a51ff",
          8830 => x"9f8f3f7f",
          8831 => x"5680587d",
          8832 => x"832e0981",
          8833 => x"069a38f8",
          8834 => x"527a51ff",
          8835 => x"9ea93fff",
          8836 => x"52841b51",
          8837 => x"ff9ea03f",
          8838 => x"f00a5288",
          8839 => x"1b519139",
          8840 => x"87fffff8",
          8841 => x"557d812e",
          8842 => x"8338f855",
          8843 => x"74527a51",
          8844 => x"ff9e843f",
          8845 => x"7c556157",
          8846 => x"74622683",
          8847 => x"38745776",
          8848 => x"5475537a",
          8849 => x"527e51ff",
          8850 => x"99fe3f82",
          8851 => x"bb980882",
          8852 => x"87388480",
          8853 => x"5382bb98",
          8854 => x"08527a51",
          8855 => x"ff9eaa3f",
          8856 => x"76167578",
          8857 => x"31565674",
          8858 => x"cd388118",
          8859 => x"5877802e",
          8860 => x"ff8d3879",
          8861 => x"557d832e",
          8862 => x"83386355",
          8863 => x"61577462",
          8864 => x"26833874",
          8865 => x"57765475",
          8866 => x"537a527e",
          8867 => x"51ff99b8",
          8868 => x"3f82bb98",
          8869 => x"0881c138",
          8870 => x"76167578",
          8871 => x"31565674",
          8872 => x"db388c56",
          8873 => x"7d832e93",
          8874 => x"38865666",
          8875 => x"83ffff26",
          8876 => x"8a388456",
          8877 => x"7d822e83",
          8878 => x"38815664",
          8879 => x"81065877",
          8880 => x"80fe3884",
          8881 => x"80537752",
          8882 => x"7a51ff9d",
          8883 => x"bc3f82d4",
          8884 => x"d5527851",
          8885 => x"ff9cc23f",
          8886 => x"83be1b55",
          8887 => x"77753481",
          8888 => x"0b811634",
          8889 => x"810b8216",
          8890 => x"34778316",
          8891 => x"34758416",
          8892 => x"34606705",
          8893 => x"5680fdc1",
          8894 => x"527551fe",
          8895 => x"bca53ffe",
          8896 => x"0b851634",
          8897 => x"82bb9808",
          8898 => x"822abf07",
          8899 => x"56758616",
          8900 => x"3482bb98",
          8901 => x"08871634",
          8902 => x"605283c6",
          8903 => x"1b51ff9c",
          8904 => x"963f6652",
          8905 => x"83ca1b51",
          8906 => x"ff9c8c3f",
          8907 => x"81547753",
          8908 => x"7a527e51",
          8909 => x"ff98913f",
          8910 => x"815682bb",
          8911 => x"9808a238",
          8912 => x"80538052",
          8913 => x"7e51ff99",
          8914 => x"e33f8156",
          8915 => x"82bb9808",
          8916 => x"90388939",
          8917 => x"8e568a39",
          8918 => x"81568639",
          8919 => x"82bb9808",
          8920 => x"567582bb",
          8921 => x"980c993d",
          8922 => x"0d04f53d",
          8923 => x"0d7d605b",
          8924 => x"59807960",
          8925 => x"ff055a57",
          8926 => x"57767825",
          8927 => x"b4388d3d",
          8928 => x"f8115555",
          8929 => x"8153fc15",
          8930 => x"527951c9",
          8931 => x"dc3f7a81",
          8932 => x"2e098106",
          8933 => x"9c388c3d",
          8934 => x"3355748d",
          8935 => x"2edb3874",
          8936 => x"76708105",
          8937 => x"58348117",
          8938 => x"57748a2e",
          8939 => x"098106c9",
          8940 => x"38807634",
          8941 => x"78557683",
          8942 => x"38765574",
          8943 => x"82bb980c",
          8944 => x"8d3d0d04",
          8945 => x"f73d0d7b",
          8946 => x"028405b3",
          8947 => x"05335957",
          8948 => x"778a2e09",
          8949 => x"81068738",
          8950 => x"8d527651",
          8951 => x"e73f8417",
          8952 => x"08568076",
          8953 => x"24be3888",
          8954 => x"17087717",
          8955 => x"8c055659",
          8956 => x"77753481",
          8957 => x"1656bb76",
          8958 => x"25a1388b",
          8959 => x"3dfc0554",
          8960 => x"75538c17",
          8961 => x"52760851",
          8962 => x"cbdc3f79",
          8963 => x"76327030",
          8964 => x"7072079f",
          8965 => x"2a703053",
          8966 => x"51565675",
          8967 => x"84180c81",
          8968 => x"1988180c",
          8969 => x"8b3d0d04",
          8970 => x"f93d0d79",
          8971 => x"84110856",
          8972 => x"56807524",
          8973 => x"a738893d",
          8974 => x"fc055474",
          8975 => x"538c1652",
          8976 => x"750851cb",
          8977 => x"a13f82bb",
          8978 => x"98089138",
          8979 => x"84160878",
          8980 => x"2e098106",
          8981 => x"87388816",
          8982 => x"08558339",
          8983 => x"ff557482",
          8984 => x"bb980c89",
          8985 => x"3d0d04fd",
          8986 => x"3d0d7554",
          8987 => x"80cc5380",
          8988 => x"527351ff",
          8989 => x"9a933f76",
          8990 => x"740c853d",
          8991 => x"0d04ea3d",
          8992 => x"0d0280e3",
          8993 => x"05336a53",
          8994 => x"863d7053",
          8995 => x"5454d83f",
          8996 => x"73527251",
          8997 => x"feae3f72",
          8998 => x"51ff8d3f",
          8999 => x"983d0d04",
          9000 => x"00ffffff",
          9001 => x"ff00ffff",
          9002 => x"ffff00ff",
          9003 => x"ffffff00",
          9004 => x"00002ba8",
          9005 => x"00002b2c",
          9006 => x"00002b33",
          9007 => x"00002b3a",
          9008 => x"00002b41",
          9009 => x"00002b48",
          9010 => x"00002b4f",
          9011 => x"00002b56",
          9012 => x"00002b5d",
          9013 => x"00002b64",
          9014 => x"00002b6b",
          9015 => x"00002b72",
          9016 => x"00002b78",
          9017 => x"00002b7e",
          9018 => x"00002b84",
          9019 => x"00002b8a",
          9020 => x"00002b90",
          9021 => x"00002b96",
          9022 => x"00002b9c",
          9023 => x"00002ba2",
          9024 => x"0000436a",
          9025 => x"00004370",
          9026 => x"00004376",
          9027 => x"0000437c",
          9028 => x"00004382",
          9029 => x"00004993",
          9030 => x"00004a89",
          9031 => x"00004b81",
          9032 => x"00004dbb",
          9033 => x"00004a71",
          9034 => x"00004868",
          9035 => x"00004c35",
          9036 => x"00004d91",
          9037 => x"00004c73",
          9038 => x"00004d09",
          9039 => x"00004c8f",
          9040 => x"00004b30",
          9041 => x"00004868",
          9042 => x"00004b81",
          9043 => x"00004ba5",
          9044 => x"00004c35",
          9045 => x"00004868",
          9046 => x"00004868",
          9047 => x"00004c8f",
          9048 => x"00004d09",
          9049 => x"00004d91",
          9050 => x"00004dbb",
          9051 => x"00000e2f",
          9052 => x"00001718",
          9053 => x"00001718",
          9054 => x"00000e5e",
          9055 => x"00001718",
          9056 => x"00001718",
          9057 => x"00001718",
          9058 => x"00001718",
          9059 => x"00001718",
          9060 => x"00001718",
          9061 => x"00001718",
          9062 => x"00000e1b",
          9063 => x"00001718",
          9064 => x"00000e46",
          9065 => x"00000e76",
          9066 => x"00001718",
          9067 => x"00001718",
          9068 => x"00001718",
          9069 => x"00001718",
          9070 => x"00001718",
          9071 => x"00001718",
          9072 => x"00001718",
          9073 => x"00001718",
          9074 => x"00001718",
          9075 => x"00001718",
          9076 => x"00001718",
          9077 => x"00001718",
          9078 => x"00001718",
          9079 => x"00001718",
          9080 => x"00001718",
          9081 => x"00001718",
          9082 => x"00001718",
          9083 => x"00001718",
          9084 => x"00001718",
          9085 => x"00001718",
          9086 => x"00001718",
          9087 => x"00001718",
          9088 => x"00001718",
          9089 => x"00001718",
          9090 => x"00001718",
          9091 => x"00001718",
          9092 => x"00001718",
          9093 => x"00001718",
          9094 => x"00001718",
          9095 => x"00001718",
          9096 => x"00001718",
          9097 => x"00001718",
          9098 => x"00001718",
          9099 => x"00001718",
          9100 => x"00001718",
          9101 => x"00001718",
          9102 => x"00000fa6",
          9103 => x"00001718",
          9104 => x"00001718",
          9105 => x"00001718",
          9106 => x"00001718",
          9107 => x"00001114",
          9108 => x"00001718",
          9109 => x"00001718",
          9110 => x"00001718",
          9111 => x"00001718",
          9112 => x"00001718",
          9113 => x"00001718",
          9114 => x"00001718",
          9115 => x"00001718",
          9116 => x"00001718",
          9117 => x"00001718",
          9118 => x"00000ed6",
          9119 => x"0000103d",
          9120 => x"00000ead",
          9121 => x"00000ead",
          9122 => x"00000ead",
          9123 => x"00001718",
          9124 => x"0000103d",
          9125 => x"00001718",
          9126 => x"00001718",
          9127 => x"00000e96",
          9128 => x"00001718",
          9129 => x"00001718",
          9130 => x"000010ea",
          9131 => x"000010f5",
          9132 => x"00001718",
          9133 => x"00001718",
          9134 => x"00000f0f",
          9135 => x"00001718",
          9136 => x"0000111d",
          9137 => x"00001718",
          9138 => x"00001718",
          9139 => x"00001114",
          9140 => x"64696e69",
          9141 => x"74000000",
          9142 => x"64696f63",
          9143 => x"746c0000",
          9144 => x"66696e69",
          9145 => x"74000000",
          9146 => x"666c6f61",
          9147 => x"64000000",
          9148 => x"66657865",
          9149 => x"63000000",
          9150 => x"6d636c65",
          9151 => x"61720000",
          9152 => x"6d636f70",
          9153 => x"79000000",
          9154 => x"6d646966",
          9155 => x"66000000",
          9156 => x"6d64756d",
          9157 => x"70000000",
          9158 => x"6d656200",
          9159 => x"6d656800",
          9160 => x"6d657700",
          9161 => x"68696400",
          9162 => x"68696500",
          9163 => x"68666400",
          9164 => x"68666500",
          9165 => x"63616c6c",
          9166 => x"00000000",
          9167 => x"6a6d7000",
          9168 => x"72657374",
          9169 => x"61727400",
          9170 => x"72657365",
          9171 => x"74000000",
          9172 => x"696e666f",
          9173 => x"00000000",
          9174 => x"74657374",
          9175 => x"00000000",
          9176 => x"74626173",
          9177 => x"69630000",
          9178 => x"6d626173",
          9179 => x"69630000",
          9180 => x"6b696c6f",
          9181 => x"00000000",
          9182 => x"65640000",
          9183 => x"4469736b",
          9184 => x"20457272",
          9185 => x"6f720a00",
          9186 => x"496e7465",
          9187 => x"726e616c",
          9188 => x"20657272",
          9189 => x"6f722e0a",
          9190 => x"00000000",
          9191 => x"4469736b",
          9192 => x"206e6f74",
          9193 => x"20726561",
          9194 => x"64792e0a",
          9195 => x"00000000",
          9196 => x"4e6f2066",
          9197 => x"696c6520",
          9198 => x"666f756e",
          9199 => x"642e0a00",
          9200 => x"4e6f2070",
          9201 => x"61746820",
          9202 => x"666f756e",
          9203 => x"642e0a00",
          9204 => x"496e7661",
          9205 => x"6c696420",
          9206 => x"66696c65",
          9207 => x"6e616d65",
          9208 => x"2e0a0000",
          9209 => x"41636365",
          9210 => x"73732064",
          9211 => x"656e6965",
          9212 => x"642e0a00",
          9213 => x"46696c65",
          9214 => x"20616c72",
          9215 => x"65616479",
          9216 => x"20657869",
          9217 => x"7374732e",
          9218 => x"0a000000",
          9219 => x"46696c65",
          9220 => x"2068616e",
          9221 => x"646c6520",
          9222 => x"696e7661",
          9223 => x"6c69642e",
          9224 => x"0a000000",
          9225 => x"53442069",
          9226 => x"73207772",
          9227 => x"69746520",
          9228 => x"70726f74",
          9229 => x"65637465",
          9230 => x"642e0a00",
          9231 => x"44726976",
          9232 => x"65206e75",
          9233 => x"6d626572",
          9234 => x"20697320",
          9235 => x"696e7661",
          9236 => x"6c69642e",
          9237 => x"0a000000",
          9238 => x"4469736b",
          9239 => x"206e6f74",
          9240 => x"20656e61",
          9241 => x"626c6564",
          9242 => x"2e0a0000",
          9243 => x"4e6f2063",
          9244 => x"6f6d7061",
          9245 => x"7469626c",
          9246 => x"65206669",
          9247 => x"6c657379",
          9248 => x"7374656d",
          9249 => x"20666f75",
          9250 => x"6e64206f",
          9251 => x"6e206469",
          9252 => x"736b2e0a",
          9253 => x"00000000",
          9254 => x"466f726d",
          9255 => x"61742061",
          9256 => x"626f7274",
          9257 => x"65642e0a",
          9258 => x"00000000",
          9259 => x"54696d65",
          9260 => x"6f75742c",
          9261 => x"206f7065",
          9262 => x"72617469",
          9263 => x"6f6e2063",
          9264 => x"616e6365",
          9265 => x"6c6c6564",
          9266 => x"2e0a0000",
          9267 => x"46696c65",
          9268 => x"20697320",
          9269 => x"6c6f636b",
          9270 => x"65642e0a",
          9271 => x"00000000",
          9272 => x"496e7375",
          9273 => x"66666963",
          9274 => x"69656e74",
          9275 => x"206d656d",
          9276 => x"6f72792e",
          9277 => x"0a000000",
          9278 => x"546f6f20",
          9279 => x"6d616e79",
          9280 => x"206f7065",
          9281 => x"6e206669",
          9282 => x"6c65732e",
          9283 => x"0a000000",
          9284 => x"50617261",
          9285 => x"6d657465",
          9286 => x"72732069",
          9287 => x"6e636f72",
          9288 => x"72656374",
          9289 => x"2e0a0000",
          9290 => x"53756363",
          9291 => x"6573732e",
          9292 => x"0a000000",
          9293 => x"556e6b6e",
          9294 => x"6f776e20",
          9295 => x"6572726f",
          9296 => x"722e0a00",
          9297 => x"0a256c75",
          9298 => x"20627974",
          9299 => x"65732025",
          9300 => x"73206174",
          9301 => x"20256c75",
          9302 => x"20627974",
          9303 => x"65732f73",
          9304 => x"65632e0a",
          9305 => x"00000000",
          9306 => x"72656164",
          9307 => x"00000000",
          9308 => x"25303858",
          9309 => x"00000000",
          9310 => x"3a202000",
          9311 => x"25303458",
          9312 => x"00000000",
          9313 => x"20202020",
          9314 => x"20202020",
          9315 => x"00000000",
          9316 => x"25303258",
          9317 => x"00000000",
          9318 => x"20200000",
          9319 => x"207c0000",
          9320 => x"7c0d0a00",
          9321 => x"5a505554",
          9322 => x"41000000",
          9323 => x"0a2a2a20",
          9324 => x"25732028",
          9325 => x"00000000",
          9326 => x"30322f30",
          9327 => x"352f3230",
          9328 => x"32300000",
          9329 => x"76312e35",
          9330 => x"32000000",
          9331 => x"205a5055",
          9332 => x"2c207265",
          9333 => x"76202530",
          9334 => x"32782920",
          9335 => x"25732025",
          9336 => x"73202a2a",
          9337 => x"0a0a0000",
          9338 => x"5a505554",
          9339 => x"4120496e",
          9340 => x"74657272",
          9341 => x"75707420",
          9342 => x"48616e64",
          9343 => x"6c65720a",
          9344 => x"00000000",
          9345 => x"54696d65",
          9346 => x"7220696e",
          9347 => x"74657272",
          9348 => x"7570740a",
          9349 => x"00000000",
          9350 => x"50533220",
          9351 => x"696e7465",
          9352 => x"72727570",
          9353 => x"740a0000",
          9354 => x"494f4354",
          9355 => x"4c205244",
          9356 => x"20696e74",
          9357 => x"65727275",
          9358 => x"70740a00",
          9359 => x"494f4354",
          9360 => x"4c205752",
          9361 => x"20696e74",
          9362 => x"65727275",
          9363 => x"70740a00",
          9364 => x"55415254",
          9365 => x"30205258",
          9366 => x"20696e74",
          9367 => x"65727275",
          9368 => x"70740a00",
          9369 => x"55415254",
          9370 => x"30205458",
          9371 => x"20696e74",
          9372 => x"65727275",
          9373 => x"70740a00",
          9374 => x"55415254",
          9375 => x"31205258",
          9376 => x"20696e74",
          9377 => x"65727275",
          9378 => x"70740a00",
          9379 => x"55415254",
          9380 => x"31205458",
          9381 => x"20696e74",
          9382 => x"65727275",
          9383 => x"70740a00",
          9384 => x"53657474",
          9385 => x"696e6720",
          9386 => x"75702074",
          9387 => x"696d6572",
          9388 => x"2e2e2e0a",
          9389 => x"00000000",
          9390 => x"456e6162",
          9391 => x"6c696e67",
          9392 => x"2074696d",
          9393 => x"65722e2e",
          9394 => x"2e0a0000",
          9395 => x"6175746f",
          9396 => x"65786563",
          9397 => x"2e626174",
          9398 => x"00000000",
          9399 => x"7a707574",
          9400 => x"612e6873",
          9401 => x"74000000",
          9402 => x"303a0000",
          9403 => x"4661696c",
          9404 => x"65642074",
          9405 => x"6f20696e",
          9406 => x"69746961",
          9407 => x"6c697365",
          9408 => x"20736420",
          9409 => x"63617264",
          9410 => x"20302c20",
          9411 => x"706c6561",
          9412 => x"73652069",
          9413 => x"6e697420",
          9414 => x"6d616e75",
          9415 => x"616c6c79",
          9416 => x"2e000000",
          9417 => x"2a200000",
          9418 => x"42616420",
          9419 => x"6469736b",
          9420 => x"20696421",
          9421 => x"00000000",
          9422 => x"496e6974",
          9423 => x"69616c69",
          9424 => x"7365642e",
          9425 => x"0a000000",
          9426 => x"4661696c",
          9427 => x"65642074",
          9428 => x"6f20696e",
          9429 => x"69746961",
          9430 => x"6c697365",
          9431 => x"2e0a0000",
          9432 => x"72633d25",
          9433 => x"640a0000",
          9434 => x"25753a00",
          9435 => x"436c6561",
          9436 => x"72696e67",
          9437 => x"2e2e2e2e",
          9438 => x"00000000",
          9439 => x"436f7079",
          9440 => x"696e672e",
          9441 => x"2e2e0000",
          9442 => x"436f6d70",
          9443 => x"6172696e",
          9444 => x"672e2e2e",
          9445 => x"00000000",
          9446 => x"2530386c",
          9447 => x"78282530",
          9448 => x"3878292d",
          9449 => x"3e253038",
          9450 => x"6c782825",
          9451 => x"30387829",
          9452 => x"0a000000",
          9453 => x"44756d70",
          9454 => x"204d656d",
          9455 => x"6f72790a",
          9456 => x"00000000",
          9457 => x"0a436f6d",
          9458 => x"706c6574",
          9459 => x"652e0a00",
          9460 => x"25303858",
          9461 => x"20253032",
          9462 => x"582d0000",
          9463 => x"3f3f3f0a",
          9464 => x"00000000",
          9465 => x"25303858",
          9466 => x"20253034",
          9467 => x"582d0000",
          9468 => x"25303858",
          9469 => x"20253038",
          9470 => x"582d0000",
          9471 => x"44697361",
          9472 => x"626c696e",
          9473 => x"6720696e",
          9474 => x"74657272",
          9475 => x"75707473",
          9476 => x"0a000000",
          9477 => x"456e6162",
          9478 => x"6c696e67",
          9479 => x"20696e74",
          9480 => x"65727275",
          9481 => x"7074730a",
          9482 => x"00000000",
          9483 => x"44697361",
          9484 => x"626c6564",
          9485 => x"20756172",
          9486 => x"74206669",
          9487 => x"666f0a00",
          9488 => x"456e6162",
          9489 => x"6c696e67",
          9490 => x"20756172",
          9491 => x"74206669",
          9492 => x"666f0a00",
          9493 => x"45786563",
          9494 => x"7574696e",
          9495 => x"6720636f",
          9496 => x"64652040",
          9497 => x"20253038",
          9498 => x"78202e2e",
          9499 => x"2e0a0000",
          9500 => x"43616c6c",
          9501 => x"696e6720",
          9502 => x"636f6465",
          9503 => x"20402025",
          9504 => x"30387820",
          9505 => x"2e2e2e0a",
          9506 => x"00000000",
          9507 => x"43616c6c",
          9508 => x"20726574",
          9509 => x"75726e65",
          9510 => x"6420636f",
          9511 => x"64652028",
          9512 => x"2564292e",
          9513 => x"0a000000",
          9514 => x"52657374",
          9515 => x"61727469",
          9516 => x"6e672061",
          9517 => x"70706c69",
          9518 => x"63617469",
          9519 => x"6f6e2e2e",
          9520 => x"2e0a0000",
          9521 => x"436f6c64",
          9522 => x"20726562",
          9523 => x"6f6f7469",
          9524 => x"6e672e2e",
          9525 => x"2e0a0000",
          9526 => x"5a505500",
          9527 => x"62696e00",
          9528 => x"25643a5c",
          9529 => x"25735c25",
          9530 => x"732e2573",
          9531 => x"00000000",
          9532 => x"25643a5c",
          9533 => x"25735c25",
          9534 => x"73000000",
          9535 => x"25643a5c",
          9536 => x"25730000",
          9537 => x"42616420",
          9538 => x"636f6d6d",
          9539 => x"616e642e",
          9540 => x"00000000",
          9541 => x"52756e6e",
          9542 => x"696e672e",
          9543 => x"2e2e0a00",
          9544 => x"456e6162",
          9545 => x"6c696e67",
          9546 => x"20696e74",
          9547 => x"65727275",
          9548 => x"7074732e",
          9549 => x"2e2e0a00",
          9550 => x"25642f25",
          9551 => x"642f2564",
          9552 => x"2025643a",
          9553 => x"25643a25",
          9554 => x"642e2564",
          9555 => x"25640a00",
          9556 => x"536f4320",
          9557 => x"436f6e66",
          9558 => x"69677572",
          9559 => x"6174696f",
          9560 => x"6e000000",
          9561 => x"20286672",
          9562 => x"6f6d2053",
          9563 => x"6f432063",
          9564 => x"6f6e6669",
          9565 => x"67290000",
          9566 => x"3a0a4465",
          9567 => x"76696365",
          9568 => x"7320696d",
          9569 => x"706c656d",
          9570 => x"656e7465",
          9571 => x"643a0a00",
          9572 => x"20202020",
          9573 => x"57422053",
          9574 => x"4452414d",
          9575 => x"20202825",
          9576 => x"3038583a",
          9577 => x"25303858",
          9578 => x"292e0a00",
          9579 => x"20202020",
          9580 => x"53445241",
          9581 => x"4d202020",
          9582 => x"20202825",
          9583 => x"3038583a",
          9584 => x"25303858",
          9585 => x"292e0a00",
          9586 => x"20202020",
          9587 => x"494e534e",
          9588 => x"20425241",
          9589 => x"4d202825",
          9590 => x"3038583a",
          9591 => x"25303858",
          9592 => x"292e0a00",
          9593 => x"20202020",
          9594 => x"4252414d",
          9595 => x"20202020",
          9596 => x"20202825",
          9597 => x"3038583a",
          9598 => x"25303858",
          9599 => x"292e0a00",
          9600 => x"20202020",
          9601 => x"52414d20",
          9602 => x"20202020",
          9603 => x"20202825",
          9604 => x"3038583a",
          9605 => x"25303858",
          9606 => x"292e0a00",
          9607 => x"20202020",
          9608 => x"53442043",
          9609 => x"41524420",
          9610 => x"20202844",
          9611 => x"65766963",
          9612 => x"6573203d",
          9613 => x"25303264",
          9614 => x"292e0a00",
          9615 => x"20202020",
          9616 => x"54494d45",
          9617 => x"52312020",
          9618 => x"20202854",
          9619 => x"696d6572",
          9620 => x"7320203d",
          9621 => x"25303264",
          9622 => x"292e0a00",
          9623 => x"20202020",
          9624 => x"494e5452",
          9625 => x"20435452",
          9626 => x"4c202843",
          9627 => x"68616e6e",
          9628 => x"656c733d",
          9629 => x"25303264",
          9630 => x"292e0a00",
          9631 => x"20202020",
          9632 => x"57495348",
          9633 => x"424f4e45",
          9634 => x"20425553",
          9635 => x"0a000000",
          9636 => x"20202020",
          9637 => x"57422049",
          9638 => x"32430a00",
          9639 => x"20202020",
          9640 => x"494f4354",
          9641 => x"4c0a0000",
          9642 => x"20202020",
          9643 => x"5053320a",
          9644 => x"00000000",
          9645 => x"20202020",
          9646 => x"5350490a",
          9647 => x"00000000",
          9648 => x"41646472",
          9649 => x"65737365",
          9650 => x"733a0a00",
          9651 => x"20202020",
          9652 => x"43505520",
          9653 => x"52657365",
          9654 => x"74205665",
          9655 => x"63746f72",
          9656 => x"20416464",
          9657 => x"72657373",
          9658 => x"203d2025",
          9659 => x"3038580a",
          9660 => x"00000000",
          9661 => x"20202020",
          9662 => x"43505520",
          9663 => x"4d656d6f",
          9664 => x"72792053",
          9665 => x"74617274",
          9666 => x"20416464",
          9667 => x"72657373",
          9668 => x"203d2025",
          9669 => x"3038580a",
          9670 => x"00000000",
          9671 => x"20202020",
          9672 => x"53746163",
          9673 => x"6b205374",
          9674 => x"61727420",
          9675 => x"41646472",
          9676 => x"65737320",
          9677 => x"20202020",
          9678 => x"203d2025",
          9679 => x"3038580a",
          9680 => x"00000000",
          9681 => x"4d697363",
          9682 => x"3a0a0000",
          9683 => x"20202020",
          9684 => x"5a505520",
          9685 => x"49642020",
          9686 => x"20202020",
          9687 => x"20202020",
          9688 => x"20202020",
          9689 => x"20202020",
          9690 => x"203d2025",
          9691 => x"3034580a",
          9692 => x"00000000",
          9693 => x"20202020",
          9694 => x"53797374",
          9695 => x"656d2043",
          9696 => x"6c6f636b",
          9697 => x"20467265",
          9698 => x"71202020",
          9699 => x"20202020",
          9700 => x"203d2025",
          9701 => x"642e2530",
          9702 => x"34644d48",
          9703 => x"7a0a0000",
          9704 => x"20202020",
          9705 => x"53445241",
          9706 => x"4d20436c",
          9707 => x"6f636b20",
          9708 => x"46726571",
          9709 => x"20202020",
          9710 => x"20202020",
          9711 => x"203d2025",
          9712 => x"642e2530",
          9713 => x"34644d48",
          9714 => x"7a0a0000",
          9715 => x"20202020",
          9716 => x"57697368",
          9717 => x"626f6e65",
          9718 => x"20534452",
          9719 => x"414d2043",
          9720 => x"6c6f636b",
          9721 => x"20467265",
          9722 => x"713d2025",
          9723 => x"642e2530",
          9724 => x"34644d48",
          9725 => x"7a0a0000",
          9726 => x"536d616c",
          9727 => x"6c000000",
          9728 => x"4d656469",
          9729 => x"756d0000",
          9730 => x"466c6578",
          9731 => x"00000000",
          9732 => x"45564f00",
          9733 => x"45564f6d",
          9734 => x"696e0000",
          9735 => x"556e6b6e",
          9736 => x"6f776e00",
          9737 => x"00009980",
          9738 => x"01000000",
          9739 => x"00000002",
          9740 => x"0000997c",
          9741 => x"01000000",
          9742 => x"00000003",
          9743 => x"00009978",
          9744 => x"01000000",
          9745 => x"00000004",
          9746 => x"00009974",
          9747 => x"01000000",
          9748 => x"00000005",
          9749 => x"00009970",
          9750 => x"01000000",
          9751 => x"00000006",
          9752 => x"0000996c",
          9753 => x"01000000",
          9754 => x"00000007",
          9755 => x"00009968",
          9756 => x"01000000",
          9757 => x"00000001",
          9758 => x"00009964",
          9759 => x"01000000",
          9760 => x"00000008",
          9761 => x"00009960",
          9762 => x"01000000",
          9763 => x"0000000b",
          9764 => x"0000995c",
          9765 => x"01000000",
          9766 => x"00000009",
          9767 => x"00009958",
          9768 => x"01000000",
          9769 => x"0000000a",
          9770 => x"00009954",
          9771 => x"04000000",
          9772 => x"0000000d",
          9773 => x"00009950",
          9774 => x"04000000",
          9775 => x"0000000c",
          9776 => x"0000994c",
          9777 => x"04000000",
          9778 => x"0000000e",
          9779 => x"00009948",
          9780 => x"03000000",
          9781 => x"0000000f",
          9782 => x"00009944",
          9783 => x"04000000",
          9784 => x"0000000f",
          9785 => x"00009940",
          9786 => x"04000000",
          9787 => x"00000010",
          9788 => x"0000993c",
          9789 => x"04000000",
          9790 => x"00000011",
          9791 => x"00009938",
          9792 => x"03000000",
          9793 => x"00000012",
          9794 => x"00009934",
          9795 => x"03000000",
          9796 => x"00000013",
          9797 => x"00009930",
          9798 => x"03000000",
          9799 => x"00000014",
          9800 => x"0000992c",
          9801 => x"03000000",
          9802 => x"00000015",
          9803 => x"1b5b4400",
          9804 => x"1b5b4300",
          9805 => x"1b5b4200",
          9806 => x"1b5b4100",
          9807 => x"1b5b367e",
          9808 => x"1b5b357e",
          9809 => x"1b5b347e",
          9810 => x"1b304600",
          9811 => x"1b5b337e",
          9812 => x"1b5b327e",
          9813 => x"1b5b317e",
          9814 => x"10000000",
          9815 => x"0e000000",
          9816 => x"0d000000",
          9817 => x"0b000000",
          9818 => x"08000000",
          9819 => x"06000000",
          9820 => x"05000000",
          9821 => x"04000000",
          9822 => x"03000000",
          9823 => x"02000000",
          9824 => x"01000000",
          9825 => x"68697374",
          9826 => x"6f727900",
          9827 => x"68697374",
          9828 => x"00000000",
          9829 => x"21000000",
          9830 => x"25303464",
          9831 => x"20202573",
          9832 => x"0a000000",
          9833 => x"4661696c",
          9834 => x"65642074",
          9835 => x"6f207265",
          9836 => x"73657420",
          9837 => x"74686520",
          9838 => x"68697374",
          9839 => x"6f727920",
          9840 => x"66696c65",
          9841 => x"20746f20",
          9842 => x"454f462e",
          9843 => x"0a000000",
          9844 => x"43616e6e",
          9845 => x"6f74206f",
          9846 => x"70656e2f",
          9847 => x"63726561",
          9848 => x"74652068",
          9849 => x"6973746f",
          9850 => x"72792066",
          9851 => x"696c652c",
          9852 => x"20646973",
          9853 => x"61626c69",
          9854 => x"6e672e00",
          9855 => x"53440000",
          9856 => x"222a2b2c",
          9857 => x"3a3b3c3d",
          9858 => x"3e3f5b5d",
          9859 => x"7c7f0000",
          9860 => x"46415400",
          9861 => x"46415433",
          9862 => x"32000000",
          9863 => x"ebfe904d",
          9864 => x"53444f53",
          9865 => x"352e3000",
          9866 => x"4e4f204e",
          9867 => x"414d4520",
          9868 => x"20202046",
          9869 => x"41543332",
          9870 => x"20202000",
          9871 => x"4e4f204e",
          9872 => x"414d4520",
          9873 => x"20202046",
          9874 => x"41542020",
          9875 => x"20202000",
          9876 => x"000099fc",
          9877 => x"00000000",
          9878 => x"00000000",
          9879 => x"00000000",
          9880 => x"809a4541",
          9881 => x"8e418f80",
          9882 => x"45454549",
          9883 => x"49498e8f",
          9884 => x"9092924f",
          9885 => x"994f5555",
          9886 => x"59999a9b",
          9887 => x"9c9d9e9f",
          9888 => x"41494f55",
          9889 => x"a5a5a6a7",
          9890 => x"a8a9aaab",
          9891 => x"acadaeaf",
          9892 => x"b0b1b2b3",
          9893 => x"b4b5b6b7",
          9894 => x"b8b9babb",
          9895 => x"bcbdbebf",
          9896 => x"c0c1c2c3",
          9897 => x"c4c5c6c7",
          9898 => x"c8c9cacb",
          9899 => x"cccdcecf",
          9900 => x"d0d1d2d3",
          9901 => x"d4d5d6d7",
          9902 => x"d8d9dadb",
          9903 => x"dcdddedf",
          9904 => x"e0e1e2e3",
          9905 => x"e4e5e6e7",
          9906 => x"e8e9eaeb",
          9907 => x"ecedeeef",
          9908 => x"f0f1f2f3",
          9909 => x"f4f5f6f7",
          9910 => x"f8f9fafb",
          9911 => x"fcfdfeff",
          9912 => x"2b2e2c3b",
          9913 => x"3d5b5d2f",
          9914 => x"5c222a3a",
          9915 => x"3c3e3f7c",
          9916 => x"7f000000",
          9917 => x"00010004",
          9918 => x"00100040",
          9919 => x"01000200",
          9920 => x"00000000",
          9921 => x"00010002",
          9922 => x"00040008",
          9923 => x"00100020",
          9924 => x"00000000",
          9925 => x"00000000",
          9926 => x"00008ed0",
          9927 => x"01020100",
          9928 => x"00000000",
          9929 => x"00000000",
          9930 => x"00008ed8",
          9931 => x"01040100",
          9932 => x"00000000",
          9933 => x"00000000",
          9934 => x"00008ee0",
          9935 => x"01140300",
          9936 => x"00000000",
          9937 => x"00000000",
          9938 => x"00008ee8",
          9939 => x"012b0300",
          9940 => x"00000000",
          9941 => x"00000000",
          9942 => x"00008ef0",
          9943 => x"01300300",
          9944 => x"00000000",
          9945 => x"00000000",
          9946 => x"00008ef8",
          9947 => x"013c0400",
          9948 => x"00000000",
          9949 => x"00000000",
          9950 => x"00008f00",
          9951 => x"013d0400",
          9952 => x"00000000",
          9953 => x"00000000",
          9954 => x"00008f08",
          9955 => x"013f0400",
          9956 => x"00000000",
          9957 => x"00000000",
          9958 => x"00008f10",
          9959 => x"01400400",
          9960 => x"00000000",
          9961 => x"00000000",
          9962 => x"00008f18",
          9963 => x"01410400",
          9964 => x"00000000",
          9965 => x"00000000",
          9966 => x"00008f1c",
          9967 => x"01420400",
          9968 => x"00000000",
          9969 => x"00000000",
          9970 => x"00008f20",
          9971 => x"01430400",
          9972 => x"00000000",
          9973 => x"00000000",
          9974 => x"00008f24",
          9975 => x"01500500",
          9976 => x"00000000",
          9977 => x"00000000",
          9978 => x"00008f28",
          9979 => x"01510500",
          9980 => x"00000000",
          9981 => x"00000000",
          9982 => x"00008f2c",
          9983 => x"01540500",
          9984 => x"00000000",
          9985 => x"00000000",
          9986 => x"00008f30",
          9987 => x"01550500",
          9988 => x"00000000",
          9989 => x"00000000",
          9990 => x"00008f34",
          9991 => x"01790700",
          9992 => x"00000000",
          9993 => x"00000000",
          9994 => x"00008f3c",
          9995 => x"01780700",
          9996 => x"00000000",
          9997 => x"00000000",
          9998 => x"00008f40",
          9999 => x"01820800",
         10000 => x"00000000",
         10001 => x"00000000",
         10002 => x"00008f48",
         10003 => x"01830800",
         10004 => x"00000000",
         10005 => x"00000000",
         10006 => x"00008f50",
         10007 => x"01850800",
         10008 => x"00000000",
         10009 => x"00000000",
         10010 => x"00008f58",
         10011 => x"01870800",
         10012 => x"00000000",
         10013 => x"00000000",
         10014 => x"00008f60",
         10015 => x"018c0900",
         10016 => x"00000000",
         10017 => x"00000000",
         10018 => x"00008f68",
         10019 => x"018d0900",
         10020 => x"00000000",
         10021 => x"00000000",
         10022 => x"00008f70",
         10023 => x"018e0900",
         10024 => x"00000000",
         10025 => x"00000000",
         10026 => x"00008f78",
         10027 => x"018f0900",
         10028 => x"00000000",
         10029 => x"00000000",
         10030 => x"00000000",
         10031 => x"00000000",
         10032 => x"00007fff",
         10033 => x"00000000",
         10034 => x"00007fff",
         10035 => x"00010000",
         10036 => x"00007fff",
         10037 => x"00010000",
         10038 => x"00810000",
         10039 => x"01000000",
         10040 => x"017fffff",
         10041 => x"00000000",
         10042 => x"00000000",
         10043 => x"00007800",
         10044 => x"00000000",
         10045 => x"05f5e100",
         10046 => x"05f5e100",
         10047 => x"05f5e100",
         10048 => x"00000000",
         10049 => x"01010101",
         10050 => x"01010101",
         10051 => x"01011001",
         10052 => x"01000000",
         10053 => x"00000000",
         10054 => x"00000000",
         10055 => x"00000000",
         10056 => x"00000000",
         10057 => x"00000000",
         10058 => x"00000000",
         10059 => x"00000000",
         10060 => x"00000000",
         10061 => x"00000000",
         10062 => x"00000000",
         10063 => x"00000000",
         10064 => x"00000000",
         10065 => x"00000000",
         10066 => x"00000000",
         10067 => x"00000000",
         10068 => x"00000000",
         10069 => x"00000000",
         10070 => x"00000000",
         10071 => x"00000000",
         10072 => x"00000000",
         10073 => x"00000000",
         10074 => x"00000000",
         10075 => x"00000000",
         10076 => x"00000000",
         10077 => x"00009984",
         10078 => x"01000000",
         10079 => x"0000998c",
         10080 => x"01000000",
         10081 => x"00009994",
         10082 => x"02000000",
         10083 => x"00000000",
         10084 => x"00000000",
         10085 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

