-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b83ff",
          2049 => x"f80d0b0b",
          2050 => x"0b93b904",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b93",
          2121 => x"9d040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b9380",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b829a",
          2210 => x"8c738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"93850400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b80c3",
          2219 => x"f42d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b80c5",
          2227 => x"e02d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"95040b0b",
          2317 => x"0b8ca404",
          2318 => x"0b0b0b8c",
          2319 => x"b3040b0b",
          2320 => x"0b8cc204",
          2321 => x"0b0b0b8c",
          2322 => x"d1040b0b",
          2323 => x"0b8ce004",
          2324 => x"0b0b0b8c",
          2325 => x"f0040b0b",
          2326 => x"0b8d8004",
          2327 => x"0b0b0b8d",
          2328 => x"8f040b0b",
          2329 => x"0b8d9e04",
          2330 => x"0b0b0b8d",
          2331 => x"ad040b0b",
          2332 => x"0b8dbd04",
          2333 => x"0b0b0b8d",
          2334 => x"cd040b0b",
          2335 => x"0b8ddd04",
          2336 => x"0b0b0b8d",
          2337 => x"ed040b0b",
          2338 => x"0b8dfd04",
          2339 => x"0b0b0b8e",
          2340 => x"8d040b0b",
          2341 => x"0b8e9d04",
          2342 => x"0b0b0b8e",
          2343 => x"ad040b0b",
          2344 => x"0b8ebd04",
          2345 => x"0b0b0b8e",
          2346 => x"cd040b0b",
          2347 => x"0b8edd04",
          2348 => x"0b0b0b8e",
          2349 => x"ed040b0b",
          2350 => x"0b8efd04",
          2351 => x"0b0b0b8f",
          2352 => x"8d040b0b",
          2353 => x"0b8f9d04",
          2354 => x"0b0b0b8f",
          2355 => x"ad040b0b",
          2356 => x"0b8fbd04",
          2357 => x"0b0b0b8f",
          2358 => x"cd040b0b",
          2359 => x"0b8fdd04",
          2360 => x"0b0b0b8f",
          2361 => x"ed040b0b",
          2362 => x"0b8ffd04",
          2363 => x"0b0b0b90",
          2364 => x"8d040b0b",
          2365 => x"0b909d04",
          2366 => x"0b0b0b90",
          2367 => x"ad040b0b",
          2368 => x"0b90bd04",
          2369 => x"0b0b0b90",
          2370 => x"cd040b0b",
          2371 => x"0b90dd04",
          2372 => x"0b0b0b90",
          2373 => x"ed040b0b",
          2374 => x"0b90fd04",
          2375 => x"0b0b0b91",
          2376 => x"8d040b0b",
          2377 => x"0b919d04",
          2378 => x"0b0b0b91",
          2379 => x"ad040b0b",
          2380 => x"0b91bd04",
          2381 => x"0b0b0b91",
          2382 => x"cd040b0b",
          2383 => x"0b91dd04",
          2384 => x"0b0b0b91",
          2385 => x"ed040b0b",
          2386 => x"0b91fd04",
          2387 => x"0b0b0b92",
          2388 => x"8d040b0b",
          2389 => x"0b929d04",
          2390 => x"0b0b0b92",
          2391 => x"ad040b0b",
          2392 => x"0b92bd04",
          2393 => x"0b0b0b92",
          2394 => x"cd04ffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0482bbe8",
          2434 => x"0c80f98d",
          2435 => x"2d82bbe8",
          2436 => x"0882d890",
          2437 => x"0482bbe8",
          2438 => x"0cb3b22d",
          2439 => x"82bbe808",
          2440 => x"82d89004",
          2441 => x"82bbe80c",
          2442 => x"afe32d82",
          2443 => x"bbe80882",
          2444 => x"d8900482",
          2445 => x"bbe80caf",
          2446 => x"ad2d82bb",
          2447 => x"e80882d8",
          2448 => x"900482bb",
          2449 => x"e80c94ad",
          2450 => x"2d82bbe8",
          2451 => x"0882d890",
          2452 => x"0482bbe8",
          2453 => x"0cb1c22d",
          2454 => x"82bbe808",
          2455 => x"82d89004",
          2456 => x"82bbe80c",
          2457 => x"80cfcc2d",
          2458 => x"82bbe808",
          2459 => x"82d89004",
          2460 => x"82bbe80c",
          2461 => x"80c9fb2d",
          2462 => x"82bbe808",
          2463 => x"82d89004",
          2464 => x"82bbe80c",
          2465 => x"93d82d82",
          2466 => x"bbe80882",
          2467 => x"d8900482",
          2468 => x"bbe80c96",
          2469 => x"c02d82bb",
          2470 => x"e80882d8",
          2471 => x"900482bb",
          2472 => x"e80c97cd",
          2473 => x"2d82bbe8",
          2474 => x"0882d890",
          2475 => x"0482bbe8",
          2476 => x"0c80fcb7",
          2477 => x"2d82bbe8",
          2478 => x"0882d890",
          2479 => x"0482bbe8",
          2480 => x"0c80fd95",
          2481 => x"2d82bbe8",
          2482 => x"0882d890",
          2483 => x"0482bbe8",
          2484 => x"0c80f4d2",
          2485 => x"2d82bbe8",
          2486 => x"0882d890",
          2487 => x"0482bbe8",
          2488 => x"0c80f6c9",
          2489 => x"2d82bbe8",
          2490 => x"0882d890",
          2491 => x"0482bbe8",
          2492 => x"0c80f7fc",
          2493 => x"2d82bbe8",
          2494 => x"0882d890",
          2495 => x"0482bbe8",
          2496 => x"0c81dcf0",
          2497 => x"2d82bbe8",
          2498 => x"0882d890",
          2499 => x"0482bbe8",
          2500 => x"0c81e9e1",
          2501 => x"2d82bbe8",
          2502 => x"0882d890",
          2503 => x"0482bbe8",
          2504 => x"0c81e1d5",
          2505 => x"2d82bbe8",
          2506 => x"0882d890",
          2507 => x"0482bbe8",
          2508 => x"0c81e4d2",
          2509 => x"2d82bbe8",
          2510 => x"0882d890",
          2511 => x"0482bbe8",
          2512 => x"0c81eef0",
          2513 => x"2d82bbe8",
          2514 => x"0882d890",
          2515 => x"0482bbe8",
          2516 => x"0c81f7d0",
          2517 => x"2d82bbe8",
          2518 => x"0882d890",
          2519 => x"0482bbe8",
          2520 => x"0c81e8c3",
          2521 => x"2d82bbe8",
          2522 => x"0882d890",
          2523 => x"0482bbe8",
          2524 => x"0c81f28f",
          2525 => x"2d82bbe8",
          2526 => x"0882d890",
          2527 => x"0482bbe8",
          2528 => x"0c81f3ae",
          2529 => x"2d82bbe8",
          2530 => x"0882d890",
          2531 => x"0482bbe8",
          2532 => x"0c81f3cd",
          2533 => x"2d82bbe8",
          2534 => x"0882d890",
          2535 => x"0482bbe8",
          2536 => x"0c81fbb7",
          2537 => x"2d82bbe8",
          2538 => x"0882d890",
          2539 => x"0482bbe8",
          2540 => x"0c81f99d",
          2541 => x"2d82bbe8",
          2542 => x"0882d890",
          2543 => x"0482bbe8",
          2544 => x"0c81fe8b",
          2545 => x"2d82bbe8",
          2546 => x"0882d890",
          2547 => x"0482bbe8",
          2548 => x"0c81f4d1",
          2549 => x"2d82bbe8",
          2550 => x"0882d890",
          2551 => x"0482bbe8",
          2552 => x"0c82818b",
          2553 => x"2d82bbe8",
          2554 => x"0882d890",
          2555 => x"0482bbe8",
          2556 => x"0c82828c",
          2557 => x"2d82bbe8",
          2558 => x"0882d890",
          2559 => x"0482bbe8",
          2560 => x"0c81eac1",
          2561 => x"2d82bbe8",
          2562 => x"0882d890",
          2563 => x"0482bbe8",
          2564 => x"0c81ea9a",
          2565 => x"2d82bbe8",
          2566 => x"0882d890",
          2567 => x"0482bbe8",
          2568 => x"0c81ebc5",
          2569 => x"2d82bbe8",
          2570 => x"0882d890",
          2571 => x"0482bbe8",
          2572 => x"0c81f5a8",
          2573 => x"2d82bbe8",
          2574 => x"0882d890",
          2575 => x"0482bbe8",
          2576 => x"0c8282fd",
          2577 => x"2d82bbe8",
          2578 => x"0882d890",
          2579 => x"0482bbe8",
          2580 => x"0c828587",
          2581 => x"2d82bbe8",
          2582 => x"0882d890",
          2583 => x"0482bbe8",
          2584 => x"0c8288c9",
          2585 => x"2d82bbe8",
          2586 => x"0882d890",
          2587 => x"0482bbe8",
          2588 => x"0c81dc8f",
          2589 => x"2d82bbe8",
          2590 => x"0882d890",
          2591 => x"0482bbe8",
          2592 => x"0c828bb5",
          2593 => x"2d82bbe8",
          2594 => x"0882d890",
          2595 => x"0482bbe8",
          2596 => x"0c8299ea",
          2597 => x"2d82bbe8",
          2598 => x"0882d890",
          2599 => x"0482bbe8",
          2600 => x"0c8297d6",
          2601 => x"2d82bbe8",
          2602 => x"0882d890",
          2603 => x"0482bbe8",
          2604 => x"0c81adca",
          2605 => x"2d82bbe8",
          2606 => x"0882d890",
          2607 => x"0482bbe8",
          2608 => x"0c81afb4",
          2609 => x"2d82bbe8",
          2610 => x"0882d890",
          2611 => x"0482bbe8",
          2612 => x"0c81b198",
          2613 => x"2d82bbe8",
          2614 => x"0882d890",
          2615 => x"0482bbe8",
          2616 => x"0c80f4fb",
          2617 => x"2d82bbe8",
          2618 => x"0882d890",
          2619 => x"0482bbe8",
          2620 => x"0c80f69f",
          2621 => x"2d82bbe8",
          2622 => x"0882d890",
          2623 => x"0482bbe8",
          2624 => x"0c80fa82",
          2625 => x"2d82bbe8",
          2626 => x"0882d890",
          2627 => x"0482bbe8",
          2628 => x"0c80d698",
          2629 => x"2d82bbe8",
          2630 => x"0882d890",
          2631 => x"0482bbe8",
          2632 => x"0c81a7de",
          2633 => x"2d82bbe8",
          2634 => x"0882d890",
          2635 => x"0482bbe8",
          2636 => x"0c81a886",
          2637 => x"2d82bbe8",
          2638 => x"0882d890",
          2639 => x"0482bbe8",
          2640 => x"0c81abfe",
          2641 => x"2d82bbe8",
          2642 => x"0882d890",
          2643 => x"0482bbe8",
          2644 => x"0c81a4c8",
          2645 => x"2d82bbe8",
          2646 => x"0882d890",
          2647 => x"043c0400",
          2648 => x"00101010",
          2649 => x"10101010",
          2650 => x"10101010",
          2651 => x"10101010",
          2652 => x"10101010",
          2653 => x"10101010",
          2654 => x"10101010",
          2655 => x"10101010",
          2656 => x"53510400",
          2657 => x"007381ff",
          2658 => x"06738306",
          2659 => x"09810583",
          2660 => x"05101010",
          2661 => x"2b0772fc",
          2662 => x"060c5151",
          2663 => x"04727280",
          2664 => x"728106ff",
          2665 => x"05097206",
          2666 => x"05711052",
          2667 => x"720a100a",
          2668 => x"5372ed38",
          2669 => x"51515351",
          2670 => x"0482bbdc",
          2671 => x"7082d3b8",
          2672 => x"278e3880",
          2673 => x"71708405",
          2674 => x"530c0b0b",
          2675 => x"0b93bc04",
          2676 => x"8c815180",
          2677 => x"f3950400",
          2678 => x"82bbe808",
          2679 => x"0282bbe8",
          2680 => x"0cfb3d0d",
          2681 => x"82bbe808",
          2682 => x"8c057082",
          2683 => x"bbe808fc",
          2684 => x"050c82bb",
          2685 => x"e808fc05",
          2686 => x"085482bb",
          2687 => x"e8088805",
          2688 => x"085382d3",
          2689 => x"b0085254",
          2690 => x"849a3f82",
          2691 => x"bbdc0870",
          2692 => x"82bbe808",
          2693 => x"f8050c82",
          2694 => x"bbe808f8",
          2695 => x"05087082",
          2696 => x"bbdc0c51",
          2697 => x"54873d0d",
          2698 => x"82bbe80c",
          2699 => x"0482bbe8",
          2700 => x"080282bb",
          2701 => x"e80cfb3d",
          2702 => x"0d82bbe8",
          2703 => x"08900508",
          2704 => x"85113370",
          2705 => x"81327081",
          2706 => x"06515151",
          2707 => x"52718f38",
          2708 => x"800b82bb",
          2709 => x"e8088c05",
          2710 => x"08258338",
          2711 => x"8d39800b",
          2712 => x"82bbe808",
          2713 => x"f4050c81",
          2714 => x"c43982bb",
          2715 => x"e8088c05",
          2716 => x"08ff0582",
          2717 => x"bbe8088c",
          2718 => x"050c800b",
          2719 => x"82bbe808",
          2720 => x"f8050c82",
          2721 => x"bbe80888",
          2722 => x"050882bb",
          2723 => x"e808fc05",
          2724 => x"0c82bbe8",
          2725 => x"08f80508",
          2726 => x"8a2e80f6",
          2727 => x"38800b82",
          2728 => x"bbe8088c",
          2729 => x"05082580",
          2730 => x"e93882bb",
          2731 => x"e8089005",
          2732 => x"0851a090",
          2733 => x"3f82bbdc",
          2734 => x"087082bb",
          2735 => x"e808f805",
          2736 => x"0c5282bb",
          2737 => x"e808f805",
          2738 => x"08ff2e09",
          2739 => x"81068d38",
          2740 => x"800b82bb",
          2741 => x"e808f405",
          2742 => x"0c80d239",
          2743 => x"82bbe808",
          2744 => x"fc050882",
          2745 => x"bbe808f8",
          2746 => x"05085353",
          2747 => x"71733482",
          2748 => x"bbe8088c",
          2749 => x"0508ff05",
          2750 => x"82bbe808",
          2751 => x"8c050c82",
          2752 => x"bbe808fc",
          2753 => x"05088105",
          2754 => x"82bbe808",
          2755 => x"fc050cff",
          2756 => x"803982bb",
          2757 => x"e808fc05",
          2758 => x"08528072",
          2759 => x"3482bbe8",
          2760 => x"08880508",
          2761 => x"7082bbe8",
          2762 => x"08f4050c",
          2763 => x"5282bbe8",
          2764 => x"08f40508",
          2765 => x"82bbdc0c",
          2766 => x"873d0d82",
          2767 => x"bbe80c04",
          2768 => x"82bbe808",
          2769 => x"0282bbe8",
          2770 => x"0cf43d0d",
          2771 => x"860b82bb",
          2772 => x"e808e505",
          2773 => x"3482bbe8",
          2774 => x"08880508",
          2775 => x"82bbe808",
          2776 => x"e0050cfe",
          2777 => x"0a0b82bb",
          2778 => x"e808e805",
          2779 => x"0c82bbe8",
          2780 => x"08900570",
          2781 => x"82bbe808",
          2782 => x"fc050c82",
          2783 => x"bbe808fc",
          2784 => x"05085482",
          2785 => x"bbe8088c",
          2786 => x"05085382",
          2787 => x"bbe808e0",
          2788 => x"05705351",
          2789 => x"54818d3f",
          2790 => x"82bbdc08",
          2791 => x"7082bbe8",
          2792 => x"08dc050c",
          2793 => x"82bbe808",
          2794 => x"ec050882",
          2795 => x"bbe80888",
          2796 => x"05080551",
          2797 => x"54807434",
          2798 => x"82bbe808",
          2799 => x"dc050870",
          2800 => x"82bbdc0c",
          2801 => x"548e3d0d",
          2802 => x"82bbe80c",
          2803 => x"0482bbe8",
          2804 => x"080282bb",
          2805 => x"e80cfb3d",
          2806 => x"0d82bbe8",
          2807 => x"08900570",
          2808 => x"82bbe808",
          2809 => x"fc050c82",
          2810 => x"bbe808fc",
          2811 => x"05085482",
          2812 => x"bbe8088c",
          2813 => x"05085382",
          2814 => x"bbe80888",
          2815 => x"05085254",
          2816 => x"a33f82bb",
          2817 => x"dc087082",
          2818 => x"bbe808f8",
          2819 => x"050c82bb",
          2820 => x"e808f805",
          2821 => x"087082bb",
          2822 => x"dc0c5154",
          2823 => x"873d0d82",
          2824 => x"bbe80c04",
          2825 => x"82bbe808",
          2826 => x"0282bbe8",
          2827 => x"0ced3d0d",
          2828 => x"800b82bb",
          2829 => x"e808e405",
          2830 => x"2382bbe8",
          2831 => x"08880508",
          2832 => x"53800b8c",
          2833 => x"140c82bb",
          2834 => x"e8088805",
          2835 => x"08851133",
          2836 => x"70812a70",
          2837 => x"81327081",
          2838 => x"06515151",
          2839 => x"51537280",
          2840 => x"2e8d38ff",
          2841 => x"0b82bbe8",
          2842 => x"08e0050c",
          2843 => x"96ac3982",
          2844 => x"bbe8088c",
          2845 => x"05085372",
          2846 => x"33537282",
          2847 => x"bbe808f8",
          2848 => x"05347281",
          2849 => x"ff065372",
          2850 => x"802e95fa",
          2851 => x"3882bbe8",
          2852 => x"088c0508",
          2853 => x"810582bb",
          2854 => x"e8088c05",
          2855 => x"0c82bbe8",
          2856 => x"08e40522",
          2857 => x"70810651",
          2858 => x"5372802e",
          2859 => x"958b3882",
          2860 => x"bbe808f8",
          2861 => x"053353af",
          2862 => x"732781fc",
          2863 => x"3882bbe8",
          2864 => x"08f80533",
          2865 => x"5372b926",
          2866 => x"81ee3882",
          2867 => x"bbe808f8",
          2868 => x"05335372",
          2869 => x"b02e0981",
          2870 => x"0680c538",
          2871 => x"82bbe808",
          2872 => x"e8053370",
          2873 => x"982b7098",
          2874 => x"2c515153",
          2875 => x"72b23882",
          2876 => x"bbe808e4",
          2877 => x"05227083",
          2878 => x"2a708132",
          2879 => x"70810651",
          2880 => x"51515372",
          2881 => x"802e9938",
          2882 => x"82bbe808",
          2883 => x"e4052270",
          2884 => x"82800751",
          2885 => x"537282bb",
          2886 => x"e808e405",
          2887 => x"23fed039",
          2888 => x"82bbe808",
          2889 => x"e8053370",
          2890 => x"982b7098",
          2891 => x"2c707083",
          2892 => x"2b721173",
          2893 => x"11515151",
          2894 => x"53515553",
          2895 => x"7282bbe8",
          2896 => x"08e80534",
          2897 => x"82bbe808",
          2898 => x"e8053354",
          2899 => x"82bbe808",
          2900 => x"f8053370",
          2901 => x"15d01151",
          2902 => x"51537282",
          2903 => x"bbe808e8",
          2904 => x"053482bb",
          2905 => x"e808e805",
          2906 => x"3370982b",
          2907 => x"70982c51",
          2908 => x"51537280",
          2909 => x"258b3880",
          2910 => x"ff0b82bb",
          2911 => x"e808e805",
          2912 => x"3482bbe8",
          2913 => x"08e40522",
          2914 => x"70832a70",
          2915 => x"81065151",
          2916 => x"5372fddb",
          2917 => x"3882bbe8",
          2918 => x"08e80533",
          2919 => x"70882b70",
          2920 => x"902b7090",
          2921 => x"2c70882c",
          2922 => x"51515151",
          2923 => x"537282bb",
          2924 => x"e808ec05",
          2925 => x"23fdb839",
          2926 => x"82bbe808",
          2927 => x"e4052270",
          2928 => x"832a7081",
          2929 => x"06515153",
          2930 => x"72802e9d",
          2931 => x"3882bbe8",
          2932 => x"08e80533",
          2933 => x"70982b70",
          2934 => x"982c5151",
          2935 => x"53728a38",
          2936 => x"810b82bb",
          2937 => x"e808e805",
          2938 => x"3482bbe8",
          2939 => x"08f80533",
          2940 => x"e01182bb",
          2941 => x"e808c405",
          2942 => x"0c5382bb",
          2943 => x"e808c405",
          2944 => x"0880d826",
          2945 => x"92943882",
          2946 => x"bbe808c4",
          2947 => x"05087082",
          2948 => x"2b829bd8",
          2949 => x"11700851",
          2950 => x"51515372",
          2951 => x"0482bbe8",
          2952 => x"08e40522",
          2953 => x"70900751",
          2954 => x"537282bb",
          2955 => x"e808e405",
          2956 => x"2382bbe8",
          2957 => x"08e40522",
          2958 => x"70a00751",
          2959 => x"537282bb",
          2960 => x"e808e405",
          2961 => x"23fca839",
          2962 => x"82bbe808",
          2963 => x"e4052270",
          2964 => x"81800751",
          2965 => x"537282bb",
          2966 => x"e808e405",
          2967 => x"23fc9039",
          2968 => x"82bbe808",
          2969 => x"e4052270",
          2970 => x"80c00751",
          2971 => x"537282bb",
          2972 => x"e808e405",
          2973 => x"23fbf839",
          2974 => x"82bbe808",
          2975 => x"e4052270",
          2976 => x"88075153",
          2977 => x"7282bbe8",
          2978 => x"08e40523",
          2979 => x"800b82bb",
          2980 => x"e808e805",
          2981 => x"34fbd839",
          2982 => x"82bbe808",
          2983 => x"e4052270",
          2984 => x"84075153",
          2985 => x"7282bbe8",
          2986 => x"08e40523",
          2987 => x"fbc139bf",
          2988 => x"0b82bbe8",
          2989 => x"08fc0534",
          2990 => x"82bbe808",
          2991 => x"ec0522ff",
          2992 => x"11515372",
          2993 => x"82bbe808",
          2994 => x"ec052380",
          2995 => x"e30b82bb",
          2996 => x"e808f805",
          2997 => x"348da839",
          2998 => x"82bbe808",
          2999 => x"90050882",
          3000 => x"bbe80890",
          3001 => x"05088405",
          3002 => x"82bbe808",
          3003 => x"90050c70",
          3004 => x"08515372",
          3005 => x"82bbe808",
          3006 => x"fc053482",
          3007 => x"bbe808ec",
          3008 => x"0522ff11",
          3009 => x"51537282",
          3010 => x"bbe808ec",
          3011 => x"05238cef",
          3012 => x"3982bbe8",
          3013 => x"08900508",
          3014 => x"82bbe808",
          3015 => x"90050884",
          3016 => x"0582bbe8",
          3017 => x"0890050c",
          3018 => x"700882bb",
          3019 => x"e808fc05",
          3020 => x"0c82bbe8",
          3021 => x"08e40522",
          3022 => x"70832a70",
          3023 => x"81065151",
          3024 => x"51537280",
          3025 => x"2eab3882",
          3026 => x"bbe808e8",
          3027 => x"05337098",
          3028 => x"2b537298",
          3029 => x"2c5382bb",
          3030 => x"e808fc05",
          3031 => x"085253a2",
          3032 => x"d83f82bb",
          3033 => x"dc085372",
          3034 => x"82bbe808",
          3035 => x"f4052399",
          3036 => x"3982bbe8",
          3037 => x"08fc0508",
          3038 => x"519d8a3f",
          3039 => x"82bbdc08",
          3040 => x"537282bb",
          3041 => x"e808f405",
          3042 => x"2382bbe8",
          3043 => x"08ec0522",
          3044 => x"5382bbe8",
          3045 => x"08f40522",
          3046 => x"73713154",
          3047 => x"547282bb",
          3048 => x"e808ec05",
          3049 => x"238bd839",
          3050 => x"82bbe808",
          3051 => x"90050882",
          3052 => x"bbe80890",
          3053 => x"05088405",
          3054 => x"82bbe808",
          3055 => x"90050c70",
          3056 => x"0882bbe8",
          3057 => x"08fc050c",
          3058 => x"82bbe808",
          3059 => x"e4052270",
          3060 => x"832a7081",
          3061 => x"06515151",
          3062 => x"5372802e",
          3063 => x"ab3882bb",
          3064 => x"e808e805",
          3065 => x"3370982b",
          3066 => x"5372982c",
          3067 => x"5382bbe8",
          3068 => x"08fc0508",
          3069 => x"5253a1c1",
          3070 => x"3f82bbdc",
          3071 => x"08537282",
          3072 => x"bbe808f4",
          3073 => x"05239939",
          3074 => x"82bbe808",
          3075 => x"fc050851",
          3076 => x"9bf33f82",
          3077 => x"bbdc0853",
          3078 => x"7282bbe8",
          3079 => x"08f40523",
          3080 => x"82bbe808",
          3081 => x"ec052253",
          3082 => x"82bbe808",
          3083 => x"f4052273",
          3084 => x"71315454",
          3085 => x"7282bbe8",
          3086 => x"08ec0523",
          3087 => x"8ac13982",
          3088 => x"bbe808e4",
          3089 => x"05227082",
          3090 => x"2a708106",
          3091 => x"51515372",
          3092 => x"802ea438",
          3093 => x"82bbe808",
          3094 => x"90050882",
          3095 => x"bbe80890",
          3096 => x"05088405",
          3097 => x"82bbe808",
          3098 => x"90050c70",
          3099 => x"0882bbe8",
          3100 => x"08dc050c",
          3101 => x"53a23982",
          3102 => x"bbe80890",
          3103 => x"050882bb",
          3104 => x"e8089005",
          3105 => x"08840582",
          3106 => x"bbe80890",
          3107 => x"050c7008",
          3108 => x"82bbe808",
          3109 => x"dc050c53",
          3110 => x"82bbe808",
          3111 => x"dc050882",
          3112 => x"bbe808fc",
          3113 => x"050c82bb",
          3114 => x"e808fc05",
          3115 => x"088025a4",
          3116 => x"3882bbe8",
          3117 => x"08e40522",
          3118 => x"70820751",
          3119 => x"537282bb",
          3120 => x"e808e405",
          3121 => x"2382bbe8",
          3122 => x"08fc0508",
          3123 => x"3082bbe8",
          3124 => x"08fc050c",
          3125 => x"82bbe808",
          3126 => x"e4052270",
          3127 => x"ffbf0651",
          3128 => x"537282bb",
          3129 => x"e808e405",
          3130 => x"2381af39",
          3131 => x"880b82bb",
          3132 => x"e808f405",
          3133 => x"23a93982",
          3134 => x"bbe808e4",
          3135 => x"05227080",
          3136 => x"c0075153",
          3137 => x"7282bbe8",
          3138 => x"08e40523",
          3139 => x"80f80b82",
          3140 => x"bbe808f8",
          3141 => x"0534900b",
          3142 => x"82bbe808",
          3143 => x"f4052382",
          3144 => x"bbe808e4",
          3145 => x"05227082",
          3146 => x"2a708106",
          3147 => x"51515372",
          3148 => x"802ea438",
          3149 => x"82bbe808",
          3150 => x"90050882",
          3151 => x"bbe80890",
          3152 => x"05088405",
          3153 => x"82bbe808",
          3154 => x"90050c70",
          3155 => x"0882bbe8",
          3156 => x"08d8050c",
          3157 => x"53a23982",
          3158 => x"bbe80890",
          3159 => x"050882bb",
          3160 => x"e8089005",
          3161 => x"08840582",
          3162 => x"bbe80890",
          3163 => x"050c7008",
          3164 => x"82bbe808",
          3165 => x"d8050c53",
          3166 => x"82bbe808",
          3167 => x"d8050882",
          3168 => x"bbe808fc",
          3169 => x"050c82bb",
          3170 => x"e808e405",
          3171 => x"2270cf06",
          3172 => x"51537282",
          3173 => x"bbe808e4",
          3174 => x"052382bb",
          3175 => x"ec0b82bb",
          3176 => x"e808f005",
          3177 => x"0c82bbe8",
          3178 => x"08f00508",
          3179 => x"82bbe808",
          3180 => x"f4052282",
          3181 => x"bbe808fc",
          3182 => x"05087155",
          3183 => x"70545654",
          3184 => x"55a3f33f",
          3185 => x"82bbdc08",
          3186 => x"53727534",
          3187 => x"82bbe808",
          3188 => x"f0050882",
          3189 => x"bbe808d4",
          3190 => x"050c82bb",
          3191 => x"e808f005",
          3192 => x"08703351",
          3193 => x"53897327",
          3194 => x"a43882bb",
          3195 => x"e808f005",
          3196 => x"08537233",
          3197 => x"5482bbe8",
          3198 => x"08f80533",
          3199 => x"7015df11",
          3200 => x"51515372",
          3201 => x"82bbe808",
          3202 => x"d0053497",
          3203 => x"3982bbe8",
          3204 => x"08f00508",
          3205 => x"537233b0",
          3206 => x"11515372",
          3207 => x"82bbe808",
          3208 => x"d0053482",
          3209 => x"bbe808d4",
          3210 => x"05085382",
          3211 => x"bbe808d0",
          3212 => x"05337334",
          3213 => x"82bbe808",
          3214 => x"f0050881",
          3215 => x"0582bbe8",
          3216 => x"08f0050c",
          3217 => x"82bbe808",
          3218 => x"f4052270",
          3219 => x"5382bbe8",
          3220 => x"08fc0508",
          3221 => x"5253a2ab",
          3222 => x"3f82bbdc",
          3223 => x"087082bb",
          3224 => x"e808fc05",
          3225 => x"0c5382bb",
          3226 => x"e808fc05",
          3227 => x"08802e84",
          3228 => x"38feb239",
          3229 => x"82bbe808",
          3230 => x"f0050882",
          3231 => x"bbec5455",
          3232 => x"72547470",
          3233 => x"75315153",
          3234 => x"7282bbe8",
          3235 => x"08fc0534",
          3236 => x"82bbe808",
          3237 => x"e4052270",
          3238 => x"b2065153",
          3239 => x"72802e94",
          3240 => x"3882bbe8",
          3241 => x"08ec0522",
          3242 => x"ff115153",
          3243 => x"7282bbe8",
          3244 => x"08ec0523",
          3245 => x"82bbe808",
          3246 => x"e4052270",
          3247 => x"862a7081",
          3248 => x"06515153",
          3249 => x"72802e80",
          3250 => x"e73882bb",
          3251 => x"e808ec05",
          3252 => x"2270902b",
          3253 => x"82bbe808",
          3254 => x"cc050c82",
          3255 => x"bbe808cc",
          3256 => x"0508902c",
          3257 => x"82bbe808",
          3258 => x"cc050c82",
          3259 => x"bbe808f4",
          3260 => x"05225153",
          3261 => x"72902e09",
          3262 => x"81069538",
          3263 => x"82bbe808",
          3264 => x"cc0508fe",
          3265 => x"05537282",
          3266 => x"bbe808c8",
          3267 => x"05239339",
          3268 => x"82bbe808",
          3269 => x"cc0508ff",
          3270 => x"05537282",
          3271 => x"bbe808c8",
          3272 => x"052382bb",
          3273 => x"e808c805",
          3274 => x"2282bbe8",
          3275 => x"08ec0523",
          3276 => x"82bbe808",
          3277 => x"e4052270",
          3278 => x"832a7081",
          3279 => x"06515153",
          3280 => x"72802e80",
          3281 => x"d03882bb",
          3282 => x"e808e805",
          3283 => x"3370982b",
          3284 => x"70982c82",
          3285 => x"bbe808fc",
          3286 => x"05335751",
          3287 => x"51537274",
          3288 => x"24973882",
          3289 => x"bbe808e4",
          3290 => x"052270f7",
          3291 => x"06515372",
          3292 => x"82bbe808",
          3293 => x"e405239d",
          3294 => x"3982bbe8",
          3295 => x"08e80533",
          3296 => x"5382bbe8",
          3297 => x"08fc0533",
          3298 => x"73713154",
          3299 => x"547282bb",
          3300 => x"e808e805",
          3301 => x"3482bbe8",
          3302 => x"08e40522",
          3303 => x"70832a70",
          3304 => x"81065151",
          3305 => x"5372802e",
          3306 => x"b13882bb",
          3307 => x"e808e805",
          3308 => x"3370882b",
          3309 => x"70902b70",
          3310 => x"902c7088",
          3311 => x"2c515151",
          3312 => x"51537254",
          3313 => x"82bbe808",
          3314 => x"ec052270",
          3315 => x"75315153",
          3316 => x"7282bbe8",
          3317 => x"08ec0523",
          3318 => x"af3982bb",
          3319 => x"e808fc05",
          3320 => x"3370882b",
          3321 => x"70902b70",
          3322 => x"902c7088",
          3323 => x"2c515151",
          3324 => x"51537254",
          3325 => x"82bbe808",
          3326 => x"ec052270",
          3327 => x"75315153",
          3328 => x"7282bbe8",
          3329 => x"08ec0523",
          3330 => x"82bbe808",
          3331 => x"e4052270",
          3332 => x"83800651",
          3333 => x"5372b038",
          3334 => x"82bbe808",
          3335 => x"ec0522ff",
          3336 => x"11545472",
          3337 => x"82bbe808",
          3338 => x"ec052373",
          3339 => x"902b7090",
          3340 => x"2c515380",
          3341 => x"73259038",
          3342 => x"82bbe808",
          3343 => x"88050852",
          3344 => x"a0518aee",
          3345 => x"3fd23982",
          3346 => x"bbe808e4",
          3347 => x"05227081",
          3348 => x"2a708106",
          3349 => x"51515372",
          3350 => x"802e9138",
          3351 => x"82bbe808",
          3352 => x"88050852",
          3353 => x"ad518aca",
          3354 => x"3f80c739",
          3355 => x"82bbe808",
          3356 => x"e4052270",
          3357 => x"842a7081",
          3358 => x"06515153",
          3359 => x"72802e90",
          3360 => x"3882bbe8",
          3361 => x"08880508",
          3362 => x"52ab518a",
          3363 => x"a53fa339",
          3364 => x"82bbe808",
          3365 => x"e4052270",
          3366 => x"852a7081",
          3367 => x"06515153",
          3368 => x"72802e8e",
          3369 => x"3882bbe8",
          3370 => x"08880508",
          3371 => x"52a0518a",
          3372 => x"813f82bb",
          3373 => x"e808e405",
          3374 => x"2270862a",
          3375 => x"70810651",
          3376 => x"51537280",
          3377 => x"2eb13882",
          3378 => x"bbe80888",
          3379 => x"050852b0",
          3380 => x"5189df3f",
          3381 => x"82bbe808",
          3382 => x"f4052253",
          3383 => x"72902e09",
          3384 => x"81069438",
          3385 => x"82bbe808",
          3386 => x"88050852",
          3387 => x"82bbe808",
          3388 => x"f8053351",
          3389 => x"89bc3f82",
          3390 => x"bbe808e4",
          3391 => x"05227088",
          3392 => x"2a708106",
          3393 => x"51515372",
          3394 => x"802eb038",
          3395 => x"82bbe808",
          3396 => x"ec0522ff",
          3397 => x"11545472",
          3398 => x"82bbe808",
          3399 => x"ec052373",
          3400 => x"902b7090",
          3401 => x"2c515380",
          3402 => x"73259038",
          3403 => x"82bbe808",
          3404 => x"88050852",
          3405 => x"b05188fa",
          3406 => x"3fd23982",
          3407 => x"bbe808e4",
          3408 => x"05227083",
          3409 => x"2a708106",
          3410 => x"51515372",
          3411 => x"802eb038",
          3412 => x"82bbe808",
          3413 => x"e80533ff",
          3414 => x"11545472",
          3415 => x"82bbe808",
          3416 => x"e8053473",
          3417 => x"982b7098",
          3418 => x"2c515380",
          3419 => x"73259038",
          3420 => x"82bbe808",
          3421 => x"88050852",
          3422 => x"b05188b6",
          3423 => x"3fd23982",
          3424 => x"bbe808e4",
          3425 => x"05227087",
          3426 => x"2a708106",
          3427 => x"51515372",
          3428 => x"b03882bb",
          3429 => x"e808ec05",
          3430 => x"22ff1154",
          3431 => x"547282bb",
          3432 => x"e808ec05",
          3433 => x"2373902b",
          3434 => x"70902c51",
          3435 => x"53807325",
          3436 => x"903882bb",
          3437 => x"e8088805",
          3438 => x"0852a051",
          3439 => x"87f43fd2",
          3440 => x"3982bbe8",
          3441 => x"08f80533",
          3442 => x"537280e3",
          3443 => x"2e098106",
          3444 => x"973882bb",
          3445 => x"e8088805",
          3446 => x"085282bb",
          3447 => x"e808fc05",
          3448 => x"335187ce",
          3449 => x"3f81ee39",
          3450 => x"82bbe808",
          3451 => x"f8053353",
          3452 => x"7280f32e",
          3453 => x"09810680",
          3454 => x"cb3882bb",
          3455 => x"e808f405",
          3456 => x"22ff1151",
          3457 => x"537282bb",
          3458 => x"e808f405",
          3459 => x"237283ff",
          3460 => x"ff065372",
          3461 => x"83ffff2e",
          3462 => x"81bb3882",
          3463 => x"bbe80888",
          3464 => x"05085282",
          3465 => x"bbe808fc",
          3466 => x"05087033",
          3467 => x"5282bbe8",
          3468 => x"08fc0508",
          3469 => x"810582bb",
          3470 => x"e808fc05",
          3471 => x"0c5386f2",
          3472 => x"3fffb739",
          3473 => x"82bbe808",
          3474 => x"f8053353",
          3475 => x"7280d32e",
          3476 => x"09810680",
          3477 => x"cb3882bb",
          3478 => x"e808f405",
          3479 => x"22ff1151",
          3480 => x"537282bb",
          3481 => x"e808f405",
          3482 => x"237283ff",
          3483 => x"ff065372",
          3484 => x"83ffff2e",
          3485 => x"80df3882",
          3486 => x"bbe80888",
          3487 => x"05085282",
          3488 => x"bbe808fc",
          3489 => x"05087033",
          3490 => x"525386a6",
          3491 => x"3f82bbe8",
          3492 => x"08fc0508",
          3493 => x"810582bb",
          3494 => x"e808fc05",
          3495 => x"0cffb739",
          3496 => x"82bbe808",
          3497 => x"f0050882",
          3498 => x"bbec2ea9",
          3499 => x"3882bbe8",
          3500 => x"08880508",
          3501 => x"5282bbe8",
          3502 => x"08f00508",
          3503 => x"ff0582bb",
          3504 => x"e808f005",
          3505 => x"0c82bbe8",
          3506 => x"08f00508",
          3507 => x"70335253",
          3508 => x"85e03fcc",
          3509 => x"3982bbe8",
          3510 => x"08e40522",
          3511 => x"70872a70",
          3512 => x"81065151",
          3513 => x"5372802e",
          3514 => x"80c33882",
          3515 => x"bbe808ec",
          3516 => x"0522ff11",
          3517 => x"54547282",
          3518 => x"bbe808ec",
          3519 => x"05237390",
          3520 => x"2b70902c",
          3521 => x"51538073",
          3522 => x"25a33882",
          3523 => x"bbe80888",
          3524 => x"050852a0",
          3525 => x"51859b3f",
          3526 => x"d23982bb",
          3527 => x"e8088805",
          3528 => x"085282bb",
          3529 => x"e808f805",
          3530 => x"33518586",
          3531 => x"3f800b82",
          3532 => x"bbe808e4",
          3533 => x"0523eab7",
          3534 => x"3982bbe8",
          3535 => x"08f80533",
          3536 => x"5372a52e",
          3537 => x"098106a8",
          3538 => x"38810b82",
          3539 => x"bbe808e4",
          3540 => x"0523800b",
          3541 => x"82bbe808",
          3542 => x"ec052380",
          3543 => x"0b82bbe8",
          3544 => x"08e80534",
          3545 => x"8a0b82bb",
          3546 => x"e808f405",
          3547 => x"23ea8039",
          3548 => x"82bbe808",
          3549 => x"88050852",
          3550 => x"82bbe808",
          3551 => x"f8053351",
          3552 => x"84b03fe9",
          3553 => x"ea3982bb",
          3554 => x"e8088805",
          3555 => x"088c1108",
          3556 => x"7082bbe8",
          3557 => x"08e0050c",
          3558 => x"515382bb",
          3559 => x"e808e005",
          3560 => x"0882bbdc",
          3561 => x"0c953d0d",
          3562 => x"82bbe80c",
          3563 => x"0482bbe8",
          3564 => x"080282bb",
          3565 => x"e80cfd3d",
          3566 => x"0d82d3ac",
          3567 => x"085382bb",
          3568 => x"e8088c05",
          3569 => x"085282bb",
          3570 => x"e8088805",
          3571 => x"0851e4dd",
          3572 => x"3f82bbdc",
          3573 => x"087082bb",
          3574 => x"dc0c5485",
          3575 => x"3d0d82bb",
          3576 => x"e80c0482",
          3577 => x"bbe80802",
          3578 => x"82bbe80c",
          3579 => x"fb3d0d80",
          3580 => x"0b82bbe8",
          3581 => x"08f8050c",
          3582 => x"82d3b008",
          3583 => x"85113370",
          3584 => x"812a7081",
          3585 => x"32708106",
          3586 => x"51515151",
          3587 => x"5372802e",
          3588 => x"8d38ff0b",
          3589 => x"82bbe808",
          3590 => x"f4050c81",
          3591 => x"923982bb",
          3592 => x"e8088805",
          3593 => x"08537233",
          3594 => x"82bbe808",
          3595 => x"88050881",
          3596 => x"0582bbe8",
          3597 => x"0888050c",
          3598 => x"537282bb",
          3599 => x"e808fc05",
          3600 => x"347281ff",
          3601 => x"06537280",
          3602 => x"2eb03882",
          3603 => x"d3b00882",
          3604 => x"d3b00853",
          3605 => x"82bbe808",
          3606 => x"fc053352",
          3607 => x"90110851",
          3608 => x"53722d82",
          3609 => x"bbdc0853",
          3610 => x"72802eff",
          3611 => x"b138ff0b",
          3612 => x"82bbe808",
          3613 => x"f8050cff",
          3614 => x"a53982d3",
          3615 => x"b00882d3",
          3616 => x"b0085353",
          3617 => x"8a519013",
          3618 => x"0853722d",
          3619 => x"82bbdc08",
          3620 => x"5372802e",
          3621 => x"8a38ff0b",
          3622 => x"82bbe808",
          3623 => x"f8050c82",
          3624 => x"bbe808f8",
          3625 => x"05087082",
          3626 => x"bbe808f4",
          3627 => x"050c5382",
          3628 => x"bbe808f4",
          3629 => x"050882bb",
          3630 => x"dc0c873d",
          3631 => x"0d82bbe8",
          3632 => x"0c0482bb",
          3633 => x"e8080282",
          3634 => x"bbe80cfb",
          3635 => x"3d0d800b",
          3636 => x"82bbe808",
          3637 => x"f8050c82",
          3638 => x"bbe8088c",
          3639 => x"05088511",
          3640 => x"3370812a",
          3641 => x"70813270",
          3642 => x"81065151",
          3643 => x"51515372",
          3644 => x"802e8d38",
          3645 => x"ff0b82bb",
          3646 => x"e808f405",
          3647 => x"0c80f339",
          3648 => x"82bbe808",
          3649 => x"88050853",
          3650 => x"723382bb",
          3651 => x"e8088805",
          3652 => x"08810582",
          3653 => x"bbe80888",
          3654 => x"050c5372",
          3655 => x"82bbe808",
          3656 => x"fc053472",
          3657 => x"81ff0653",
          3658 => x"72802eb6",
          3659 => x"3882bbe8",
          3660 => x"088c0508",
          3661 => x"82bbe808",
          3662 => x"8c050853",
          3663 => x"82bbe808",
          3664 => x"fc053352",
          3665 => x"90110851",
          3666 => x"53722d82",
          3667 => x"bbdc0853",
          3668 => x"72802eff",
          3669 => x"ab38ff0b",
          3670 => x"82bbe808",
          3671 => x"f8050cff",
          3672 => x"9f3982bb",
          3673 => x"e808f805",
          3674 => x"087082bb",
          3675 => x"e808f405",
          3676 => x"0c5382bb",
          3677 => x"e808f405",
          3678 => x"0882bbdc",
          3679 => x"0c873d0d",
          3680 => x"82bbe80c",
          3681 => x"0482bbe8",
          3682 => x"080282bb",
          3683 => x"e80cfe3d",
          3684 => x"0d82d3b0",
          3685 => x"085282bb",
          3686 => x"e8088805",
          3687 => x"0851933f",
          3688 => x"82bbdc08",
          3689 => x"7082bbdc",
          3690 => x"0c53843d",
          3691 => x"0d82bbe8",
          3692 => x"0c0482bb",
          3693 => x"e8080282",
          3694 => x"bbe80cfb",
          3695 => x"3d0d82bb",
          3696 => x"e8088c05",
          3697 => x"08851133",
          3698 => x"70812a70",
          3699 => x"81327081",
          3700 => x"06515151",
          3701 => x"51537280",
          3702 => x"2e8d38ff",
          3703 => x"0b82bbe8",
          3704 => x"08fc050c",
          3705 => x"81cb3982",
          3706 => x"bbe8088c",
          3707 => x"05088511",
          3708 => x"3370822a",
          3709 => x"70810651",
          3710 => x"51515372",
          3711 => x"802e80db",
          3712 => x"3882bbe8",
          3713 => x"088c0508",
          3714 => x"82bbe808",
          3715 => x"8c050854",
          3716 => x"548c1408",
          3717 => x"88140825",
          3718 => x"9f3882bb",
          3719 => x"e8088c05",
          3720 => x"08700870",
          3721 => x"82bbe808",
          3722 => x"88050852",
          3723 => x"57545472",
          3724 => x"75347308",
          3725 => x"8105740c",
          3726 => x"82bbe808",
          3727 => x"8c05088c",
          3728 => x"11088105",
          3729 => x"8c120c82",
          3730 => x"bbe80888",
          3731 => x"05087082",
          3732 => x"bbe808fc",
          3733 => x"050c5153",
          3734 => x"80d73982",
          3735 => x"bbe8088c",
          3736 => x"050882bb",
          3737 => x"e8088c05",
          3738 => x"085382bb",
          3739 => x"e8088805",
          3740 => x"087081ff",
          3741 => x"06539012",
          3742 => x"08515454",
          3743 => x"722d82bb",
          3744 => x"dc085372",
          3745 => x"a33882bb",
          3746 => x"e8088c05",
          3747 => x"088c1108",
          3748 => x"81058c12",
          3749 => x"0c82bbe8",
          3750 => x"08880508",
          3751 => x"7082bbe8",
          3752 => x"08fc050c",
          3753 => x"51538a39",
          3754 => x"ff0b82bb",
          3755 => x"e808fc05",
          3756 => x"0c82bbe8",
          3757 => x"08fc0508",
          3758 => x"82bbdc0c",
          3759 => x"873d0d82",
          3760 => x"bbe80c04",
          3761 => x"82bbe808",
          3762 => x"0282bbe8",
          3763 => x"0cf93d0d",
          3764 => x"82bbe808",
          3765 => x"88050885",
          3766 => x"11337081",
          3767 => x"32708106",
          3768 => x"51515152",
          3769 => x"71802e8d",
          3770 => x"38ff0b82",
          3771 => x"bbe808f8",
          3772 => x"050c8394",
          3773 => x"3982bbe8",
          3774 => x"08880508",
          3775 => x"85113370",
          3776 => x"862a7081",
          3777 => x"06515151",
          3778 => x"5271802e",
          3779 => x"80c53882",
          3780 => x"bbe80888",
          3781 => x"050882bb",
          3782 => x"e8088805",
          3783 => x"08535385",
          3784 => x"123370ff",
          3785 => x"bf065152",
          3786 => x"71851434",
          3787 => x"82bbe808",
          3788 => x"8805088c",
          3789 => x"11088105",
          3790 => x"8c120c82",
          3791 => x"bbe80888",
          3792 => x"05088411",
          3793 => x"337082bb",
          3794 => x"e808f805",
          3795 => x"0c515152",
          3796 => x"82b63982",
          3797 => x"bbe80888",
          3798 => x"05088511",
          3799 => x"3370822a",
          3800 => x"70810651",
          3801 => x"51515271",
          3802 => x"802e80d7",
          3803 => x"3882bbe8",
          3804 => x"08880508",
          3805 => x"70087033",
          3806 => x"82bbe808",
          3807 => x"fc050c51",
          3808 => x"5282bbe8",
          3809 => x"08fc0508",
          3810 => x"a93882bb",
          3811 => x"e8088805",
          3812 => x"0882bbe8",
          3813 => x"08880508",
          3814 => x"53538512",
          3815 => x"3370a007",
          3816 => x"51527185",
          3817 => x"1434ff0b",
          3818 => x"82bbe808",
          3819 => x"f8050c81",
          3820 => x"d73982bb",
          3821 => x"e8088805",
          3822 => x"08700881",
          3823 => x"05710c52",
          3824 => x"81a13982",
          3825 => x"bbe80888",
          3826 => x"050882bb",
          3827 => x"e8088805",
          3828 => x"08529411",
          3829 => x"08515271",
          3830 => x"2d82bbdc",
          3831 => x"087082bb",
          3832 => x"e808fc05",
          3833 => x"0c5282bb",
          3834 => x"e808fc05",
          3835 => x"08802580",
          3836 => x"f23882bb",
          3837 => x"e8088805",
          3838 => x"0882bbe8",
          3839 => x"08f4050c",
          3840 => x"82bbe808",
          3841 => x"88050885",
          3842 => x"113382bb",
          3843 => x"e808f005",
          3844 => x"0c5282bb",
          3845 => x"e808fc05",
          3846 => x"08ff2e09",
          3847 => x"81069538",
          3848 => x"82bbe808",
          3849 => x"f0050890",
          3850 => x"07527182",
          3851 => x"bbe808ec",
          3852 => x"05349339",
          3853 => x"82bbe808",
          3854 => x"f00508a0",
          3855 => x"07527182",
          3856 => x"bbe808ec",
          3857 => x"053482bb",
          3858 => x"e808f405",
          3859 => x"085282bb",
          3860 => x"e808ec05",
          3861 => x"33851334",
          3862 => x"ff0b82bb",
          3863 => x"e808f805",
          3864 => x"0ca63982",
          3865 => x"bbe80888",
          3866 => x"05088c11",
          3867 => x"0881058c",
          3868 => x"120c82bb",
          3869 => x"e808fc05",
          3870 => x"087081ff",
          3871 => x"067082bb",
          3872 => x"e808f805",
          3873 => x"0c515152",
          3874 => x"82bbe808",
          3875 => x"f8050882",
          3876 => x"bbdc0c89",
          3877 => x"3d0d82bb",
          3878 => x"e80c0482",
          3879 => x"bbe80802",
          3880 => x"82bbe80c",
          3881 => x"fd3d0d82",
          3882 => x"bbe80888",
          3883 => x"050882bb",
          3884 => x"e808fc05",
          3885 => x"0c82bbe8",
          3886 => x"088c0508",
          3887 => x"82bbe808",
          3888 => x"f8050c82",
          3889 => x"bbe80890",
          3890 => x"0508802e",
          3891 => x"82a23882",
          3892 => x"bbe808f8",
          3893 => x"050882bb",
          3894 => x"e808fc05",
          3895 => x"082681ac",
          3896 => x"3882bbe8",
          3897 => x"08f80508",
          3898 => x"82bbe808",
          3899 => x"90050805",
          3900 => x"5182bbe8",
          3901 => x"08fc0508",
          3902 => x"71278190",
          3903 => x"3882bbe8",
          3904 => x"08fc0508",
          3905 => x"82bbe808",
          3906 => x"90050805",
          3907 => x"82bbe808",
          3908 => x"fc050c82",
          3909 => x"bbe808f8",
          3910 => x"050882bb",
          3911 => x"e8089005",
          3912 => x"080582bb",
          3913 => x"e808f805",
          3914 => x"0c82bbe8",
          3915 => x"08900508",
          3916 => x"810582bb",
          3917 => x"e8089005",
          3918 => x"0c82bbe8",
          3919 => x"08900508",
          3920 => x"ff0582bb",
          3921 => x"e8089005",
          3922 => x"0c82bbe8",
          3923 => x"08900508",
          3924 => x"802e819c",
          3925 => x"3882bbe8",
          3926 => x"08fc0508",
          3927 => x"ff0582bb",
          3928 => x"e808fc05",
          3929 => x"0c82bbe8",
          3930 => x"08f80508",
          3931 => x"ff0582bb",
          3932 => x"e808f805",
          3933 => x"0c82bbe8",
          3934 => x"08fc0508",
          3935 => x"82bbe808",
          3936 => x"f8050853",
          3937 => x"51713371",
          3938 => x"34ffae39",
          3939 => x"82bbe808",
          3940 => x"90050881",
          3941 => x"0582bbe8",
          3942 => x"0890050c",
          3943 => x"82bbe808",
          3944 => x"900508ff",
          3945 => x"0582bbe8",
          3946 => x"0890050c",
          3947 => x"82bbe808",
          3948 => x"90050880",
          3949 => x"2eba3882",
          3950 => x"bbe808f8",
          3951 => x"05085170",
          3952 => x"3382bbe8",
          3953 => x"08f80508",
          3954 => x"810582bb",
          3955 => x"e808f805",
          3956 => x"0c82bbe8",
          3957 => x"08fc0508",
          3958 => x"52527171",
          3959 => x"3482bbe8",
          3960 => x"08fc0508",
          3961 => x"810582bb",
          3962 => x"e808fc05",
          3963 => x"0cffad39",
          3964 => x"82bbe808",
          3965 => x"88050870",
          3966 => x"82bbdc0c",
          3967 => x"51853d0d",
          3968 => x"82bbe80c",
          3969 => x"0482bbe8",
          3970 => x"080282bb",
          3971 => x"e80cfe3d",
          3972 => x"0d82bbe8",
          3973 => x"08880508",
          3974 => x"82bbe808",
          3975 => x"fc050c82",
          3976 => x"bbe808fc",
          3977 => x"05085271",
          3978 => x"3382bbe8",
          3979 => x"08fc0508",
          3980 => x"810582bb",
          3981 => x"e808fc05",
          3982 => x"0c7081ff",
          3983 => x"06515170",
          3984 => x"802e8338",
          3985 => x"da3982bb",
          3986 => x"e808fc05",
          3987 => x"08ff0582",
          3988 => x"bbe808fc",
          3989 => x"050c82bb",
          3990 => x"e808fc05",
          3991 => x"0882bbe8",
          3992 => x"08880508",
          3993 => x"317082bb",
          3994 => x"dc0c5184",
          3995 => x"3d0d82bb",
          3996 => x"e80c0482",
          3997 => x"bbe80802",
          3998 => x"82bbe80c",
          3999 => x"fe3d0d82",
          4000 => x"bbe80888",
          4001 => x"050882bb",
          4002 => x"e808fc05",
          4003 => x"0c82bbe8",
          4004 => x"088c0508",
          4005 => x"52713382",
          4006 => x"bbe8088c",
          4007 => x"05088105",
          4008 => x"82bbe808",
          4009 => x"8c050c82",
          4010 => x"bbe808fc",
          4011 => x"05085351",
          4012 => x"70723482",
          4013 => x"bbe808fc",
          4014 => x"05088105",
          4015 => x"82bbe808",
          4016 => x"fc050c70",
          4017 => x"81ff0651",
          4018 => x"70802e84",
          4019 => x"38ffbe39",
          4020 => x"82bbe808",
          4021 => x"88050870",
          4022 => x"82bbdc0c",
          4023 => x"51843d0d",
          4024 => x"82bbe80c",
          4025 => x"0482bbe8",
          4026 => x"080282bb",
          4027 => x"e80cfd3d",
          4028 => x"0d82bbe8",
          4029 => x"08880508",
          4030 => x"82bbe808",
          4031 => x"fc050c82",
          4032 => x"bbe8088c",
          4033 => x"050882bb",
          4034 => x"e808f805",
          4035 => x"0c82bbe8",
          4036 => x"08900508",
          4037 => x"802e80e5",
          4038 => x"3882bbe8",
          4039 => x"08900508",
          4040 => x"810582bb",
          4041 => x"e8089005",
          4042 => x"0c82bbe8",
          4043 => x"08900508",
          4044 => x"ff0582bb",
          4045 => x"e8089005",
          4046 => x"0c82bbe8",
          4047 => x"08900508",
          4048 => x"802eba38",
          4049 => x"82bbe808",
          4050 => x"f8050851",
          4051 => x"703382bb",
          4052 => x"e808f805",
          4053 => x"08810582",
          4054 => x"bbe808f8",
          4055 => x"050c82bb",
          4056 => x"e808fc05",
          4057 => x"08525271",
          4058 => x"713482bb",
          4059 => x"e808fc05",
          4060 => x"08810582",
          4061 => x"bbe808fc",
          4062 => x"050cffad",
          4063 => x"3982bbe8",
          4064 => x"08880508",
          4065 => x"7082bbdc",
          4066 => x"0c51853d",
          4067 => x"0d82bbe8",
          4068 => x"0c0482bb",
          4069 => x"e8080282",
          4070 => x"bbe80cfd",
          4071 => x"3d0d82bb",
          4072 => x"e8089005",
          4073 => x"08802e81",
          4074 => x"f43882bb",
          4075 => x"e8088c05",
          4076 => x"08527133",
          4077 => x"82bbe808",
          4078 => x"8c050881",
          4079 => x"0582bbe8",
          4080 => x"088c050c",
          4081 => x"82bbe808",
          4082 => x"88050870",
          4083 => x"337281ff",
          4084 => x"06535454",
          4085 => x"5171712e",
          4086 => x"843880ce",
          4087 => x"3982bbe8",
          4088 => x"08880508",
          4089 => x"52713382",
          4090 => x"bbe80888",
          4091 => x"05088105",
          4092 => x"82bbe808",
          4093 => x"88050c70",
          4094 => x"81ff0651",
          4095 => x"51708d38",
          4096 => x"800b82bb",
          4097 => x"e808fc05",
          4098 => x"0c819b39",
          4099 => x"82bbe808",
          4100 => x"900508ff",
          4101 => x"0582bbe8",
          4102 => x"0890050c",
          4103 => x"82bbe808",
          4104 => x"90050880",
          4105 => x"2e8438ff",
          4106 => x"813982bb",
          4107 => x"e8089005",
          4108 => x"08802e80",
          4109 => x"e83882bb",
          4110 => x"e8088805",
          4111 => x"08703352",
          4112 => x"53708d38",
          4113 => x"ff0b82bb",
          4114 => x"e808fc05",
          4115 => x"0c80d739",
          4116 => x"82bbe808",
          4117 => x"8c0508ff",
          4118 => x"0582bbe8",
          4119 => x"088c050c",
          4120 => x"82bbe808",
          4121 => x"8c050870",
          4122 => x"33525270",
          4123 => x"8c38810b",
          4124 => x"82bbe808",
          4125 => x"fc050cae",
          4126 => x"3982bbe8",
          4127 => x"08880508",
          4128 => x"703382bb",
          4129 => x"e8088c05",
          4130 => x"08703372",
          4131 => x"71317082",
          4132 => x"bbe808fc",
          4133 => x"050c5355",
          4134 => x"5252538a",
          4135 => x"39800b82",
          4136 => x"bbe808fc",
          4137 => x"050c82bb",
          4138 => x"e808fc05",
          4139 => x"0882bbdc",
          4140 => x"0c853d0d",
          4141 => x"82bbe80c",
          4142 => x"0482bbe8",
          4143 => x"080282bb",
          4144 => x"e80cfd3d",
          4145 => x"0d82bbe8",
          4146 => x"08880508",
          4147 => x"82bbe808",
          4148 => x"f8050c82",
          4149 => x"bbe8088c",
          4150 => x"05088d38",
          4151 => x"800b82bb",
          4152 => x"e808fc05",
          4153 => x"0c80ec39",
          4154 => x"82bbe808",
          4155 => x"f8050852",
          4156 => x"713382bb",
          4157 => x"e808f805",
          4158 => x"08810582",
          4159 => x"bbe808f8",
          4160 => x"050c7081",
          4161 => x"ff065151",
          4162 => x"70802e9f",
          4163 => x"3882bbe8",
          4164 => x"088c0508",
          4165 => x"ff0582bb",
          4166 => x"e8088c05",
          4167 => x"0c82bbe8",
          4168 => x"088c0508",
          4169 => x"ff2e8438",
          4170 => x"ffbe3982",
          4171 => x"bbe808f8",
          4172 => x"0508ff05",
          4173 => x"82bbe808",
          4174 => x"f8050c82",
          4175 => x"bbe808f8",
          4176 => x"050882bb",
          4177 => x"e8088805",
          4178 => x"08317082",
          4179 => x"bbe808fc",
          4180 => x"050c5182",
          4181 => x"bbe808fc",
          4182 => x"050882bb",
          4183 => x"dc0c853d",
          4184 => x"0d82bbe8",
          4185 => x"0c0482bb",
          4186 => x"e8080282",
          4187 => x"bbe80cfe",
          4188 => x"3d0d82bb",
          4189 => x"e8088805",
          4190 => x"0882bbe8",
          4191 => x"08fc050c",
          4192 => x"82bbe808",
          4193 => x"90050880",
          4194 => x"2e80d438",
          4195 => x"82bbe808",
          4196 => x"90050881",
          4197 => x"0582bbe8",
          4198 => x"0890050c",
          4199 => x"82bbe808",
          4200 => x"900508ff",
          4201 => x"0582bbe8",
          4202 => x"0890050c",
          4203 => x"82bbe808",
          4204 => x"90050880",
          4205 => x"2ea93882",
          4206 => x"bbe8088c",
          4207 => x"05085170",
          4208 => x"82bbe808",
          4209 => x"fc050852",
          4210 => x"52717134",
          4211 => x"82bbe808",
          4212 => x"fc050881",
          4213 => x"0582bbe8",
          4214 => x"08fc050c",
          4215 => x"ffbe3982",
          4216 => x"bbe80888",
          4217 => x"05087082",
          4218 => x"bbdc0c51",
          4219 => x"843d0d82",
          4220 => x"bbe80c04",
          4221 => x"82bbe808",
          4222 => x"0282bbe8",
          4223 => x"0cf93d0d",
          4224 => x"800b82bb",
          4225 => x"e808fc05",
          4226 => x"0c82bbe8",
          4227 => x"08880508",
          4228 => x"8025b938",
          4229 => x"82bbe808",
          4230 => x"88050830",
          4231 => x"82bbe808",
          4232 => x"88050c80",
          4233 => x"0b82bbe8",
          4234 => x"08f4050c",
          4235 => x"82bbe808",
          4236 => x"fc05088a",
          4237 => x"38810b82",
          4238 => x"bbe808f4",
          4239 => x"050c82bb",
          4240 => x"e808f405",
          4241 => x"0882bbe8",
          4242 => x"08fc050c",
          4243 => x"82bbe808",
          4244 => x"8c050880",
          4245 => x"25b93882",
          4246 => x"bbe8088c",
          4247 => x"05083082",
          4248 => x"bbe8088c",
          4249 => x"050c800b",
          4250 => x"82bbe808",
          4251 => x"f0050c82",
          4252 => x"bbe808fc",
          4253 => x"05088a38",
          4254 => x"810b82bb",
          4255 => x"e808f005",
          4256 => x"0c82bbe8",
          4257 => x"08f00508",
          4258 => x"82bbe808",
          4259 => x"fc050c80",
          4260 => x"5382bbe8",
          4261 => x"088c0508",
          4262 => x"5282bbe8",
          4263 => x"08880508",
          4264 => x"5182c53f",
          4265 => x"82bbdc08",
          4266 => x"7082bbe8",
          4267 => x"08f8050c",
          4268 => x"5482bbe8",
          4269 => x"08fc0508",
          4270 => x"802e9038",
          4271 => x"82bbe808",
          4272 => x"f8050830",
          4273 => x"82bbe808",
          4274 => x"f8050c82",
          4275 => x"bbe808f8",
          4276 => x"05087082",
          4277 => x"bbdc0c54",
          4278 => x"893d0d82",
          4279 => x"bbe80c04",
          4280 => x"82bbe808",
          4281 => x"0282bbe8",
          4282 => x"0cfb3d0d",
          4283 => x"800b82bb",
          4284 => x"e808fc05",
          4285 => x"0c82bbe8",
          4286 => x"08880508",
          4287 => x"80259938",
          4288 => x"82bbe808",
          4289 => x"88050830",
          4290 => x"82bbe808",
          4291 => x"88050c81",
          4292 => x"0b82bbe8",
          4293 => x"08fc050c",
          4294 => x"82bbe808",
          4295 => x"8c050880",
          4296 => x"25903882",
          4297 => x"bbe8088c",
          4298 => x"05083082",
          4299 => x"bbe8088c",
          4300 => x"050c8153",
          4301 => x"82bbe808",
          4302 => x"8c050852",
          4303 => x"82bbe808",
          4304 => x"88050851",
          4305 => x"81a23f82",
          4306 => x"bbdc0870",
          4307 => x"82bbe808",
          4308 => x"f8050c54",
          4309 => x"82bbe808",
          4310 => x"fc050880",
          4311 => x"2e903882",
          4312 => x"bbe808f8",
          4313 => x"05083082",
          4314 => x"bbe808f8",
          4315 => x"050c82bb",
          4316 => x"e808f805",
          4317 => x"087082bb",
          4318 => x"dc0c5487",
          4319 => x"3d0d82bb",
          4320 => x"e80c0482",
          4321 => x"bbe80802",
          4322 => x"82bbe80c",
          4323 => x"fd3d0d80",
          4324 => x"5382bbe8",
          4325 => x"088c0508",
          4326 => x"5282bbe8",
          4327 => x"08880508",
          4328 => x"5180c53f",
          4329 => x"82bbdc08",
          4330 => x"7082bbdc",
          4331 => x"0c54853d",
          4332 => x"0d82bbe8",
          4333 => x"0c0482bb",
          4334 => x"e8080282",
          4335 => x"bbe80cfd",
          4336 => x"3d0d8153",
          4337 => x"82bbe808",
          4338 => x"8c050852",
          4339 => x"82bbe808",
          4340 => x"88050851",
          4341 => x"933f82bb",
          4342 => x"dc087082",
          4343 => x"bbdc0c54",
          4344 => x"853d0d82",
          4345 => x"bbe80c04",
          4346 => x"82bbe808",
          4347 => x"0282bbe8",
          4348 => x"0cfd3d0d",
          4349 => x"810b82bb",
          4350 => x"e808fc05",
          4351 => x"0c800b82",
          4352 => x"bbe808f8",
          4353 => x"050c82bb",
          4354 => x"e8088c05",
          4355 => x"0882bbe8",
          4356 => x"08880508",
          4357 => x"27b93882",
          4358 => x"bbe808fc",
          4359 => x"0508802e",
          4360 => x"ae38800b",
          4361 => x"82bbe808",
          4362 => x"8c050824",
          4363 => x"a23882bb",
          4364 => x"e8088c05",
          4365 => x"081082bb",
          4366 => x"e8088c05",
          4367 => x"0c82bbe8",
          4368 => x"08fc0508",
          4369 => x"1082bbe8",
          4370 => x"08fc050c",
          4371 => x"ffb83982",
          4372 => x"bbe808fc",
          4373 => x"0508802e",
          4374 => x"80e13882",
          4375 => x"bbe8088c",
          4376 => x"050882bb",
          4377 => x"e8088805",
          4378 => x"0826ad38",
          4379 => x"82bbe808",
          4380 => x"88050882",
          4381 => x"bbe8088c",
          4382 => x"05083182",
          4383 => x"bbe80888",
          4384 => x"050c82bb",
          4385 => x"e808f805",
          4386 => x"0882bbe8",
          4387 => x"08fc0508",
          4388 => x"0782bbe8",
          4389 => x"08f8050c",
          4390 => x"82bbe808",
          4391 => x"fc050881",
          4392 => x"2a82bbe8",
          4393 => x"08fc050c",
          4394 => x"82bbe808",
          4395 => x"8c050881",
          4396 => x"2a82bbe8",
          4397 => x"088c050c",
          4398 => x"ff953982",
          4399 => x"bbe80890",
          4400 => x"0508802e",
          4401 => x"933882bb",
          4402 => x"e8088805",
          4403 => x"087082bb",
          4404 => x"e808f405",
          4405 => x"0c519139",
          4406 => x"82bbe808",
          4407 => x"f8050870",
          4408 => x"82bbe808",
          4409 => x"f4050c51",
          4410 => x"82bbe808",
          4411 => x"f4050882",
          4412 => x"bbdc0c85",
          4413 => x"3d0d82bb",
          4414 => x"e80c0482",
          4415 => x"bbe80802",
          4416 => x"82bbe80c",
          4417 => x"f73d0d80",
          4418 => x"0b82bbe8",
          4419 => x"08f00534",
          4420 => x"82bbe808",
          4421 => x"8c050853",
          4422 => x"80730c82",
          4423 => x"bbe80888",
          4424 => x"05087008",
          4425 => x"51537233",
          4426 => x"537282bb",
          4427 => x"e808f805",
          4428 => x"347281ff",
          4429 => x"065372a0",
          4430 => x"2e098106",
          4431 => x"913882bb",
          4432 => x"e8088805",
          4433 => x"08700881",
          4434 => x"05710c53",
          4435 => x"ce3982bb",
          4436 => x"e808f805",
          4437 => x"335372ad",
          4438 => x"2e098106",
          4439 => x"a438810b",
          4440 => x"82bbe808",
          4441 => x"f0053482",
          4442 => x"bbe80888",
          4443 => x"05087008",
          4444 => x"8105710c",
          4445 => x"70085153",
          4446 => x"723382bb",
          4447 => x"e808f805",
          4448 => x"3482bbe8",
          4449 => x"08f80533",
          4450 => x"5372b02e",
          4451 => x"09810681",
          4452 => x"dc3882bb",
          4453 => x"e8088805",
          4454 => x"08700881",
          4455 => x"05710c70",
          4456 => x"08515372",
          4457 => x"3382bbe8",
          4458 => x"08f80534",
          4459 => x"82bbe808",
          4460 => x"f8053382",
          4461 => x"bbe808e8",
          4462 => x"050c82bb",
          4463 => x"e808e805",
          4464 => x"0880e22e",
          4465 => x"b63882bb",
          4466 => x"e808e805",
          4467 => x"0880f82e",
          4468 => x"843880cd",
          4469 => x"39900b82",
          4470 => x"bbe808f4",
          4471 => x"053482bb",
          4472 => x"e8088805",
          4473 => x"08700881",
          4474 => x"05710c70",
          4475 => x"08515372",
          4476 => x"3382bbe8",
          4477 => x"08f80534",
          4478 => x"81a43982",
          4479 => x"0b82bbe8",
          4480 => x"08f40534",
          4481 => x"82bbe808",
          4482 => x"88050870",
          4483 => x"08810571",
          4484 => x"0c700851",
          4485 => x"53723382",
          4486 => x"bbe808f8",
          4487 => x"053480fe",
          4488 => x"3982bbe8",
          4489 => x"08f80533",
          4490 => x"5372a026",
          4491 => x"8d38810b",
          4492 => x"82bbe808",
          4493 => x"ec050c83",
          4494 => x"803982bb",
          4495 => x"e808f805",
          4496 => x"3353af73",
          4497 => x"27903882",
          4498 => x"bbe808f8",
          4499 => x"05335372",
          4500 => x"b9268338",
          4501 => x"8d39800b",
          4502 => x"82bbe808",
          4503 => x"ec050c82",
          4504 => x"d839880b",
          4505 => x"82bbe808",
          4506 => x"f40534b2",
          4507 => x"3982bbe8",
          4508 => x"08f80533",
          4509 => x"53af7327",
          4510 => x"903882bb",
          4511 => x"e808f805",
          4512 => x"335372b9",
          4513 => x"2683388d",
          4514 => x"39800b82",
          4515 => x"bbe808ec",
          4516 => x"050c82a5",
          4517 => x"398a0b82",
          4518 => x"bbe808f4",
          4519 => x"0534800b",
          4520 => x"82bbe808",
          4521 => x"fc050c82",
          4522 => x"bbe808f8",
          4523 => x"053353a0",
          4524 => x"732781cf",
          4525 => x"3882bbe8",
          4526 => x"08f80533",
          4527 => x"5380e073",
          4528 => x"27943882",
          4529 => x"bbe808f8",
          4530 => x"0533e011",
          4531 => x"51537282",
          4532 => x"bbe808f8",
          4533 => x"053482bb",
          4534 => x"e808f805",
          4535 => x"33d01151",
          4536 => x"537282bb",
          4537 => x"e808f805",
          4538 => x"3482bbe8",
          4539 => x"08f80533",
          4540 => x"53907327",
          4541 => x"ad3882bb",
          4542 => x"e808f805",
          4543 => x"33f91151",
          4544 => x"537282bb",
          4545 => x"e808f805",
          4546 => x"3482bbe8",
          4547 => x"08f80533",
          4548 => x"53728926",
          4549 => x"8d38800b",
          4550 => x"82bbe808",
          4551 => x"ec050c81",
          4552 => x"983982bb",
          4553 => x"e808f805",
          4554 => x"3382bbe8",
          4555 => x"08f40533",
          4556 => x"54547274",
          4557 => x"268d3880",
          4558 => x"0b82bbe8",
          4559 => x"08ec050c",
          4560 => x"80f73982",
          4561 => x"bbe808f4",
          4562 => x"05337082",
          4563 => x"bbe808fc",
          4564 => x"05082982",
          4565 => x"bbe808f8",
          4566 => x"05337012",
          4567 => x"82bbe808",
          4568 => x"fc050c82",
          4569 => x"bbe80888",
          4570 => x"05087008",
          4571 => x"8105710c",
          4572 => x"70085151",
          4573 => x"52555372",
          4574 => x"3382bbe8",
          4575 => x"08f80534",
          4576 => x"fea53982",
          4577 => x"bbe808f0",
          4578 => x"05335372",
          4579 => x"802e9038",
          4580 => x"82bbe808",
          4581 => x"fc050830",
          4582 => x"82bbe808",
          4583 => x"fc050c82",
          4584 => x"bbe8088c",
          4585 => x"050882bb",
          4586 => x"e808fc05",
          4587 => x"08710c53",
          4588 => x"810b82bb",
          4589 => x"e808ec05",
          4590 => x"0c82bbe8",
          4591 => x"08ec0508",
          4592 => x"82bbdc0c",
          4593 => x"8b3d0d82",
          4594 => x"bbe80c04",
          4595 => x"82bbe808",
          4596 => x"0282bbe8",
          4597 => x"0cf73d0d",
          4598 => x"800b82bb",
          4599 => x"e808f005",
          4600 => x"3482bbe8",
          4601 => x"088c0508",
          4602 => x"5380730c",
          4603 => x"82bbe808",
          4604 => x"88050870",
          4605 => x"08515372",
          4606 => x"33537282",
          4607 => x"bbe808f8",
          4608 => x"05347281",
          4609 => x"ff065372",
          4610 => x"a02e0981",
          4611 => x"06913882",
          4612 => x"bbe80888",
          4613 => x"05087008",
          4614 => x"8105710c",
          4615 => x"53ce3982",
          4616 => x"bbe808f8",
          4617 => x"05335372",
          4618 => x"ad2e0981",
          4619 => x"06a43881",
          4620 => x"0b82bbe8",
          4621 => x"08f00534",
          4622 => x"82bbe808",
          4623 => x"88050870",
          4624 => x"08810571",
          4625 => x"0c700851",
          4626 => x"53723382",
          4627 => x"bbe808f8",
          4628 => x"053482bb",
          4629 => x"e808f805",
          4630 => x"335372b0",
          4631 => x"2e098106",
          4632 => x"81dc3882",
          4633 => x"bbe80888",
          4634 => x"05087008",
          4635 => x"8105710c",
          4636 => x"70085153",
          4637 => x"723382bb",
          4638 => x"e808f805",
          4639 => x"3482bbe8",
          4640 => x"08f80533",
          4641 => x"82bbe808",
          4642 => x"e8050c82",
          4643 => x"bbe808e8",
          4644 => x"050880e2",
          4645 => x"2eb63882",
          4646 => x"bbe808e8",
          4647 => x"050880f8",
          4648 => x"2e843880",
          4649 => x"cd39900b",
          4650 => x"82bbe808",
          4651 => x"f4053482",
          4652 => x"bbe80888",
          4653 => x"05087008",
          4654 => x"8105710c",
          4655 => x"70085153",
          4656 => x"723382bb",
          4657 => x"e808f805",
          4658 => x"3481a439",
          4659 => x"820b82bb",
          4660 => x"e808f405",
          4661 => x"3482bbe8",
          4662 => x"08880508",
          4663 => x"70088105",
          4664 => x"710c7008",
          4665 => x"51537233",
          4666 => x"82bbe808",
          4667 => x"f8053480",
          4668 => x"fe3982bb",
          4669 => x"e808f805",
          4670 => x"335372a0",
          4671 => x"268d3881",
          4672 => x"0b82bbe8",
          4673 => x"08ec050c",
          4674 => x"83803982",
          4675 => x"bbe808f8",
          4676 => x"053353af",
          4677 => x"73279038",
          4678 => x"82bbe808",
          4679 => x"f8053353",
          4680 => x"72b92683",
          4681 => x"388d3980",
          4682 => x"0b82bbe8",
          4683 => x"08ec050c",
          4684 => x"82d83988",
          4685 => x"0b82bbe8",
          4686 => x"08f40534",
          4687 => x"b23982bb",
          4688 => x"e808f805",
          4689 => x"3353af73",
          4690 => x"27903882",
          4691 => x"bbe808f8",
          4692 => x"05335372",
          4693 => x"b9268338",
          4694 => x"8d39800b",
          4695 => x"82bbe808",
          4696 => x"ec050c82",
          4697 => x"a5398a0b",
          4698 => x"82bbe808",
          4699 => x"f4053480",
          4700 => x"0b82bbe8",
          4701 => x"08fc050c",
          4702 => x"82bbe808",
          4703 => x"f8053353",
          4704 => x"a0732781",
          4705 => x"cf3882bb",
          4706 => x"e808f805",
          4707 => x"335380e0",
          4708 => x"73279438",
          4709 => x"82bbe808",
          4710 => x"f80533e0",
          4711 => x"11515372",
          4712 => x"82bbe808",
          4713 => x"f8053482",
          4714 => x"bbe808f8",
          4715 => x"0533d011",
          4716 => x"51537282",
          4717 => x"bbe808f8",
          4718 => x"053482bb",
          4719 => x"e808f805",
          4720 => x"33539073",
          4721 => x"27ad3882",
          4722 => x"bbe808f8",
          4723 => x"0533f911",
          4724 => x"51537282",
          4725 => x"bbe808f8",
          4726 => x"053482bb",
          4727 => x"e808f805",
          4728 => x"33537289",
          4729 => x"268d3880",
          4730 => x"0b82bbe8",
          4731 => x"08ec050c",
          4732 => x"81983982",
          4733 => x"bbe808f8",
          4734 => x"053382bb",
          4735 => x"e808f405",
          4736 => x"33545472",
          4737 => x"74268d38",
          4738 => x"800b82bb",
          4739 => x"e808ec05",
          4740 => x"0c80f739",
          4741 => x"82bbe808",
          4742 => x"f4053370",
          4743 => x"82bbe808",
          4744 => x"fc050829",
          4745 => x"82bbe808",
          4746 => x"f8053370",
          4747 => x"1282bbe8",
          4748 => x"08fc050c",
          4749 => x"82bbe808",
          4750 => x"88050870",
          4751 => x"08810571",
          4752 => x"0c700851",
          4753 => x"51525553",
          4754 => x"723382bb",
          4755 => x"e808f805",
          4756 => x"34fea539",
          4757 => x"82bbe808",
          4758 => x"f0053353",
          4759 => x"72802e90",
          4760 => x"3882bbe8",
          4761 => x"08fc0508",
          4762 => x"3082bbe8",
          4763 => x"08fc050c",
          4764 => x"82bbe808",
          4765 => x"8c050882",
          4766 => x"bbe808fc",
          4767 => x"0508710c",
          4768 => x"53810b82",
          4769 => x"bbe808ec",
          4770 => x"050c82bb",
          4771 => x"e808ec05",
          4772 => x"0882bbdc",
          4773 => x"0c8b3d0d",
          4774 => x"82bbe80c",
          4775 => x"04f93d0d",
          4776 => x"79700870",
          4777 => x"56565874",
          4778 => x"802e80e3",
          4779 => x"38953975",
          4780 => x"0851e6d1",
          4781 => x"3f82bbdc",
          4782 => x"0815780c",
          4783 => x"85163354",
          4784 => x"80cd3974",
          4785 => x"335473a0",
          4786 => x"2e098106",
          4787 => x"86388115",
          4788 => x"55f13980",
          4789 => x"57769029",
          4790 => x"82b6dc05",
          4791 => x"70085256",
          4792 => x"e6a33f82",
          4793 => x"bbdc0853",
          4794 => x"74527508",
          4795 => x"51e9a33f",
          4796 => x"82bbdc08",
          4797 => x"8b388416",
          4798 => x"33547381",
          4799 => x"2effb038",
          4800 => x"81177081",
          4801 => x"ff065854",
          4802 => x"997727c9",
          4803 => x"38ff5473",
          4804 => x"82bbdc0c",
          4805 => x"893d0d04",
          4806 => x"ff3d0d73",
          4807 => x"52719326",
          4808 => x"818e3871",
          4809 => x"8429829a",
          4810 => x"9c055271",
          4811 => x"0804829f",
          4812 => x"e8518180",
          4813 => x"39829ff4",
          4814 => x"5180f939",
          4815 => x"82a08451",
          4816 => x"80f23982",
          4817 => x"a0945180",
          4818 => x"eb3982a0",
          4819 => x"a45180e4",
          4820 => x"3982a0b4",
          4821 => x"5180dd39",
          4822 => x"82a0c851",
          4823 => x"80d63982",
          4824 => x"a0d85180",
          4825 => x"cf3982a0",
          4826 => x"f05180c8",
          4827 => x"3982a188",
          4828 => x"5180c139",
          4829 => x"82a1a051",
          4830 => x"bb3982a1",
          4831 => x"bc51b539",
          4832 => x"82a1d051",
          4833 => x"af3982a1",
          4834 => x"f851a939",
          4835 => x"82a28851",
          4836 => x"a33982a2",
          4837 => x"a8519d39",
          4838 => x"82a2b851",
          4839 => x"973982a2",
          4840 => x"d0519139",
          4841 => x"82a2e851",
          4842 => x"8b3982a3",
          4843 => x"80518539",
          4844 => x"82a38c51",
          4845 => x"d8ad3f83",
          4846 => x"3d0d04fb",
          4847 => x"3d0d7779",
          4848 => x"56567487",
          4849 => x"e7268a38",
          4850 => x"74527587",
          4851 => x"e8295190",
          4852 => x"3987e852",
          4853 => x"7451efab",
          4854 => x"3f82bbdc",
          4855 => x"08527551",
          4856 => x"efa13f82",
          4857 => x"bbdc0854",
          4858 => x"79537552",
          4859 => x"82a39c51",
          4860 => x"ffbbe53f",
          4861 => x"873d0d04",
          4862 => x"ec3d0d66",
          4863 => x"02840580",
          4864 => x"e305335b",
          4865 => x"57806878",
          4866 => x"30707a07",
          4867 => x"73255157",
          4868 => x"59597856",
          4869 => x"7787ff26",
          4870 => x"83388156",
          4871 => x"74760770",
          4872 => x"81ff0651",
          4873 => x"55935674",
          4874 => x"81823881",
          4875 => x"5376528c",
          4876 => x"3d705256",
          4877 => x"8184b93f",
          4878 => x"82bbdc08",
          4879 => x"5782bbdc",
          4880 => x"08b93882",
          4881 => x"bbdc0887",
          4882 => x"c098880c",
          4883 => x"82bbdc08",
          4884 => x"59963dd4",
          4885 => x"05548480",
          4886 => x"53775275",
          4887 => x"518188f5",
          4888 => x"3f82bbdc",
          4889 => x"085782bb",
          4890 => x"dc089038",
          4891 => x"7a557480",
          4892 => x"2e893874",
          4893 => x"19751959",
          4894 => x"59d73996",
          4895 => x"3dd80551",
          4896 => x"8190de3f",
          4897 => x"76307078",
          4898 => x"0780257b",
          4899 => x"30709f2a",
          4900 => x"72065157",
          4901 => x"51567480",
          4902 => x"2e903882",
          4903 => x"a3c05387",
          4904 => x"c0988808",
          4905 => x"527851fe",
          4906 => x"923f7656",
          4907 => x"7582bbdc",
          4908 => x"0c963d0d",
          4909 => x"04f83d0d",
          4910 => x"7c028405",
          4911 => x"b7053358",
          4912 => x"59ff5880",
          4913 => x"537b527a",
          4914 => x"51fead3f",
          4915 => x"82bbdc08",
          4916 => x"a8387680",
          4917 => x"2e883876",
          4918 => x"812e9c38",
          4919 => x"9c3982d3",
          4920 => x"ac566155",
          4921 => x"605482bb",
          4922 => x"dc537f52",
          4923 => x"7e51782d",
          4924 => x"82bbdc08",
          4925 => x"58833978",
          4926 => x"047782bb",
          4927 => x"dc0c8a3d",
          4928 => x"0d04f33d",
          4929 => x"0d7f6163",
          4930 => x"028c0580",
          4931 => x"cf053373",
          4932 => x"73156841",
          4933 => x"5f5c5c5e",
          4934 => x"5e5e7a52",
          4935 => x"82a3c851",
          4936 => x"ffb9b53f",
          4937 => x"82a3d051",
          4938 => x"ffb9ad3f",
          4939 => x"80557479",
          4940 => x"27818038",
          4941 => x"7b902e89",
          4942 => x"387ba02e",
          4943 => x"a73880c6",
          4944 => x"39741853",
          4945 => x"727a278e",
          4946 => x"38722252",
          4947 => x"82a3d451",
          4948 => x"ffb9853f",
          4949 => x"893982a3",
          4950 => x"e051ffb8",
          4951 => x"fb3f8215",
          4952 => x"5580c339",
          4953 => x"74185372",
          4954 => x"7a278e38",
          4955 => x"72085282",
          4956 => x"a3c851ff",
          4957 => x"b8e23f89",
          4958 => x"3982a3dc",
          4959 => x"51ffb8d8",
          4960 => x"3f841555",
          4961 => x"a1397418",
          4962 => x"53727a27",
          4963 => x"8e387233",
          4964 => x"5282a3e8",
          4965 => x"51ffb8c0",
          4966 => x"3f893982",
          4967 => x"a3f051ff",
          4968 => x"b8b63f81",
          4969 => x"155582d3",
          4970 => x"b00852a0",
          4971 => x"51d8833f",
          4972 => x"fefc3982",
          4973 => x"a3f451ff",
          4974 => x"b89e3f80",
          4975 => x"55747927",
          4976 => x"80c63874",
          4977 => x"18703355",
          4978 => x"53805672",
          4979 => x"7a278338",
          4980 => x"81568053",
          4981 => x"9f742783",
          4982 => x"38815375",
          4983 => x"73067081",
          4984 => x"ff065153",
          4985 => x"72802e90",
          4986 => x"387380fe",
          4987 => x"268a3882",
          4988 => x"d3b00852",
          4989 => x"73518839",
          4990 => x"82d3b008",
          4991 => x"52a051d7",
          4992 => x"b13f8115",
          4993 => x"55ffb639",
          4994 => x"82a3f851",
          4995 => x"d3d53f78",
          4996 => x"18791c5c",
          4997 => x"58a0fe3f",
          4998 => x"82bbdc08",
          4999 => x"982b7098",
          5000 => x"2c515776",
          5001 => x"a02e0981",
          5002 => x"06aa38a0",
          5003 => x"e83f82bb",
          5004 => x"dc08982b",
          5005 => x"70982c70",
          5006 => x"a0327030",
          5007 => x"729b3270",
          5008 => x"30707207",
          5009 => x"73750706",
          5010 => x"51585859",
          5011 => x"57515780",
          5012 => x"7324d838",
          5013 => x"769b2e09",
          5014 => x"81068538",
          5015 => x"80538c39",
          5016 => x"7c1e5372",
          5017 => x"7826fdb2",
          5018 => x"38ff5372",
          5019 => x"82bbdc0c",
          5020 => x"8f3d0d04",
          5021 => x"fc3d0d02",
          5022 => x"9b053382",
          5023 => x"a3fc5382",
          5024 => x"a4845255",
          5025 => x"ffb6d13f",
          5026 => x"82bab422",
          5027 => x"51a9d93f",
          5028 => x"82a49054",
          5029 => x"82a49c53",
          5030 => x"82bab533",
          5031 => x"5282a4a4",
          5032 => x"51ffb6b4",
          5033 => x"3f74802e",
          5034 => x"8438a58b",
          5035 => x"3f863d0d",
          5036 => x"04fe3d0d",
          5037 => x"87c09680",
          5038 => x"0853aab6",
          5039 => x"3f81519c",
          5040 => x"c13f82a4",
          5041 => x"c0519dd6",
          5042 => x"3f80519c",
          5043 => x"b53f7281",
          5044 => x"2a708106",
          5045 => x"51527180",
          5046 => x"2e923881",
          5047 => x"519ca33f",
          5048 => x"82a4d851",
          5049 => x"9db83f80",
          5050 => x"519c973f",
          5051 => x"72822a70",
          5052 => x"81065152",
          5053 => x"71802e92",
          5054 => x"3881519c",
          5055 => x"853f82a4",
          5056 => x"e8519d9a",
          5057 => x"3f80519b",
          5058 => x"f93f7283",
          5059 => x"2a708106",
          5060 => x"51527180",
          5061 => x"2e923881",
          5062 => x"519be73f",
          5063 => x"82a4f851",
          5064 => x"9cfc3f80",
          5065 => x"519bdb3f",
          5066 => x"72842a70",
          5067 => x"81065152",
          5068 => x"71802e92",
          5069 => x"3881519b",
          5070 => x"c93f82a5",
          5071 => x"8c519cde",
          5072 => x"3f80519b",
          5073 => x"bd3f7285",
          5074 => x"2a708106",
          5075 => x"51527180",
          5076 => x"2e923881",
          5077 => x"519bab3f",
          5078 => x"82a5a051",
          5079 => x"9cc03f80",
          5080 => x"519b9f3f",
          5081 => x"72862a70",
          5082 => x"81065152",
          5083 => x"71802e92",
          5084 => x"3881519b",
          5085 => x"8d3f82a5",
          5086 => x"b4519ca2",
          5087 => x"3f80519b",
          5088 => x"813f7287",
          5089 => x"2a708106",
          5090 => x"51527180",
          5091 => x"2e923881",
          5092 => x"519aef3f",
          5093 => x"82a5c851",
          5094 => x"9c843f80",
          5095 => x"519ae33f",
          5096 => x"72882a70",
          5097 => x"81065152",
          5098 => x"71802e92",
          5099 => x"3881519a",
          5100 => x"d13f82a5",
          5101 => x"dc519be6",
          5102 => x"3f80519a",
          5103 => x"c53fa8ba",
          5104 => x"3f843d0d",
          5105 => x"04fb3d0d",
          5106 => x"77028405",
          5107 => x"a3053370",
          5108 => x"55565680",
          5109 => x"527551e3",
          5110 => x"8d3f0b0b",
          5111 => x"82b6d833",
          5112 => x"5473a938",
          5113 => x"815382a6",
          5114 => x"985282d2",
          5115 => x"dc5180fc",
          5116 => x"ff3f82bb",
          5117 => x"dc083070",
          5118 => x"82bbdc08",
          5119 => x"07802582",
          5120 => x"71315151",
          5121 => x"54730b0b",
          5122 => x"82b6d834",
          5123 => x"0b0b82b6",
          5124 => x"d8335473",
          5125 => x"812e0981",
          5126 => x"06af3882",
          5127 => x"d2dc5374",
          5128 => x"52755181",
          5129 => x"b7b03f82",
          5130 => x"bbdc0880",
          5131 => x"2e8b3882",
          5132 => x"bbdc0851",
          5133 => x"cfad3f91",
          5134 => x"3982d2dc",
          5135 => x"518189a1",
          5136 => x"3f820b0b",
          5137 => x"0b82b6d8",
          5138 => x"340b0b82",
          5139 => x"b6d83354",
          5140 => x"73822e09",
          5141 => x"81068c38",
          5142 => x"82a6a853",
          5143 => x"74527551",
          5144 => x"aeb23f80",
          5145 => x"0b82bbdc",
          5146 => x"0c873d0d",
          5147 => x"04ce3d0d",
          5148 => x"80707182",
          5149 => x"d2d80c5f",
          5150 => x"5d81527c",
          5151 => x"5180cbcb",
          5152 => x"3f82bbdc",
          5153 => x"0881ff06",
          5154 => x"59787d2e",
          5155 => x"098106a3",
          5156 => x"38963d59",
          5157 => x"835382a6",
          5158 => x"b4527851",
          5159 => x"dcc73f7c",
          5160 => x"53785282",
          5161 => x"bd885180",
          5162 => x"fae53f82",
          5163 => x"bbdc087d",
          5164 => x"2e883882",
          5165 => x"a6b85191",
          5166 => x"d5398170",
          5167 => x"5f5d82a6",
          5168 => x"f051ffb2",
          5169 => x"933f963d",
          5170 => x"70465a80",
          5171 => x"f8527951",
          5172 => x"fdf33fb4",
          5173 => x"3dff8405",
          5174 => x"51f3c23f",
          5175 => x"82bbdc08",
          5176 => x"902b7090",
          5177 => x"2c515978",
          5178 => x"80c12e89",
          5179 => x"d4387880",
          5180 => x"c12480d9",
          5181 => x"3878ab2e",
          5182 => x"83b93878",
          5183 => x"ab24a438",
          5184 => x"78822e81",
          5185 => x"b3387882",
          5186 => x"248a3878",
          5187 => x"802effae",
          5188 => x"388f8039",
          5189 => x"78842e82",
          5190 => x"83387894",
          5191 => x"2e82ad38",
          5192 => x"8ef13978",
          5193 => x"bd2e84fc",
          5194 => x"3878bd24",
          5195 => x"903878b0",
          5196 => x"2e83a638",
          5197 => x"78bc2e84",
          5198 => x"84388ed7",
          5199 => x"3978bf2e",
          5200 => x"85c43878",
          5201 => x"80c02e86",
          5202 => x"bd388ec7",
          5203 => x"397880d5",
          5204 => x"2e8da038",
          5205 => x"7880d524",
          5206 => x"b0387880",
          5207 => x"d02e8cd9",
          5208 => x"387880d0",
          5209 => x"24923878",
          5210 => x"80c22e89",
          5211 => x"fc387880",
          5212 => x"c32e8ba5",
          5213 => x"388e9c39",
          5214 => x"7880d12e",
          5215 => x"8cca3878",
          5216 => x"80d42e8c",
          5217 => x"d2388e8b",
          5218 => x"39788182",
          5219 => x"2e8de238",
          5220 => x"78818224",
          5221 => x"92387880",
          5222 => x"f82e8cf4",
          5223 => x"387880f9",
          5224 => x"2e8d9138",
          5225 => x"8ded3978",
          5226 => x"81832e8d",
          5227 => x"d3387881",
          5228 => x"852e8dd9",
          5229 => x"388ddc39",
          5230 => x"b43dff80",
          5231 => x"1153ff84",
          5232 => x"0551ec88",
          5233 => x"3f82bbdc",
          5234 => x"08883882",
          5235 => x"a6f4518f",
          5236 => x"bd39b43d",
          5237 => x"fefc1153",
          5238 => x"ff840551",
          5239 => x"ebee3f82",
          5240 => x"bbdc0880",
          5241 => x"2e883881",
          5242 => x"63258338",
          5243 => x"80430280",
          5244 => x"cb053352",
          5245 => x"0280cf05",
          5246 => x"335180c8",
          5247 => x"ce3f82bb",
          5248 => x"dc0881ff",
          5249 => x"0659788d",
          5250 => x"3882a784",
          5251 => x"51cbd43f",
          5252 => x"815efdaa",
          5253 => x"3982a794",
          5254 => x"518ef339",
          5255 => x"b43dff80",
          5256 => x"1153ff84",
          5257 => x"0551eba4",
          5258 => x"3f82bbdc",
          5259 => x"08802efd",
          5260 => x"8d388053",
          5261 => x"80520280",
          5262 => x"cf053351",
          5263 => x"80ccd93f",
          5264 => x"82bbdc08",
          5265 => x"5282a7ac",
          5266 => x"518c9f39",
          5267 => x"b43dff80",
          5268 => x"1153ff84",
          5269 => x"0551eaf4",
          5270 => x"3f82bbdc",
          5271 => x"08802e87",
          5272 => x"38638926",
          5273 => x"fcd838b4",
          5274 => x"3dfefc11",
          5275 => x"53ff8405",
          5276 => x"51ead93f",
          5277 => x"82bbdc08",
          5278 => x"863882bb",
          5279 => x"dc084363",
          5280 => x"5382a7b4",
          5281 => x"527951ff",
          5282 => x"b1b63f02",
          5283 => x"80cb0533",
          5284 => x"53795263",
          5285 => x"84b42982",
          5286 => x"bd880551",
          5287 => x"80f6f03f",
          5288 => x"82bbdc08",
          5289 => x"818c3882",
          5290 => x"a78451ca",
          5291 => x"b63f815d",
          5292 => x"fc8c39b4",
          5293 => x"3dff8405",
          5294 => x"518fc03f",
          5295 => x"82bbdc08",
          5296 => x"b53dff84",
          5297 => x"05525b90",
          5298 => x"d63f8153",
          5299 => x"82bbdc08",
          5300 => x"527a51f2",
          5301 => x"a33f80d1",
          5302 => x"39b43dff",
          5303 => x"8405518f",
          5304 => x"9a3f82bb",
          5305 => x"dc08b53d",
          5306 => x"ff840552",
          5307 => x"5b90b03f",
          5308 => x"82bbdc08",
          5309 => x"b53dff84",
          5310 => x"05525a90",
          5311 => x"a23f82bb",
          5312 => x"dc08b53d",
          5313 => x"ff840552",
          5314 => x"5990943f",
          5315 => x"82ba8058",
          5316 => x"82bc8c57",
          5317 => x"80568055",
          5318 => x"82bbdc08",
          5319 => x"81ff0654",
          5320 => x"78537952",
          5321 => x"7a51f38d",
          5322 => x"3f82bbdc",
          5323 => x"08802efb",
          5324 => x"8d3882bb",
          5325 => x"dc0851ef",
          5326 => x"df3ffb82",
          5327 => x"39b43dff",
          5328 => x"801153ff",
          5329 => x"840551e9",
          5330 => x"833f82bb",
          5331 => x"dc08802e",
          5332 => x"faec38b4",
          5333 => x"3dfefc11",
          5334 => x"53ff8405",
          5335 => x"51e8ed3f",
          5336 => x"82bbdc08",
          5337 => x"802efad6",
          5338 => x"38b43dfe",
          5339 => x"f81153ff",
          5340 => x"840551e8",
          5341 => x"d73f82bb",
          5342 => x"dc088638",
          5343 => x"82bbdc08",
          5344 => x"4282a7b8",
          5345 => x"51ffacd0",
          5346 => x"3f63635c",
          5347 => x"5a797b27",
          5348 => x"81ec3861",
          5349 => x"59787a70",
          5350 => x"84055c0c",
          5351 => x"7a7a26f5",
          5352 => x"3881db39",
          5353 => x"b43dff80",
          5354 => x"1153ff84",
          5355 => x"0551e89c",
          5356 => x"3f82bbdc",
          5357 => x"08802efa",
          5358 => x"8538b43d",
          5359 => x"fefc1153",
          5360 => x"ff840551",
          5361 => x"e8863f82",
          5362 => x"bbdc0880",
          5363 => x"2ef9ef38",
          5364 => x"b43dfef8",
          5365 => x"1153ff84",
          5366 => x"0551e7f0",
          5367 => x"3f82bbdc",
          5368 => x"08802ef9",
          5369 => x"d93882a7",
          5370 => x"c851ffab",
          5371 => x"eb3f635a",
          5372 => x"79632781",
          5373 => x"89386159",
          5374 => x"79708105",
          5375 => x"5b337934",
          5376 => x"61810542",
          5377 => x"eb39b43d",
          5378 => x"ff801153",
          5379 => x"ff840551",
          5380 => x"e7ba3f82",
          5381 => x"bbdc0880",
          5382 => x"2ef9a338",
          5383 => x"b43dfefc",
          5384 => x"1153ff84",
          5385 => x"0551e7a4",
          5386 => x"3f82bbdc",
          5387 => x"08802ef9",
          5388 => x"8d38b43d",
          5389 => x"fef81153",
          5390 => x"ff840551",
          5391 => x"e78e3f82",
          5392 => x"bbdc0880",
          5393 => x"2ef8f738",
          5394 => x"82a7d451",
          5395 => x"ffab893f",
          5396 => x"635a7963",
          5397 => x"27a83861",
          5398 => x"70337b33",
          5399 => x"5e5a5b78",
          5400 => x"7c2e9238",
          5401 => x"78557a54",
          5402 => x"79335379",
          5403 => x"5282a7e4",
          5404 => x"51ffaae4",
          5405 => x"3f811a62",
          5406 => x"8105435a",
          5407 => x"d5398a51",
          5408 => x"ca833ff8",
          5409 => x"b939b43d",
          5410 => x"ff801153",
          5411 => x"ff840551",
          5412 => x"e6ba3f82",
          5413 => x"bbdc0880",
          5414 => x"df3882ba",
          5415 => x"c8335978",
          5416 => x"802e8938",
          5417 => x"82ba8008",
          5418 => x"4480cd39",
          5419 => x"82bac933",
          5420 => x"5978802e",
          5421 => x"883882ba",
          5422 => x"880844bc",
          5423 => x"3982baca",
          5424 => x"33597880",
          5425 => x"2e883882",
          5426 => x"ba900844",
          5427 => x"ab3982ba",
          5428 => x"cb335978",
          5429 => x"802e8838",
          5430 => x"82ba9808",
          5431 => x"449a3982",
          5432 => x"bac63359",
          5433 => x"78802e88",
          5434 => x"3882baa0",
          5435 => x"08448939",
          5436 => x"82bab008",
          5437 => x"fc800544",
          5438 => x"b43dfefc",
          5439 => x"1153ff84",
          5440 => x"0551e5c8",
          5441 => x"3f82bbdc",
          5442 => x"0880de38",
          5443 => x"82bac833",
          5444 => x"5978802e",
          5445 => x"893882ba",
          5446 => x"84084380",
          5447 => x"cc3982ba",
          5448 => x"c9335978",
          5449 => x"802e8838",
          5450 => x"82ba8c08",
          5451 => x"43bb3982",
          5452 => x"baca3359",
          5453 => x"78802e88",
          5454 => x"3882ba94",
          5455 => x"0843aa39",
          5456 => x"82bacb33",
          5457 => x"5978802e",
          5458 => x"883882ba",
          5459 => x"9c084399",
          5460 => x"3982bac6",
          5461 => x"33597880",
          5462 => x"2e883882",
          5463 => x"baa40843",
          5464 => x"883982ba",
          5465 => x"b0088805",
          5466 => x"43b43dfe",
          5467 => x"f81153ff",
          5468 => x"840551e4",
          5469 => x"d73f82bb",
          5470 => x"dc08802e",
          5471 => x"a7388062",
          5472 => x"5c5c7a88",
          5473 => x"2e833881",
          5474 => x"5c7a9032",
          5475 => x"70307072",
          5476 => x"079f2a70",
          5477 => x"7f065151",
          5478 => x"5a5a7880",
          5479 => x"2e88387a",
          5480 => x"a02e8338",
          5481 => x"884282a8",
          5482 => x"8051c4b7",
          5483 => x"3fa05563",
          5484 => x"54615362",
          5485 => x"526351ee",
          5486 => x"c93f82a8",
          5487 => x"8c5187ce",
          5488 => x"39b43dff",
          5489 => x"801153ff",
          5490 => x"840551e3",
          5491 => x"ff3f82bb",
          5492 => x"dc08802e",
          5493 => x"f5e838b4",
          5494 => x"3dfefc11",
          5495 => x"53ff8405",
          5496 => x"51e3e93f",
          5497 => x"82bbdc08",
          5498 => x"802ea438",
          5499 => x"63590280",
          5500 => x"cb053379",
          5501 => x"34638105",
          5502 => x"44b43dfe",
          5503 => x"fc1153ff",
          5504 => x"840551e3",
          5505 => x"c73f82bb",
          5506 => x"dc08e138",
          5507 => x"f5b03963",
          5508 => x"70335452",
          5509 => x"82a89851",
          5510 => x"ffa7bd3f",
          5511 => x"82d3ac08",
          5512 => x"5380f852",
          5513 => x"7951ffa8",
          5514 => x"843f7945",
          5515 => x"79335978",
          5516 => x"ae2ef58a",
          5517 => x"389f7927",
          5518 => x"9f38b43d",
          5519 => x"fefc1153",
          5520 => x"ff840551",
          5521 => x"e3863f82",
          5522 => x"bbdc0880",
          5523 => x"2e913863",
          5524 => x"590280cb",
          5525 => x"05337934",
          5526 => x"63810544",
          5527 => x"ffb13982",
          5528 => x"a8a451c2",
          5529 => x"fe3fffa7",
          5530 => x"39b43dfe",
          5531 => x"f41153ff",
          5532 => x"840551dd",
          5533 => x"863f82bb",
          5534 => x"dc08802e",
          5535 => x"f4c038b4",
          5536 => x"3dfef011",
          5537 => x"53ff8405",
          5538 => x"51dcf03f",
          5539 => x"82bbdc08",
          5540 => x"802ea538",
          5541 => x"605902be",
          5542 => x"05227970",
          5543 => x"82055b23",
          5544 => x"7841b43d",
          5545 => x"fef01153",
          5546 => x"ff840551",
          5547 => x"dccd3f82",
          5548 => x"bbdc08e0",
          5549 => x"38f48739",
          5550 => x"60702254",
          5551 => x"5282a8a8",
          5552 => x"51ffa694",
          5553 => x"3f82d3ac",
          5554 => x"085380f8",
          5555 => x"527951ff",
          5556 => x"a6db3f79",
          5557 => x"45793359",
          5558 => x"78ae2ef3",
          5559 => x"e138789f",
          5560 => x"26873860",
          5561 => x"820541d0",
          5562 => x"39b43dfe",
          5563 => x"f01153ff",
          5564 => x"840551dc",
          5565 => x"863f82bb",
          5566 => x"dc08802e",
          5567 => x"92386059",
          5568 => x"02be0522",
          5569 => x"79708205",
          5570 => x"5b237841",
          5571 => x"ffaa3982",
          5572 => x"a8a451c1",
          5573 => x"ce3fffa0",
          5574 => x"39b43dfe",
          5575 => x"f41153ff",
          5576 => x"840551db",
          5577 => x"d63f82bb",
          5578 => x"dc08802e",
          5579 => x"f39038b4",
          5580 => x"3dfef011",
          5581 => x"53ff8405",
          5582 => x"51dbc03f",
          5583 => x"82bbdc08",
          5584 => x"802ea038",
          5585 => x"6060710c",
          5586 => x"59608405",
          5587 => x"41b43dfe",
          5588 => x"f01153ff",
          5589 => x"840551db",
          5590 => x"a23f82bb",
          5591 => x"dc08e538",
          5592 => x"f2dc3960",
          5593 => x"70085452",
          5594 => x"82a8b451",
          5595 => x"ffa4e93f",
          5596 => x"82d3ac08",
          5597 => x"5380f852",
          5598 => x"7951ffa5",
          5599 => x"b03f7945",
          5600 => x"79335978",
          5601 => x"ae2ef2b6",
          5602 => x"389f7927",
          5603 => x"9b38b43d",
          5604 => x"fef01153",
          5605 => x"ff840551",
          5606 => x"dae13f82",
          5607 => x"bbdc0880",
          5608 => x"2e8d3860",
          5609 => x"60710c59",
          5610 => x"60840541",
          5611 => x"ffb53982",
          5612 => x"a8a451c0",
          5613 => x"ae3fffab",
          5614 => x"3982a8c4",
          5615 => x"51c0a43f",
          5616 => x"82519889",
          5617 => x"3ff1f739",
          5618 => x"82a8dc51",
          5619 => x"c0953fa2",
          5620 => x"5197de3f",
          5621 => x"f1e83982",
          5622 => x"a8f051c0",
          5623 => x"863f8480",
          5624 => x"810b87c0",
          5625 => x"94840c84",
          5626 => x"80810b87",
          5627 => x"c094940c",
          5628 => x"f1cc3982",
          5629 => x"a98451ff",
          5630 => x"bfe93f8c",
          5631 => x"80830b87",
          5632 => x"c094840c",
          5633 => x"8c80830b",
          5634 => x"87c09494",
          5635 => x"0cf1af39",
          5636 => x"b43dff80",
          5637 => x"1153ff84",
          5638 => x"0551dfb0",
          5639 => x"3f82bbdc",
          5640 => x"08802ef1",
          5641 => x"99386352",
          5642 => x"82a99851",
          5643 => x"ffa3a93f",
          5644 => x"63597804",
          5645 => x"b43dff80",
          5646 => x"1153ff84",
          5647 => x"0551df8c",
          5648 => x"3f82bbdc",
          5649 => x"08802ef0",
          5650 => x"f5386352",
          5651 => x"82a9b451",
          5652 => x"ffa3853f",
          5653 => x"6359782d",
          5654 => x"82bbdc08",
          5655 => x"802ef0de",
          5656 => x"3882bbdc",
          5657 => x"085282a9",
          5658 => x"d051ffa2",
          5659 => x"eb3ff0ce",
          5660 => x"3982a9ec",
          5661 => x"51ffbeeb",
          5662 => x"3fffa2bd",
          5663 => x"3ff0bf39",
          5664 => x"82aa8851",
          5665 => x"ffbedc3f",
          5666 => x"8059ffa6",
          5667 => x"3991a83f",
          5668 => x"f0ac3979",
          5669 => x"45793359",
          5670 => x"78802ef0",
          5671 => x"a1387d7d",
          5672 => x"06597880",
          5673 => x"2e81cf38",
          5674 => x"b43dff84",
          5675 => x"055183cb",
          5676 => x"3f82bbdc",
          5677 => x"085b815c",
          5678 => x"7b822eb2",
          5679 => x"387b8224",
          5680 => x"89387b81",
          5681 => x"2e8c3880",
          5682 => x"ca397b83",
          5683 => x"2ead3880",
          5684 => x"c23982aa",
          5685 => x"9c567a55",
          5686 => x"82aaa054",
          5687 => x"805382aa",
          5688 => x"a452b43d",
          5689 => x"ffb00551",
          5690 => x"ffa4d53f",
          5691 => x"b8397a52",
          5692 => x"b43dffb0",
          5693 => x"0551cafb",
          5694 => x"3fab397a",
          5695 => x"5582aaa0",
          5696 => x"54805382",
          5697 => x"aab452b4",
          5698 => x"3dffb005",
          5699 => x"51ffa4b0",
          5700 => x"3f93397a",
          5701 => x"54805382",
          5702 => x"aac052b4",
          5703 => x"3dffb005",
          5704 => x"51ffa49c",
          5705 => x"3f82ba80",
          5706 => x"5882bc8c",
          5707 => x"57805664",
          5708 => x"55805482",
          5709 => x"d8805382",
          5710 => x"d88052b4",
          5711 => x"3dffb005",
          5712 => x"51e6f23f",
          5713 => x"82bbdc08",
          5714 => x"82bbdc08",
          5715 => x"09703070",
          5716 => x"72078025",
          5717 => x"515b5b5f",
          5718 => x"805a7b83",
          5719 => x"26833881",
          5720 => x"5a787a06",
          5721 => x"5978802e",
          5722 => x"8d38811c",
          5723 => x"7081ff06",
          5724 => x"5d597bfe",
          5725 => x"c3387d81",
          5726 => x"327d8132",
          5727 => x"0759788a",
          5728 => x"387eff2e",
          5729 => x"098106ee",
          5730 => x"b53882aa",
          5731 => x"c851ffbc",
          5732 => x"d23feeaa",
          5733 => x"39f53d0d",
          5734 => x"800b82bc",
          5735 => x"8c3487c0",
          5736 => x"948c7008",
          5737 => x"54558784",
          5738 => x"80527251",
          5739 => x"d3d53f82",
          5740 => x"bbdc0890",
          5741 => x"2b750855",
          5742 => x"53878480",
          5743 => x"527351d3",
          5744 => x"c23f7282",
          5745 => x"bbdc0807",
          5746 => x"750c87c0",
          5747 => x"949c7008",
          5748 => x"54558784",
          5749 => x"80527251",
          5750 => x"d3a93f82",
          5751 => x"bbdc0890",
          5752 => x"2b750855",
          5753 => x"53878480",
          5754 => x"527351d3",
          5755 => x"963f7282",
          5756 => x"bbdc0807",
          5757 => x"750c8c80",
          5758 => x"830b87c0",
          5759 => x"94840c8c",
          5760 => x"80830b87",
          5761 => x"c094940c",
          5762 => x"80fa9a5a",
          5763 => x"80fd865b",
          5764 => x"83028405",
          5765 => x"99053480",
          5766 => x"5c82d3ac",
          5767 => x"0b873d70",
          5768 => x"88130c70",
          5769 => x"720c82d3",
          5770 => x"b00c5489",
          5771 => x"be3f93c2",
          5772 => x"3f82aad8",
          5773 => x"51ffbbab",
          5774 => x"3f82aae4",
          5775 => x"51ffbba3",
          5776 => x"3f80ddb1",
          5777 => x"5192e53f",
          5778 => x"8151e8a8",
          5779 => x"3fec9e3f",
          5780 => x"8004fe3d",
          5781 => x"0d805283",
          5782 => x"5371882b",
          5783 => x"5287d83f",
          5784 => x"82bbdc08",
          5785 => x"81ff0672",
          5786 => x"07ff1454",
          5787 => x"52728025",
          5788 => x"e8387182",
          5789 => x"bbdc0c84",
          5790 => x"3d0d04fc",
          5791 => x"3d0d7670",
          5792 => x"08545580",
          5793 => x"73525472",
          5794 => x"742e818a",
          5795 => x"38723351",
          5796 => x"70a02e09",
          5797 => x"81068638",
          5798 => x"811353f1",
          5799 => x"39723351",
          5800 => x"70a22e09",
          5801 => x"81068638",
          5802 => x"81135381",
          5803 => x"54725273",
          5804 => x"812e0981",
          5805 => x"069f3884",
          5806 => x"39811252",
          5807 => x"80723352",
          5808 => x"5470a22e",
          5809 => x"83388154",
          5810 => x"70802e9d",
          5811 => x"3873ea38",
          5812 => x"98398112",
          5813 => x"52807233",
          5814 => x"525470a0",
          5815 => x"2e833881",
          5816 => x"5470802e",
          5817 => x"843873ea",
          5818 => x"38807233",
          5819 => x"525470a0",
          5820 => x"2e098106",
          5821 => x"83388154",
          5822 => x"70a23270",
          5823 => x"30708025",
          5824 => x"76075151",
          5825 => x"5170802e",
          5826 => x"88388072",
          5827 => x"70810554",
          5828 => x"3471750c",
          5829 => x"72517082",
          5830 => x"bbdc0c86",
          5831 => x"3d0d04fc",
          5832 => x"3d0d7653",
          5833 => x"7208802e",
          5834 => x"9138863d",
          5835 => x"fc055272",
          5836 => x"51d3c83f",
          5837 => x"82bbdc08",
          5838 => x"85388053",
          5839 => x"83397453",
          5840 => x"7282bbdc",
          5841 => x"0c863d0d",
          5842 => x"04fc3d0d",
          5843 => x"76821133",
          5844 => x"ff055253",
          5845 => x"8152708b",
          5846 => x"26819838",
          5847 => x"831333ff",
          5848 => x"05518252",
          5849 => x"709e2681",
          5850 => x"8a388413",
          5851 => x"33518352",
          5852 => x"70972680",
          5853 => x"fe388513",
          5854 => x"33518452",
          5855 => x"70bb2680",
          5856 => x"f2388613",
          5857 => x"33518552",
          5858 => x"70bb2680",
          5859 => x"e6388813",
          5860 => x"22558652",
          5861 => x"7487e726",
          5862 => x"80d9388a",
          5863 => x"13225487",
          5864 => x"527387e7",
          5865 => x"2680cc38",
          5866 => x"810b87c0",
          5867 => x"989c0c72",
          5868 => x"2287c098",
          5869 => x"bc0c8213",
          5870 => x"3387c098",
          5871 => x"b80c8313",
          5872 => x"3387c098",
          5873 => x"b40c8413",
          5874 => x"3387c098",
          5875 => x"b00c8513",
          5876 => x"3387c098",
          5877 => x"ac0c8613",
          5878 => x"3387c098",
          5879 => x"a80c7487",
          5880 => x"c098a40c",
          5881 => x"7387c098",
          5882 => x"a00c800b",
          5883 => x"87c0989c",
          5884 => x"0c805271",
          5885 => x"82bbdc0c",
          5886 => x"863d0d04",
          5887 => x"f33d0d7f",
          5888 => x"5b87c098",
          5889 => x"9c5d817d",
          5890 => x"0c87c098",
          5891 => x"bc085e7d",
          5892 => x"7b2387c0",
          5893 => x"98b8085a",
          5894 => x"79821c34",
          5895 => x"87c098b4",
          5896 => x"085a7983",
          5897 => x"1c3487c0",
          5898 => x"98b0085a",
          5899 => x"79841c34",
          5900 => x"87c098ac",
          5901 => x"085a7985",
          5902 => x"1c3487c0",
          5903 => x"98a8085a",
          5904 => x"79861c34",
          5905 => x"87c098a4",
          5906 => x"085c7b88",
          5907 => x"1c2387c0",
          5908 => x"98a0085a",
          5909 => x"798a1c23",
          5910 => x"807d0c79",
          5911 => x"83ffff06",
          5912 => x"597b83ff",
          5913 => x"ff065886",
          5914 => x"1b335785",
          5915 => x"1b335684",
          5916 => x"1b335583",
          5917 => x"1b335482",
          5918 => x"1b33537d",
          5919 => x"83ffff06",
          5920 => x"5282aafc",
          5921 => x"51ff9ad0",
          5922 => x"3f8f3d0d",
          5923 => x"04fb3d0d",
          5924 => x"029f0533",
          5925 => x"82b9fc33",
          5926 => x"7081ff06",
          5927 => x"58555587",
          5928 => x"c0948451",
          5929 => x"75802e86",
          5930 => x"3887c094",
          5931 => x"94517008",
          5932 => x"70962a70",
          5933 => x"81065354",
          5934 => x"5270802e",
          5935 => x"8c387191",
          5936 => x"2a708106",
          5937 => x"515170d7",
          5938 => x"38728132",
          5939 => x"70810651",
          5940 => x"5170802e",
          5941 => x"8d387193",
          5942 => x"2a708106",
          5943 => x"515170ff",
          5944 => x"be387381",
          5945 => x"ff065187",
          5946 => x"c0948052",
          5947 => x"70802e86",
          5948 => x"3887c094",
          5949 => x"90527472",
          5950 => x"0c7482bb",
          5951 => x"dc0c873d",
          5952 => x"0d04ff3d",
          5953 => x"0d028f05",
          5954 => x"33703070",
          5955 => x"9f2a5152",
          5956 => x"527082b9",
          5957 => x"fc34833d",
          5958 => x"0d04f93d",
          5959 => x"0d02a705",
          5960 => x"3358778a",
          5961 => x"2e098106",
          5962 => x"87387a52",
          5963 => x"8d51eb3f",
          5964 => x"82b9fc33",
          5965 => x"7081ff06",
          5966 => x"585687c0",
          5967 => x"94845376",
          5968 => x"802e8638",
          5969 => x"87c09494",
          5970 => x"53720870",
          5971 => x"962a7081",
          5972 => x"06555654",
          5973 => x"72802e8c",
          5974 => x"3873912a",
          5975 => x"70810651",
          5976 => x"5372d738",
          5977 => x"74813270",
          5978 => x"81065153",
          5979 => x"72802e8d",
          5980 => x"3873932a",
          5981 => x"70810651",
          5982 => x"5372ffbe",
          5983 => x"387581ff",
          5984 => x"065387c0",
          5985 => x"94805472",
          5986 => x"802e8638",
          5987 => x"87c09490",
          5988 => x"5477740c",
          5989 => x"800b82bb",
          5990 => x"dc0c893d",
          5991 => x"0d04f93d",
          5992 => x"0d795480",
          5993 => x"74337081",
          5994 => x"ff065353",
          5995 => x"5770772e",
          5996 => x"80fc3871",
          5997 => x"81ff0681",
          5998 => x"1582b9fc",
          5999 => x"337081ff",
          6000 => x"06595755",
          6001 => x"5887c094",
          6002 => x"84517580",
          6003 => x"2e863887",
          6004 => x"c0949451",
          6005 => x"70087096",
          6006 => x"2a708106",
          6007 => x"53545270",
          6008 => x"802e8c38",
          6009 => x"71912a70",
          6010 => x"81065151",
          6011 => x"70d73872",
          6012 => x"81327081",
          6013 => x"06515170",
          6014 => x"802e8d38",
          6015 => x"71932a70",
          6016 => x"81065151",
          6017 => x"70ffbe38",
          6018 => x"7481ff06",
          6019 => x"5187c094",
          6020 => x"80527080",
          6021 => x"2e863887",
          6022 => x"c0949052",
          6023 => x"77720c81",
          6024 => x"17743370",
          6025 => x"81ff0653",
          6026 => x"535770ff",
          6027 => x"86387682",
          6028 => x"bbdc0c89",
          6029 => x"3d0d04fe",
          6030 => x"3d0d82b9",
          6031 => x"fc337081",
          6032 => x"ff065452",
          6033 => x"87c09484",
          6034 => x"5172802e",
          6035 => x"863887c0",
          6036 => x"94945170",
          6037 => x"0870822a",
          6038 => x"70810651",
          6039 => x"51517080",
          6040 => x"2ee23871",
          6041 => x"81ff0651",
          6042 => x"87c09480",
          6043 => x"5270802e",
          6044 => x"863887c0",
          6045 => x"94905271",
          6046 => x"087081ff",
          6047 => x"0682bbdc",
          6048 => x"0c51843d",
          6049 => x"0d04ffaf",
          6050 => x"3f82bbdc",
          6051 => x"0881ff06",
          6052 => x"82bbdc0c",
          6053 => x"04fe3d0d",
          6054 => x"82b9fc33",
          6055 => x"7081ff06",
          6056 => x"525387c0",
          6057 => x"94845270",
          6058 => x"802e8638",
          6059 => x"87c09494",
          6060 => x"52710870",
          6061 => x"822a7081",
          6062 => x"06515151",
          6063 => x"ff527080",
          6064 => x"2ea03872",
          6065 => x"81ff0651",
          6066 => x"87c09480",
          6067 => x"5270802e",
          6068 => x"863887c0",
          6069 => x"94905271",
          6070 => x"0870982b",
          6071 => x"70982c51",
          6072 => x"53517182",
          6073 => x"bbdc0c84",
          6074 => x"3d0d04ff",
          6075 => x"3d0d87c0",
          6076 => x"9e800870",
          6077 => x"9c2a8a06",
          6078 => x"51517080",
          6079 => x"2e84b438",
          6080 => x"87c09ea4",
          6081 => x"0882ba80",
          6082 => x"0c87c09e",
          6083 => x"a80882ba",
          6084 => x"840c87c0",
          6085 => x"9e940882",
          6086 => x"ba880c87",
          6087 => x"c09e9808",
          6088 => x"82ba8c0c",
          6089 => x"87c09e9c",
          6090 => x"0882ba90",
          6091 => x"0c87c09e",
          6092 => x"a00882ba",
          6093 => x"940c87c0",
          6094 => x"9eac0882",
          6095 => x"ba980c87",
          6096 => x"c09eb008",
          6097 => x"82ba9c0c",
          6098 => x"87c09eb4",
          6099 => x"0882baa0",
          6100 => x"0c87c09e",
          6101 => x"b80882ba",
          6102 => x"a40c87c0",
          6103 => x"9ebc0882",
          6104 => x"baa80c87",
          6105 => x"c09ec008",
          6106 => x"82baac0c",
          6107 => x"87c09ec4",
          6108 => x"0882bab0",
          6109 => x"0c87c09e",
          6110 => x"80085170",
          6111 => x"82bab423",
          6112 => x"87c09e84",
          6113 => x"0882bab8",
          6114 => x"0c87c09e",
          6115 => x"880882ba",
          6116 => x"bc0c87c0",
          6117 => x"9e8c0882",
          6118 => x"bac00c81",
          6119 => x"0b82bac4",
          6120 => x"34800b87",
          6121 => x"c09e9008",
          6122 => x"7084800a",
          6123 => x"06515252",
          6124 => x"70802e83",
          6125 => x"38815271",
          6126 => x"82bac534",
          6127 => x"800b87c0",
          6128 => x"9e900870",
          6129 => x"88800a06",
          6130 => x"51525270",
          6131 => x"802e8338",
          6132 => x"81527182",
          6133 => x"bac63480",
          6134 => x"0b87c09e",
          6135 => x"90087090",
          6136 => x"800a0651",
          6137 => x"52527080",
          6138 => x"2e833881",
          6139 => x"527182ba",
          6140 => x"c734800b",
          6141 => x"87c09e90",
          6142 => x"08708880",
          6143 => x"80065152",
          6144 => x"5270802e",
          6145 => x"83388152",
          6146 => x"7182bac8",
          6147 => x"34800b87",
          6148 => x"c09e9008",
          6149 => x"70a08080",
          6150 => x"06515252",
          6151 => x"70802e83",
          6152 => x"38815271",
          6153 => x"82bac934",
          6154 => x"800b87c0",
          6155 => x"9e900870",
          6156 => x"90808006",
          6157 => x"51525270",
          6158 => x"802e8338",
          6159 => x"81527182",
          6160 => x"baca3480",
          6161 => x"0b87c09e",
          6162 => x"90087084",
          6163 => x"80800651",
          6164 => x"52527080",
          6165 => x"2e833881",
          6166 => x"527182ba",
          6167 => x"cb34800b",
          6168 => x"87c09e90",
          6169 => x"08708280",
          6170 => x"80065152",
          6171 => x"5270802e",
          6172 => x"83388152",
          6173 => x"7182bacc",
          6174 => x"34800b87",
          6175 => x"c09e9008",
          6176 => x"70818080",
          6177 => x"06515252",
          6178 => x"70802e83",
          6179 => x"38815271",
          6180 => x"82bacd34",
          6181 => x"800b87c0",
          6182 => x"9e900870",
          6183 => x"80c08006",
          6184 => x"51525270",
          6185 => x"802e8338",
          6186 => x"81527182",
          6187 => x"bace3480",
          6188 => x"0b87c09e",
          6189 => x"900870a0",
          6190 => x"80065152",
          6191 => x"5270802e",
          6192 => x"83388152",
          6193 => x"7182bacf",
          6194 => x"3487c09e",
          6195 => x"90087098",
          6196 => x"8006708a",
          6197 => x"2a515151",
          6198 => x"7082bad0",
          6199 => x"34800b87",
          6200 => x"c09e9008",
          6201 => x"70848006",
          6202 => x"51525270",
          6203 => x"802e8338",
          6204 => x"81527182",
          6205 => x"bad13487",
          6206 => x"c09e9008",
          6207 => x"7083f006",
          6208 => x"70842a51",
          6209 => x"51517082",
          6210 => x"bad23480",
          6211 => x"0b87c09e",
          6212 => x"90087088",
          6213 => x"06515252",
          6214 => x"70802e83",
          6215 => x"38815271",
          6216 => x"82bad334",
          6217 => x"87c09e90",
          6218 => x"08708706",
          6219 => x"51517082",
          6220 => x"bad43483",
          6221 => x"3d0d04fb",
          6222 => x"3d0d82ab",
          6223 => x"9451ffad",
          6224 => x"a23f82ba",
          6225 => x"c4335473",
          6226 => x"802e8938",
          6227 => x"82aba851",
          6228 => x"ffad903f",
          6229 => x"82abbc51",
          6230 => x"ffad883f",
          6231 => x"82bac633",
          6232 => x"5473802e",
          6233 => x"943882ba",
          6234 => x"a00882ba",
          6235 => x"a4081154",
          6236 => x"5282abd4",
          6237 => x"51ff90e0",
          6238 => x"3f82bacb",
          6239 => x"33547380",
          6240 => x"2e943882",
          6241 => x"ba980882",
          6242 => x"ba9c0811",
          6243 => x"545282ab",
          6244 => x"f051ff90",
          6245 => x"c33f82ba",
          6246 => x"c8335473",
          6247 => x"802e9438",
          6248 => x"82ba8008",
          6249 => x"82ba8408",
          6250 => x"11545282",
          6251 => x"ac8c51ff",
          6252 => x"90a63f82",
          6253 => x"bac93354",
          6254 => x"73802e94",
          6255 => x"3882ba88",
          6256 => x"0882ba8c",
          6257 => x"08115452",
          6258 => x"82aca851",
          6259 => x"ff90893f",
          6260 => x"82baca33",
          6261 => x"5473802e",
          6262 => x"943882ba",
          6263 => x"900882ba",
          6264 => x"94081154",
          6265 => x"5282acc4",
          6266 => x"51ff8fec",
          6267 => x"3f82bacf",
          6268 => x"33547380",
          6269 => x"2e8e3882",
          6270 => x"bad03352",
          6271 => x"82ace051",
          6272 => x"ff8fd53f",
          6273 => x"82bad333",
          6274 => x"5473802e",
          6275 => x"8e3882ba",
          6276 => x"d4335282",
          6277 => x"ad8051ff",
          6278 => x"8fbe3f82",
          6279 => x"bad13354",
          6280 => x"73802e8e",
          6281 => x"3882bad2",
          6282 => x"335282ad",
          6283 => x"a051ff8f",
          6284 => x"a73f82ba",
          6285 => x"c5335473",
          6286 => x"802e8938",
          6287 => x"82adc051",
          6288 => x"ffaba03f",
          6289 => x"82bac733",
          6290 => x"5473802e",
          6291 => x"893882ad",
          6292 => x"d451ffab",
          6293 => x"8e3f82ba",
          6294 => x"cc335473",
          6295 => x"802e8938",
          6296 => x"82ade051",
          6297 => x"ffaafc3f",
          6298 => x"82bacd33",
          6299 => x"5473802e",
          6300 => x"893882ad",
          6301 => x"ec51ffaa",
          6302 => x"ea3f82ba",
          6303 => x"ce335473",
          6304 => x"802e8938",
          6305 => x"82adf851",
          6306 => x"ffaad83f",
          6307 => x"82ae8451",
          6308 => x"ffaad03f",
          6309 => x"82baa808",
          6310 => x"5282ae90",
          6311 => x"51ff8eb8",
          6312 => x"3f82baac",
          6313 => x"085282ae",
          6314 => x"b851ff8e",
          6315 => x"ab3f82ba",
          6316 => x"b0085282",
          6317 => x"aee051ff",
          6318 => x"8e9e3f82",
          6319 => x"af8851ff",
          6320 => x"aaa13f82",
          6321 => x"bab42252",
          6322 => x"82af9051",
          6323 => x"ff8e893f",
          6324 => x"82bab808",
          6325 => x"56bd84c0",
          6326 => x"527551c1",
          6327 => x"a63f82bb",
          6328 => x"dc08bd84",
          6329 => x"c0297671",
          6330 => x"31545482",
          6331 => x"bbdc0852",
          6332 => x"82afb851",
          6333 => x"ff8de13f",
          6334 => x"82bacb33",
          6335 => x"5473802e",
          6336 => x"a93882ba",
          6337 => x"bc0856bd",
          6338 => x"84c05275",
          6339 => x"51c0f43f",
          6340 => x"82bbdc08",
          6341 => x"bd84c029",
          6342 => x"76713154",
          6343 => x"5482bbdc",
          6344 => x"085282af",
          6345 => x"e451ff8d",
          6346 => x"af3f82ba",
          6347 => x"c6335473",
          6348 => x"802ea938",
          6349 => x"82bac008",
          6350 => x"56bd84c0",
          6351 => x"527551c0",
          6352 => x"c23f82bb",
          6353 => x"dc08bd84",
          6354 => x"c0297671",
          6355 => x"31545482",
          6356 => x"bbdc0852",
          6357 => x"82b09051",
          6358 => x"ff8cfd3f",
          6359 => x"82a7fc51",
          6360 => x"ffa9803f",
          6361 => x"873d0d04",
          6362 => x"fe3d0d02",
          6363 => x"920533ff",
          6364 => x"05527184",
          6365 => x"26aa3871",
          6366 => x"8429829a",
          6367 => x"ec055271",
          6368 => x"080482b0",
          6369 => x"bc519d39",
          6370 => x"82b0c451",
          6371 => x"973982b0",
          6372 => x"cc519139",
          6373 => x"82b0d451",
          6374 => x"8b3982b0",
          6375 => x"d8518539",
          6376 => x"82b0e051",
          6377 => x"ffa8bc3f",
          6378 => x"843d0d04",
          6379 => x"7188800c",
          6380 => x"04ff3d0d",
          6381 => x"87c09684",
          6382 => x"70085252",
          6383 => x"80720c70",
          6384 => x"74077082",
          6385 => x"bad80c72",
          6386 => x"0c833d0d",
          6387 => x"04ff3d0d",
          6388 => x"87c09684",
          6389 => x"700882ba",
          6390 => x"d80c5280",
          6391 => x"720c7309",
          6392 => x"7082bad8",
          6393 => x"08067082",
          6394 => x"bad80c73",
          6395 => x"0c51833d",
          6396 => x"0d04800b",
          6397 => x"87c09684",
          6398 => x"0c0482ba",
          6399 => x"d80887c0",
          6400 => x"96840c04",
          6401 => x"fd3d0d76",
          6402 => x"982b7098",
          6403 => x"2c79982b",
          6404 => x"70982c72",
          6405 => x"10137082",
          6406 => x"2b515351",
          6407 => x"54515180",
          6408 => x"0b82b0ec",
          6409 => x"12335553",
          6410 => x"7174259c",
          6411 => x"3882b0e8",
          6412 => x"11081202",
          6413 => x"84059705",
          6414 => x"33713352",
          6415 => x"52527072",
          6416 => x"2e098106",
          6417 => x"83388153",
          6418 => x"7282bbdc",
          6419 => x"0c853d0d",
          6420 => x"04fb3d0d",
          6421 => x"79028405",
          6422 => x"a3053371",
          6423 => x"33555654",
          6424 => x"72802eb1",
          6425 => x"3882d3b0",
          6426 => x"08528851",
          6427 => x"ffaac33f",
          6428 => x"82d3b008",
          6429 => x"52a051ff",
          6430 => x"aab83f82",
          6431 => x"d3b00852",
          6432 => x"8851ffaa",
          6433 => x"ad3f7333",
          6434 => x"ff055372",
          6435 => x"74347281",
          6436 => x"ff0653cc",
          6437 => x"397751ff",
          6438 => x"8abe3f74",
          6439 => x"7434873d",
          6440 => x"0d04f63d",
          6441 => x"0d7c0284",
          6442 => x"05b70533",
          6443 => x"028805bb",
          6444 => x"053382bb",
          6445 => x"b4337084",
          6446 => x"2982badc",
          6447 => x"05700851",
          6448 => x"59595a58",
          6449 => x"5974802e",
          6450 => x"86387451",
          6451 => x"9afa3f82",
          6452 => x"bbb43370",
          6453 => x"842982ba",
          6454 => x"dc058119",
          6455 => x"70545856",
          6456 => x"5a9dfb3f",
          6457 => x"82bbdc08",
          6458 => x"750c82bb",
          6459 => x"b4337084",
          6460 => x"2982badc",
          6461 => x"05700851",
          6462 => x"565a7480",
          6463 => x"2ea73875",
          6464 => x"53785274",
          6465 => x"51ffb3dd",
          6466 => x"3f82bbb4",
          6467 => x"33810555",
          6468 => x"7482bbb4",
          6469 => x"347481ff",
          6470 => x"06559375",
          6471 => x"27873880",
          6472 => x"0b82bbb4",
          6473 => x"3477802e",
          6474 => x"b63882bb",
          6475 => x"b0085675",
          6476 => x"802eac38",
          6477 => x"82bbac33",
          6478 => x"5574a438",
          6479 => x"8c3dfc05",
          6480 => x"54765378",
          6481 => x"52755180",
          6482 => x"da883f82",
          6483 => x"bbb00852",
          6484 => x"8a51818f",
          6485 => x"953f82bb",
          6486 => x"b0085180",
          6487 => x"dde53f8c",
          6488 => x"3d0d04fd",
          6489 => x"3d0d82ba",
          6490 => x"dc539354",
          6491 => x"72085271",
          6492 => x"802e8938",
          6493 => x"715199d0",
          6494 => x"3f80730c",
          6495 => x"ff148414",
          6496 => x"54547380",
          6497 => x"25e63880",
          6498 => x"0b82bbb4",
          6499 => x"3482bbb0",
          6500 => x"08527180",
          6501 => x"2e953871",
          6502 => x"5180dec5",
          6503 => x"3f82bbb0",
          6504 => x"085199a4",
          6505 => x"3f800b82",
          6506 => x"bbb00c85",
          6507 => x"3d0d04dc",
          6508 => x"3d0d8157",
          6509 => x"805282bb",
          6510 => x"b0085180",
          6511 => x"e3b23f82",
          6512 => x"bbdc0880",
          6513 => x"d33882bb",
          6514 => x"b0085380",
          6515 => x"f852883d",
          6516 => x"70525681",
          6517 => x"8c803f82",
          6518 => x"bbdc0880",
          6519 => x"2eba3875",
          6520 => x"51ffb0a1",
          6521 => x"3f82bbdc",
          6522 => x"0855800b",
          6523 => x"82bbdc08",
          6524 => x"259d3882",
          6525 => x"bbdc08ff",
          6526 => x"05701755",
          6527 => x"55807434",
          6528 => x"75537652",
          6529 => x"811782b3",
          6530 => x"dc5257ff",
          6531 => x"87ca3f74",
          6532 => x"ff2e0981",
          6533 => x"06ffaf38",
          6534 => x"a63d0d04",
          6535 => x"d93d0daa",
          6536 => x"3d08ad3d",
          6537 => x"085a5a81",
          6538 => x"70585880",
          6539 => x"5282bbb0",
          6540 => x"085180e2",
          6541 => x"bb3f82bb",
          6542 => x"dc088195",
          6543 => x"38ff0b82",
          6544 => x"bbb00854",
          6545 => x"5580f852",
          6546 => x"8b3d7052",
          6547 => x"56818b86",
          6548 => x"3f82bbdc",
          6549 => x"08802ea5",
          6550 => x"387551ff",
          6551 => x"afa73f82",
          6552 => x"bbdc0881",
          6553 => x"18585580",
          6554 => x"0b82bbdc",
          6555 => x"08258e38",
          6556 => x"82bbdc08",
          6557 => x"ff057017",
          6558 => x"55558074",
          6559 => x"34740970",
          6560 => x"30707207",
          6561 => x"9f2a5155",
          6562 => x"5578772e",
          6563 => x"853873ff",
          6564 => x"ac3882bb",
          6565 => x"b0088c11",
          6566 => x"08535180",
          6567 => x"e1d23f82",
          6568 => x"bbdc0880",
          6569 => x"2e893882",
          6570 => x"b3e851ff",
          6571 => x"86aa3f78",
          6572 => x"772e0981",
          6573 => x"069b3875",
          6574 => x"527951ff",
          6575 => x"afb53f79",
          6576 => x"51ffaec1",
          6577 => x"3fab3d08",
          6578 => x"5482bbdc",
          6579 => x"08743480",
          6580 => x"587782bb",
          6581 => x"dc0ca93d",
          6582 => x"0d04f63d",
          6583 => x"0d7c7e71",
          6584 => x"5c717233",
          6585 => x"57595a58",
          6586 => x"73a02e09",
          6587 => x"8106a238",
          6588 => x"78337805",
          6589 => x"56777627",
          6590 => x"98388117",
          6591 => x"705b7071",
          6592 => x"33565855",
          6593 => x"73a02e09",
          6594 => x"81068638",
          6595 => x"757526ea",
          6596 => x"38805473",
          6597 => x"882982bb",
          6598 => x"b8057008",
          6599 => x"5255ffad",
          6600 => x"e43f82bb",
          6601 => x"dc085379",
          6602 => x"52740851",
          6603 => x"ffb0e33f",
          6604 => x"82bbdc08",
          6605 => x"80c53884",
          6606 => x"15335574",
          6607 => x"812e8838",
          6608 => x"74822e88",
          6609 => x"38b539fc",
          6610 => x"e63fac39",
          6611 => x"811a5a8c",
          6612 => x"3dfc1153",
          6613 => x"f80551c0",
          6614 => x"f33f82bb",
          6615 => x"dc08802e",
          6616 => x"9a38ff1b",
          6617 => x"53785277",
          6618 => x"51fdb13f",
          6619 => x"82bbdc08",
          6620 => x"81ff0655",
          6621 => x"74853874",
          6622 => x"54913981",
          6623 => x"147081ff",
          6624 => x"06515482",
          6625 => x"7427ff8b",
          6626 => x"38805473",
          6627 => x"82bbdc0c",
          6628 => x"8c3d0d04",
          6629 => x"d33d0db0",
          6630 => x"3d08b23d",
          6631 => x"08b43d08",
          6632 => x"595f5a80",
          6633 => x"0baf3d34",
          6634 => x"82bbb433",
          6635 => x"82bbb008",
          6636 => x"555b7381",
          6637 => x"cb387382",
          6638 => x"bbac3355",
          6639 => x"55738338",
          6640 => x"81557680",
          6641 => x"2e81bc38",
          6642 => x"81707606",
          6643 => x"55567380",
          6644 => x"2e81ad38",
          6645 => x"a8519886",
          6646 => x"3f82bbdc",
          6647 => x"0882bbb0",
          6648 => x"0c82bbdc",
          6649 => x"08802e81",
          6650 => x"92389353",
          6651 => x"765282bb",
          6652 => x"dc085180",
          6653 => x"ccfa3f82",
          6654 => x"bbdc0880",
          6655 => x"2e8c3882",
          6656 => x"b49451ff",
          6657 => x"9fdd3f80",
          6658 => x"f73982bb",
          6659 => x"dc085b82",
          6660 => x"bbb00853",
          6661 => x"80f85290",
          6662 => x"3d705254",
          6663 => x"8187b73f",
          6664 => x"82bbdc08",
          6665 => x"5682bbdc",
          6666 => x"08742e09",
          6667 => x"810680d0",
          6668 => x"3882bbdc",
          6669 => x"0851ffab",
          6670 => x"cc3f82bb",
          6671 => x"dc085580",
          6672 => x"0b82bbdc",
          6673 => x"0825a938",
          6674 => x"82bbdc08",
          6675 => x"ff057017",
          6676 => x"55558074",
          6677 => x"34805374",
          6678 => x"81ff0652",
          6679 => x"7551f8c2",
          6680 => x"3f811b70",
          6681 => x"81ff065c",
          6682 => x"54937b27",
          6683 => x"8338805b",
          6684 => x"74ff2e09",
          6685 => x"8106ff97",
          6686 => x"38863975",
          6687 => x"82bbac34",
          6688 => x"768c3882",
          6689 => x"bbb00880",
          6690 => x"2e8438f9",
          6691 => x"d63f8f3d",
          6692 => x"5dec823f",
          6693 => x"82bbdc08",
          6694 => x"982b7098",
          6695 => x"2c515978",
          6696 => x"ff2eee38",
          6697 => x"7881ff06",
          6698 => x"82d38833",
          6699 => x"70982b70",
          6700 => x"982c82d3",
          6701 => x"84337098",
          6702 => x"2b70972c",
          6703 => x"71982c05",
          6704 => x"70842982",
          6705 => x"b0e80570",
          6706 => x"08157033",
          6707 => x"51515151",
          6708 => x"59595159",
          6709 => x"5d588156",
          6710 => x"73782e80",
          6711 => x"e9387774",
          6712 => x"27b43874",
          6713 => x"81800a29",
          6714 => x"81ff0a05",
          6715 => x"70982c51",
          6716 => x"55807524",
          6717 => x"80ce3876",
          6718 => x"53745277",
          6719 => x"51f6853f",
          6720 => x"82bbdc08",
          6721 => x"81ff0654",
          6722 => x"73802ed7",
          6723 => x"387482d3",
          6724 => x"84348156",
          6725 => x"b1397481",
          6726 => x"800a2981",
          6727 => x"800a0570",
          6728 => x"982c7081",
          6729 => x"ff065651",
          6730 => x"55739526",
          6731 => x"97387653",
          6732 => x"74527751",
          6733 => x"f5ce3f82",
          6734 => x"bbdc0881",
          6735 => x"ff065473",
          6736 => x"cc38d339",
          6737 => x"80567580",
          6738 => x"2e80ca38",
          6739 => x"811c5574",
          6740 => x"82d38834",
          6741 => x"74982b70",
          6742 => x"982c82d3",
          6743 => x"84337098",
          6744 => x"2b70982c",
          6745 => x"70101170",
          6746 => x"822b82b0",
          6747 => x"ec11335e",
          6748 => x"51515157",
          6749 => x"58515574",
          6750 => x"772e0981",
          6751 => x"06fe9238",
          6752 => x"82b0f014",
          6753 => x"087d0c80",
          6754 => x"0b82d388",
          6755 => x"34800b82",
          6756 => x"d3843492",
          6757 => x"397582d3",
          6758 => x"88347582",
          6759 => x"d3843478",
          6760 => x"af3d3475",
          6761 => x"7d0c7e54",
          6762 => x"739526fd",
          6763 => x"e1387384",
          6764 => x"29829b80",
          6765 => x"05547308",
          6766 => x"0482d390",
          6767 => x"3354737e",
          6768 => x"2efdcb38",
          6769 => x"82d38c33",
          6770 => x"55737527",
          6771 => x"ab387498",
          6772 => x"2b70982c",
          6773 => x"51557375",
          6774 => x"249e3874",
          6775 => x"1a547333",
          6776 => x"81153474",
          6777 => x"81800a29",
          6778 => x"81ff0a05",
          6779 => x"70982c82",
          6780 => x"d3903356",
          6781 => x"5155df39",
          6782 => x"82d39033",
          6783 => x"81115654",
          6784 => x"7482d390",
          6785 => x"34731a54",
          6786 => x"ae3d3374",
          6787 => x"3482d38c",
          6788 => x"3354737e",
          6789 => x"25893881",
          6790 => x"14547382",
          6791 => x"d38c3482",
          6792 => x"d3903370",
          6793 => x"81800a29",
          6794 => x"81ff0a05",
          6795 => x"70982c82",
          6796 => x"d38c335a",
          6797 => x"51565674",
          6798 => x"7725a838",
          6799 => x"82d3b008",
          6800 => x"52741a70",
          6801 => x"335254ff",
          6802 => x"9ee83f74",
          6803 => x"81800a29",
          6804 => x"81800a05",
          6805 => x"70982c82",
          6806 => x"d38c3356",
          6807 => x"51557375",
          6808 => x"24da3882",
          6809 => x"d3903370",
          6810 => x"982b7098",
          6811 => x"2c82d38c",
          6812 => x"335a5156",
          6813 => x"56747725",
          6814 => x"fc943882",
          6815 => x"d3b00852",
          6816 => x"8851ff9e",
          6817 => x"ad3f7481",
          6818 => x"800a2981",
          6819 => x"800a0570",
          6820 => x"982c82d3",
          6821 => x"8c335651",
          6822 => x"55737524",
          6823 => x"de38fbee",
          6824 => x"39837a34",
          6825 => x"800b811b",
          6826 => x"3482d390",
          6827 => x"53805282",
          6828 => x"a3bc51f3",
          6829 => x"9c3f81fd",
          6830 => x"3982d390",
          6831 => x"337081ff",
          6832 => x"06555573",
          6833 => x"802efbc6",
          6834 => x"3882d38c",
          6835 => x"33ff0554",
          6836 => x"7382d38c",
          6837 => x"34ff1554",
          6838 => x"7382d390",
          6839 => x"3482d3b0",
          6840 => x"08528851",
          6841 => x"ff9dcb3f",
          6842 => x"82d39033",
          6843 => x"70982b70",
          6844 => x"982c82d3",
          6845 => x"8c335751",
          6846 => x"56577474",
          6847 => x"25ad3874",
          6848 => x"1a548114",
          6849 => x"33743482",
          6850 => x"d3b00852",
          6851 => x"733351ff",
          6852 => x"9da03f74",
          6853 => x"81800a29",
          6854 => x"81800a05",
          6855 => x"70982c82",
          6856 => x"d38c3358",
          6857 => x"51557575",
          6858 => x"24d53882",
          6859 => x"d3b00852",
          6860 => x"a051ff9c",
          6861 => x"fd3f82d3",
          6862 => x"90337098",
          6863 => x"2b70982c",
          6864 => x"82d38c33",
          6865 => x"57515657",
          6866 => x"747424fa",
          6867 => x"c13882d3",
          6868 => x"b0085288",
          6869 => x"51ff9cda",
          6870 => x"3f748180",
          6871 => x"0a298180",
          6872 => x"0a057098",
          6873 => x"2c82d38c",
          6874 => x"33585155",
          6875 => x"757525de",
          6876 => x"38fa9b39",
          6877 => x"82d38c33",
          6878 => x"7a055480",
          6879 => x"743482d3",
          6880 => x"b008528a",
          6881 => x"51ff9caa",
          6882 => x"3f82d38c",
          6883 => x"527951f6",
          6884 => x"c93f82bb",
          6885 => x"dc0881ff",
          6886 => x"06547396",
          6887 => x"3882d38c",
          6888 => x"33547380",
          6889 => x"2e8f3881",
          6890 => x"53735279",
          6891 => x"51f1f33f",
          6892 => x"8439807a",
          6893 => x"34800b82",
          6894 => x"d3903480",
          6895 => x"0b82d38c",
          6896 => x"347982bb",
          6897 => x"dc0caf3d",
          6898 => x"0d0482d3",
          6899 => x"90335473",
          6900 => x"802ef9ba",
          6901 => x"3882d3b0",
          6902 => x"08528851",
          6903 => x"ff9bd33f",
          6904 => x"82d39033",
          6905 => x"ff055473",
          6906 => x"82d39034",
          6907 => x"7381ff06",
          6908 => x"54dd3982",
          6909 => x"d3903382",
          6910 => x"d38c3355",
          6911 => x"5573752e",
          6912 => x"f98c38ff",
          6913 => x"14547382",
          6914 => x"d38c3474",
          6915 => x"982b7098",
          6916 => x"2c7581ff",
          6917 => x"06565155",
          6918 => x"747425ad",
          6919 => x"38741a54",
          6920 => x"81143374",
          6921 => x"3482d3b0",
          6922 => x"08527333",
          6923 => x"51ff9b82",
          6924 => x"3f748180",
          6925 => x"0a298180",
          6926 => x"0a057098",
          6927 => x"2c82d38c",
          6928 => x"33585155",
          6929 => x"757524d5",
          6930 => x"3882d3b0",
          6931 => x"0852a051",
          6932 => x"ff9adf3f",
          6933 => x"82d39033",
          6934 => x"70982b70",
          6935 => x"982c82d3",
          6936 => x"8c335751",
          6937 => x"56577474",
          6938 => x"24f8a338",
          6939 => x"82d3b008",
          6940 => x"528851ff",
          6941 => x"9abc3f74",
          6942 => x"81800a29",
          6943 => x"81800a05",
          6944 => x"70982c82",
          6945 => x"d38c3358",
          6946 => x"51557575",
          6947 => x"25de38f7",
          6948 => x"fd3982d3",
          6949 => x"90337081",
          6950 => x"ff0682d3",
          6951 => x"8c335956",
          6952 => x"54747727",
          6953 => x"f7e83882",
          6954 => x"d3b00852",
          6955 => x"81145473",
          6956 => x"82d39034",
          6957 => x"741a7033",
          6958 => x"5254ff99",
          6959 => x"f53f82d3",
          6960 => x"90337081",
          6961 => x"ff0682d3",
          6962 => x"8c335856",
          6963 => x"54757526",
          6964 => x"d638f7ba",
          6965 => x"3982d390",
          6966 => x"53805282",
          6967 => x"a3bc51ee",
          6968 => x"f03f800b",
          6969 => x"82d39034",
          6970 => x"800b82d3",
          6971 => x"8c34f79e",
          6972 => x"397ab038",
          6973 => x"82bba808",
          6974 => x"5574802e",
          6975 => x"a6387451",
          6976 => x"ffa2823f",
          6977 => x"82bbdc08",
          6978 => x"82d38c34",
          6979 => x"82bbdc08",
          6980 => x"81ff0681",
          6981 => x"05537452",
          6982 => x"7951ffa3",
          6983 => x"c83f935b",
          6984 => x"81c0397a",
          6985 => x"842982ba",
          6986 => x"dc05fc11",
          6987 => x"08565474",
          6988 => x"802ea738",
          6989 => x"7451ffa1",
          6990 => x"cc3f82bb",
          6991 => x"dc0882d3",
          6992 => x"8c3482bb",
          6993 => x"dc0881ff",
          6994 => x"06810553",
          6995 => x"74527951",
          6996 => x"ffa3923f",
          6997 => x"ff1b5480",
          6998 => x"fa397308",
          6999 => x"5574802e",
          7000 => x"f6ac3874",
          7001 => x"51ffa19d",
          7002 => x"3f99397a",
          7003 => x"932e0981",
          7004 => x"06ae3882",
          7005 => x"badc0855",
          7006 => x"74802ea4",
          7007 => x"387451ff",
          7008 => x"a1833f82",
          7009 => x"bbdc0882",
          7010 => x"d38c3482",
          7011 => x"bbdc0881",
          7012 => x"ff068105",
          7013 => x"53745279",
          7014 => x"51ffa2c9",
          7015 => x"3f80c339",
          7016 => x"7a842982",
          7017 => x"bae00570",
          7018 => x"08565474",
          7019 => x"802eab38",
          7020 => x"7451ffa0",
          7021 => x"d03f82bb",
          7022 => x"dc0882d3",
          7023 => x"8c3482bb",
          7024 => x"dc0881ff",
          7025 => x"06810553",
          7026 => x"74527951",
          7027 => x"ffa2963f",
          7028 => x"811b5473",
          7029 => x"81ff065b",
          7030 => x"89397482",
          7031 => x"d38c3474",
          7032 => x"7a3482d3",
          7033 => x"905382d3",
          7034 => x"8c335279",
          7035 => x"51ece23f",
          7036 => x"f59c3982",
          7037 => x"d3903370",
          7038 => x"81ff0682",
          7039 => x"d38c3359",
          7040 => x"56547477",
          7041 => x"27f58738",
          7042 => x"82d3b008",
          7043 => x"52811454",
          7044 => x"7382d390",
          7045 => x"34741a70",
          7046 => x"335254ff",
          7047 => x"97943ff4",
          7048 => x"ed3982d3",
          7049 => x"90335473",
          7050 => x"802ef4e2",
          7051 => x"3882d3b0",
          7052 => x"08528851",
          7053 => x"ff96fb3f",
          7054 => x"82d39033",
          7055 => x"ff055473",
          7056 => x"82d39034",
          7057 => x"f4c839f9",
          7058 => x"3d0d83c0",
          7059 => x"800b82bb",
          7060 => x"d40c8480",
          7061 => x"0b82bbd0",
          7062 => x"23a08053",
          7063 => x"805283c0",
          7064 => x"8051ffa6",
          7065 => x"813f82bb",
          7066 => x"d4085480",
          7067 => x"58777434",
          7068 => x"81577681",
          7069 => x"153482bb",
          7070 => x"d4085477",
          7071 => x"84153476",
          7072 => x"85153482",
          7073 => x"bbd40854",
          7074 => x"77861534",
          7075 => x"76871534",
          7076 => x"82bbd408",
          7077 => x"82bbd022",
          7078 => x"ff05fe80",
          7079 => x"80077083",
          7080 => x"ffff0670",
          7081 => x"882a5851",
          7082 => x"55567488",
          7083 => x"17347389",
          7084 => x"173482bb",
          7085 => x"d0227088",
          7086 => x"2982bbd4",
          7087 => x"0805f811",
          7088 => x"51555577",
          7089 => x"82153476",
          7090 => x"83153489",
          7091 => x"3d0d04ff",
          7092 => x"3d0d7352",
          7093 => x"81518472",
          7094 => x"278f38fb",
          7095 => x"12832a82",
          7096 => x"117083ff",
          7097 => x"ff065151",
          7098 => x"517082bb",
          7099 => x"dc0c833d",
          7100 => x"0d04f93d",
          7101 => x"0d02a605",
          7102 => x"22028405",
          7103 => x"aa052271",
          7104 => x"0582bbd4",
          7105 => x"0871832b",
          7106 => x"71117483",
          7107 => x"2b731170",
          7108 => x"33811233",
          7109 => x"71882b07",
          7110 => x"02a405ae",
          7111 => x"05227181",
          7112 => x"ffff0607",
          7113 => x"70882a53",
          7114 => x"51525954",
          7115 => x"5b5b5753",
          7116 => x"54557177",
          7117 => x"34708118",
          7118 => x"3482bbd4",
          7119 => x"08147588",
          7120 => x"2a525470",
          7121 => x"82153474",
          7122 => x"83153482",
          7123 => x"bbd40870",
          7124 => x"17703381",
          7125 => x"12337188",
          7126 => x"2b077083",
          7127 => x"2b8ffff8",
          7128 => x"06515256",
          7129 => x"52710573",
          7130 => x"83ffff06",
          7131 => x"70882a54",
          7132 => x"54517182",
          7133 => x"12347281",
          7134 => x"ff065372",
          7135 => x"83123482",
          7136 => x"bbd40816",
          7137 => x"56717634",
          7138 => x"72811734",
          7139 => x"893d0d04",
          7140 => x"fb3d0d82",
          7141 => x"bbd40802",
          7142 => x"84059e05",
          7143 => x"2270832b",
          7144 => x"72118611",
          7145 => x"33871233",
          7146 => x"718b2b71",
          7147 => x"832b0758",
          7148 => x"5b595255",
          7149 => x"52720584",
          7150 => x"12338513",
          7151 => x"3371882b",
          7152 => x"0770882a",
          7153 => x"54565652",
          7154 => x"70841334",
          7155 => x"73851334",
          7156 => x"82bbd408",
          7157 => x"70148411",
          7158 => x"33851233",
          7159 => x"718b2b71",
          7160 => x"832b0756",
          7161 => x"59575272",
          7162 => x"05861233",
          7163 => x"87133371",
          7164 => x"882b0770",
          7165 => x"882a5456",
          7166 => x"56527086",
          7167 => x"13347387",
          7168 => x"133482bb",
          7169 => x"d4081370",
          7170 => x"33811233",
          7171 => x"71882b07",
          7172 => x"7081ffff",
          7173 => x"0670882a",
          7174 => x"53515353",
          7175 => x"53717334",
          7176 => x"70811434",
          7177 => x"873d0d04",
          7178 => x"fa3d0d02",
          7179 => x"a2052282",
          7180 => x"bbd40871",
          7181 => x"832b7111",
          7182 => x"70338112",
          7183 => x"3371882b",
          7184 => x"07708829",
          7185 => x"15703381",
          7186 => x"12337198",
          7187 => x"2b71902b",
          7188 => x"07535f53",
          7189 => x"55525a56",
          7190 => x"57535471",
          7191 => x"802580f6",
          7192 => x"387251fe",
          7193 => x"ab3f82bb",
          7194 => x"d4087016",
          7195 => x"70338112",
          7196 => x"33718b2b",
          7197 => x"71832b07",
          7198 => x"74117033",
          7199 => x"81123371",
          7200 => x"882b0770",
          7201 => x"832b8fff",
          7202 => x"f8065152",
          7203 => x"5451535a",
          7204 => x"58537205",
          7205 => x"74882a54",
          7206 => x"52728213",
          7207 => x"34738313",
          7208 => x"3482bbd4",
          7209 => x"08701670",
          7210 => x"33811233",
          7211 => x"718b2b71",
          7212 => x"832b0756",
          7213 => x"59575572",
          7214 => x"05703381",
          7215 => x"12337188",
          7216 => x"2b077081",
          7217 => x"ffff0670",
          7218 => x"882a5751",
          7219 => x"52585272",
          7220 => x"74347181",
          7221 => x"1534883d",
          7222 => x"0d04fb3d",
          7223 => x"0d82bbd4",
          7224 => x"08028405",
          7225 => x"9e052270",
          7226 => x"832b7211",
          7227 => x"82113383",
          7228 => x"1233718b",
          7229 => x"2b71832b",
          7230 => x"07595b59",
          7231 => x"52565273",
          7232 => x"05713381",
          7233 => x"13337188",
          7234 => x"2b07028c",
          7235 => x"05a20522",
          7236 => x"71077088",
          7237 => x"2a535153",
          7238 => x"53537173",
          7239 => x"34708114",
          7240 => x"3482bbd4",
          7241 => x"08701570",
          7242 => x"33811233",
          7243 => x"718b2b71",
          7244 => x"832b0756",
          7245 => x"59575272",
          7246 => x"05821233",
          7247 => x"83133371",
          7248 => x"882b0770",
          7249 => x"882a5455",
          7250 => x"56527082",
          7251 => x"13347283",
          7252 => x"133482bb",
          7253 => x"d4081482",
          7254 => x"11338312",
          7255 => x"3371882b",
          7256 => x"0782bbdc",
          7257 => x"0c525487",
          7258 => x"3d0d04f7",
          7259 => x"3d0d7b82",
          7260 => x"bbd40831",
          7261 => x"832a7083",
          7262 => x"ffff0670",
          7263 => x"535753fd",
          7264 => x"a73f82bb",
          7265 => x"d4087683",
          7266 => x"2b711182",
          7267 => x"11338312",
          7268 => x"33718b2b",
          7269 => x"71832b07",
          7270 => x"75117033",
          7271 => x"81123371",
          7272 => x"982b7190",
          7273 => x"2b075342",
          7274 => x"4051535b",
          7275 => x"58555954",
          7276 => x"7280258d",
          7277 => x"38828080",
          7278 => x"527551fe",
          7279 => x"9d3f8184",
          7280 => x"39841433",
          7281 => x"85153371",
          7282 => x"8b2b7183",
          7283 => x"2b077611",
          7284 => x"79882a53",
          7285 => x"51555855",
          7286 => x"76861434",
          7287 => x"7581ff06",
          7288 => x"56758714",
          7289 => x"3482bbd4",
          7290 => x"08701984",
          7291 => x"12338513",
          7292 => x"3371882b",
          7293 => x"0770882a",
          7294 => x"54575b56",
          7295 => x"53728416",
          7296 => x"34738516",
          7297 => x"3482bbd4",
          7298 => x"08185380",
          7299 => x"0b861434",
          7300 => x"800b8714",
          7301 => x"3482bbd4",
          7302 => x"08537684",
          7303 => x"14347585",
          7304 => x"143482bb",
          7305 => x"d4081870",
          7306 => x"33811233",
          7307 => x"71882b07",
          7308 => x"70828080",
          7309 => x"0770882a",
          7310 => x"53515556",
          7311 => x"54747434",
          7312 => x"72811534",
          7313 => x"8b3d0d04",
          7314 => x"ff3d0d73",
          7315 => x"5282bbd4",
          7316 => x"088438f7",
          7317 => x"f23f7180",
          7318 => x"2e863871",
          7319 => x"51fe8c3f",
          7320 => x"833d0d04",
          7321 => x"f53d0d80",
          7322 => x"7e5258f8",
          7323 => x"e23f82bb",
          7324 => x"dc0883ff",
          7325 => x"ff0682bb",
          7326 => x"d4088411",
          7327 => x"33851233",
          7328 => x"71882b07",
          7329 => x"705f5956",
          7330 => x"585a81ff",
          7331 => x"ff597578",
          7332 => x"2e80cb38",
          7333 => x"75882917",
          7334 => x"70338112",
          7335 => x"3371882b",
          7336 => x"077081ff",
          7337 => x"ff067931",
          7338 => x"7083ffff",
          7339 => x"06707f27",
          7340 => x"52535156",
          7341 => x"59557779",
          7342 => x"278a3873",
          7343 => x"802e8538",
          7344 => x"75785a5b",
          7345 => x"84153385",
          7346 => x"16337188",
          7347 => x"2b075754",
          7348 => x"75c23878",
          7349 => x"81ffff2e",
          7350 => x"85387a79",
          7351 => x"59568076",
          7352 => x"832b82bb",
          7353 => x"d4081170",
          7354 => x"33811233",
          7355 => x"71882b07",
          7356 => x"7081ffff",
          7357 => x"0651525a",
          7358 => x"565c5573",
          7359 => x"752e8338",
          7360 => x"81558054",
          7361 => x"79782681",
          7362 => x"cc387454",
          7363 => x"74802e81",
          7364 => x"c438777a",
          7365 => x"2e098106",
          7366 => x"89387551",
          7367 => x"f8f23f81",
          7368 => x"ac398280",
          7369 => x"80537952",
          7370 => x"7551f7c6",
          7371 => x"3f82bbd4",
          7372 => x"08701c86",
          7373 => x"11338712",
          7374 => x"33718b2b",
          7375 => x"71832b07",
          7376 => x"535a5e55",
          7377 => x"74057a17",
          7378 => x"7083ffff",
          7379 => x"0670882a",
          7380 => x"5c595654",
          7381 => x"78841534",
          7382 => x"7681ff06",
          7383 => x"57768515",
          7384 => x"3482bbd4",
          7385 => x"0875832b",
          7386 => x"7111721e",
          7387 => x"86113387",
          7388 => x"12337188",
          7389 => x"2b077088",
          7390 => x"2a535b5e",
          7391 => x"535a5654",
          7392 => x"73861934",
          7393 => x"75871934",
          7394 => x"82bbd408",
          7395 => x"701c8411",
          7396 => x"33851233",
          7397 => x"718b2b71",
          7398 => x"832b0753",
          7399 => x"5d5a5574",
          7400 => x"05547886",
          7401 => x"15347687",
          7402 => x"153482bb",
          7403 => x"d4087016",
          7404 => x"711d8411",
          7405 => x"33851233",
          7406 => x"71882b07",
          7407 => x"70882a53",
          7408 => x"5a5f5256",
          7409 => x"54738416",
          7410 => x"34758516",
          7411 => x"3482bbd4",
          7412 => x"081b8405",
          7413 => x"547382bb",
          7414 => x"dc0c8d3d",
          7415 => x"0d04fe3d",
          7416 => x"0d745282",
          7417 => x"bbd40884",
          7418 => x"38f4dc3f",
          7419 => x"71537180",
          7420 => x"2e8b3871",
          7421 => x"51fced3f",
          7422 => x"82bbdc08",
          7423 => x"537282bb",
          7424 => x"dc0c843d",
          7425 => x"0d04ee3d",
          7426 => x"0d646640",
          7427 => x"5c807042",
          7428 => x"4082bbd4",
          7429 => x"08602e09",
          7430 => x"81068438",
          7431 => x"f4a93f7b",
          7432 => x"8e387e51",
          7433 => x"ffb83f82",
          7434 => x"bbdc0854",
          7435 => x"83c7397e",
          7436 => x"8b387b51",
          7437 => x"fc923f7e",
          7438 => x"5483ba39",
          7439 => x"7e51f58f",
          7440 => x"3f82bbdc",
          7441 => x"0883ffff",
          7442 => x"0682bbd4",
          7443 => x"087d7131",
          7444 => x"832a7083",
          7445 => x"ffff0670",
          7446 => x"832b7311",
          7447 => x"70338112",
          7448 => x"3371882b",
          7449 => x"07707531",
          7450 => x"7083ffff",
          7451 => x"06708829",
          7452 => x"fc057388",
          7453 => x"291a7033",
          7454 => x"81123371",
          7455 => x"882b0770",
          7456 => x"902b5344",
          7457 => x"4e534841",
          7458 => x"525c545b",
          7459 => x"415c565b",
          7460 => x"5b738025",
          7461 => x"8f387681",
          7462 => x"ffff0675",
          7463 => x"317083ff",
          7464 => x"ff064254",
          7465 => x"82163383",
          7466 => x"17337188",
          7467 => x"2b077088",
          7468 => x"291c7033",
          7469 => x"81123371",
          7470 => x"982b7190",
          7471 => x"2b075347",
          7472 => x"45525654",
          7473 => x"7380258b",
          7474 => x"38787531",
          7475 => x"7083ffff",
          7476 => x"06415477",
          7477 => x"7b2781fe",
          7478 => x"38601854",
          7479 => x"737b2e09",
          7480 => x"81068f38",
          7481 => x"7851f6c0",
          7482 => x"3f7a83ff",
          7483 => x"ff065881",
          7484 => x"e5397f8e",
          7485 => x"387a7424",
          7486 => x"89387851",
          7487 => x"f6aa3f81",
          7488 => x"a5397f18",
          7489 => x"557a7524",
          7490 => x"80c83879",
          7491 => x"1d821133",
          7492 => x"83123371",
          7493 => x"882b0753",
          7494 => x"5754f4f4",
          7495 => x"3f805278",
          7496 => x"51f7b73f",
          7497 => x"82bbdc08",
          7498 => x"83ffff06",
          7499 => x"7e547c53",
          7500 => x"70832b82",
          7501 => x"bbd40811",
          7502 => x"84055355",
          7503 => x"59ff8edb",
          7504 => x"3f82bbd4",
          7505 => x"08148405",
          7506 => x"7583ffff",
          7507 => x"06595c81",
          7508 => x"85396015",
          7509 => x"547a7424",
          7510 => x"80d43878",
          7511 => x"51f5c93f",
          7512 => x"82bbd408",
          7513 => x"1d821133",
          7514 => x"83123371",
          7515 => x"882b0753",
          7516 => x"4354f49c",
          7517 => x"3f805278",
          7518 => x"51f6df3f",
          7519 => x"82bbdc08",
          7520 => x"83ffff06",
          7521 => x"7e547c53",
          7522 => x"70832b82",
          7523 => x"bbd40811",
          7524 => x"84055355",
          7525 => x"59ff8e83",
          7526 => x"3f82bbd4",
          7527 => x"08148405",
          7528 => x"60620519",
          7529 => x"555c7383",
          7530 => x"ffff0658",
          7531 => x"a9397b7f",
          7532 => x"5254f9b0",
          7533 => x"3f82bbdc",
          7534 => x"085c82bb",
          7535 => x"dc08802e",
          7536 => x"93387d53",
          7537 => x"735282bb",
          7538 => x"dc0851ff",
          7539 => x"92973f73",
          7540 => x"51f7983f",
          7541 => x"7a587a78",
          7542 => x"27993880",
          7543 => x"537a5278",
          7544 => x"51f28f3f",
          7545 => x"7a19832b",
          7546 => x"82bbd408",
          7547 => x"05840551",
          7548 => x"f6f93f7b",
          7549 => x"547382bb",
          7550 => x"dc0c943d",
          7551 => x"0d04fc3d",
          7552 => x"0d777729",
          7553 => x"705254fb",
          7554 => x"d53f82bb",
          7555 => x"dc085582",
          7556 => x"bbdc0880",
          7557 => x"2e8e3873",
          7558 => x"53805282",
          7559 => x"bbdc0851",
          7560 => x"ff96c33f",
          7561 => x"7482bbdc",
          7562 => x"0c863d0d",
          7563 => x"04ff3d0d",
          7564 => x"028f0533",
          7565 => x"51815270",
          7566 => x"72268738",
          7567 => x"82bbd811",
          7568 => x"33527182",
          7569 => x"bbdc0c83",
          7570 => x"3d0d04fc",
          7571 => x"3d0d029b",
          7572 => x"05330284",
          7573 => x"059f0533",
          7574 => x"56538351",
          7575 => x"72812680",
          7576 => x"e0387284",
          7577 => x"2b87c092",
          7578 => x"8c115351",
          7579 => x"88547480",
          7580 => x"2e843881",
          7581 => x"88547372",
          7582 => x"0c87c092",
          7583 => x"8c115181",
          7584 => x"710c850b",
          7585 => x"87c0988c",
          7586 => x"0c705271",
          7587 => x"08708206",
          7588 => x"51517080",
          7589 => x"2e8a3887",
          7590 => x"c0988c08",
          7591 => x"5170ec38",
          7592 => x"7108fc80",
          7593 => x"80065271",
          7594 => x"923887c0",
          7595 => x"988c0851",
          7596 => x"70802e87",
          7597 => x"387182bb",
          7598 => x"d8143482",
          7599 => x"bbd81333",
          7600 => x"517082bb",
          7601 => x"dc0c863d",
          7602 => x"0d04f33d",
          7603 => x"0d606264",
          7604 => x"028c05bf",
          7605 => x"05335740",
          7606 => x"585b8374",
          7607 => x"525afecd",
          7608 => x"3f82bbdc",
          7609 => x"0881067a",
          7610 => x"54527181",
          7611 => x"be387172",
          7612 => x"75842b87",
          7613 => x"c0928011",
          7614 => x"87c0928c",
          7615 => x"1287c092",
          7616 => x"8413415a",
          7617 => x"40575a58",
          7618 => x"850b87c0",
          7619 => x"988c0c76",
          7620 => x"7d0c8476",
          7621 => x"0c750870",
          7622 => x"852a7081",
          7623 => x"06515354",
          7624 => x"71802e8e",
          7625 => x"387b0852",
          7626 => x"717b7081",
          7627 => x"055d3481",
          7628 => x"19598074",
          7629 => x"a2065353",
          7630 => x"71732e83",
          7631 => x"38815378",
          7632 => x"83ff268f",
          7633 => x"3872802e",
          7634 => x"8a3887c0",
          7635 => x"988c0852",
          7636 => x"71c33887",
          7637 => x"c0988c08",
          7638 => x"5271802e",
          7639 => x"87387884",
          7640 => x"802e9938",
          7641 => x"81760c87",
          7642 => x"c0928c15",
          7643 => x"53720870",
          7644 => x"82065152",
          7645 => x"71f738ff",
          7646 => x"1a5a8d39",
          7647 => x"84801781",
          7648 => x"197081ff",
          7649 => x"065a5357",
          7650 => x"79802e90",
          7651 => x"3873fc80",
          7652 => x"80065271",
          7653 => x"87387d78",
          7654 => x"26feed38",
          7655 => x"73fc8080",
          7656 => x"06527180",
          7657 => x"2e833881",
          7658 => x"52715372",
          7659 => x"82bbdc0c",
          7660 => x"8f3d0d04",
          7661 => x"f33d0d60",
          7662 => x"6264028c",
          7663 => x"05bf0533",
          7664 => x"5740585b",
          7665 => x"83598074",
          7666 => x"5258fce1",
          7667 => x"3f82bbdc",
          7668 => x"08810679",
          7669 => x"54527178",
          7670 => x"2e098106",
          7671 => x"81b13877",
          7672 => x"74842b87",
          7673 => x"c0928011",
          7674 => x"87c0928c",
          7675 => x"1287c092",
          7676 => x"84134059",
          7677 => x"5f565a85",
          7678 => x"0b87c098",
          7679 => x"8c0c767d",
          7680 => x"0c82760c",
          7681 => x"80587508",
          7682 => x"70842a70",
          7683 => x"81065153",
          7684 => x"5471802e",
          7685 => x"8c387a70",
          7686 => x"81055c33",
          7687 => x"7c0c8118",
          7688 => x"5873812a",
          7689 => x"70810651",
          7690 => x"5271802e",
          7691 => x"8a3887c0",
          7692 => x"988c0852",
          7693 => x"71d03887",
          7694 => x"c0988c08",
          7695 => x"5271802e",
          7696 => x"87387784",
          7697 => x"802e9938",
          7698 => x"81760c87",
          7699 => x"c0928c15",
          7700 => x"53720870",
          7701 => x"82065152",
          7702 => x"71f738ff",
          7703 => x"19598d39",
          7704 => x"811a7081",
          7705 => x"ff068480",
          7706 => x"19595b52",
          7707 => x"78802e90",
          7708 => x"3873fc80",
          7709 => x"80065271",
          7710 => x"87387d7a",
          7711 => x"26fef838",
          7712 => x"73fc8080",
          7713 => x"06527180",
          7714 => x"2e833881",
          7715 => x"52715372",
          7716 => x"82bbdc0c",
          7717 => x"8f3d0d04",
          7718 => x"fa3d0d7a",
          7719 => x"028405a3",
          7720 => x"05330288",
          7721 => x"05a70533",
          7722 => x"71545456",
          7723 => x"57fafe3f",
          7724 => x"82bbdc08",
          7725 => x"81065383",
          7726 => x"547280fe",
          7727 => x"38850b87",
          7728 => x"c0988c0c",
          7729 => x"81567176",
          7730 => x"2e80dc38",
          7731 => x"71762493",
          7732 => x"3874842b",
          7733 => x"87c0928c",
          7734 => x"11545471",
          7735 => x"802e8d38",
          7736 => x"80d43971",
          7737 => x"832e80c6",
          7738 => x"3880cb39",
          7739 => x"72087081",
          7740 => x"2a708106",
          7741 => x"51515271",
          7742 => x"802e8a38",
          7743 => x"87c0988c",
          7744 => x"085271e8",
          7745 => x"3887c098",
          7746 => x"8c085271",
          7747 => x"96388173",
          7748 => x"0c87c092",
          7749 => x"8c145372",
          7750 => x"08708206",
          7751 => x"515271f7",
          7752 => x"38963980",
          7753 => x"56923988",
          7754 => x"800a770c",
          7755 => x"85398180",
          7756 => x"770c7256",
          7757 => x"83398456",
          7758 => x"75547382",
          7759 => x"bbdc0c88",
          7760 => x"3d0d04fe",
          7761 => x"3d0d7481",
          7762 => x"11337133",
          7763 => x"71882b07",
          7764 => x"82bbdc0c",
          7765 => x"5351843d",
          7766 => x"0d04fd3d",
          7767 => x"0d758311",
          7768 => x"33821233",
          7769 => x"71902b71",
          7770 => x"882b0781",
          7771 => x"14337072",
          7772 => x"07882b75",
          7773 => x"33710782",
          7774 => x"bbdc0c52",
          7775 => x"53545654",
          7776 => x"52853d0d",
          7777 => x"04ff3d0d",
          7778 => x"73028405",
          7779 => x"92052252",
          7780 => x"52707270",
          7781 => x"81055434",
          7782 => x"70882a51",
          7783 => x"70723483",
          7784 => x"3d0d04ff",
          7785 => x"3d0d7375",
          7786 => x"52527072",
          7787 => x"70810554",
          7788 => x"3470882a",
          7789 => x"51707270",
          7790 => x"81055434",
          7791 => x"70882a51",
          7792 => x"70727081",
          7793 => x"05543470",
          7794 => x"882a5170",
          7795 => x"7234833d",
          7796 => x"0d04fe3d",
          7797 => x"0d767577",
          7798 => x"54545170",
          7799 => x"802e9238",
          7800 => x"71708105",
          7801 => x"53337370",
          7802 => x"81055534",
          7803 => x"ff1151eb",
          7804 => x"39843d0d",
          7805 => x"04fe3d0d",
          7806 => x"75777654",
          7807 => x"52537272",
          7808 => x"70810554",
          7809 => x"34ff1151",
          7810 => x"70f43884",
          7811 => x"3d0d04fc",
          7812 => x"3d0d7877",
          7813 => x"79565653",
          7814 => x"74708105",
          7815 => x"56337470",
          7816 => x"81055633",
          7817 => x"717131ff",
          7818 => x"16565252",
          7819 => x"5272802e",
          7820 => x"86387180",
          7821 => x"2ee23871",
          7822 => x"82bbdc0c",
          7823 => x"863d0d04",
          7824 => x"fe3d0d74",
          7825 => x"76545189",
          7826 => x"3971732e",
          7827 => x"8a388111",
          7828 => x"51703352",
          7829 => x"71f33870",
          7830 => x"3382bbdc",
          7831 => x"0c843d0d",
          7832 => x"04800b82",
          7833 => x"bbdc0c04",
          7834 => x"800b82bb",
          7835 => x"dc0c04f7",
          7836 => x"3d0d7b56",
          7837 => x"800b8317",
          7838 => x"33565a74",
          7839 => x"7a2e80d6",
          7840 => x"388154b0",
          7841 => x"160853b4",
          7842 => x"16705381",
          7843 => x"17335259",
          7844 => x"faa23f82",
          7845 => x"bbdc087a",
          7846 => x"2e098106",
          7847 => x"b73882bb",
          7848 => x"dc088317",
          7849 => x"34b01608",
          7850 => x"70a41808",
          7851 => x"319c1808",
          7852 => x"59565874",
          7853 => x"77279f38",
          7854 => x"82163355",
          7855 => x"74822e09",
          7856 => x"81069338",
          7857 => x"81547618",
          7858 => x"53785281",
          7859 => x"163351f9",
          7860 => x"e33f8339",
          7861 => x"815a7982",
          7862 => x"bbdc0c8b",
          7863 => x"3d0d04fa",
          7864 => x"3d0d787a",
          7865 => x"56568057",
          7866 => x"74b01708",
          7867 => x"2eaf3875",
          7868 => x"51fefc3f",
          7869 => x"82bbdc08",
          7870 => x"5782bbdc",
          7871 => x"089f3881",
          7872 => x"547453b4",
          7873 => x"16528116",
          7874 => x"3351f7be",
          7875 => x"3f82bbdc",
          7876 => x"08802e85",
          7877 => x"38ff5581",
          7878 => x"5774b017",
          7879 => x"0c7682bb",
          7880 => x"dc0c883d",
          7881 => x"0d04f83d",
          7882 => x"0d7a7052",
          7883 => x"57fec03f",
          7884 => x"82bbdc08",
          7885 => x"5882bbdc",
          7886 => x"08819138",
          7887 => x"76335574",
          7888 => x"832e0981",
          7889 => x"0680f038",
          7890 => x"84173359",
          7891 => x"78812e09",
          7892 => x"810680e3",
          7893 => x"38848053",
          7894 => x"82bbdc08",
          7895 => x"52b41770",
          7896 => x"5256fd91",
          7897 => x"3f82d4d5",
          7898 => x"5284b217",
          7899 => x"51fc963f",
          7900 => x"848b85a4",
          7901 => x"d2527551",
          7902 => x"fca93f86",
          7903 => x"8a85e4f2",
          7904 => x"52849817",
          7905 => x"51fc9c3f",
          7906 => x"90170852",
          7907 => x"849c1751",
          7908 => x"fc913f8c",
          7909 => x"17085284",
          7910 => x"a01751fc",
          7911 => x"863fa017",
          7912 => x"08810570",
          7913 => x"b0190c79",
          7914 => x"55537552",
          7915 => x"81173351",
          7916 => x"f8823f77",
          7917 => x"84183480",
          7918 => x"53805281",
          7919 => x"173351f9",
          7920 => x"d73f82bb",
          7921 => x"dc08802e",
          7922 => x"83388158",
          7923 => x"7782bbdc",
          7924 => x"0c8a3d0d",
          7925 => x"04fb3d0d",
          7926 => x"77fe1a98",
          7927 => x"1208fe05",
          7928 => x"55565480",
          7929 => x"56747327",
          7930 => x"8d388a14",
          7931 => x"22757129",
          7932 => x"ac160805",
          7933 => x"57537582",
          7934 => x"bbdc0c87",
          7935 => x"3d0d04f9",
          7936 => x"3d0d7a7a",
          7937 => x"70085654",
          7938 => x"57817727",
          7939 => x"81df3876",
          7940 => x"98150827",
          7941 => x"81d738ff",
          7942 => x"74335458",
          7943 => x"72822e80",
          7944 => x"f5387282",
          7945 => x"24893872",
          7946 => x"812e8d38",
          7947 => x"81bf3972",
          7948 => x"832e818e",
          7949 => x"3881b639",
          7950 => x"76812a17",
          7951 => x"70892aa4",
          7952 => x"16080553",
          7953 => x"745255fd",
          7954 => x"963f82bb",
          7955 => x"dc08819f",
          7956 => x"387483ff",
          7957 => x"0614b411",
          7958 => x"33811770",
          7959 => x"892aa418",
          7960 => x"08055576",
          7961 => x"54575753",
          7962 => x"fcf53f82",
          7963 => x"bbdc0880",
          7964 => x"fe387483",
          7965 => x"ff0614b4",
          7966 => x"11337088",
          7967 => x"2b780779",
          7968 => x"81067184",
          7969 => x"2a5c5258",
          7970 => x"51537280",
          7971 => x"e238759f",
          7972 => x"ff065880",
          7973 => x"da397688",
          7974 => x"2aa41508",
          7975 => x"05527351",
          7976 => x"fcbd3f82",
          7977 => x"bbdc0880",
          7978 => x"c6387610",
          7979 => x"83fe0674",
          7980 => x"05b40551",
          7981 => x"f98d3f82",
          7982 => x"bbdc0883",
          7983 => x"ffff0658",
          7984 => x"ae397687",
          7985 => x"2aa41508",
          7986 => x"05527351",
          7987 => x"fc913f82",
          7988 => x"bbdc089b",
          7989 => x"3876822b",
          7990 => x"83fc0674",
          7991 => x"05b40551",
          7992 => x"f8f83f82",
          7993 => x"bbdc08f0",
          7994 => x"0a065883",
          7995 => x"39815877",
          7996 => x"82bbdc0c",
          7997 => x"893d0d04",
          7998 => x"f83d0d7a",
          7999 => x"7c7e5a58",
          8000 => x"56825981",
          8001 => x"7727829e",
          8002 => x"38769817",
          8003 => x"08278296",
          8004 => x"38753353",
          8005 => x"72792e81",
          8006 => x"9d387279",
          8007 => x"24893872",
          8008 => x"812e8d38",
          8009 => x"82803972",
          8010 => x"832e81b8",
          8011 => x"3881f739",
          8012 => x"76812a17",
          8013 => x"70892aa4",
          8014 => x"18080553",
          8015 => x"765255fb",
          8016 => x"9e3f82bb",
          8017 => x"dc085982",
          8018 => x"bbdc0881",
          8019 => x"d9387483",
          8020 => x"ff0616b4",
          8021 => x"05811678",
          8022 => x"81065956",
          8023 => x"54775376",
          8024 => x"802e8f38",
          8025 => x"77842b9f",
          8026 => x"f0067433",
          8027 => x"8f067107",
          8028 => x"51537274",
          8029 => x"34810b83",
          8030 => x"17347489",
          8031 => x"2aa41708",
          8032 => x"05527551",
          8033 => x"fad93f82",
          8034 => x"bbdc0859",
          8035 => x"82bbdc08",
          8036 => x"81943874",
          8037 => x"83ff0616",
          8038 => x"b4057884",
          8039 => x"2a545476",
          8040 => x"8f387788",
          8041 => x"2a743381",
          8042 => x"f006718f",
          8043 => x"06075153",
          8044 => x"72743480",
          8045 => x"ec397688",
          8046 => x"2aa41708",
          8047 => x"05527551",
          8048 => x"fa9d3f82",
          8049 => x"bbdc0859",
          8050 => x"82bbdc08",
          8051 => x"80d83877",
          8052 => x"83ffff06",
          8053 => x"52761083",
          8054 => x"fe067605",
          8055 => x"b40551f7",
          8056 => x"a43fbe39",
          8057 => x"76872aa4",
          8058 => x"17080552",
          8059 => x"7551f9ef",
          8060 => x"3f82bbdc",
          8061 => x"085982bb",
          8062 => x"dc08ab38",
          8063 => x"77f00a06",
          8064 => x"77822b83",
          8065 => x"fc067018",
          8066 => x"b4057054",
          8067 => x"515454f6",
          8068 => x"c93f82bb",
          8069 => x"dc088f0a",
          8070 => x"06740752",
          8071 => x"7251f783",
          8072 => x"3f810b83",
          8073 => x"17347882",
          8074 => x"bbdc0c8a",
          8075 => x"3d0d04f8",
          8076 => x"3d0d7a7c",
          8077 => x"7e720859",
          8078 => x"56565981",
          8079 => x"7527a438",
          8080 => x"74981708",
          8081 => x"279d3873",
          8082 => x"802eaa38",
          8083 => x"ff537352",
          8084 => x"7551fda4",
          8085 => x"3f82bbdc",
          8086 => x"085482bb",
          8087 => x"dc0880f2",
          8088 => x"38933982",
          8089 => x"5480eb39",
          8090 => x"815480e6",
          8091 => x"3982bbdc",
          8092 => x"085480de",
          8093 => x"39745278",
          8094 => x"51fb843f",
          8095 => x"82bbdc08",
          8096 => x"5882bbdc",
          8097 => x"08802e80",
          8098 => x"c73882bb",
          8099 => x"dc08812e",
          8100 => x"d23882bb",
          8101 => x"dc08ff2e",
          8102 => x"cf388053",
          8103 => x"74527551",
          8104 => x"fcd63f82",
          8105 => x"bbdc08c5",
          8106 => x"38981608",
          8107 => x"fe119018",
          8108 => x"08575557",
          8109 => x"74742790",
          8110 => x"38811590",
          8111 => x"170c8416",
          8112 => x"33810754",
          8113 => x"73841734",
          8114 => x"77557678",
          8115 => x"26ffa638",
          8116 => x"80547382",
          8117 => x"bbdc0c8a",
          8118 => x"3d0d04f6",
          8119 => x"3d0d7c7e",
          8120 => x"7108595b",
          8121 => x"5b799538",
          8122 => x"8c170858",
          8123 => x"77802e88",
          8124 => x"38981708",
          8125 => x"7826b238",
          8126 => x"8158ae39",
          8127 => x"79527a51",
          8128 => x"f9fd3f81",
          8129 => x"557482bb",
          8130 => x"dc082782",
          8131 => x"e03882bb",
          8132 => x"dc085582",
          8133 => x"bbdc08ff",
          8134 => x"2e82d238",
          8135 => x"98170882",
          8136 => x"bbdc0826",
          8137 => x"82c73879",
          8138 => x"58901708",
          8139 => x"70565473",
          8140 => x"802e82b9",
          8141 => x"38777a2e",
          8142 => x"09810680",
          8143 => x"e238811a",
          8144 => x"56981708",
          8145 => x"76268338",
          8146 => x"82567552",
          8147 => x"7a51f9af",
          8148 => x"3f805982",
          8149 => x"bbdc0881",
          8150 => x"2e098106",
          8151 => x"863882bb",
          8152 => x"dc085982",
          8153 => x"bbdc0809",
          8154 => x"70307072",
          8155 => x"07802570",
          8156 => x"7c0782bb",
          8157 => x"dc085451",
          8158 => x"51555573",
          8159 => x"81ef3882",
          8160 => x"bbdc0880",
          8161 => x"2e95388c",
          8162 => x"17085481",
          8163 => x"74279038",
          8164 => x"73981808",
          8165 => x"27893873",
          8166 => x"58853975",
          8167 => x"80db3877",
          8168 => x"56811656",
          8169 => x"98170876",
          8170 => x"26893882",
          8171 => x"56757826",
          8172 => x"81ac3875",
          8173 => x"527a51f8",
          8174 => x"c63f82bb",
          8175 => x"dc08802e",
          8176 => x"b8388059",
          8177 => x"82bbdc08",
          8178 => x"812e0981",
          8179 => x"06863882",
          8180 => x"bbdc0859",
          8181 => x"82bbdc08",
          8182 => x"09703070",
          8183 => x"72078025",
          8184 => x"707c0751",
          8185 => x"51555573",
          8186 => x"80f83875",
          8187 => x"782e0981",
          8188 => x"06ffae38",
          8189 => x"735580f5",
          8190 => x"39ff5375",
          8191 => x"527651f9",
          8192 => x"f73f82bb",
          8193 => x"dc0882bb",
          8194 => x"dc083070",
          8195 => x"82bbdc08",
          8196 => x"07802551",
          8197 => x"55557980",
          8198 => x"2e943873",
          8199 => x"802e8f38",
          8200 => x"75537952",
          8201 => x"7651f9d0",
          8202 => x"3f82bbdc",
          8203 => x"085574a5",
          8204 => x"38758c18",
          8205 => x"0c981708",
          8206 => x"fe059018",
          8207 => x"08565474",
          8208 => x"74268638",
          8209 => x"ff159018",
          8210 => x"0c841733",
          8211 => x"81075473",
          8212 => x"84183497",
          8213 => x"39ff5674",
          8214 => x"812e9038",
          8215 => x"8c398055",
          8216 => x"8c3982bb",
          8217 => x"dc085585",
          8218 => x"39815675",
          8219 => x"557482bb",
          8220 => x"dc0c8c3d",
          8221 => x"0d04f83d",
          8222 => x"0d7a7052",
          8223 => x"55f3f03f",
          8224 => x"82bbdc08",
          8225 => x"58815682",
          8226 => x"bbdc0880",
          8227 => x"d8387b52",
          8228 => x"7451f6c1",
          8229 => x"3f82bbdc",
          8230 => x"0882bbdc",
          8231 => x"08b0170c",
          8232 => x"59848053",
          8233 => x"7752b415",
          8234 => x"705257f2",
          8235 => x"c83f7756",
          8236 => x"84398116",
          8237 => x"568a1522",
          8238 => x"58757827",
          8239 => x"97388154",
          8240 => x"75195376",
          8241 => x"52811533",
          8242 => x"51ede93f",
          8243 => x"82bbdc08",
          8244 => x"802edf38",
          8245 => x"8a152276",
          8246 => x"32703070",
          8247 => x"7207709f",
          8248 => x"2a535156",
          8249 => x"567582bb",
          8250 => x"dc0c8a3d",
          8251 => x"0d04f83d",
          8252 => x"0d7a7c71",
          8253 => x"08585657",
          8254 => x"74f0800a",
          8255 => x"2680f138",
          8256 => x"749f0653",
          8257 => x"7280e938",
          8258 => x"7490180c",
          8259 => x"88170854",
          8260 => x"73aa3875",
          8261 => x"33538273",
          8262 => x"278838a8",
          8263 => x"16085473",
          8264 => x"9b387485",
          8265 => x"2a53820b",
          8266 => x"8817225a",
          8267 => x"58727927",
          8268 => x"80fe38a8",
          8269 => x"16089818",
          8270 => x"0c80cd39",
          8271 => x"8a162270",
          8272 => x"892b5458",
          8273 => x"727526b2",
          8274 => x"38735276",
          8275 => x"51f5b03f",
          8276 => x"82bbdc08",
          8277 => x"5482bbdc",
          8278 => x"08ff2ebd",
          8279 => x"38810b82",
          8280 => x"bbdc0827",
          8281 => x"8b389816",
          8282 => x"0882bbdc",
          8283 => x"08268538",
          8284 => x"8258bd39",
          8285 => x"74733155",
          8286 => x"cb397352",
          8287 => x"7551f4d5",
          8288 => x"3f82bbdc",
          8289 => x"0898180c",
          8290 => x"7394180c",
          8291 => x"98170853",
          8292 => x"82587280",
          8293 => x"2e9a3885",
          8294 => x"39815894",
          8295 => x"3974892a",
          8296 => x"1398180c",
          8297 => x"7483ff06",
          8298 => x"16b4059c",
          8299 => x"180c8058",
          8300 => x"7782bbdc",
          8301 => x"0c8a3d0d",
          8302 => x"04f83d0d",
          8303 => x"7a700890",
          8304 => x"1208a005",
          8305 => x"595754f0",
          8306 => x"800a7727",
          8307 => x"8638800b",
          8308 => x"98150c98",
          8309 => x"14085384",
          8310 => x"5572802e",
          8311 => x"81cb3876",
          8312 => x"83ff0658",
          8313 => x"7781b538",
          8314 => x"81139815",
          8315 => x"0c941408",
          8316 => x"55749238",
          8317 => x"76852a88",
          8318 => x"17225653",
          8319 => x"74732681",
          8320 => x"9b3880c0",
          8321 => x"398a1622",
          8322 => x"ff057789",
          8323 => x"2a065372",
          8324 => x"818a3874",
          8325 => x"527351f3",
          8326 => x"e63f82bb",
          8327 => x"dc085382",
          8328 => x"55810b82",
          8329 => x"bbdc0827",
          8330 => x"80ff3881",
          8331 => x"5582bbdc",
          8332 => x"08ff2e80",
          8333 => x"f4389816",
          8334 => x"0882bbdc",
          8335 => x"082680ca",
          8336 => x"387b8a38",
          8337 => x"7798150c",
          8338 => x"845580dd",
          8339 => x"39941408",
          8340 => x"527351f9",
          8341 => x"863f82bb",
          8342 => x"dc085387",
          8343 => x"5582bbdc",
          8344 => x"08802e80",
          8345 => x"c4388255",
          8346 => x"82bbdc08",
          8347 => x"812eba38",
          8348 => x"815582bb",
          8349 => x"dc08ff2e",
          8350 => x"b03882bb",
          8351 => x"dc085275",
          8352 => x"51fbf33f",
          8353 => x"82bbdc08",
          8354 => x"a0387294",
          8355 => x"150c7252",
          8356 => x"7551f2c1",
          8357 => x"3f82bbdc",
          8358 => x"0898150c",
          8359 => x"7690150c",
          8360 => x"7716b405",
          8361 => x"9c150c80",
          8362 => x"557482bb",
          8363 => x"dc0c8a3d",
          8364 => x"0d04f73d",
          8365 => x"0d7b7d71",
          8366 => x"085b5b57",
          8367 => x"80527651",
          8368 => x"fcac3f82",
          8369 => x"bbdc0854",
          8370 => x"82bbdc08",
          8371 => x"80ec3882",
          8372 => x"bbdc0856",
          8373 => x"98170852",
          8374 => x"7851f083",
          8375 => x"3f82bbdc",
          8376 => x"085482bb",
          8377 => x"dc0880d2",
          8378 => x"3882bbdc",
          8379 => x"089c1808",
          8380 => x"70335154",
          8381 => x"587281e5",
          8382 => x"2e098106",
          8383 => x"83388158",
          8384 => x"82bbdc08",
          8385 => x"55728338",
          8386 => x"81557775",
          8387 => x"07537280",
          8388 => x"2e8e3881",
          8389 => x"1656757a",
          8390 => x"2e098106",
          8391 => x"8838a539",
          8392 => x"82bbdc08",
          8393 => x"56815276",
          8394 => x"51fd8e3f",
          8395 => x"82bbdc08",
          8396 => x"5482bbdc",
          8397 => x"08802eff",
          8398 => x"9b387384",
          8399 => x"2e098106",
          8400 => x"83388754",
          8401 => x"7382bbdc",
          8402 => x"0c8b3d0d",
          8403 => x"04fd3d0d",
          8404 => x"769a1152",
          8405 => x"54ebec3f",
          8406 => x"82bbdc08",
          8407 => x"83ffff06",
          8408 => x"76703351",
          8409 => x"53537183",
          8410 => x"2e098106",
          8411 => x"90389414",
          8412 => x"51ebd03f",
          8413 => x"82bbdc08",
          8414 => x"902b7307",
          8415 => x"537282bb",
          8416 => x"dc0c853d",
          8417 => x"0d04fc3d",
          8418 => x"0d777970",
          8419 => x"83ffff06",
          8420 => x"549a1253",
          8421 => x"5555ebed",
          8422 => x"3f767033",
          8423 => x"51537283",
          8424 => x"2e098106",
          8425 => x"8b387390",
          8426 => x"2a529415",
          8427 => x"51ebd63f",
          8428 => x"863d0d04",
          8429 => x"f73d0d7b",
          8430 => x"7d5b5584",
          8431 => x"75085a58",
          8432 => x"98150880",
          8433 => x"2e818a38",
          8434 => x"98150852",
          8435 => x"7851ee8f",
          8436 => x"3f82bbdc",
          8437 => x"085882bb",
          8438 => x"dc0880f5",
          8439 => x"389c1508",
          8440 => x"70335553",
          8441 => x"73863884",
          8442 => x"5880e639",
          8443 => x"8b133370",
          8444 => x"bf067081",
          8445 => x"ff065851",
          8446 => x"53728616",
          8447 => x"3482bbdc",
          8448 => x"08537381",
          8449 => x"e52e8338",
          8450 => x"815373ae",
          8451 => x"2ea93881",
          8452 => x"70740654",
          8453 => x"5772802e",
          8454 => x"9e38758f",
          8455 => x"2e993882",
          8456 => x"bbdc0876",
          8457 => x"df065454",
          8458 => x"72882e09",
          8459 => x"81068338",
          8460 => x"7654737a",
          8461 => x"2ea03880",
          8462 => x"527451fa",
          8463 => x"fc3f82bb",
          8464 => x"dc085882",
          8465 => x"bbdc0889",
          8466 => x"38981508",
          8467 => x"fefa3886",
          8468 => x"39800b98",
          8469 => x"160c7782",
          8470 => x"bbdc0c8b",
          8471 => x"3d0d04fb",
          8472 => x"3d0d7770",
          8473 => x"08575481",
          8474 => x"527351fc",
          8475 => x"c53f82bb",
          8476 => x"dc085582",
          8477 => x"bbdc08b4",
          8478 => x"38981408",
          8479 => x"527551ec",
          8480 => x"de3f82bb",
          8481 => x"dc085582",
          8482 => x"bbdc08a0",
          8483 => x"38a05382",
          8484 => x"bbdc0852",
          8485 => x"9c140851",
          8486 => x"eadb3f8b",
          8487 => x"53a01452",
          8488 => x"9c140851",
          8489 => x"eaac3f81",
          8490 => x"0b831734",
          8491 => x"7482bbdc",
          8492 => x"0c873d0d",
          8493 => x"04fd3d0d",
          8494 => x"75700898",
          8495 => x"12085470",
          8496 => x"535553ec",
          8497 => x"9a3f82bb",
          8498 => x"dc088d38",
          8499 => x"9c130853",
          8500 => x"e5733481",
          8501 => x"0b831534",
          8502 => x"853d0d04",
          8503 => x"fa3d0d78",
          8504 => x"7a575780",
          8505 => x"0b891734",
          8506 => x"98170880",
          8507 => x"2e818238",
          8508 => x"80708918",
          8509 => x"5555559c",
          8510 => x"17081470",
          8511 => x"33811656",
          8512 => x"515271a0",
          8513 => x"2ea83871",
          8514 => x"852e0981",
          8515 => x"06843881",
          8516 => x"e5527389",
          8517 => x"2e098106",
          8518 => x"8b38ae73",
          8519 => x"70810555",
          8520 => x"34811555",
          8521 => x"71737081",
          8522 => x"05553481",
          8523 => x"15558a74",
          8524 => x"27c53875",
          8525 => x"15880552",
          8526 => x"800b8113",
          8527 => x"349c1708",
          8528 => x"528b1233",
          8529 => x"8817349c",
          8530 => x"17089c11",
          8531 => x"5252e88a",
          8532 => x"3f82bbdc",
          8533 => x"08760c96",
          8534 => x"1251e7e7",
          8535 => x"3f82bbdc",
          8536 => x"08861723",
          8537 => x"981251e7",
          8538 => x"da3f82bb",
          8539 => x"dc088417",
          8540 => x"23883d0d",
          8541 => x"04f33d0d",
          8542 => x"7f70085e",
          8543 => x"5b806170",
          8544 => x"33515555",
          8545 => x"73af2e83",
          8546 => x"38815573",
          8547 => x"80dc2e91",
          8548 => x"3874802e",
          8549 => x"8c38941d",
          8550 => x"08881c0c",
          8551 => x"aa398115",
          8552 => x"41806170",
          8553 => x"33565656",
          8554 => x"73af2e09",
          8555 => x"81068338",
          8556 => x"81567380",
          8557 => x"dc327030",
          8558 => x"70802578",
          8559 => x"07515154",
          8560 => x"73dc3873",
          8561 => x"881c0c60",
          8562 => x"70335154",
          8563 => x"739f2696",
          8564 => x"38ff800b",
          8565 => x"ab1c3480",
          8566 => x"527a51f6",
          8567 => x"913f82bb",
          8568 => x"dc085585",
          8569 => x"9839913d",
          8570 => x"61a01d5c",
          8571 => x"5a5e8b53",
          8572 => x"a0527951",
          8573 => x"e7ff3f80",
          8574 => x"70595788",
          8575 => x"7933555c",
          8576 => x"73ae2e09",
          8577 => x"810680d4",
          8578 => x"38781870",
          8579 => x"33811a71",
          8580 => x"ae327030",
          8581 => x"709f2a73",
          8582 => x"82260751",
          8583 => x"51535a57",
          8584 => x"54738c38",
          8585 => x"79175475",
          8586 => x"74348117",
          8587 => x"57db3975",
          8588 => x"af327030",
          8589 => x"709f2a51",
          8590 => x"51547580",
          8591 => x"dc2e8c38",
          8592 => x"73802e87",
          8593 => x"3875a026",
          8594 => x"82bd3877",
          8595 => x"197e0ca4",
          8596 => x"54a07627",
          8597 => x"82bd38a0",
          8598 => x"5482b839",
          8599 => x"78187033",
          8600 => x"811a5a57",
          8601 => x"54a07627",
          8602 => x"81fc3875",
          8603 => x"af327030",
          8604 => x"7780dc32",
          8605 => x"70307280",
          8606 => x"25718025",
          8607 => x"07515156",
          8608 => x"51557380",
          8609 => x"2eac3884",
          8610 => x"39811858",
          8611 => x"80781a70",
          8612 => x"33515555",
          8613 => x"73af2e09",
          8614 => x"81068338",
          8615 => x"81557380",
          8616 => x"dc327030",
          8617 => x"70802577",
          8618 => x"07515154",
          8619 => x"73db3881",
          8620 => x"b53975ae",
          8621 => x"2e098106",
          8622 => x"83388154",
          8623 => x"767c2774",
          8624 => x"07547380",
          8625 => x"2ea2387b",
          8626 => x"8b327030",
          8627 => x"77ae3270",
          8628 => x"30728025",
          8629 => x"719f2a07",
          8630 => x"53515651",
          8631 => x"557481a7",
          8632 => x"3888578b",
          8633 => x"5cfef539",
          8634 => x"75982b54",
          8635 => x"7380258c",
          8636 => x"387580ff",
          8637 => x"0682b5a4",
          8638 => x"11335754",
          8639 => x"7551e6e1",
          8640 => x"3f82bbdc",
          8641 => x"08802eb2",
          8642 => x"38781870",
          8643 => x"33811a71",
          8644 => x"545a5654",
          8645 => x"e6d23f82",
          8646 => x"bbdc0880",
          8647 => x"2e80e838",
          8648 => x"ff1c5476",
          8649 => x"742780df",
          8650 => x"38791754",
          8651 => x"75743481",
          8652 => x"177a1155",
          8653 => x"57747434",
          8654 => x"a7397552",
          8655 => x"82b4c451",
          8656 => x"e5fe3f82",
          8657 => x"bbdc08bf",
          8658 => x"38ff9f16",
          8659 => x"54739926",
          8660 => x"8938e016",
          8661 => x"7081ff06",
          8662 => x"57547917",
          8663 => x"54757434",
          8664 => x"811757fd",
          8665 => x"f7397719",
          8666 => x"7e0c7680",
          8667 => x"2e993879",
          8668 => x"33547381",
          8669 => x"e52e0981",
          8670 => x"06843885",
          8671 => x"7a348454",
          8672 => x"a076278f",
          8673 => x"388b3986",
          8674 => x"5581f239",
          8675 => x"845680f3",
          8676 => x"39805473",
          8677 => x"8b1b3480",
          8678 => x"7b085852",
          8679 => x"7a51f2ce",
          8680 => x"3f82bbdc",
          8681 => x"085682bb",
          8682 => x"dc0880d7",
          8683 => x"38981b08",
          8684 => x"527651e6",
          8685 => x"aa3f82bb",
          8686 => x"dc085682",
          8687 => x"bbdc0880",
          8688 => x"c2389c1b",
          8689 => x"08703355",
          8690 => x"5573802e",
          8691 => x"ffbe388b",
          8692 => x"1533bf06",
          8693 => x"5473861c",
          8694 => x"348b1533",
          8695 => x"70832a70",
          8696 => x"81065155",
          8697 => x"58739238",
          8698 => x"8b537952",
          8699 => x"7451e49f",
          8700 => x"3f82bbdc",
          8701 => x"08802e8b",
          8702 => x"3875527a",
          8703 => x"51f3ba3f",
          8704 => x"ff9f3975",
          8705 => x"ab1c3357",
          8706 => x"5574802e",
          8707 => x"bb387484",
          8708 => x"2e098106",
          8709 => x"80e73875",
          8710 => x"852a7081",
          8711 => x"0677822a",
          8712 => x"58515473",
          8713 => x"802e9638",
          8714 => x"75810654",
          8715 => x"73802efb",
          8716 => x"b538ff80",
          8717 => x"0bab1c34",
          8718 => x"805580c1",
          8719 => x"39758106",
          8720 => x"5473ba38",
          8721 => x"8555b639",
          8722 => x"75822a70",
          8723 => x"81065154",
          8724 => x"73ab3886",
          8725 => x"1b337084",
          8726 => x"2a708106",
          8727 => x"51555573",
          8728 => x"802ee138",
          8729 => x"901b0883",
          8730 => x"ff061db4",
          8731 => x"05527c51",
          8732 => x"f5db3f82",
          8733 => x"bbdc0888",
          8734 => x"1c0cfaea",
          8735 => x"397482bb",
          8736 => x"dc0c8f3d",
          8737 => x"0d04f63d",
          8738 => x"0d7c5bff",
          8739 => x"7b087071",
          8740 => x"7355595c",
          8741 => x"55597380",
          8742 => x"2e81c638",
          8743 => x"75708105",
          8744 => x"573370a0",
          8745 => x"26525271",
          8746 => x"ba2e8d38",
          8747 => x"70ee3871",
          8748 => x"ba2e0981",
          8749 => x"0681a538",
          8750 => x"7333d011",
          8751 => x"7081ff06",
          8752 => x"51525370",
          8753 => x"89269138",
          8754 => x"82147381",
          8755 => x"ff06d005",
          8756 => x"56527176",
          8757 => x"2e80f738",
          8758 => x"800b82b5",
          8759 => x"94595577",
          8760 => x"087a5557",
          8761 => x"76708105",
          8762 => x"58337470",
          8763 => x"81055633",
          8764 => x"ff9f1253",
          8765 => x"53537099",
          8766 => x"268938e0",
          8767 => x"137081ff",
          8768 => x"065451ff",
          8769 => x"9f125170",
          8770 => x"99268938",
          8771 => x"e0127081",
          8772 => x"ff065351",
          8773 => x"7230709f",
          8774 => x"2a515172",
          8775 => x"722e0981",
          8776 => x"06853870",
          8777 => x"ffbe3872",
          8778 => x"30747732",
          8779 => x"70307072",
          8780 => x"079f2a73",
          8781 => x"9f2a0753",
          8782 => x"54545170",
          8783 => x"802e8f38",
          8784 => x"81158419",
          8785 => x"59558375",
          8786 => x"25ff9438",
          8787 => x"8b397483",
          8788 => x"24863874",
          8789 => x"767c0c59",
          8790 => x"78518639",
          8791 => x"82d3a833",
          8792 => x"517082bb",
          8793 => x"dc0c8c3d",
          8794 => x"0d04fa3d",
          8795 => x"0d785680",
          8796 => x"0b831734",
          8797 => x"ff0bb017",
          8798 => x"0c795275",
          8799 => x"51e2e03f",
          8800 => x"845582bb",
          8801 => x"dc088180",
          8802 => x"3884b216",
          8803 => x"51dfb43f",
          8804 => x"82bbdc08",
          8805 => x"83ffff06",
          8806 => x"54835573",
          8807 => x"82d4d52e",
          8808 => x"09810680",
          8809 => x"e338800b",
          8810 => x"b4173356",
          8811 => x"577481e9",
          8812 => x"2e098106",
          8813 => x"83388157",
          8814 => x"7481eb32",
          8815 => x"70307080",
          8816 => x"25790751",
          8817 => x"5154738a",
          8818 => x"387481e8",
          8819 => x"2e098106",
          8820 => x"b5388353",
          8821 => x"82b4d452",
          8822 => x"80ea1651",
          8823 => x"e0b13f82",
          8824 => x"bbdc0855",
          8825 => x"82bbdc08",
          8826 => x"802e9d38",
          8827 => x"855382b4",
          8828 => x"d8528186",
          8829 => x"1651e097",
          8830 => x"3f82bbdc",
          8831 => x"085582bb",
          8832 => x"dc08802e",
          8833 => x"83388255",
          8834 => x"7482bbdc",
          8835 => x"0c883d0d",
          8836 => x"04f23d0d",
          8837 => x"61028405",
          8838 => x"80cb0533",
          8839 => x"58558075",
          8840 => x"0c6051fc",
          8841 => x"e13f82bb",
          8842 => x"dc08588b",
          8843 => x"56800b82",
          8844 => x"bbdc0824",
          8845 => x"86fc3882",
          8846 => x"bbdc0884",
          8847 => x"2982d394",
          8848 => x"05700855",
          8849 => x"538c5673",
          8850 => x"802e86e6",
          8851 => x"3873750c",
          8852 => x"7681fe06",
          8853 => x"74335457",
          8854 => x"72802eae",
          8855 => x"38811433",
          8856 => x"51d7ca3f",
          8857 => x"82bbdc08",
          8858 => x"81ff0670",
          8859 => x"81065455",
          8860 => x"72983876",
          8861 => x"802e86b8",
          8862 => x"3874822a",
          8863 => x"70810651",
          8864 => x"538a5672",
          8865 => x"86ac3886",
          8866 => x"a7398074",
          8867 => x"34778115",
          8868 => x"34815281",
          8869 => x"143351d7",
          8870 => x"b23f82bb",
          8871 => x"dc0881ff",
          8872 => x"06708106",
          8873 => x"54558356",
          8874 => x"72868738",
          8875 => x"76802e8f",
          8876 => x"3874822a",
          8877 => x"70810651",
          8878 => x"538a5672",
          8879 => x"85f43880",
          8880 => x"70537452",
          8881 => x"5bfda33f",
          8882 => x"82bbdc08",
          8883 => x"81ff0657",
          8884 => x"76822e09",
          8885 => x"810680e2",
          8886 => x"388c3d74",
          8887 => x"56588356",
          8888 => x"83f61533",
          8889 => x"70585372",
          8890 => x"802e8d38",
          8891 => x"83fa1551",
          8892 => x"dce83f82",
          8893 => x"bbdc0857",
          8894 => x"76787084",
          8895 => x"055a0cff",
          8896 => x"16901656",
          8897 => x"56758025",
          8898 => x"d738800b",
          8899 => x"8d3d5456",
          8900 => x"72708405",
          8901 => x"54085b83",
          8902 => x"577a802e",
          8903 => x"95387a52",
          8904 => x"7351fcc6",
          8905 => x"3f82bbdc",
          8906 => x"0881ff06",
          8907 => x"57817727",
          8908 => x"89388116",
          8909 => x"56837627",
          8910 => x"d7388156",
          8911 => x"76842e84",
          8912 => x"f1388d56",
          8913 => x"76812684",
          8914 => x"e938bf14",
          8915 => x"51dbf43f",
          8916 => x"82bbdc08",
          8917 => x"83ffff06",
          8918 => x"53728480",
          8919 => x"2e098106",
          8920 => x"84d03880",
          8921 => x"ca1451db",
          8922 => x"da3f82bb",
          8923 => x"dc0883ff",
          8924 => x"ff065877",
          8925 => x"8d3880d8",
          8926 => x"1451dbde",
          8927 => x"3f82bbdc",
          8928 => x"0858779c",
          8929 => x"150c80c4",
          8930 => x"14338215",
          8931 => x"3480c414",
          8932 => x"33ff1170",
          8933 => x"81ff0651",
          8934 => x"54558d56",
          8935 => x"72812684",
          8936 => x"91387481",
          8937 => x"ff067871",
          8938 => x"2980c116",
          8939 => x"33525953",
          8940 => x"728a1523",
          8941 => x"72802e8b",
          8942 => x"38ff1373",
          8943 => x"06537280",
          8944 => x"2e86388d",
          8945 => x"5683eb39",
          8946 => x"80c51451",
          8947 => x"daf53f82",
          8948 => x"bbdc0853",
          8949 => x"82bbdc08",
          8950 => x"88152372",
          8951 => x"8f06578d",
          8952 => x"567683ce",
          8953 => x"3880c714",
          8954 => x"51dad83f",
          8955 => x"82bbdc08",
          8956 => x"83ffff06",
          8957 => x"55748d38",
          8958 => x"80d41451",
          8959 => x"dadc3f82",
          8960 => x"bbdc0855",
          8961 => x"80c21451",
          8962 => x"dab93f82",
          8963 => x"bbdc0883",
          8964 => x"ffff0653",
          8965 => x"8d567280",
          8966 => x"2e839738",
          8967 => x"88142278",
          8968 => x"1471842a",
          8969 => x"055a5a78",
          8970 => x"75268386",
          8971 => x"388a1422",
          8972 => x"52747931",
          8973 => x"51feeecb",
          8974 => x"3f82bbdc",
          8975 => x"085582bb",
          8976 => x"dc08802e",
          8977 => x"82ec3882",
          8978 => x"bbdc0880",
          8979 => x"fffffff5",
          8980 => x"26833883",
          8981 => x"577483ff",
          8982 => x"f5268338",
          8983 => x"8257749f",
          8984 => x"f5268538",
          8985 => x"81578939",
          8986 => x"8d567680",
          8987 => x"2e82c338",
          8988 => x"82157098",
          8989 => x"160c7ba0",
          8990 => x"160c731c",
          8991 => x"70a4170c",
          8992 => x"7a1dac17",
          8993 => x"0c545576",
          8994 => x"832e0981",
          8995 => x"06af3880",
          8996 => x"de1451d9",
          8997 => x"ae3f82bb",
          8998 => x"dc0883ff",
          8999 => x"ff06538d",
          9000 => x"5672828e",
          9001 => x"3879828a",
          9002 => x"3880e014",
          9003 => x"51d9ab3f",
          9004 => x"82bbdc08",
          9005 => x"a8150c74",
          9006 => x"822b53a2",
          9007 => x"398d5679",
          9008 => x"802e81ee",
          9009 => x"387713a8",
          9010 => x"150c7415",
          9011 => x"5376822e",
          9012 => x"8d387410",
          9013 => x"1570812a",
          9014 => x"76810605",
          9015 => x"515383ff",
          9016 => x"13892a53",
          9017 => x"8d56729c",
          9018 => x"15082681",
          9019 => x"c538ff0b",
          9020 => x"90150cff",
          9021 => x"0b8c150c",
          9022 => x"ff800b84",
          9023 => x"15347683",
          9024 => x"2e098106",
          9025 => x"81923880",
          9026 => x"e41451d8",
          9027 => x"b63f82bb",
          9028 => x"dc0883ff",
          9029 => x"ff065372",
          9030 => x"812e0981",
          9031 => x"0680f938",
          9032 => x"811b5273",
          9033 => x"51dbb83f",
          9034 => x"82bbdc08",
          9035 => x"80ea3882",
          9036 => x"bbdc0884",
          9037 => x"153484b2",
          9038 => x"1451d887",
          9039 => x"3f82bbdc",
          9040 => x"0883ffff",
          9041 => x"06537282",
          9042 => x"d4d52e09",
          9043 => x"810680c8",
          9044 => x"38b41451",
          9045 => x"d8843f82",
          9046 => x"bbdc0884",
          9047 => x"8b85a4d2",
          9048 => x"2e098106",
          9049 => x"b3388498",
          9050 => x"1451d7ee",
          9051 => x"3f82bbdc",
          9052 => x"08868a85",
          9053 => x"e4f22e09",
          9054 => x"81069d38",
          9055 => x"849c1451",
          9056 => x"d7d83f82",
          9057 => x"bbdc0890",
          9058 => x"150c84a0",
          9059 => x"1451d7ca",
          9060 => x"3f82bbdc",
          9061 => x"088c150c",
          9062 => x"76743482",
          9063 => x"d3a42281",
          9064 => x"05537282",
          9065 => x"d3a42372",
          9066 => x"86152380",
          9067 => x"0b94150c",
          9068 => x"80567582",
          9069 => x"bbdc0c90",
          9070 => x"3d0d04fb",
          9071 => x"3d0d7754",
          9072 => x"89557380",
          9073 => x"2eb93873",
          9074 => x"08537280",
          9075 => x"2eb13872",
          9076 => x"33527180",
          9077 => x"2ea93886",
          9078 => x"13228415",
          9079 => x"22575271",
          9080 => x"762e0981",
          9081 => x"06993881",
          9082 => x"133351d0",
          9083 => x"c03f82bb",
          9084 => x"dc088106",
          9085 => x"52718838",
          9086 => x"71740854",
          9087 => x"55833980",
          9088 => x"53787371",
          9089 => x"0c527482",
          9090 => x"bbdc0c87",
          9091 => x"3d0d04fa",
          9092 => x"3d0d02ab",
          9093 => x"05337a58",
          9094 => x"893dfc05",
          9095 => x"5256f4e6",
          9096 => x"3f8b5480",
          9097 => x"0b82bbdc",
          9098 => x"0824bc38",
          9099 => x"82bbdc08",
          9100 => x"842982d3",
          9101 => x"94057008",
          9102 => x"55557380",
          9103 => x"2e843880",
          9104 => x"74347854",
          9105 => x"73802e84",
          9106 => x"38807434",
          9107 => x"78750c75",
          9108 => x"5475802e",
          9109 => x"92388053",
          9110 => x"893d7053",
          9111 => x"840551f7",
          9112 => x"b03f82bb",
          9113 => x"dc085473",
          9114 => x"82bbdc0c",
          9115 => x"883d0d04",
          9116 => x"eb3d0d67",
          9117 => x"02840580",
          9118 => x"e7053359",
          9119 => x"59895478",
          9120 => x"802e84c8",
          9121 => x"3877bf06",
          9122 => x"7054983d",
          9123 => x"d0055399",
          9124 => x"3d840552",
          9125 => x"58f6fa3f",
          9126 => x"82bbdc08",
          9127 => x"5582bbdc",
          9128 => x"0884a438",
          9129 => x"7a5c6852",
          9130 => x"8c3d7052",
          9131 => x"56edc63f",
          9132 => x"82bbdc08",
          9133 => x"5582bbdc",
          9134 => x"08923802",
          9135 => x"80d70533",
          9136 => x"70982b55",
          9137 => x"57738025",
          9138 => x"83388655",
          9139 => x"779c0654",
          9140 => x"73802e81",
          9141 => x"ab387480",
          9142 => x"2e953874",
          9143 => x"842e0981",
          9144 => x"06aa3875",
          9145 => x"51eaf83f",
          9146 => x"82bbdc08",
          9147 => x"559e3902",
          9148 => x"b2053391",
          9149 => x"06547381",
          9150 => x"b8387782",
          9151 => x"2a708106",
          9152 => x"51547380",
          9153 => x"2e8e3888",
          9154 => x"5583bc39",
          9155 => x"77880758",
          9156 => x"7483b438",
          9157 => x"77832a70",
          9158 => x"81065154",
          9159 => x"73802e81",
          9160 => x"af386252",
          9161 => x"7a51e8a5",
          9162 => x"3f82bbdc",
          9163 => x"08568288",
          9164 => x"b20a5262",
          9165 => x"8e0551d4",
          9166 => x"ea3f6254",
          9167 => x"a00b8b15",
          9168 => x"34805362",
          9169 => x"527a51e8",
          9170 => x"bd3f8052",
          9171 => x"629c0551",
          9172 => x"d4d13f7a",
          9173 => x"54810b83",
          9174 => x"15347580",
          9175 => x"2e80f138",
          9176 => x"7ab01108",
          9177 => x"51548053",
          9178 => x"7552973d",
          9179 => x"d40551dd",
          9180 => x"be3f82bb",
          9181 => x"dc085582",
          9182 => x"bbdc0882",
          9183 => x"ca38b739",
          9184 => x"7482c438",
          9185 => x"02b20533",
          9186 => x"70842a70",
          9187 => x"81065155",
          9188 => x"5673802e",
          9189 => x"86388455",
          9190 => x"82ad3977",
          9191 => x"812a7081",
          9192 => x"06515473",
          9193 => x"802ea938",
          9194 => x"75810654",
          9195 => x"73802ea0",
          9196 => x"38875582",
          9197 => x"92397352",
          9198 => x"7a51d6a3",
          9199 => x"3f82bbdc",
          9200 => x"087bff18",
          9201 => x"8c120c55",
          9202 => x"5582bbdc",
          9203 => x"0881f838",
          9204 => x"77832a70",
          9205 => x"81065154",
          9206 => x"73802e86",
          9207 => x"387780c0",
          9208 => x"07587ab0",
          9209 => x"1108a01b",
          9210 => x"0c63a41b",
          9211 => x"0c635370",
          9212 => x"5257e6d9",
          9213 => x"3f82bbdc",
          9214 => x"0882bbdc",
          9215 => x"08881b0c",
          9216 => x"639c0552",
          9217 => x"5ad2d33f",
          9218 => x"82bbdc08",
          9219 => x"82bbdc08",
          9220 => x"8c1b0c77",
          9221 => x"7a0c5686",
          9222 => x"1722841a",
          9223 => x"2377901a",
          9224 => x"34800b91",
          9225 => x"1a34800b",
          9226 => x"9c1a0c80",
          9227 => x"0b941a0c",
          9228 => x"77852a70",
          9229 => x"81065154",
          9230 => x"73802e81",
          9231 => x"8d3882bb",
          9232 => x"dc08802e",
          9233 => x"81843882",
          9234 => x"bbdc0894",
          9235 => x"1a0c8a17",
          9236 => x"2270892b",
          9237 => x"7b525957",
          9238 => x"a8397652",
          9239 => x"7851d79f",
          9240 => x"3f82bbdc",
          9241 => x"085782bb",
          9242 => x"dc088126",
          9243 => x"83388255",
          9244 => x"82bbdc08",
          9245 => x"ff2e0981",
          9246 => x"06833879",
          9247 => x"55757831",
          9248 => x"56743070",
          9249 => x"76078025",
          9250 => x"51547776",
          9251 => x"278a3881",
          9252 => x"70750655",
          9253 => x"5a73c338",
          9254 => x"76981a0c",
          9255 => x"74a93875",
          9256 => x"83ff0654",
          9257 => x"73802ea2",
          9258 => x"3876527a",
          9259 => x"51d6a63f",
          9260 => x"82bbdc08",
          9261 => x"85388255",
          9262 => x"8e397589",
          9263 => x"2a82bbdc",
          9264 => x"08059c1a",
          9265 => x"0c843980",
          9266 => x"790c7454",
          9267 => x"7382bbdc",
          9268 => x"0c973d0d",
          9269 => x"04f23d0d",
          9270 => x"60636564",
          9271 => x"40405d59",
          9272 => x"807e0c90",
          9273 => x"3dfc0552",
          9274 => x"7851f9cf",
          9275 => x"3f82bbdc",
          9276 => x"085582bb",
          9277 => x"dc088a38",
          9278 => x"91193355",
          9279 => x"74802e86",
          9280 => x"38745682",
          9281 => x"c4399019",
          9282 => x"33810655",
          9283 => x"87567480",
          9284 => x"2e82b638",
          9285 => x"9539820b",
          9286 => x"911a3482",
          9287 => x"5682aa39",
          9288 => x"810b911a",
          9289 => x"34815682",
          9290 => x"a0398c19",
          9291 => x"08941a08",
          9292 => x"3155747c",
          9293 => x"27833874",
          9294 => x"5c7b802e",
          9295 => x"82893894",
          9296 => x"19087083",
          9297 => x"ff065656",
          9298 => x"7481b238",
          9299 => x"7e8a1122",
          9300 => x"ff057789",
          9301 => x"2a065b55",
          9302 => x"79a83875",
          9303 => x"87388819",
          9304 => x"08558f39",
          9305 => x"98190852",
          9306 => x"7851d593",
          9307 => x"3f82bbdc",
          9308 => x"08558175",
          9309 => x"27ff9f38",
          9310 => x"74ff2eff",
          9311 => x"a3387498",
          9312 => x"1a0c9819",
          9313 => x"08527e51",
          9314 => x"d4cb3f82",
          9315 => x"bbdc0880",
          9316 => x"2eff8338",
          9317 => x"82bbdc08",
          9318 => x"1a7c892a",
          9319 => x"59577780",
          9320 => x"2e80d638",
          9321 => x"771a7f8a",
          9322 => x"1122585c",
          9323 => x"55757527",
          9324 => x"8538757a",
          9325 => x"31587754",
          9326 => x"76537c52",
          9327 => x"811b3351",
          9328 => x"ca883f82",
          9329 => x"bbdc08fe",
          9330 => x"d7387e83",
          9331 => x"11335656",
          9332 => x"74802e9f",
          9333 => x"38b01608",
          9334 => x"77315574",
          9335 => x"78279438",
          9336 => x"848053b4",
          9337 => x"1652b016",
          9338 => x"08773189",
          9339 => x"2b7d0551",
          9340 => x"cfe03f77",
          9341 => x"892b56b9",
          9342 => x"39769c1a",
          9343 => x"0c941908",
          9344 => x"83ff0684",
          9345 => x"80713157",
          9346 => x"557b7627",
          9347 => x"83387b56",
          9348 => x"9c190852",
          9349 => x"7e51d1c7",
          9350 => x"3f82bbdc",
          9351 => x"08fe8138",
          9352 => x"75539419",
          9353 => x"0883ff06",
          9354 => x"1fb40552",
          9355 => x"7c51cfa2",
          9356 => x"3f7b7631",
          9357 => x"7e08177f",
          9358 => x"0c761e94",
          9359 => x"1b081894",
          9360 => x"1c0c5e5c",
          9361 => x"fdf33980",
          9362 => x"567582bb",
          9363 => x"dc0c903d",
          9364 => x"0d04f23d",
          9365 => x"0d606365",
          9366 => x"6440405d",
          9367 => x"58807e0c",
          9368 => x"903dfc05",
          9369 => x"527751f6",
          9370 => x"d23f82bb",
          9371 => x"dc085582",
          9372 => x"bbdc088a",
          9373 => x"38911833",
          9374 => x"5574802e",
          9375 => x"86387456",
          9376 => x"83b83990",
          9377 => x"18337081",
          9378 => x"2a708106",
          9379 => x"51565687",
          9380 => x"5674802e",
          9381 => x"83a43895",
          9382 => x"39820b91",
          9383 => x"19348256",
          9384 => x"83983981",
          9385 => x"0b911934",
          9386 => x"8156838e",
          9387 => x"39941808",
          9388 => x"7c115656",
          9389 => x"74762784",
          9390 => x"3875095c",
          9391 => x"7b802e82",
          9392 => x"ec389418",
          9393 => x"087083ff",
          9394 => x"06565674",
          9395 => x"81fd387e",
          9396 => x"8a1122ff",
          9397 => x"0577892a",
          9398 => x"065c557a",
          9399 => x"bf38758c",
          9400 => x"38881808",
          9401 => x"55749c38",
          9402 => x"7a528539",
          9403 => x"98180852",
          9404 => x"7751d7e7",
          9405 => x"3f82bbdc",
          9406 => x"085582bb",
          9407 => x"dc08802e",
          9408 => x"82ab3874",
          9409 => x"812eff91",
          9410 => x"3874ff2e",
          9411 => x"ff953874",
          9412 => x"98190c88",
          9413 => x"18088538",
          9414 => x"7488190c",
          9415 => x"7e55b015",
          9416 => x"089c1908",
          9417 => x"2e098106",
          9418 => x"8d387451",
          9419 => x"cec13f82",
          9420 => x"bbdc08fe",
          9421 => x"ee389818",
          9422 => x"08527e51",
          9423 => x"d1973f82",
          9424 => x"bbdc0880",
          9425 => x"2efed238",
          9426 => x"82bbdc08",
          9427 => x"1b7c892a",
          9428 => x"5a577880",
          9429 => x"2e80d538",
          9430 => x"781b7f8a",
          9431 => x"1122585b",
          9432 => x"55757527",
          9433 => x"8538757b",
          9434 => x"31597854",
          9435 => x"76537c52",
          9436 => x"811a3351",
          9437 => x"c8be3f82",
          9438 => x"bbdc08fe",
          9439 => x"a6387eb0",
          9440 => x"11087831",
          9441 => x"56567479",
          9442 => x"279b3884",
          9443 => x"8053b016",
          9444 => x"08773189",
          9445 => x"2b7d0552",
          9446 => x"b41651cc",
          9447 => x"b53f7e55",
          9448 => x"800b8316",
          9449 => x"3478892b",
          9450 => x"5680db39",
          9451 => x"8c180894",
          9452 => x"19082693",
          9453 => x"387e51cd",
          9454 => x"b63f82bb",
          9455 => x"dc08fde3",
          9456 => x"387e77b0",
          9457 => x"120c5576",
          9458 => x"9c190c94",
          9459 => x"180883ff",
          9460 => x"06848071",
          9461 => x"3157557b",
          9462 => x"76278338",
          9463 => x"7b569c18",
          9464 => x"08527e51",
          9465 => x"cdf93f82",
          9466 => x"bbdc08fd",
          9467 => x"b6387553",
          9468 => x"7c529418",
          9469 => x"0883ff06",
          9470 => x"1fb40551",
          9471 => x"cbd43f7e",
          9472 => x"55810b83",
          9473 => x"16347b76",
          9474 => x"317e0817",
          9475 => x"7f0c761e",
          9476 => x"941a0818",
          9477 => x"70941c0c",
          9478 => x"8c1b0858",
          9479 => x"585e5c74",
          9480 => x"76278338",
          9481 => x"7555748c",
          9482 => x"190cfd90",
          9483 => x"39901833",
          9484 => x"80c00755",
          9485 => x"74901934",
          9486 => x"80567582",
          9487 => x"bbdc0c90",
          9488 => x"3d0d04f8",
          9489 => x"3d0d7a8b",
          9490 => x"3dfc0553",
          9491 => x"705256f2",
          9492 => x"ea3f82bb",
          9493 => x"dc085782",
          9494 => x"bbdc0880",
          9495 => x"fb389016",
          9496 => x"3370862a",
          9497 => x"70810651",
          9498 => x"55557380",
          9499 => x"2e80e938",
          9500 => x"a0160852",
          9501 => x"7851cce7",
          9502 => x"3f82bbdc",
          9503 => x"085782bb",
          9504 => x"dc0880d4",
          9505 => x"38a41608",
          9506 => x"8b1133a0",
          9507 => x"07555573",
          9508 => x"8b163488",
          9509 => x"16085374",
          9510 => x"52750851",
          9511 => x"dde83f8c",
          9512 => x"1608529c",
          9513 => x"1551c9fb",
          9514 => x"3f8288b2",
          9515 => x"0a529615",
          9516 => x"51c9f03f",
          9517 => x"76529215",
          9518 => x"51c9ca3f",
          9519 => x"7854810b",
          9520 => x"83153478",
          9521 => x"51ccdf3f",
          9522 => x"82bbdc08",
          9523 => x"90173381",
          9524 => x"bf065557",
          9525 => x"73901734",
          9526 => x"7682bbdc",
          9527 => x"0c8a3d0d",
          9528 => x"04fc3d0d",
          9529 => x"76705254",
          9530 => x"fed93f82",
          9531 => x"bbdc0853",
          9532 => x"82bbdc08",
          9533 => x"9c38863d",
          9534 => x"fc055273",
          9535 => x"51f1bc3f",
          9536 => x"82bbdc08",
          9537 => x"5382bbdc",
          9538 => x"08873882",
          9539 => x"bbdc0874",
          9540 => x"0c7282bb",
          9541 => x"dc0c863d",
          9542 => x"0d04ff3d",
          9543 => x"0d843d51",
          9544 => x"e6e43f8b",
          9545 => x"52800b82",
          9546 => x"bbdc0824",
          9547 => x"8b3882bb",
          9548 => x"dc0882d3",
          9549 => x"a8348052",
          9550 => x"7182bbdc",
          9551 => x"0c833d0d",
          9552 => x"04ef3d0d",
          9553 => x"8053933d",
          9554 => x"d0055294",
          9555 => x"3d51e9c1",
          9556 => x"3f82bbdc",
          9557 => x"085582bb",
          9558 => x"dc0880e0",
          9559 => x"38765863",
          9560 => x"52933dd4",
          9561 => x"0551e08d",
          9562 => x"3f82bbdc",
          9563 => x"085582bb",
          9564 => x"dc08bc38",
          9565 => x"0280c705",
          9566 => x"3370982b",
          9567 => x"55567380",
          9568 => x"25893876",
          9569 => x"7a94120c",
          9570 => x"54b23902",
          9571 => x"a2053370",
          9572 => x"842a7081",
          9573 => x"06515556",
          9574 => x"73802e9e",
          9575 => x"38767f53",
          9576 => x"705254db",
          9577 => x"a83f82bb",
          9578 => x"dc089415",
          9579 => x"0c8e3982",
          9580 => x"bbdc0884",
          9581 => x"2e098106",
          9582 => x"83388555",
          9583 => x"7482bbdc",
          9584 => x"0c933d0d",
          9585 => x"04e43d0d",
          9586 => x"6f6f5b5b",
          9587 => x"807a3480",
          9588 => x"539e3dff",
          9589 => x"b805529f",
          9590 => x"3d51e8b5",
          9591 => x"3f82bbdc",
          9592 => x"085782bb",
          9593 => x"dc0882fc",
          9594 => x"387b437a",
          9595 => x"7c941108",
          9596 => x"47555864",
          9597 => x"5473802e",
          9598 => x"81ed38a0",
          9599 => x"52933d70",
          9600 => x"5255d5ea",
          9601 => x"3f82bbdc",
          9602 => x"085782bb",
          9603 => x"dc0882d4",
          9604 => x"3868527b",
          9605 => x"51c9c83f",
          9606 => x"82bbdc08",
          9607 => x"5782bbdc",
          9608 => x"0882c138",
          9609 => x"69527b51",
          9610 => x"daa33f82",
          9611 => x"bbdc0845",
          9612 => x"76527451",
          9613 => x"d5b83f82",
          9614 => x"bbdc0857",
          9615 => x"82bbdc08",
          9616 => x"82a23880",
          9617 => x"527451da",
          9618 => x"eb3f82bb",
          9619 => x"dc085782",
          9620 => x"bbdc08a4",
          9621 => x"3869527b",
          9622 => x"51d9f23f",
          9623 => x"7382bbdc",
          9624 => x"082ea638",
          9625 => x"76527451",
          9626 => x"d6cf3f82",
          9627 => x"bbdc0857",
          9628 => x"82bbdc08",
          9629 => x"802ecc38",
          9630 => x"76842e09",
          9631 => x"81068638",
          9632 => x"825781e0",
          9633 => x"397681dc",
          9634 => x"389e3dff",
          9635 => x"bc055274",
          9636 => x"51dcc93f",
          9637 => x"76903d78",
          9638 => x"11811133",
          9639 => x"51565a56",
          9640 => x"73802e91",
          9641 => x"3802b905",
          9642 => x"55811681",
          9643 => x"16703356",
          9644 => x"565673f5",
          9645 => x"38811654",
          9646 => x"73782681",
          9647 => x"90387580",
          9648 => x"2e993878",
          9649 => x"16810555",
          9650 => x"ff186f11",
          9651 => x"ff18ff18",
          9652 => x"58585558",
          9653 => x"74337434",
          9654 => x"75ee38ff",
          9655 => x"186f1155",
          9656 => x"58af7434",
          9657 => x"fe8d3977",
          9658 => x"7b2e0981",
          9659 => x"068a38ff",
          9660 => x"186f1155",
          9661 => x"58af7434",
          9662 => x"800b82d3",
          9663 => x"a8337084",
          9664 => x"2982b594",
          9665 => x"05700870",
          9666 => x"33525c56",
          9667 => x"56567376",
          9668 => x"2e8d3881",
          9669 => x"16701a70",
          9670 => x"33515556",
          9671 => x"73f53882",
          9672 => x"16547378",
          9673 => x"26a73880",
          9674 => x"55747627",
          9675 => x"91387419",
          9676 => x"5473337a",
          9677 => x"7081055c",
          9678 => x"34811555",
          9679 => x"ec39ba7a",
          9680 => x"7081055c",
          9681 => x"3474ff2e",
          9682 => x"09810685",
          9683 => x"38915794",
          9684 => x"396e1881",
          9685 => x"19595473",
          9686 => x"337a7081",
          9687 => x"055c347a",
          9688 => x"7826ee38",
          9689 => x"807a3476",
          9690 => x"82bbdc0c",
          9691 => x"9e3d0d04",
          9692 => x"f73d0d7b",
          9693 => x"7d8d3dfc",
          9694 => x"05547153",
          9695 => x"5755ecbb",
          9696 => x"3f82bbdc",
          9697 => x"085382bb",
          9698 => x"dc0882fa",
          9699 => x"38911533",
          9700 => x"537282f2",
          9701 => x"388c1508",
          9702 => x"54737627",
          9703 => x"92389015",
          9704 => x"3370812a",
          9705 => x"70810651",
          9706 => x"54577283",
          9707 => x"38735694",
          9708 => x"15085480",
          9709 => x"7094170c",
          9710 => x"5875782e",
          9711 => x"82973879",
          9712 => x"8a112270",
          9713 => x"892b5951",
          9714 => x"5373782e",
          9715 => x"b7387652",
          9716 => x"ff1651fe",
          9717 => x"d7ad3f82",
          9718 => x"bbdc08ff",
          9719 => x"15785470",
          9720 => x"535553fe",
          9721 => x"d79d3f82",
          9722 => x"bbdc0873",
          9723 => x"26963876",
          9724 => x"30707506",
          9725 => x"7094180c",
          9726 => x"77713198",
          9727 => x"18085758",
          9728 => x"5153b139",
          9729 => x"88150854",
          9730 => x"73a63873",
          9731 => x"527451cd",
          9732 => x"ca3f82bb",
          9733 => x"dc085482",
          9734 => x"bbdc0881",
          9735 => x"2e819a38",
          9736 => x"82bbdc08",
          9737 => x"ff2e819b",
          9738 => x"3882bbdc",
          9739 => x"0888160c",
          9740 => x"7398160c",
          9741 => x"73802e81",
          9742 => x"9c387676",
          9743 => x"2780dc38",
          9744 => x"75773194",
          9745 => x"16081894",
          9746 => x"170c9016",
          9747 => x"3370812a",
          9748 => x"70810651",
          9749 => x"555a5672",
          9750 => x"802e9a38",
          9751 => x"73527451",
          9752 => x"ccf93f82",
          9753 => x"bbdc0854",
          9754 => x"82bbdc08",
          9755 => x"943882bb",
          9756 => x"dc0856a7",
          9757 => x"39735274",
          9758 => x"51c7843f",
          9759 => x"82bbdc08",
          9760 => x"5473ff2e",
          9761 => x"be388174",
          9762 => x"27af3879",
          9763 => x"53739814",
          9764 => x"0827a638",
          9765 => x"7398160c",
          9766 => x"ffa03994",
          9767 => x"15081694",
          9768 => x"160c7583",
          9769 => x"ff065372",
          9770 => x"802eaa38",
          9771 => x"73527951",
          9772 => x"c6a33f82",
          9773 => x"bbdc0894",
          9774 => x"38820b91",
          9775 => x"16348253",
          9776 => x"80c43981",
          9777 => x"0b911634",
          9778 => x"8153bb39",
          9779 => x"75892a82",
          9780 => x"bbdc0805",
          9781 => x"58941508",
          9782 => x"548c1508",
          9783 => x"74279038",
          9784 => x"738c160c",
          9785 => x"90153380",
          9786 => x"c0075372",
          9787 => x"90163473",
          9788 => x"83ff0653",
          9789 => x"72802e8c",
          9790 => x"38779c16",
          9791 => x"082e8538",
          9792 => x"779c160c",
          9793 => x"80537282",
          9794 => x"bbdc0c8b",
          9795 => x"3d0d04f9",
          9796 => x"3d0d7956",
          9797 => x"89547580",
          9798 => x"2e818a38",
          9799 => x"8053893d",
          9800 => x"fc05528a",
          9801 => x"3d840551",
          9802 => x"e1e73f82",
          9803 => x"bbdc0855",
          9804 => x"82bbdc08",
          9805 => x"80ea3877",
          9806 => x"760c7a52",
          9807 => x"7551d8b5",
          9808 => x"3f82bbdc",
          9809 => x"085582bb",
          9810 => x"dc0880c3",
          9811 => x"38ab1633",
          9812 => x"70982b55",
          9813 => x"57807424",
          9814 => x"a2388616",
          9815 => x"3370842a",
          9816 => x"70810651",
          9817 => x"55577380",
          9818 => x"2ead389c",
          9819 => x"16085277",
          9820 => x"51d3da3f",
          9821 => x"82bbdc08",
          9822 => x"88170c77",
          9823 => x"54861422",
          9824 => x"84172374",
          9825 => x"527551ce",
          9826 => x"e53f82bb",
          9827 => x"dc085574",
          9828 => x"842e0981",
          9829 => x"06853885",
          9830 => x"55863974",
          9831 => x"802e8438",
          9832 => x"80760c74",
          9833 => x"547382bb",
          9834 => x"dc0c893d",
          9835 => x"0d04fc3d",
          9836 => x"0d76873d",
          9837 => x"fc055370",
          9838 => x"5253e7ff",
          9839 => x"3f82bbdc",
          9840 => x"08873882",
          9841 => x"bbdc0873",
          9842 => x"0c863d0d",
          9843 => x"04fb3d0d",
          9844 => x"7779893d",
          9845 => x"fc055471",
          9846 => x"535654e7",
          9847 => x"de3f82bb",
          9848 => x"dc085382",
          9849 => x"bbdc0880",
          9850 => x"df387493",
          9851 => x"3882bbdc",
          9852 => x"08527351",
          9853 => x"cdf83f82",
          9854 => x"bbdc0853",
          9855 => x"80ca3982",
          9856 => x"bbdc0852",
          9857 => x"7351d3ac",
          9858 => x"3f82bbdc",
          9859 => x"085382bb",
          9860 => x"dc08842e",
          9861 => x"09810685",
          9862 => x"38805387",
          9863 => x"3982bbdc",
          9864 => x"08a63874",
          9865 => x"527351d5",
          9866 => x"b33f7252",
          9867 => x"7351cf89",
          9868 => x"3f82bbdc",
          9869 => x"08843270",
          9870 => x"30707207",
          9871 => x"9f2c7082",
          9872 => x"bbdc0806",
          9873 => x"51515454",
          9874 => x"7282bbdc",
          9875 => x"0c873d0d",
          9876 => x"04ee3d0d",
          9877 => x"65578053",
          9878 => x"893d7053",
          9879 => x"963d5256",
          9880 => x"dfaf3f82",
          9881 => x"bbdc0855",
          9882 => x"82bbdc08",
          9883 => x"b2386452",
          9884 => x"7551d681",
          9885 => x"3f82bbdc",
          9886 => x"085582bb",
          9887 => x"dc08a038",
          9888 => x"0280cb05",
          9889 => x"3370982b",
          9890 => x"55587380",
          9891 => x"25853886",
          9892 => x"558d3976",
          9893 => x"802e8838",
          9894 => x"76527551",
          9895 => x"d4be3f74",
          9896 => x"82bbdc0c",
          9897 => x"943d0d04",
          9898 => x"f03d0d63",
          9899 => x"65555c80",
          9900 => x"53923dec",
          9901 => x"0552933d",
          9902 => x"51ded63f",
          9903 => x"82bbdc08",
          9904 => x"5b82bbdc",
          9905 => x"08828038",
          9906 => x"7c740c73",
          9907 => x"08981108",
          9908 => x"fe119013",
          9909 => x"08595658",
          9910 => x"55757426",
          9911 => x"9138757c",
          9912 => x"0c81e439",
          9913 => x"815b81cc",
          9914 => x"39825b81",
          9915 => x"c73982bb",
          9916 => x"dc087533",
          9917 => x"55597381",
          9918 => x"2e098106",
          9919 => x"bf388275",
          9920 => x"5f577652",
          9921 => x"923df005",
          9922 => x"51c1f43f",
          9923 => x"82bbdc08",
          9924 => x"ff2ed138",
          9925 => x"82bbdc08",
          9926 => x"812ece38",
          9927 => x"82bbdc08",
          9928 => x"307082bb",
          9929 => x"dc080780",
          9930 => x"257a0581",
          9931 => x"197f5359",
          9932 => x"5a549814",
          9933 => x"087726ca",
          9934 => x"3880f939",
          9935 => x"a4150882",
          9936 => x"bbdc0857",
          9937 => x"58759838",
          9938 => x"77528118",
          9939 => x"7d5258ff",
          9940 => x"bf8d3f82",
          9941 => x"bbdc085b",
          9942 => x"82bbdc08",
          9943 => x"80d6387c",
          9944 => x"70337712",
          9945 => x"ff1a5d52",
          9946 => x"56547482",
          9947 => x"2e098106",
          9948 => x"9e38b414",
          9949 => x"51ffbbcb",
          9950 => x"3f82bbdc",
          9951 => x"0883ffff",
          9952 => x"06703070",
          9953 => x"80251b82",
          9954 => x"19595b51",
          9955 => x"549b39b4",
          9956 => x"1451ffbb",
          9957 => x"c53f82bb",
          9958 => x"dc08f00a",
          9959 => x"06703070",
          9960 => x"80251b84",
          9961 => x"19595b51",
          9962 => x"547583ff",
          9963 => x"067a5856",
          9964 => x"79ff9238",
          9965 => x"787c0c7c",
          9966 => x"7990120c",
          9967 => x"84113381",
          9968 => x"07565474",
          9969 => x"8415347a",
          9970 => x"82bbdc0c",
          9971 => x"923d0d04",
          9972 => x"f93d0d79",
          9973 => x"8a3dfc05",
          9974 => x"53705257",
          9975 => x"e3dd3f82",
          9976 => x"bbdc0856",
          9977 => x"82bbdc08",
          9978 => x"81a83891",
          9979 => x"17335675",
          9980 => x"81a03890",
          9981 => x"17337081",
          9982 => x"2a708106",
          9983 => x"51555587",
          9984 => x"5573802e",
          9985 => x"818e3894",
          9986 => x"17085473",
          9987 => x"8c180827",
          9988 => x"81803873",
          9989 => x"9b3882bb",
          9990 => x"dc085388",
          9991 => x"17085276",
          9992 => x"51c48c3f",
          9993 => x"82bbdc08",
          9994 => x"7488190c",
          9995 => x"5680c939",
          9996 => x"98170852",
          9997 => x"7651ffbf",
          9998 => x"c63f82bb",
          9999 => x"dc08ff2e",
         10000 => x"09810683",
         10001 => x"38815682",
         10002 => x"bbdc0881",
         10003 => x"2e098106",
         10004 => x"85388256",
         10005 => x"a33975a0",
         10006 => x"38775482",
         10007 => x"bbdc0898",
         10008 => x"15082794",
         10009 => x"38981708",
         10010 => x"5382bbdc",
         10011 => x"08527651",
         10012 => x"c3bd3f82",
         10013 => x"bbdc0856",
         10014 => x"9417088c",
         10015 => x"180c9017",
         10016 => x"3380c007",
         10017 => x"54739018",
         10018 => x"3475802e",
         10019 => x"85387591",
         10020 => x"18347555",
         10021 => x"7482bbdc",
         10022 => x"0c893d0d",
         10023 => x"04e23d0d",
         10024 => x"8253a03d",
         10025 => x"ffa40552",
         10026 => x"a13d51da",
         10027 => x"e43f82bb",
         10028 => x"dc085582",
         10029 => x"bbdc0881",
         10030 => x"f5387845",
         10031 => x"a13d0852",
         10032 => x"953d7052",
         10033 => x"58d1ae3f",
         10034 => x"82bbdc08",
         10035 => x"5582bbdc",
         10036 => x"0881db38",
         10037 => x"0280fb05",
         10038 => x"3370852a",
         10039 => x"70810651",
         10040 => x"55568655",
         10041 => x"7381c738",
         10042 => x"75982b54",
         10043 => x"80742481",
         10044 => x"bd380280",
         10045 => x"d6053370",
         10046 => x"81065854",
         10047 => x"87557681",
         10048 => x"ad386b52",
         10049 => x"7851ccc5",
         10050 => x"3f82bbdc",
         10051 => x"0874842a",
         10052 => x"70810651",
         10053 => x"55567380",
         10054 => x"2e80d438",
         10055 => x"785482bb",
         10056 => x"dc089415",
         10057 => x"082e8186",
         10058 => x"38735a82",
         10059 => x"bbdc085c",
         10060 => x"76528a3d",
         10061 => x"705254c7",
         10062 => x"b53f82bb",
         10063 => x"dc085582",
         10064 => x"bbdc0880",
         10065 => x"e93882bb",
         10066 => x"dc085273",
         10067 => x"51cce53f",
         10068 => x"82bbdc08",
         10069 => x"5582bbdc",
         10070 => x"08863887",
         10071 => x"5580cf39",
         10072 => x"82bbdc08",
         10073 => x"842e8838",
         10074 => x"82bbdc08",
         10075 => x"80c03877",
         10076 => x"51cec23f",
         10077 => x"82bbdc08",
         10078 => x"82bbdc08",
         10079 => x"307082bb",
         10080 => x"dc080780",
         10081 => x"25515555",
         10082 => x"75802e94",
         10083 => x"3873802e",
         10084 => x"8f388053",
         10085 => x"75527751",
         10086 => x"c1953f82",
         10087 => x"bbdc0855",
         10088 => x"748c3878",
         10089 => x"51ffbafe",
         10090 => x"3f82bbdc",
         10091 => x"08557482",
         10092 => x"bbdc0ca0",
         10093 => x"3d0d04e9",
         10094 => x"3d0d8253",
         10095 => x"993dc005",
         10096 => x"529a3d51",
         10097 => x"d8cb3f82",
         10098 => x"bbdc0854",
         10099 => x"82bbdc08",
         10100 => x"82b03878",
         10101 => x"5e69528e",
         10102 => x"3d705258",
         10103 => x"cf973f82",
         10104 => x"bbdc0854",
         10105 => x"82bbdc08",
         10106 => x"86388854",
         10107 => x"82943982",
         10108 => x"bbdc0884",
         10109 => x"2e098106",
         10110 => x"82883802",
         10111 => x"80df0533",
         10112 => x"70852a81",
         10113 => x"06515586",
         10114 => x"547481f6",
         10115 => x"38785a74",
         10116 => x"528a3d70",
         10117 => x"5257c1c3",
         10118 => x"3f82bbdc",
         10119 => x"08755556",
         10120 => x"82bbdc08",
         10121 => x"83388754",
         10122 => x"82bbdc08",
         10123 => x"812e0981",
         10124 => x"06833882",
         10125 => x"5482bbdc",
         10126 => x"08ff2e09",
         10127 => x"81068638",
         10128 => x"815481b4",
         10129 => x"397381b0",
         10130 => x"3882bbdc",
         10131 => x"08527851",
         10132 => x"c4a43f82",
         10133 => x"bbdc0854",
         10134 => x"82bbdc08",
         10135 => x"819a388b",
         10136 => x"53a052b4",
         10137 => x"1951ffb7",
         10138 => x"8c3f7854",
         10139 => x"ae0bb415",
         10140 => x"34785490",
         10141 => x"0bbf1534",
         10142 => x"8288b20a",
         10143 => x"5280ca19",
         10144 => x"51ffb69f",
         10145 => x"3f755378",
         10146 => x"b4115351",
         10147 => x"c9f83fa0",
         10148 => x"5378b411",
         10149 => x"5380d405",
         10150 => x"51ffb6b6",
         10151 => x"3f7854ae",
         10152 => x"0b80d515",
         10153 => x"347f5378",
         10154 => x"80d41153",
         10155 => x"51c9d73f",
         10156 => x"7854810b",
         10157 => x"83153477",
         10158 => x"51cba43f",
         10159 => x"82bbdc08",
         10160 => x"5482bbdc",
         10161 => x"08b23882",
         10162 => x"88b20a52",
         10163 => x"64960551",
         10164 => x"ffb5d03f",
         10165 => x"75536452",
         10166 => x"7851c9aa",
         10167 => x"3f645490",
         10168 => x"0b8b1534",
         10169 => x"7854810b",
         10170 => x"83153478",
         10171 => x"51ffb8b6",
         10172 => x"3f82bbdc",
         10173 => x"08548b39",
         10174 => x"80537552",
         10175 => x"7651ffbe",
         10176 => x"ae3f7382",
         10177 => x"bbdc0c99",
         10178 => x"3d0d04da",
         10179 => x"3d0da93d",
         10180 => x"840551d2",
         10181 => x"f13f8253",
         10182 => x"a83dff84",
         10183 => x"0552a93d",
         10184 => x"51d5ee3f",
         10185 => x"82bbdc08",
         10186 => x"5582bbdc",
         10187 => x"0882d338",
         10188 => x"784da93d",
         10189 => x"08529d3d",
         10190 => x"705258cc",
         10191 => x"b83f82bb",
         10192 => x"dc085582",
         10193 => x"bbdc0882",
         10194 => x"b9380281",
         10195 => x"9b053381",
         10196 => x"a0065486",
         10197 => x"557382aa",
         10198 => x"38a053a4",
         10199 => x"3d0852a8",
         10200 => x"3dff8805",
         10201 => x"51ffb4ea",
         10202 => x"3fac5377",
         10203 => x"52923d70",
         10204 => x"5254ffb4",
         10205 => x"dd3faa3d",
         10206 => x"08527351",
         10207 => x"cbf73f82",
         10208 => x"bbdc0855",
         10209 => x"82bbdc08",
         10210 => x"9538636f",
         10211 => x"2e098106",
         10212 => x"883865a2",
         10213 => x"3d082e92",
         10214 => x"38885581",
         10215 => x"e53982bb",
         10216 => x"dc08842e",
         10217 => x"09810681",
         10218 => x"b8387351",
         10219 => x"c9b13f82",
         10220 => x"bbdc0855",
         10221 => x"82bbdc08",
         10222 => x"81c83868",
         10223 => x"569353a8",
         10224 => x"3dff9505",
         10225 => x"528d1651",
         10226 => x"ffb4873f",
         10227 => x"02af0533",
         10228 => x"8b17348b",
         10229 => x"16337084",
         10230 => x"2a708106",
         10231 => x"51555573",
         10232 => x"893874a0",
         10233 => x"0754738b",
         10234 => x"17347854",
         10235 => x"810b8315",
         10236 => x"348b1633",
         10237 => x"70842a70",
         10238 => x"81065155",
         10239 => x"5573802e",
         10240 => x"80e5386e",
         10241 => x"642e80df",
         10242 => x"38755278",
         10243 => x"51c6be3f",
         10244 => x"82bbdc08",
         10245 => x"527851ff",
         10246 => x"b7bb3f82",
         10247 => x"5582bbdc",
         10248 => x"08802e80",
         10249 => x"dd3882bb",
         10250 => x"dc085278",
         10251 => x"51ffb5af",
         10252 => x"3f82bbdc",
         10253 => x"087980d4",
         10254 => x"11585855",
         10255 => x"82bbdc08",
         10256 => x"80c03881",
         10257 => x"16335473",
         10258 => x"ae2e0981",
         10259 => x"06993863",
         10260 => x"53755276",
         10261 => x"51c6af3f",
         10262 => x"7854810b",
         10263 => x"83153487",
         10264 => x"3982bbdc",
         10265 => x"089c3877",
         10266 => x"51c8ca3f",
         10267 => x"82bbdc08",
         10268 => x"5582bbdc",
         10269 => x"088c3878",
         10270 => x"51ffb5aa",
         10271 => x"3f82bbdc",
         10272 => x"08557482",
         10273 => x"bbdc0ca8",
         10274 => x"3d0d04ed",
         10275 => x"3d0d0280",
         10276 => x"db053302",
         10277 => x"840580df",
         10278 => x"05335757",
         10279 => x"8253953d",
         10280 => x"d0055296",
         10281 => x"3d51d2e9",
         10282 => x"3f82bbdc",
         10283 => x"085582bb",
         10284 => x"dc0880cf",
         10285 => x"38785a65",
         10286 => x"52953dd4",
         10287 => x"0551c9b5",
         10288 => x"3f82bbdc",
         10289 => x"085582bb",
         10290 => x"dc08b838",
         10291 => x"0280cf05",
         10292 => x"3381a006",
         10293 => x"54865573",
         10294 => x"aa3875a7",
         10295 => x"06617109",
         10296 => x"8b123371",
         10297 => x"067a7406",
         10298 => x"07515755",
         10299 => x"56748b15",
         10300 => x"34785481",
         10301 => x"0b831534",
         10302 => x"7851ffb4",
         10303 => x"a93f82bb",
         10304 => x"dc085574",
         10305 => x"82bbdc0c",
         10306 => x"953d0d04",
         10307 => x"ef3d0d64",
         10308 => x"56825393",
         10309 => x"3dd00552",
         10310 => x"943d51d1",
         10311 => x"f43f82bb",
         10312 => x"dc085582",
         10313 => x"bbdc0880",
         10314 => x"cb387658",
         10315 => x"6352933d",
         10316 => x"d40551c8",
         10317 => x"c03f82bb",
         10318 => x"dc085582",
         10319 => x"bbdc08b4",
         10320 => x"380280c7",
         10321 => x"053381a0",
         10322 => x"06548655",
         10323 => x"73a63884",
         10324 => x"16228617",
         10325 => x"2271902b",
         10326 => x"07535496",
         10327 => x"1f51ffb0",
         10328 => x"c23f7654",
         10329 => x"810b8315",
         10330 => x"347651ff",
         10331 => x"b3b83f82",
         10332 => x"bbdc0855",
         10333 => x"7482bbdc",
         10334 => x"0c933d0d",
         10335 => x"04ea3d0d",
         10336 => x"696b5c5a",
         10337 => x"8053983d",
         10338 => x"d0055299",
         10339 => x"3d51d181",
         10340 => x"3f82bbdc",
         10341 => x"0882bbdc",
         10342 => x"08307082",
         10343 => x"bbdc0807",
         10344 => x"80255155",
         10345 => x"5779802e",
         10346 => x"81853881",
         10347 => x"70750655",
         10348 => x"5573802e",
         10349 => x"80f9387b",
         10350 => x"5d805f80",
         10351 => x"528d3d70",
         10352 => x"5254ffbe",
         10353 => x"a93f82bb",
         10354 => x"dc085782",
         10355 => x"bbdc0880",
         10356 => x"d1387452",
         10357 => x"7351c3dc",
         10358 => x"3f82bbdc",
         10359 => x"085782bb",
         10360 => x"dc08bf38",
         10361 => x"82bbdc08",
         10362 => x"82bbdc08",
         10363 => x"655b5956",
         10364 => x"78188119",
         10365 => x"7b185659",
         10366 => x"55743374",
         10367 => x"34811656",
         10368 => x"8a7827ec",
         10369 => x"388b5675",
         10370 => x"1a548074",
         10371 => x"3475802e",
         10372 => x"9e38ff16",
         10373 => x"701b7033",
         10374 => x"51555673",
         10375 => x"a02ee838",
         10376 => x"8e397684",
         10377 => x"2e098106",
         10378 => x"8638807a",
         10379 => x"34805776",
         10380 => x"30707807",
         10381 => x"80255154",
         10382 => x"7a802e80",
         10383 => x"c1387380",
         10384 => x"2ebc387b",
         10385 => x"a0110853",
         10386 => x"51ffb193",
         10387 => x"3f82bbdc",
         10388 => x"085782bb",
         10389 => x"dc08a738",
         10390 => x"7b703355",
         10391 => x"5580c356",
         10392 => x"73832e8b",
         10393 => x"3880e456",
         10394 => x"73842e83",
         10395 => x"38a75675",
         10396 => x"15b40551",
         10397 => x"ffade33f",
         10398 => x"82bbdc08",
         10399 => x"7b0c7682",
         10400 => x"bbdc0c98",
         10401 => x"3d0d04e6",
         10402 => x"3d0d8253",
         10403 => x"9c3dffb8",
         10404 => x"05529d3d",
         10405 => x"51cefa3f",
         10406 => x"82bbdc08",
         10407 => x"82bbdc08",
         10408 => x"565482bb",
         10409 => x"dc088398",
         10410 => x"388b53a0",
         10411 => x"528b3d70",
         10412 => x"5259ffae",
         10413 => x"c03f736d",
         10414 => x"70337081",
         10415 => x"ff065257",
         10416 => x"55579f74",
         10417 => x"2781bc38",
         10418 => x"78587481",
         10419 => x"ff066d81",
         10420 => x"054e7052",
         10421 => x"55ffaf89",
         10422 => x"3f82bbdc",
         10423 => x"08802ea5",
         10424 => x"386c7033",
         10425 => x"70535754",
         10426 => x"ffaefd3f",
         10427 => x"82bbdc08",
         10428 => x"802e8d38",
         10429 => x"74882b76",
         10430 => x"076d8105",
         10431 => x"4e558639",
         10432 => x"82bbdc08",
         10433 => x"55ff9f15",
         10434 => x"7083ffff",
         10435 => x"06515473",
         10436 => x"99268a38",
         10437 => x"e0157083",
         10438 => x"ffff0656",
         10439 => x"5480ff75",
         10440 => x"27873882",
         10441 => x"b4a41533",
         10442 => x"5574802e",
         10443 => x"a3387452",
         10444 => x"82b6a451",
         10445 => x"ffae893f",
         10446 => x"82bbdc08",
         10447 => x"933881ff",
         10448 => x"75278838",
         10449 => x"76892688",
         10450 => x"388b398a",
         10451 => x"77278638",
         10452 => x"865581ec",
         10453 => x"3981ff75",
         10454 => x"278f3874",
         10455 => x"882a5473",
         10456 => x"78708105",
         10457 => x"5a348117",
         10458 => x"57747870",
         10459 => x"81055a34",
         10460 => x"81176d70",
         10461 => x"337081ff",
         10462 => x"06525755",
         10463 => x"57739f26",
         10464 => x"fec8388b",
         10465 => x"3d335486",
         10466 => x"557381e5",
         10467 => x"2e81b138",
         10468 => x"76802e99",
         10469 => x"3802a705",
         10470 => x"55761570",
         10471 => x"33515473",
         10472 => x"a02e0981",
         10473 => x"068738ff",
         10474 => x"175776ed",
         10475 => x"38794180",
         10476 => x"43805291",
         10477 => x"3d705255",
         10478 => x"ffbab33f",
         10479 => x"82bbdc08",
         10480 => x"5482bbdc",
         10481 => x"0880f738",
         10482 => x"81527451",
         10483 => x"ffbfe53f",
         10484 => x"82bbdc08",
         10485 => x"5482bbdc",
         10486 => x"088d3876",
         10487 => x"80c43867",
         10488 => x"54e57434",
         10489 => x"80c63982",
         10490 => x"bbdc0884",
         10491 => x"2e098106",
         10492 => x"80cc3880",
         10493 => x"5476742e",
         10494 => x"80c43881",
         10495 => x"527451ff",
         10496 => x"bdb03f82",
         10497 => x"bbdc0854",
         10498 => x"82bbdc08",
         10499 => x"b138a053",
         10500 => x"82bbdc08",
         10501 => x"526751ff",
         10502 => x"abdb3f67",
         10503 => x"54880b8b",
         10504 => x"15348b53",
         10505 => x"78526751",
         10506 => x"ffaba73f",
         10507 => x"7954810b",
         10508 => x"83153479",
         10509 => x"51ffadee",
         10510 => x"3f82bbdc",
         10511 => x"08547355",
         10512 => x"7482bbdc",
         10513 => x"0c9c3d0d",
         10514 => x"04f23d0d",
         10515 => x"60620288",
         10516 => x"0580cb05",
         10517 => x"33933dfc",
         10518 => x"05557254",
         10519 => x"405e5ad2",
         10520 => x"da3f82bb",
         10521 => x"dc085882",
         10522 => x"bbdc0882",
         10523 => x"bd38911a",
         10524 => x"33587782",
         10525 => x"b5387c80",
         10526 => x"2e97388c",
         10527 => x"1a085978",
         10528 => x"9038901a",
         10529 => x"3370812a",
         10530 => x"70810651",
         10531 => x"55557390",
         10532 => x"38875482",
         10533 => x"97398258",
         10534 => x"82903981",
         10535 => x"58828b39",
         10536 => x"7e8a1122",
         10537 => x"70892b70",
         10538 => x"557f5456",
         10539 => x"5656febd",
         10540 => x"d23fff14",
         10541 => x"7d067030",
         10542 => x"7072079f",
         10543 => x"2a82bbdc",
         10544 => x"08058c19",
         10545 => x"087c405a",
         10546 => x"5d555581",
         10547 => x"77278838",
         10548 => x"98160877",
         10549 => x"26833882",
         10550 => x"57767756",
         10551 => x"59805674",
         10552 => x"527951ff",
         10553 => x"ae993f81",
         10554 => x"157f5555",
         10555 => x"98140875",
         10556 => x"26833882",
         10557 => x"5582bbdc",
         10558 => x"08812eff",
         10559 => x"993882bb",
         10560 => x"dc08ff2e",
         10561 => x"ff953882",
         10562 => x"bbdc088e",
         10563 => x"38811656",
         10564 => x"757b2e09",
         10565 => x"81068738",
         10566 => x"93397459",
         10567 => x"80567477",
         10568 => x"2e098106",
         10569 => x"ffb93887",
         10570 => x"5880ff39",
         10571 => x"7d802eba",
         10572 => x"38787b55",
         10573 => x"557a802e",
         10574 => x"b4388115",
         10575 => x"5673812e",
         10576 => x"09810683",
         10577 => x"38ff5675",
         10578 => x"5374527e",
         10579 => x"51ffafa8",
         10580 => x"3f82bbdc",
         10581 => x"085882bb",
         10582 => x"dc0880ce",
         10583 => x"38748116",
         10584 => x"ff165656",
         10585 => x"5c73d338",
         10586 => x"8439ff19",
         10587 => x"5c7e7c8c",
         10588 => x"120c557d",
         10589 => x"802eb338",
         10590 => x"78881b0c",
         10591 => x"7c8c1b0c",
         10592 => x"901a3380",
         10593 => x"c0075473",
         10594 => x"901b3498",
         10595 => x"1508fe05",
         10596 => x"90160857",
         10597 => x"54757426",
         10598 => x"9138757b",
         10599 => x"3190160c",
         10600 => x"84153381",
         10601 => x"07547384",
         10602 => x"16347754",
         10603 => x"7382bbdc",
         10604 => x"0c903d0d",
         10605 => x"04e93d0d",
         10606 => x"6b6d0288",
         10607 => x"0580eb05",
         10608 => x"339d3d54",
         10609 => x"5a5c59c5",
         10610 => x"bd3f8b56",
         10611 => x"800b82bb",
         10612 => x"dc08248b",
         10613 => x"f83882bb",
         10614 => x"dc088429",
         10615 => x"82d39405",
         10616 => x"70085155",
         10617 => x"74802e84",
         10618 => x"38807534",
         10619 => x"82bbdc08",
         10620 => x"81ff065f",
         10621 => x"81527e51",
         10622 => x"ffa0d03f",
         10623 => x"82bbdc08",
         10624 => x"81ff0670",
         10625 => x"81065657",
         10626 => x"8356748b",
         10627 => x"c0387682",
         10628 => x"2a708106",
         10629 => x"51558a56",
         10630 => x"748bb238",
         10631 => x"993dfc05",
         10632 => x"5383527e",
         10633 => x"51ffa4f0",
         10634 => x"3f82bbdc",
         10635 => x"08993867",
         10636 => x"5574802e",
         10637 => x"92387482",
         10638 => x"8080268b",
         10639 => x"38ff1575",
         10640 => x"06557480",
         10641 => x"2e833881",
         10642 => x"4878802e",
         10643 => x"87388480",
         10644 => x"79269238",
         10645 => x"7881800a",
         10646 => x"268b38ff",
         10647 => x"19790655",
         10648 => x"74802e86",
         10649 => x"3893568a",
         10650 => x"e4397889",
         10651 => x"2a6e892a",
         10652 => x"70892b77",
         10653 => x"59484359",
         10654 => x"7a833881",
         10655 => x"56613070",
         10656 => x"80257707",
         10657 => x"51559156",
         10658 => x"748ac238",
         10659 => x"993df805",
         10660 => x"5381527e",
         10661 => x"51ffa480",
         10662 => x"3f815682",
         10663 => x"bbdc088a",
         10664 => x"ac387783",
         10665 => x"2a707706",
         10666 => x"82bbdc08",
         10667 => x"43564574",
         10668 => x"8338bf41",
         10669 => x"66558e56",
         10670 => x"6075268a",
         10671 => x"90387461",
         10672 => x"31704855",
         10673 => x"80ff7527",
         10674 => x"8a833893",
         10675 => x"56788180",
         10676 => x"2689fa38",
         10677 => x"77812a70",
         10678 => x"81065643",
         10679 => x"74802e95",
         10680 => x"38778706",
         10681 => x"5574822e",
         10682 => x"838d3877",
         10683 => x"81065574",
         10684 => x"802e8383",
         10685 => x"38778106",
         10686 => x"55935682",
         10687 => x"5e74802e",
         10688 => x"89cb3878",
         10689 => x"5a7d832e",
         10690 => x"09810680",
         10691 => x"e13878ae",
         10692 => x"3866912a",
         10693 => x"57810b82",
         10694 => x"b6c82256",
         10695 => x"5a74802e",
         10696 => x"9d387477",
         10697 => x"26983882",
         10698 => x"b6c85679",
         10699 => x"10821770",
         10700 => x"2257575a",
         10701 => x"74802e86",
         10702 => x"38767527",
         10703 => x"ee387952",
         10704 => x"6651feb8",
         10705 => x"be3f82bb",
         10706 => x"dc088429",
         10707 => x"84870570",
         10708 => x"892a5e55",
         10709 => x"a05c800b",
         10710 => x"82bbdc08",
         10711 => x"fc808a05",
         10712 => x"5644fdff",
         10713 => x"f00a7527",
         10714 => x"80ec3888",
         10715 => x"d33978ae",
         10716 => x"38668c2a",
         10717 => x"57810b82",
         10718 => x"b6b82256",
         10719 => x"5a74802e",
         10720 => x"9d387477",
         10721 => x"26983882",
         10722 => x"b6b85679",
         10723 => x"10821770",
         10724 => x"2257575a",
         10725 => x"74802e86",
         10726 => x"38767527",
         10727 => x"ee387952",
         10728 => x"6651feb7",
         10729 => x"de3f82bb",
         10730 => x"dc081084",
         10731 => x"055782bb",
         10732 => x"dc089ff5",
         10733 => x"26963881",
         10734 => x"0b82bbdc",
         10735 => x"081082bb",
         10736 => x"dc080571",
         10737 => x"11722a83",
         10738 => x"0559565e",
         10739 => x"83ff1789",
         10740 => x"2a5d815c",
         10741 => x"a044601c",
         10742 => x"7d116505",
         10743 => x"697012ff",
         10744 => x"05713070",
         10745 => x"72067431",
         10746 => x"5c525957",
         10747 => x"59407d83",
         10748 => x"2e098106",
         10749 => x"8938761c",
         10750 => x"6018415c",
         10751 => x"8439761d",
         10752 => x"5d799029",
         10753 => x"18706231",
         10754 => x"68585155",
         10755 => x"74762687",
         10756 => x"af38757c",
         10757 => x"317d317a",
         10758 => x"53706531",
         10759 => x"5255feb6",
         10760 => x"e23f82bb",
         10761 => x"dc08587d",
         10762 => x"832e0981",
         10763 => x"069b3882",
         10764 => x"bbdc0883",
         10765 => x"fff52680",
         10766 => x"dd387887",
         10767 => x"83387981",
         10768 => x"2a5978fd",
         10769 => x"be3886f8",
         10770 => x"397d822e",
         10771 => x"09810680",
         10772 => x"c53883ff",
         10773 => x"f50b82bb",
         10774 => x"dc0827a0",
         10775 => x"38788f38",
         10776 => x"791a5574",
         10777 => x"80c02686",
         10778 => x"387459fd",
         10779 => x"96396281",
         10780 => x"06557480",
         10781 => x"2e8f3883",
         10782 => x"5efd8839",
         10783 => x"82bbdc08",
         10784 => x"9ff52692",
         10785 => x"387886b8",
         10786 => x"38791a59",
         10787 => x"81807927",
         10788 => x"fcf13886",
         10789 => x"ab398055",
         10790 => x"7d812e09",
         10791 => x"81068338",
         10792 => x"7d559ff5",
         10793 => x"78278b38",
         10794 => x"74810655",
         10795 => x"8e567486",
         10796 => x"9c388480",
         10797 => x"5380527a",
         10798 => x"51ffa2b9",
         10799 => x"3f8b5382",
         10800 => x"b4e0527a",
         10801 => x"51ffa28a",
         10802 => x"3f848052",
         10803 => x"8b1b51ff",
         10804 => x"a1b33f79",
         10805 => x"8d1c347b",
         10806 => x"83ffff06",
         10807 => x"528e1b51",
         10808 => x"ffa1a23f",
         10809 => x"810b901c",
         10810 => x"347d8332",
         10811 => x"70307096",
         10812 => x"2a848006",
         10813 => x"54515591",
         10814 => x"1b51ffa1",
         10815 => x"883f6655",
         10816 => x"7483ffff",
         10817 => x"26903874",
         10818 => x"83ffff06",
         10819 => x"52931b51",
         10820 => x"ffa0f23f",
         10821 => x"8a397452",
         10822 => x"a01b51ff",
         10823 => x"a1853ff8",
         10824 => x"0b951c34",
         10825 => x"bf52981b",
         10826 => x"51ffa0d9",
         10827 => x"3f81ff52",
         10828 => x"9a1b51ff",
         10829 => x"a0cf3f60",
         10830 => x"529c1b51",
         10831 => x"ffa0e43f",
         10832 => x"7d832e09",
         10833 => x"810680cb",
         10834 => x"388288b2",
         10835 => x"0a5280c3",
         10836 => x"1b51ffa0",
         10837 => x"ce3f7c52",
         10838 => x"a41b51ff",
         10839 => x"a0c53f82",
         10840 => x"52ac1b51",
         10841 => x"ffa0bc3f",
         10842 => x"8152b01b",
         10843 => x"51ffa095",
         10844 => x"3f8652b2",
         10845 => x"1b51ffa0",
         10846 => x"8c3fff80",
         10847 => x"0b80c01c",
         10848 => x"34a90b80",
         10849 => x"c21c3493",
         10850 => x"5382b4ec",
         10851 => x"5280c71b",
         10852 => x"51ae3982",
         10853 => x"88b20a52",
         10854 => x"a71b51ff",
         10855 => x"a0853f7c",
         10856 => x"83ffff06",
         10857 => x"52961b51",
         10858 => x"ff9fda3f",
         10859 => x"ff800ba4",
         10860 => x"1c34a90b",
         10861 => x"a61c3493",
         10862 => x"5382b580",
         10863 => x"52ab1b51",
         10864 => x"ffa08f3f",
         10865 => x"82d4d552",
         10866 => x"83fe1b70",
         10867 => x"5259ff9f",
         10868 => x"b43f8154",
         10869 => x"60537a52",
         10870 => x"7e51ff9b",
         10871 => x"d73f8156",
         10872 => x"82bbdc08",
         10873 => x"83e7387d",
         10874 => x"832e0981",
         10875 => x"0680ee38",
         10876 => x"75546086",
         10877 => x"05537a52",
         10878 => x"7e51ff9b",
         10879 => x"b73f8480",
         10880 => x"5380527a",
         10881 => x"51ff9fed",
         10882 => x"3f848b85",
         10883 => x"a4d2527a",
         10884 => x"51ff9f8f",
         10885 => x"3f868a85",
         10886 => x"e4f25283",
         10887 => x"e41b51ff",
         10888 => x"9f813fff",
         10889 => x"185283e8",
         10890 => x"1b51ff9e",
         10891 => x"f63f8252",
         10892 => x"83ec1b51",
         10893 => x"ff9eec3f",
         10894 => x"82d4d552",
         10895 => x"7851ff9e",
         10896 => x"c43f7554",
         10897 => x"60870553",
         10898 => x"7a527e51",
         10899 => x"ff9ae53f",
         10900 => x"75546016",
         10901 => x"537a527e",
         10902 => x"51ff9ad8",
         10903 => x"3f655380",
         10904 => x"527a51ff",
         10905 => x"9f8f3f7f",
         10906 => x"5680587d",
         10907 => x"832e0981",
         10908 => x"069a38f8",
         10909 => x"527a51ff",
         10910 => x"9ea93fff",
         10911 => x"52841b51",
         10912 => x"ff9ea03f",
         10913 => x"f00a5288",
         10914 => x"1b519139",
         10915 => x"87fffff8",
         10916 => x"557d812e",
         10917 => x"8338f855",
         10918 => x"74527a51",
         10919 => x"ff9e843f",
         10920 => x"7c556157",
         10921 => x"74622683",
         10922 => x"38745776",
         10923 => x"5475537a",
         10924 => x"527e51ff",
         10925 => x"99fe3f82",
         10926 => x"bbdc0882",
         10927 => x"87388480",
         10928 => x"5382bbdc",
         10929 => x"08527a51",
         10930 => x"ff9eaa3f",
         10931 => x"76167578",
         10932 => x"31565674",
         10933 => x"cd388118",
         10934 => x"5877802e",
         10935 => x"ff8d3879",
         10936 => x"557d832e",
         10937 => x"83386355",
         10938 => x"61577462",
         10939 => x"26833874",
         10940 => x"57765475",
         10941 => x"537a527e",
         10942 => x"51ff99b8",
         10943 => x"3f82bbdc",
         10944 => x"0881c138",
         10945 => x"76167578",
         10946 => x"31565674",
         10947 => x"db388c56",
         10948 => x"7d832e93",
         10949 => x"38865666",
         10950 => x"83ffff26",
         10951 => x"8a388456",
         10952 => x"7d822e83",
         10953 => x"38815664",
         10954 => x"81065877",
         10955 => x"80fe3884",
         10956 => x"80537752",
         10957 => x"7a51ff9d",
         10958 => x"bc3f82d4",
         10959 => x"d5527851",
         10960 => x"ff9cc23f",
         10961 => x"83be1b55",
         10962 => x"77753481",
         10963 => x"0b811634",
         10964 => x"810b8216",
         10965 => x"34778316",
         10966 => x"34758416",
         10967 => x"34606705",
         10968 => x"5680fdc1",
         10969 => x"527551fe",
         10970 => x"b0993ffe",
         10971 => x"0b851634",
         10972 => x"82bbdc08",
         10973 => x"822abf07",
         10974 => x"56758616",
         10975 => x"3482bbdc",
         10976 => x"08871634",
         10977 => x"605283c6",
         10978 => x"1b51ff9c",
         10979 => x"963f6652",
         10980 => x"83ca1b51",
         10981 => x"ff9c8c3f",
         10982 => x"81547753",
         10983 => x"7a527e51",
         10984 => x"ff98913f",
         10985 => x"815682bb",
         10986 => x"dc08a238",
         10987 => x"80538052",
         10988 => x"7e51ff99",
         10989 => x"e33f8156",
         10990 => x"82bbdc08",
         10991 => x"90388939",
         10992 => x"8e568a39",
         10993 => x"81568639",
         10994 => x"82bbdc08",
         10995 => x"567582bb",
         10996 => x"dc0c993d",
         10997 => x"0d04f53d",
         10998 => x"0d7d605b",
         10999 => x"59807960",
         11000 => x"ff055a57",
         11001 => x"57767825",
         11002 => x"b4388d3d",
         11003 => x"f8115555",
         11004 => x"8153fc15",
         11005 => x"527951c9",
         11006 => x"dc3f7a81",
         11007 => x"2e098106",
         11008 => x"9c388c3d",
         11009 => x"3355748d",
         11010 => x"2edb3874",
         11011 => x"76708105",
         11012 => x"58348117",
         11013 => x"57748a2e",
         11014 => x"098106c9",
         11015 => x"38807634",
         11016 => x"78557683",
         11017 => x"38765574",
         11018 => x"82bbdc0c",
         11019 => x"8d3d0d04",
         11020 => x"f73d0d7b",
         11021 => x"028405b3",
         11022 => x"05335957",
         11023 => x"778a2e09",
         11024 => x"81068738",
         11025 => x"8d527651",
         11026 => x"e73f8417",
         11027 => x"08568076",
         11028 => x"24be3888",
         11029 => x"17087717",
         11030 => x"8c055659",
         11031 => x"77753481",
         11032 => x"1656bb76",
         11033 => x"25a1388b",
         11034 => x"3dfc0554",
         11035 => x"75538c17",
         11036 => x"52760851",
         11037 => x"cbdc3f79",
         11038 => x"76327030",
         11039 => x"7072079f",
         11040 => x"2a703053",
         11041 => x"51565675",
         11042 => x"84180c81",
         11043 => x"1988180c",
         11044 => x"8b3d0d04",
         11045 => x"f93d0d79",
         11046 => x"84110856",
         11047 => x"56807524",
         11048 => x"a738893d",
         11049 => x"fc055474",
         11050 => x"538c1652",
         11051 => x"750851cb",
         11052 => x"a13f82bb",
         11053 => x"dc089138",
         11054 => x"84160878",
         11055 => x"2e098106",
         11056 => x"87388816",
         11057 => x"08558339",
         11058 => x"ff557482",
         11059 => x"bbdc0c89",
         11060 => x"3d0d04fd",
         11061 => x"3d0d7554",
         11062 => x"80cc5380",
         11063 => x"527351ff",
         11064 => x"9a933f76",
         11065 => x"740c853d",
         11066 => x"0d04ea3d",
         11067 => x"0d0280e3",
         11068 => x"05336a53",
         11069 => x"863d7053",
         11070 => x"5454d83f",
         11071 => x"73527251",
         11072 => x"feae3f72",
         11073 => x"51ff8d3f",
         11074 => x"983d0d04",
         11075 => x"00ffffff",
         11076 => x"ff00ffff",
         11077 => x"ffff00ff",
         11078 => x"ffffff00",
         11079 => x"00002baa",
         11080 => x"00002b2e",
         11081 => x"00002b35",
         11082 => x"00002b3c",
         11083 => x"00002b43",
         11084 => x"00002b4a",
         11085 => x"00002b51",
         11086 => x"00002b58",
         11087 => x"00002b5f",
         11088 => x"00002b66",
         11089 => x"00002b6d",
         11090 => x"00002b74",
         11091 => x"00002b7a",
         11092 => x"00002b80",
         11093 => x"00002b86",
         11094 => x"00002b8c",
         11095 => x"00002b92",
         11096 => x"00002b98",
         11097 => x"00002b9e",
         11098 => x"00002ba4",
         11099 => x"00004382",
         11100 => x"00004388",
         11101 => x"0000438e",
         11102 => x"00004394",
         11103 => x"0000439a",
         11104 => x"000049b9",
         11105 => x"00004ab9",
         11106 => x"00004bca",
         11107 => x"00004e22",
         11108 => x"00004aa1",
         11109 => x"0000488e",
         11110 => x"00004c92",
         11111 => x"00004df3",
         11112 => x"00004cd5",
         11113 => x"00004d6b",
         11114 => x"00004cf1",
         11115 => x"00004b74",
         11116 => x"0000488e",
         11117 => x"00004bca",
         11118 => x"00004bf3",
         11119 => x"00004c92",
         11120 => x"0000488e",
         11121 => x"0000488e",
         11122 => x"00004cf1",
         11123 => x"00004d6b",
         11124 => x"00004df3",
         11125 => x"00004e22",
         11126 => x"00000e31",
         11127 => x"0000171a",
         11128 => x"0000171a",
         11129 => x"00000e60",
         11130 => x"0000171a",
         11131 => x"0000171a",
         11132 => x"0000171a",
         11133 => x"0000171a",
         11134 => x"0000171a",
         11135 => x"0000171a",
         11136 => x"0000171a",
         11137 => x"00000e1d",
         11138 => x"0000171a",
         11139 => x"00000e48",
         11140 => x"00000e78",
         11141 => x"0000171a",
         11142 => x"0000171a",
         11143 => x"0000171a",
         11144 => x"0000171a",
         11145 => x"0000171a",
         11146 => x"0000171a",
         11147 => x"0000171a",
         11148 => x"0000171a",
         11149 => x"0000171a",
         11150 => x"0000171a",
         11151 => x"0000171a",
         11152 => x"0000171a",
         11153 => x"0000171a",
         11154 => x"0000171a",
         11155 => x"0000171a",
         11156 => x"0000171a",
         11157 => x"0000171a",
         11158 => x"0000171a",
         11159 => x"0000171a",
         11160 => x"0000171a",
         11161 => x"0000171a",
         11162 => x"0000171a",
         11163 => x"0000171a",
         11164 => x"0000171a",
         11165 => x"0000171a",
         11166 => x"0000171a",
         11167 => x"0000171a",
         11168 => x"0000171a",
         11169 => x"0000171a",
         11170 => x"0000171a",
         11171 => x"0000171a",
         11172 => x"0000171a",
         11173 => x"0000171a",
         11174 => x"0000171a",
         11175 => x"0000171a",
         11176 => x"0000171a",
         11177 => x"00000fa8",
         11178 => x"0000171a",
         11179 => x"0000171a",
         11180 => x"0000171a",
         11181 => x"0000171a",
         11182 => x"00001116",
         11183 => x"0000171a",
         11184 => x"0000171a",
         11185 => x"0000171a",
         11186 => x"0000171a",
         11187 => x"0000171a",
         11188 => x"0000171a",
         11189 => x"0000171a",
         11190 => x"0000171a",
         11191 => x"0000171a",
         11192 => x"0000171a",
         11193 => x"00000ed8",
         11194 => x"0000103f",
         11195 => x"00000eaf",
         11196 => x"00000eaf",
         11197 => x"00000eaf",
         11198 => x"0000171a",
         11199 => x"0000103f",
         11200 => x"0000171a",
         11201 => x"0000171a",
         11202 => x"00000e98",
         11203 => x"0000171a",
         11204 => x"0000171a",
         11205 => x"000010ec",
         11206 => x"000010f7",
         11207 => x"0000171a",
         11208 => x"0000171a",
         11209 => x"00000f11",
         11210 => x"0000171a",
         11211 => x"0000111f",
         11212 => x"0000171a",
         11213 => x"0000171a",
         11214 => x"00001116",
         11215 => x"64696e69",
         11216 => x"74000000",
         11217 => x"64696f63",
         11218 => x"746c0000",
         11219 => x"66696e69",
         11220 => x"74000000",
         11221 => x"666c6f61",
         11222 => x"64000000",
         11223 => x"66657865",
         11224 => x"63000000",
         11225 => x"6d636c65",
         11226 => x"61720000",
         11227 => x"6d636f70",
         11228 => x"79000000",
         11229 => x"6d646966",
         11230 => x"66000000",
         11231 => x"6d64756d",
         11232 => x"70000000",
         11233 => x"6d656200",
         11234 => x"6d656800",
         11235 => x"6d657700",
         11236 => x"68696400",
         11237 => x"68696500",
         11238 => x"68666400",
         11239 => x"68666500",
         11240 => x"63616c6c",
         11241 => x"00000000",
         11242 => x"6a6d7000",
         11243 => x"72657374",
         11244 => x"61727400",
         11245 => x"72657365",
         11246 => x"74000000",
         11247 => x"696e666f",
         11248 => x"00000000",
         11249 => x"74657374",
         11250 => x"00000000",
         11251 => x"74626173",
         11252 => x"69630000",
         11253 => x"6d626173",
         11254 => x"69630000",
         11255 => x"6b696c6f",
         11256 => x"00000000",
         11257 => x"65640000",
         11258 => x"4469736b",
         11259 => x"20457272",
         11260 => x"6f720000",
         11261 => x"496e7465",
         11262 => x"726e616c",
         11263 => x"20657272",
         11264 => x"6f722e00",
         11265 => x"4469736b",
         11266 => x"206e6f74",
         11267 => x"20726561",
         11268 => x"64792e00",
         11269 => x"4e6f2066",
         11270 => x"696c6520",
         11271 => x"666f756e",
         11272 => x"642e0000",
         11273 => x"4e6f2070",
         11274 => x"61746820",
         11275 => x"666f756e",
         11276 => x"642e0000",
         11277 => x"496e7661",
         11278 => x"6c696420",
         11279 => x"66696c65",
         11280 => x"6e616d65",
         11281 => x"2e000000",
         11282 => x"41636365",
         11283 => x"73732064",
         11284 => x"656e6965",
         11285 => x"642e0000",
         11286 => x"46696c65",
         11287 => x"20616c72",
         11288 => x"65616479",
         11289 => x"20657869",
         11290 => x"7374732e",
         11291 => x"00000000",
         11292 => x"46696c65",
         11293 => x"2068616e",
         11294 => x"646c6520",
         11295 => x"696e7661",
         11296 => x"6c69642e",
         11297 => x"00000000",
         11298 => x"53442069",
         11299 => x"73207772",
         11300 => x"69746520",
         11301 => x"70726f74",
         11302 => x"65637465",
         11303 => x"642e0000",
         11304 => x"44726976",
         11305 => x"65206e75",
         11306 => x"6d626572",
         11307 => x"20697320",
         11308 => x"696e7661",
         11309 => x"6c69642e",
         11310 => x"00000000",
         11311 => x"4469736b",
         11312 => x"206e6f74",
         11313 => x"20656e61",
         11314 => x"626c6564",
         11315 => x"2e000000",
         11316 => x"4e6f2063",
         11317 => x"6f6d7061",
         11318 => x"7469626c",
         11319 => x"65206669",
         11320 => x"6c657379",
         11321 => x"7374656d",
         11322 => x"20666f75",
         11323 => x"6e64206f",
         11324 => x"6e206469",
         11325 => x"736b2e00",
         11326 => x"466f726d",
         11327 => x"61742061",
         11328 => x"626f7274",
         11329 => x"65642e00",
         11330 => x"54696d65",
         11331 => x"6f75742c",
         11332 => x"206f7065",
         11333 => x"72617469",
         11334 => x"6f6e2063",
         11335 => x"616e6365",
         11336 => x"6c6c6564",
         11337 => x"2e000000",
         11338 => x"46696c65",
         11339 => x"20697320",
         11340 => x"6c6f636b",
         11341 => x"65642e00",
         11342 => x"496e7375",
         11343 => x"66666963",
         11344 => x"69656e74",
         11345 => x"206d656d",
         11346 => x"6f72792e",
         11347 => x"00000000",
         11348 => x"546f6f20",
         11349 => x"6d616e79",
         11350 => x"206f7065",
         11351 => x"6e206669",
         11352 => x"6c65732e",
         11353 => x"00000000",
         11354 => x"50617261",
         11355 => x"6d657465",
         11356 => x"72732069",
         11357 => x"6e636f72",
         11358 => x"72656374",
         11359 => x"2e000000",
         11360 => x"53756363",
         11361 => x"6573732e",
         11362 => x"00000000",
         11363 => x"556e6b6e",
         11364 => x"6f776e20",
         11365 => x"6572726f",
         11366 => x"722e0000",
         11367 => x"0a256c75",
         11368 => x"20627974",
         11369 => x"65732025",
         11370 => x"73206174",
         11371 => x"20256c75",
         11372 => x"20627974",
         11373 => x"65732f73",
         11374 => x"65632e0a",
         11375 => x"00000000",
         11376 => x"72656164",
         11377 => x"00000000",
         11378 => x"2530386c",
         11379 => x"58000000",
         11380 => x"3a202000",
         11381 => x"25303458",
         11382 => x"00000000",
         11383 => x"20202020",
         11384 => x"20202020",
         11385 => x"00000000",
         11386 => x"25303258",
         11387 => x"00000000",
         11388 => x"20200000",
         11389 => x"207c0000",
         11390 => x"7c000000",
         11391 => x"5a505554",
         11392 => x"41000000",
         11393 => x"0a2a2a20",
         11394 => x"25732028",
         11395 => x"00000000",
         11396 => x"30322f30",
         11397 => x"352f3230",
         11398 => x"32300000",
         11399 => x"76312e35",
         11400 => x"32000000",
         11401 => x"205a5055",
         11402 => x"2c207265",
         11403 => x"76202530",
         11404 => x"32782920",
         11405 => x"25732025",
         11406 => x"73202a2a",
         11407 => x"0a0a0000",
         11408 => x"5a505554",
         11409 => x"4120496e",
         11410 => x"74657272",
         11411 => x"75707420",
         11412 => x"48616e64",
         11413 => x"6c657200",
         11414 => x"54696d65",
         11415 => x"7220696e",
         11416 => x"74657272",
         11417 => x"75707400",
         11418 => x"50533220",
         11419 => x"696e7465",
         11420 => x"72727570",
         11421 => x"74000000",
         11422 => x"494f4354",
         11423 => x"4c205244",
         11424 => x"20696e74",
         11425 => x"65727275",
         11426 => x"70740000",
         11427 => x"494f4354",
         11428 => x"4c205752",
         11429 => x"20696e74",
         11430 => x"65727275",
         11431 => x"70740000",
         11432 => x"55415254",
         11433 => x"30205258",
         11434 => x"20696e74",
         11435 => x"65727275",
         11436 => x"70740000",
         11437 => x"55415254",
         11438 => x"30205458",
         11439 => x"20696e74",
         11440 => x"65727275",
         11441 => x"70740000",
         11442 => x"55415254",
         11443 => x"31205258",
         11444 => x"20696e74",
         11445 => x"65727275",
         11446 => x"70740000",
         11447 => x"55415254",
         11448 => x"31205458",
         11449 => x"20696e74",
         11450 => x"65727275",
         11451 => x"70740000",
         11452 => x"53657474",
         11453 => x"696e6720",
         11454 => x"75702074",
         11455 => x"696d6572",
         11456 => x"2e2e2e00",
         11457 => x"456e6162",
         11458 => x"6c696e67",
         11459 => x"2074696d",
         11460 => x"65722e2e",
         11461 => x"2e000000",
         11462 => x"6175746f",
         11463 => x"65786563",
         11464 => x"2e626174",
         11465 => x"00000000",
         11466 => x"7a707574",
         11467 => x"612e6873",
         11468 => x"74000000",
         11469 => x"303a0000",
         11470 => x"4661696c",
         11471 => x"65642074",
         11472 => x"6f20696e",
         11473 => x"69746961",
         11474 => x"6c697365",
         11475 => x"20736420",
         11476 => x"63617264",
         11477 => x"20302c20",
         11478 => x"706c6561",
         11479 => x"73652069",
         11480 => x"6e697420",
         11481 => x"6d616e75",
         11482 => x"616c6c79",
         11483 => x"2e000000",
         11484 => x"2a200000",
         11485 => x"42616420",
         11486 => x"6469736b",
         11487 => x"20696421",
         11488 => x"00000000",
         11489 => x"496e6974",
         11490 => x"69616c69",
         11491 => x"7365642e",
         11492 => x"00000000",
         11493 => x"4661696c",
         11494 => x"65642074",
         11495 => x"6f20696e",
         11496 => x"69746961",
         11497 => x"6c697365",
         11498 => x"2e000000",
         11499 => x"72633d25",
         11500 => x"640a0000",
         11501 => x"25753a00",
         11502 => x"436c6561",
         11503 => x"72696e67",
         11504 => x"2e2e2e2e",
         11505 => x"00000000",
         11506 => x"436f7079",
         11507 => x"696e672e",
         11508 => x"2e2e0000",
         11509 => x"436f6d70",
         11510 => x"6172696e",
         11511 => x"672e2e2e",
         11512 => x"00000000",
         11513 => x"2530386c",
         11514 => x"78282530",
         11515 => x"3878292d",
         11516 => x"3e253038",
         11517 => x"6c782825",
         11518 => x"30387829",
         11519 => x"0a000000",
         11520 => x"44756d70",
         11521 => x"204d656d",
         11522 => x"6f727900",
         11523 => x"0a436f6d",
         11524 => x"706c6574",
         11525 => x"652e0000",
         11526 => x"2530386c",
         11527 => x"58202530",
         11528 => x"32582d00",
         11529 => x"3f3f3f00",
         11530 => x"2530386c",
         11531 => x"58202530",
         11532 => x"34582d00",
         11533 => x"2530386c",
         11534 => x"58202530",
         11535 => x"386c582d",
         11536 => x"00000000",
         11537 => x"44697361",
         11538 => x"626c696e",
         11539 => x"6720696e",
         11540 => x"74657272",
         11541 => x"75707473",
         11542 => x"00000000",
         11543 => x"456e6162",
         11544 => x"6c696e67",
         11545 => x"20696e74",
         11546 => x"65727275",
         11547 => x"70747300",
         11548 => x"44697361",
         11549 => x"626c6564",
         11550 => x"20756172",
         11551 => x"74206669",
         11552 => x"666f0000",
         11553 => x"456e6162",
         11554 => x"6c696e67",
         11555 => x"20756172",
         11556 => x"74206669",
         11557 => x"666f0000",
         11558 => x"45786563",
         11559 => x"7574696e",
         11560 => x"6720636f",
         11561 => x"64652040",
         11562 => x"20253038",
         11563 => x"6c78202e",
         11564 => x"2e2e0a00",
         11565 => x"43616c6c",
         11566 => x"696e6720",
         11567 => x"636f6465",
         11568 => x"20402025",
         11569 => x"30386c78",
         11570 => x"202e2e2e",
         11571 => x"0a000000",
         11572 => x"43616c6c",
         11573 => x"20726574",
         11574 => x"75726e65",
         11575 => x"6420636f",
         11576 => x"64652028",
         11577 => x"2564292e",
         11578 => x"0a000000",
         11579 => x"52657374",
         11580 => x"61727469",
         11581 => x"6e672061",
         11582 => x"70706c69",
         11583 => x"63617469",
         11584 => x"6f6e2e2e",
         11585 => x"2e000000",
         11586 => x"436f6c64",
         11587 => x"20726562",
         11588 => x"6f6f7469",
         11589 => x"6e672e2e",
         11590 => x"2e000000",
         11591 => x"5a505500",
         11592 => x"62696e00",
         11593 => x"25643a5c",
         11594 => x"25735c25",
         11595 => x"732e2573",
         11596 => x"00000000",
         11597 => x"25643a5c",
         11598 => x"25735c25",
         11599 => x"73000000",
         11600 => x"25643a5c",
         11601 => x"25730000",
         11602 => x"42616420",
         11603 => x"636f6d6d",
         11604 => x"616e642e",
         11605 => x"00000000",
         11606 => x"52756e6e",
         11607 => x"696e672e",
         11608 => x"2e2e0000",
         11609 => x"456e6162",
         11610 => x"6c696e67",
         11611 => x"20696e74",
         11612 => x"65727275",
         11613 => x"7074732e",
         11614 => x"2e2e0000",
         11615 => x"25642f25",
         11616 => x"642f2564",
         11617 => x"2025643a",
         11618 => x"25643a25",
         11619 => x"642e2564",
         11620 => x"25640a00",
         11621 => x"536f4320",
         11622 => x"436f6e66",
         11623 => x"69677572",
         11624 => x"6174696f",
         11625 => x"6e000000",
         11626 => x"20286672",
         11627 => x"6f6d2053",
         11628 => x"6f432063",
         11629 => x"6f6e6669",
         11630 => x"67290000",
         11631 => x"3a0a4465",
         11632 => x"76696365",
         11633 => x"7320696d",
         11634 => x"706c656d",
         11635 => x"656e7465",
         11636 => x"643a0a00",
         11637 => x"20202020",
         11638 => x"57422053",
         11639 => x"4452414d",
         11640 => x"20202825",
         11641 => x"3038583a",
         11642 => x"25303858",
         11643 => x"292e0a00",
         11644 => x"20202020",
         11645 => x"53445241",
         11646 => x"4d202020",
         11647 => x"20202825",
         11648 => x"3038583a",
         11649 => x"25303858",
         11650 => x"292e0a00",
         11651 => x"20202020",
         11652 => x"494e534e",
         11653 => x"20425241",
         11654 => x"4d202825",
         11655 => x"3038583a",
         11656 => x"25303858",
         11657 => x"292e0a00",
         11658 => x"20202020",
         11659 => x"4252414d",
         11660 => x"20202020",
         11661 => x"20202825",
         11662 => x"3038583a",
         11663 => x"25303858",
         11664 => x"292e0a00",
         11665 => x"20202020",
         11666 => x"52414d20",
         11667 => x"20202020",
         11668 => x"20202825",
         11669 => x"3038583a",
         11670 => x"25303858",
         11671 => x"292e0a00",
         11672 => x"20202020",
         11673 => x"53442043",
         11674 => x"41524420",
         11675 => x"20202844",
         11676 => x"65766963",
         11677 => x"6573203d",
         11678 => x"25303264",
         11679 => x"292e0a00",
         11680 => x"20202020",
         11681 => x"54494d45",
         11682 => x"52312020",
         11683 => x"20202854",
         11684 => x"696d6572",
         11685 => x"7320203d",
         11686 => x"25303264",
         11687 => x"292e0a00",
         11688 => x"20202020",
         11689 => x"494e5452",
         11690 => x"20435452",
         11691 => x"4c202843",
         11692 => x"68616e6e",
         11693 => x"656c733d",
         11694 => x"25303264",
         11695 => x"292e0a00",
         11696 => x"20202020",
         11697 => x"57495348",
         11698 => x"424f4e45",
         11699 => x"20425553",
         11700 => x"0a000000",
         11701 => x"20202020",
         11702 => x"57422049",
         11703 => x"32430a00",
         11704 => x"20202020",
         11705 => x"494f4354",
         11706 => x"4c0a0000",
         11707 => x"20202020",
         11708 => x"5053320a",
         11709 => x"00000000",
         11710 => x"20202020",
         11711 => x"5350490a",
         11712 => x"00000000",
         11713 => x"41646472",
         11714 => x"65737365",
         11715 => x"733a0a00",
         11716 => x"20202020",
         11717 => x"43505520",
         11718 => x"52657365",
         11719 => x"74205665",
         11720 => x"63746f72",
         11721 => x"20416464",
         11722 => x"72657373",
         11723 => x"203d2025",
         11724 => x"3038580a",
         11725 => x"00000000",
         11726 => x"20202020",
         11727 => x"43505520",
         11728 => x"4d656d6f",
         11729 => x"72792053",
         11730 => x"74617274",
         11731 => x"20416464",
         11732 => x"72657373",
         11733 => x"203d2025",
         11734 => x"3038580a",
         11735 => x"00000000",
         11736 => x"20202020",
         11737 => x"53746163",
         11738 => x"6b205374",
         11739 => x"61727420",
         11740 => x"41646472",
         11741 => x"65737320",
         11742 => x"20202020",
         11743 => x"203d2025",
         11744 => x"3038580a",
         11745 => x"00000000",
         11746 => x"4d697363",
         11747 => x"3a0a0000",
         11748 => x"20202020",
         11749 => x"5a505520",
         11750 => x"49642020",
         11751 => x"20202020",
         11752 => x"20202020",
         11753 => x"20202020",
         11754 => x"20202020",
         11755 => x"203d2025",
         11756 => x"3034580a",
         11757 => x"00000000",
         11758 => x"20202020",
         11759 => x"53797374",
         11760 => x"656d2043",
         11761 => x"6c6f636b",
         11762 => x"20467265",
         11763 => x"71202020",
         11764 => x"20202020",
         11765 => x"203d2025",
         11766 => x"642e2530",
         11767 => x"34644d48",
         11768 => x"7a0a0000",
         11769 => x"20202020",
         11770 => x"53445241",
         11771 => x"4d20436c",
         11772 => x"6f636b20",
         11773 => x"46726571",
         11774 => x"20202020",
         11775 => x"20202020",
         11776 => x"203d2025",
         11777 => x"642e2530",
         11778 => x"34644d48",
         11779 => x"7a0a0000",
         11780 => x"20202020",
         11781 => x"57697368",
         11782 => x"626f6e65",
         11783 => x"20534452",
         11784 => x"414d2043",
         11785 => x"6c6f636b",
         11786 => x"20467265",
         11787 => x"713d2025",
         11788 => x"642e2530",
         11789 => x"34644d48",
         11790 => x"7a0a0000",
         11791 => x"536d616c",
         11792 => x"6c000000",
         11793 => x"4d656469",
         11794 => x"756d0000",
         11795 => x"466c6578",
         11796 => x"00000000",
         11797 => x"45564f00",
         11798 => x"45564f6d",
         11799 => x"696e0000",
         11800 => x"556e6b6e",
         11801 => x"6f776e00",
         11802 => x"000099c4",
         11803 => x"01000000",
         11804 => x"00000002",
         11805 => x"000099c0",
         11806 => x"01000000",
         11807 => x"00000003",
         11808 => x"000099bc",
         11809 => x"01000000",
         11810 => x"00000004",
         11811 => x"000099b8",
         11812 => x"01000000",
         11813 => x"00000005",
         11814 => x"000099b4",
         11815 => x"01000000",
         11816 => x"00000006",
         11817 => x"000099b0",
         11818 => x"01000000",
         11819 => x"00000007",
         11820 => x"000099ac",
         11821 => x"01000000",
         11822 => x"00000001",
         11823 => x"000099a8",
         11824 => x"01000000",
         11825 => x"00000008",
         11826 => x"000099a4",
         11827 => x"01000000",
         11828 => x"0000000b",
         11829 => x"000099a0",
         11830 => x"01000000",
         11831 => x"00000009",
         11832 => x"0000999c",
         11833 => x"01000000",
         11834 => x"0000000a",
         11835 => x"00009998",
         11836 => x"04000000",
         11837 => x"0000000d",
         11838 => x"00009994",
         11839 => x"04000000",
         11840 => x"0000000c",
         11841 => x"00009990",
         11842 => x"04000000",
         11843 => x"0000000e",
         11844 => x"0000998c",
         11845 => x"03000000",
         11846 => x"0000000f",
         11847 => x"00009988",
         11848 => x"04000000",
         11849 => x"0000000f",
         11850 => x"00009984",
         11851 => x"04000000",
         11852 => x"00000010",
         11853 => x"00009980",
         11854 => x"04000000",
         11855 => x"00000011",
         11856 => x"0000997c",
         11857 => x"03000000",
         11858 => x"00000012",
         11859 => x"00009978",
         11860 => x"03000000",
         11861 => x"00000013",
         11862 => x"00009974",
         11863 => x"03000000",
         11864 => x"00000014",
         11865 => x"00009970",
         11866 => x"03000000",
         11867 => x"00000015",
         11868 => x"1b5b4400",
         11869 => x"1b5b4300",
         11870 => x"1b5b4200",
         11871 => x"1b5b4100",
         11872 => x"1b5b367e",
         11873 => x"1b5b357e",
         11874 => x"1b5b347e",
         11875 => x"1b304600",
         11876 => x"1b5b337e",
         11877 => x"1b5b327e",
         11878 => x"1b5b317e",
         11879 => x"10000000",
         11880 => x"0e000000",
         11881 => x"0d000000",
         11882 => x"0b000000",
         11883 => x"08000000",
         11884 => x"06000000",
         11885 => x"05000000",
         11886 => x"04000000",
         11887 => x"03000000",
         11888 => x"02000000",
         11889 => x"01000000",
         11890 => x"68697374",
         11891 => x"6f727900",
         11892 => x"68697374",
         11893 => x"00000000",
         11894 => x"21000000",
         11895 => x"2530346c",
         11896 => x"75202025",
         11897 => x"730a0000",
         11898 => x"4661696c",
         11899 => x"65642074",
         11900 => x"6f207265",
         11901 => x"73657420",
         11902 => x"74686520",
         11903 => x"68697374",
         11904 => x"6f727920",
         11905 => x"66696c65",
         11906 => x"20746f20",
         11907 => x"454f462e",
         11908 => x"00000000",
         11909 => x"43616e6e",
         11910 => x"6f74206f",
         11911 => x"70656e2f",
         11912 => x"63726561",
         11913 => x"74652068",
         11914 => x"6973746f",
         11915 => x"72792066",
         11916 => x"696c652c",
         11917 => x"20646973",
         11918 => x"61626c69",
         11919 => x"6e672e00",
         11920 => x"53440000",
         11921 => x"222a2b2c",
         11922 => x"3a3b3c3d",
         11923 => x"3e3f5b5d",
         11924 => x"7c7f0000",
         11925 => x"46415400",
         11926 => x"46415433",
         11927 => x"32000000",
         11928 => x"ebfe904d",
         11929 => x"53444f53",
         11930 => x"352e3000",
         11931 => x"4e4f204e",
         11932 => x"414d4520",
         11933 => x"20202046",
         11934 => x"41543332",
         11935 => x"20202000",
         11936 => x"4e4f204e",
         11937 => x"414d4520",
         11938 => x"20202046",
         11939 => x"41542020",
         11940 => x"20202000",
         11941 => x"00009a40",
         11942 => x"00000000",
         11943 => x"00000000",
         11944 => x"00000000",
         11945 => x"809a4541",
         11946 => x"8e418f80",
         11947 => x"45454549",
         11948 => x"49498e8f",
         11949 => x"9092924f",
         11950 => x"994f5555",
         11951 => x"59999a9b",
         11952 => x"9c9d9e9f",
         11953 => x"41494f55",
         11954 => x"a5a5a6a7",
         11955 => x"a8a9aaab",
         11956 => x"acadaeaf",
         11957 => x"b0b1b2b3",
         11958 => x"b4b5b6b7",
         11959 => x"b8b9babb",
         11960 => x"bcbdbebf",
         11961 => x"c0c1c2c3",
         11962 => x"c4c5c6c7",
         11963 => x"c8c9cacb",
         11964 => x"cccdcecf",
         11965 => x"d0d1d2d3",
         11966 => x"d4d5d6d7",
         11967 => x"d8d9dadb",
         11968 => x"dcdddedf",
         11969 => x"e0e1e2e3",
         11970 => x"e4e5e6e7",
         11971 => x"e8e9eaeb",
         11972 => x"ecedeeef",
         11973 => x"f0f1f2f3",
         11974 => x"f4f5f6f7",
         11975 => x"f8f9fafb",
         11976 => x"fcfdfeff",
         11977 => x"2b2e2c3b",
         11978 => x"3d5b5d2f",
         11979 => x"5c222a3a",
         11980 => x"3c3e3f7c",
         11981 => x"7f000000",
         11982 => x"00010004",
         11983 => x"00100040",
         11984 => x"01000200",
         11985 => x"00000000",
         11986 => x"00010002",
         11987 => x"00040008",
         11988 => x"00100020",
         11989 => x"00000000",
         11990 => x"00000000",
         11991 => x"00008f3c",
         11992 => x"01020100",
         11993 => x"00000000",
         11994 => x"00000000",
         11995 => x"00008f44",
         11996 => x"01040100",
         11997 => x"00000000",
         11998 => x"00000000",
         11999 => x"00008f4c",
         12000 => x"01140300",
         12001 => x"00000000",
         12002 => x"00000000",
         12003 => x"00008f54",
         12004 => x"012b0300",
         12005 => x"00000000",
         12006 => x"00000000",
         12007 => x"00008f5c",
         12008 => x"01300300",
         12009 => x"00000000",
         12010 => x"00000000",
         12011 => x"00008f64",
         12012 => x"013c0400",
         12013 => x"00000000",
         12014 => x"00000000",
         12015 => x"00008f6c",
         12016 => x"013d0400",
         12017 => x"00000000",
         12018 => x"00000000",
         12019 => x"00008f74",
         12020 => x"013f0400",
         12021 => x"00000000",
         12022 => x"00000000",
         12023 => x"00008f7c",
         12024 => x"01400400",
         12025 => x"00000000",
         12026 => x"00000000",
         12027 => x"00008f84",
         12028 => x"01410400",
         12029 => x"00000000",
         12030 => x"00000000",
         12031 => x"00008f88",
         12032 => x"01420400",
         12033 => x"00000000",
         12034 => x"00000000",
         12035 => x"00008f8c",
         12036 => x"01430400",
         12037 => x"00000000",
         12038 => x"00000000",
         12039 => x"00008f90",
         12040 => x"01500500",
         12041 => x"00000000",
         12042 => x"00000000",
         12043 => x"00008f94",
         12044 => x"01510500",
         12045 => x"00000000",
         12046 => x"00000000",
         12047 => x"00008f98",
         12048 => x"01540500",
         12049 => x"00000000",
         12050 => x"00000000",
         12051 => x"00008f9c",
         12052 => x"01550500",
         12053 => x"00000000",
         12054 => x"00000000",
         12055 => x"00008fa0",
         12056 => x"01790700",
         12057 => x"00000000",
         12058 => x"00000000",
         12059 => x"00008fa8",
         12060 => x"01780700",
         12061 => x"00000000",
         12062 => x"00000000",
         12063 => x"00008fac",
         12064 => x"01820800",
         12065 => x"00000000",
         12066 => x"00000000",
         12067 => x"00008fb4",
         12068 => x"01830800",
         12069 => x"00000000",
         12070 => x"00000000",
         12071 => x"00008fbc",
         12072 => x"01850800",
         12073 => x"00000000",
         12074 => x"00000000",
         12075 => x"00008fc4",
         12076 => x"01870800",
         12077 => x"00000000",
         12078 => x"00000000",
         12079 => x"00008fcc",
         12080 => x"018c0900",
         12081 => x"00000000",
         12082 => x"00000000",
         12083 => x"00008fd4",
         12084 => x"018d0900",
         12085 => x"00000000",
         12086 => x"00000000",
         12087 => x"00008fdc",
         12088 => x"018e0900",
         12089 => x"00000000",
         12090 => x"00000000",
         12091 => x"00008fe4",
         12092 => x"018f0900",
         12093 => x"00000000",
         12094 => x"00000000",
         12095 => x"00000000",
         12096 => x"00000000",
         12097 => x"00007fff",
         12098 => x"00000000",
         12099 => x"00007fff",
         12100 => x"00010000",
         12101 => x"00007fff",
         12102 => x"00010000",
         12103 => x"00810000",
         12104 => x"01000000",
         12105 => x"017fffff",
         12106 => x"00000000",
         12107 => x"00000000",
         12108 => x"00007800",
         12109 => x"00000000",
         12110 => x"05f5e100",
         12111 => x"05f5e100",
         12112 => x"05f5e100",
         12113 => x"00000000",
         12114 => x"01010101",
         12115 => x"01010101",
         12116 => x"01011001",
         12117 => x"01000000",
         12118 => x"00000000",
         12119 => x"00000000",
         12120 => x"00000000",
         12121 => x"00000000",
         12122 => x"00000000",
         12123 => x"00000000",
         12124 => x"00000000",
         12125 => x"00000000",
         12126 => x"00000000",
         12127 => x"00000000",
         12128 => x"00000000",
         12129 => x"00000000",
         12130 => x"00000000",
         12131 => x"00000000",
         12132 => x"00000000",
         12133 => x"00000000",
         12134 => x"00000000",
         12135 => x"00000000",
         12136 => x"00000000",
         12137 => x"00000000",
         12138 => x"00000000",
         12139 => x"00000000",
         12140 => x"00000000",
         12141 => x"00000000",
         12142 => x"000099c8",
         12143 => x"01000000",
         12144 => x"000099d0",
         12145 => x"01000000",
         12146 => x"000099d8",
         12147 => x"02000000",
         12148 => x"00000000",
         12149 => x"00000000",
         12150 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

