-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b87fa",
          2049 => x"f80d0b0b",
          2050 => x"0b93e904",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b93",
          2121 => x"cd040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b93b0",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b83bd",
          2210 => x"f4738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"93b50400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b0bac",
          2219 => x"cc2d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b0bab",
          2227 => x"ab2d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"96040b0b",
          2317 => x"0b8ca604",
          2318 => x"0b0b0b8c",
          2319 => x"b6040b0b",
          2320 => x"0b8cc604",
          2321 => x"0b0b0b8c",
          2322 => x"d6040b0b",
          2323 => x"0b8ce604",
          2324 => x"0b0b0b8c",
          2325 => x"f6040b0b",
          2326 => x"0b8d8604",
          2327 => x"0b0b0b8d",
          2328 => x"96040b0b",
          2329 => x"0b8da604",
          2330 => x"0b0b0b8d",
          2331 => x"b6040b0b",
          2332 => x"0b8dc604",
          2333 => x"0b0b0b8d",
          2334 => x"d7040b0b",
          2335 => x"0b8de804",
          2336 => x"0b0b0b8d",
          2337 => x"f9040b0b",
          2338 => x"0b8e8a04",
          2339 => x"0b0b0b8e",
          2340 => x"9b040b0b",
          2341 => x"0b8eac04",
          2342 => x"0b0b0b8e",
          2343 => x"bd040b0b",
          2344 => x"0b8ece04",
          2345 => x"0b0b0b8e",
          2346 => x"df040b0b",
          2347 => x"0b8ef004",
          2348 => x"0b0b0b8f",
          2349 => x"81040b0b",
          2350 => x"0b8f9204",
          2351 => x"0b0b0b8f",
          2352 => x"a3040b0b",
          2353 => x"0b8fb404",
          2354 => x"0b0b0b8f",
          2355 => x"c5040b0b",
          2356 => x"0b8fd604",
          2357 => x"0b0b0b8f",
          2358 => x"e7040b0b",
          2359 => x"0b8ff804",
          2360 => x"0b0b0b90",
          2361 => x"89040b0b",
          2362 => x"0b909a04",
          2363 => x"0b0b0b90",
          2364 => x"ab040b0b",
          2365 => x"0b90bc04",
          2366 => x"0b0b0b90",
          2367 => x"cd040b0b",
          2368 => x"0b90de04",
          2369 => x"0b0b0b90",
          2370 => x"ef040b0b",
          2371 => x"0b918004",
          2372 => x"0b0b0b91",
          2373 => x"91040b0b",
          2374 => x"0b91a204",
          2375 => x"0b0b0b91",
          2376 => x"b3040b0b",
          2377 => x"0b91c404",
          2378 => x"0b0b0b91",
          2379 => x"d5040b0b",
          2380 => x"0b91e604",
          2381 => x"0b0b0b91",
          2382 => x"f7040b0b",
          2383 => x"0b928804",
          2384 => x"0b0b0b92",
          2385 => x"99040b0b",
          2386 => x"0b92aa04",
          2387 => x"0b0b0b92",
          2388 => x"bb040b0b",
          2389 => x"0b92cb04",
          2390 => x"0b0b0b92",
          2391 => x"dc040b0b",
          2392 => x"0b92ed04",
          2393 => x"0b0b0b92",
          2394 => x"fe04ffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0484b9d4",
          2434 => x"0c80d687",
          2435 => x"2d84b9d4",
          2436 => x"0880c080",
          2437 => x"900484b9",
          2438 => x"d40ca2ee",
          2439 => x"2d84b9d4",
          2440 => x"0880c080",
          2441 => x"900484b9",
          2442 => x"d40ca0f3",
          2443 => x"2d84b9d4",
          2444 => x"0880c080",
          2445 => x"900484b9",
          2446 => x"d40ca0e0",
          2447 => x"2d84b9d4",
          2448 => x"0880c080",
          2449 => x"900484b9",
          2450 => x"d40c94a3",
          2451 => x"2d84b9d4",
          2452 => x"0880c080",
          2453 => x"900484b9",
          2454 => x"d40ca1f6",
          2455 => x"2d84b9d4",
          2456 => x"0880c080",
          2457 => x"900484b9",
          2458 => x"d40caf86",
          2459 => x"2d84b9d4",
          2460 => x"0880c080",
          2461 => x"900484b9",
          2462 => x"d40cad82",
          2463 => x"2d84b9d4",
          2464 => x"0880c080",
          2465 => x"900484b9",
          2466 => x"d40c9488",
          2467 => x"2d84b9d4",
          2468 => x"0880c080",
          2469 => x"900484b9",
          2470 => x"d40c95a8",
          2471 => x"2d84b9d4",
          2472 => x"0880c080",
          2473 => x"900484b9",
          2474 => x"d40c95d1",
          2475 => x"2d84b9d4",
          2476 => x"0880c080",
          2477 => x"900484b9",
          2478 => x"d40cb18a",
          2479 => x"2d84b9d4",
          2480 => x"0880c080",
          2481 => x"900484b9",
          2482 => x"d40c80d4",
          2483 => x"ec2d84b9",
          2484 => x"d40880c0",
          2485 => x"80900484",
          2486 => x"b9d40c80",
          2487 => x"d5d12d84",
          2488 => x"b9d40880",
          2489 => x"c0809004",
          2490 => x"84b9d40c",
          2491 => x"80d2a82d",
          2492 => x"84b9d408",
          2493 => x"80c08090",
          2494 => x"0484b9d4",
          2495 => x"0c80d3db",
          2496 => x"2d84b9d4",
          2497 => x"0880c080",
          2498 => x"900484b9",
          2499 => x"d40c82c9",
          2500 => x"ae2d84b9",
          2501 => x"d40880c0",
          2502 => x"80900484",
          2503 => x"b9d40c82",
          2504 => x"e3802d84",
          2505 => x"b9d40880",
          2506 => x"c0809004",
          2507 => x"84b9d40c",
          2508 => x"82d29e2d",
          2509 => x"84b9d408",
          2510 => x"80c08090",
          2511 => x"0484b9d4",
          2512 => x"0c82d7c0",
          2513 => x"2d84b9d4",
          2514 => x"0880c080",
          2515 => x"900484b9",
          2516 => x"d40c82ed",
          2517 => x"9d2d84b9",
          2518 => x"d40880c0",
          2519 => x"80900484",
          2520 => x"b9d40c82",
          2521 => x"faa52d84",
          2522 => x"b9d40880",
          2523 => x"c0809004",
          2524 => x"84b9d40c",
          2525 => x"82df872d",
          2526 => x"84b9d408",
          2527 => x"80c08090",
          2528 => x"0484b9d4",
          2529 => x"0c82f1be",
          2530 => x"2d84b9d4",
          2531 => x"0880c080",
          2532 => x"900484b9",
          2533 => x"d40c82f3",
          2534 => x"8b2d84b9",
          2535 => x"d40880c0",
          2536 => x"80900484",
          2537 => x"b9d40c82",
          2538 => x"f3e02d84",
          2539 => x"b9d40880",
          2540 => x"c0809004",
          2541 => x"84b9d40c",
          2542 => x"8384a22d",
          2543 => x"84b9d408",
          2544 => x"80c08090",
          2545 => x"0484b9d4",
          2546 => x"0c82fee7",
          2547 => x"2d84b9d4",
          2548 => x"0880c080",
          2549 => x"900484b9",
          2550 => x"d40c838b",
          2551 => x"862d84b9",
          2552 => x"d40880c0",
          2553 => x"80900484",
          2554 => x"b9d40c82",
          2555 => x"f5bd2d84",
          2556 => x"b9d40880",
          2557 => x"c0809004",
          2558 => x"84b9d40c",
          2559 => x"8393fd2d",
          2560 => x"84b9d408",
          2561 => x"80c08090",
          2562 => x"0484b9d4",
          2563 => x"0c839588",
          2564 => x"2d84b9d4",
          2565 => x"0880c080",
          2566 => x"900484b9",
          2567 => x"d40c82e5",
          2568 => x"d02d84b9",
          2569 => x"d40880c0",
          2570 => x"80900484",
          2571 => x"b9d40c82",
          2572 => x"e3e72d84",
          2573 => x"b9d40880",
          2574 => x"c0809004",
          2575 => x"84b9d40c",
          2576 => x"82e78e2d",
          2577 => x"84b9d408",
          2578 => x"80c08090",
          2579 => x"0484b9d4",
          2580 => x"0c82f6a7",
          2581 => x"2d84b9d4",
          2582 => x"0880c080",
          2583 => x"900484b9",
          2584 => x"d40c8396",
          2585 => x"9a2d84b9",
          2586 => x"d40880c0",
          2587 => x"80900484",
          2588 => x"b9d40c83",
          2589 => x"99f72d84",
          2590 => x"b9d40880",
          2591 => x"c0809004",
          2592 => x"84b9d40c",
          2593 => x"83a0e92d",
          2594 => x"84b9d408",
          2595 => x"80c08090",
          2596 => x"0484b9d4",
          2597 => x"0c82c6ff",
          2598 => x"2d84b9d4",
          2599 => x"0880c080",
          2600 => x"900484b9",
          2601 => x"d40c83a4",
          2602 => x"922d84b9",
          2603 => x"d40880c0",
          2604 => x"80900484",
          2605 => x"b9d40c83",
          2606 => x"b9932d84",
          2607 => x"b9d40880",
          2608 => x"c0809004",
          2609 => x"84b9d40c",
          2610 => x"83b7c52d",
          2611 => x"84b9d408",
          2612 => x"80c08090",
          2613 => x"0484b9d4",
          2614 => x"0c81f3e3",
          2615 => x"2d84b9d4",
          2616 => x"0880c080",
          2617 => x"900484b9",
          2618 => x"d40c81f4",
          2619 => x"e22d84b9",
          2620 => x"d40880c0",
          2621 => x"80900484",
          2622 => x"b9d40c81",
          2623 => x"f5e12d84",
          2624 => x"b9d40880",
          2625 => x"c0809004",
          2626 => x"84b9d40c",
          2627 => x"80d0aa2d",
          2628 => x"84b9d408",
          2629 => x"80c08090",
          2630 => x"0484b9d4",
          2631 => x"0c80d1fa",
          2632 => x"2d84b9d4",
          2633 => x"0880c080",
          2634 => x"900484b9",
          2635 => x"d40c80d7",
          2636 => x"a52d84b9",
          2637 => x"d40880c0",
          2638 => x"80900484",
          2639 => x"b9d40cb1",
          2640 => x"9a2d84b9",
          2641 => x"d40880c0",
          2642 => x"80900484",
          2643 => x"b9d40c81",
          2644 => x"db812d84",
          2645 => x"b9d40880",
          2646 => x"c0809004",
          2647 => x"84b9d40c",
          2648 => x"81dcbc2d",
          2649 => x"84b9d408",
          2650 => x"80c08090",
          2651 => x"0484b9d4",
          2652 => x"0c81f1bd",
          2653 => x"2d84b9d4",
          2654 => x"0880c080",
          2655 => x"900484b9",
          2656 => x"d40c81d5",
          2657 => x"912d84b9",
          2658 => x"d40880c0",
          2659 => x"8090043c",
          2660 => x"04101010",
          2661 => x"10101010",
          2662 => x"10101010",
          2663 => x"10101010",
          2664 => x"10101010",
          2665 => x"10101010",
          2666 => x"10101010",
          2667 => x"10101010",
          2668 => x"53510400",
          2669 => x"007381ff",
          2670 => x"06738306",
          2671 => x"09810583",
          2672 => x"05101010",
          2673 => x"2b0772fc",
          2674 => x"060c5151",
          2675 => x"04727280",
          2676 => x"728106ff",
          2677 => x"05097206",
          2678 => x"05711052",
          2679 => x"720a100a",
          2680 => x"5372ed38",
          2681 => x"51515351",
          2682 => x"0484b9c8",
          2683 => x"7084d5b4",
          2684 => x"278e3880",
          2685 => x"71708405",
          2686 => x"530c0b0b",
          2687 => x"0b93ec04",
          2688 => x"8c815180",
          2689 => x"ceba0400",
          2690 => x"fc3d0d87",
          2691 => x"3d707084",
          2692 => x"05520856",
          2693 => x"53745284",
          2694 => x"d5ac0851",
          2695 => x"81c53f86",
          2696 => x"3d0d04fa",
          2697 => x"3d0d787a",
          2698 => x"7c851133",
          2699 => x"81328106",
          2700 => x"80732507",
          2701 => x"56585557",
          2702 => x"80527272",
          2703 => x"2e098106",
          2704 => x"80d338ff",
          2705 => x"1477748a",
          2706 => x"32703070",
          2707 => x"72079f2a",
          2708 => x"51555556",
          2709 => x"54807425",
          2710 => x"b7387180",
          2711 => x"2eb23875",
          2712 => x"518efa3f",
          2713 => x"84b9c808",
          2714 => x"5384b9c8",
          2715 => x"08ff2eae",
          2716 => x"3884b9c8",
          2717 => x"08757081",
          2718 => x"055734ff",
          2719 => x"14738a32",
          2720 => x"70307072",
          2721 => x"079f2a51",
          2722 => x"54545473",
          2723 => x"8024cb38",
          2724 => x"80753476",
          2725 => x"527184b9",
          2726 => x"c80c883d",
          2727 => x"0d04800b",
          2728 => x"84b9c80c",
          2729 => x"883d0d04",
          2730 => x"f53d0d7d",
          2731 => x"54860284",
          2732 => x"05990534",
          2733 => x"7356fe0a",
          2734 => x"588e3d88",
          2735 => x"05537e52",
          2736 => x"8d3de405",
          2737 => x"519d3f73",
          2738 => x"19548074",
          2739 => x"348d3d0d",
          2740 => x"04fd3d0d",
          2741 => x"863d8805",
          2742 => x"53765275",
          2743 => x"51853f85",
          2744 => x"3d0d04f1",
          2745 => x"3d0d6163",
          2746 => x"65425d5d",
          2747 => x"80708c1f",
          2748 => x"0c851e33",
          2749 => x"70812a81",
          2750 => x"32810655",
          2751 => x"555bff54",
          2752 => x"727b2e09",
          2753 => x"810680d2",
          2754 => x"387b3357",
          2755 => x"767b2e80",
          2756 => x"c538811c",
          2757 => x"7b810654",
          2758 => x"5c72802e",
          2759 => x"818138d0",
          2760 => x"175f7e89",
          2761 => x"2681a338",
          2762 => x"76b03270",
          2763 => x"30708025",
          2764 => x"51545578",
          2765 => x"ae387280",
          2766 => x"2ea9387a",
          2767 => x"832a7081",
          2768 => x"32810640",
          2769 => x"547e802e",
          2770 => x"9e387a82",
          2771 => x"80075b7b",
          2772 => x"335776ff",
          2773 => x"bd388c1d",
          2774 => x"08547384",
          2775 => x"b9c80c91",
          2776 => x"3d0d047a",
          2777 => x"832a5478",
          2778 => x"10101079",
          2779 => x"10057098",
          2780 => x"2b70982c",
          2781 => x"19708180",
          2782 => x"0a298b0a",
          2783 => x"0570982c",
          2784 => x"525a5b56",
          2785 => x"5f807924",
          2786 => x"81863873",
          2787 => x"81065372",
          2788 => x"ffbd3878",
          2789 => x"7c335858",
          2790 => x"76fef738",
          2791 => x"ffb83976",
          2792 => x"a52e0981",
          2793 => x"06933881",
          2794 => x"73745a5a",
          2795 => x"5b8a7c33",
          2796 => x"585a76fe",
          2797 => x"dd38ff9e",
          2798 => x"397c5276",
          2799 => x"518baf3f",
          2800 => x"7b335776",
          2801 => x"fecc38ff",
          2802 => x"8d397a83",
          2803 => x"2a708106",
          2804 => x"5455788a",
          2805 => x"38817074",
          2806 => x"0640547e",
          2807 => x"9538e017",
          2808 => x"537280d8",
          2809 => x"26973872",
          2810 => x"101083ca",
          2811 => x"84055473",
          2812 => x"080473e0",
          2813 => x"18545980",
          2814 => x"d87327eb",
          2815 => x"387c5276",
          2816 => x"518aeb3f",
          2817 => x"807c3358",
          2818 => x"5b76fe86",
          2819 => x"38fec739",
          2820 => x"80ff59fe",
          2821 => x"f639885a",
          2822 => x"7f608405",
          2823 => x"71087d83",
          2824 => x"ffcf065e",
          2825 => x"58415484",
          2826 => x"b9d85e79",
          2827 => x"52755193",
          2828 => x"9a3f84b9",
          2829 => x"c80881ff",
          2830 => x"0684b9c8",
          2831 => x"0818df05",
          2832 => x"56537289",
          2833 => x"26883884",
          2834 => x"b9c808b0",
          2835 => x"0555747e",
          2836 => x"70810540",
          2837 => x"34795275",
          2838 => x"5190ca3f",
          2839 => x"84b9c808",
          2840 => x"5684b9c8",
          2841 => x"08c5387d",
          2842 => x"84b9d831",
          2843 => x"982b7bb2",
          2844 => x"0640567e",
          2845 => x"802e8f38",
          2846 => x"77848080",
          2847 => x"29fc8080",
          2848 => x"0570902c",
          2849 => x"59557a86",
          2850 => x"2a708106",
          2851 => x"555f7380",
          2852 => x"2e9e3877",
          2853 => x"84808029",
          2854 => x"f8808005",
          2855 => x"5379902e",
          2856 => x"8b387784",
          2857 => x"808029fc",
          2858 => x"80800553",
          2859 => x"72902c58",
          2860 => x"7a832a70",
          2861 => x"81065455",
          2862 => x"72802e9e",
          2863 => x"3875982c",
          2864 => x"7081ff06",
          2865 => x"54547873",
          2866 => x"2486cc38",
          2867 => x"7a83fff7",
          2868 => x"0670832a",
          2869 => x"71862a41",
          2870 => x"565b7481",
          2871 => x"06547380",
          2872 => x"2e85f038",
          2873 => x"77793190",
          2874 => x"2b70902c",
          2875 => x"7c838006",
          2876 => x"56595373",
          2877 => x"802e8596",
          2878 => x"387a812a",
          2879 => x"81065473",
          2880 => x"85eb387a",
          2881 => x"842a8106",
          2882 => x"54738698",
          2883 => x"387a852a",
          2884 => x"81065473",
          2885 => x"8697387e",
          2886 => x"81065473",
          2887 => x"858f387a",
          2888 => x"882a8106",
          2889 => x"5f7e802e",
          2890 => x"b2387778",
          2891 => x"84808029",
          2892 => x"fc808005",
          2893 => x"70902c5a",
          2894 => x"40548074",
          2895 => x"259d387c",
          2896 => x"52b05188",
          2897 => x"a93f7778",
          2898 => x"84808029",
          2899 => x"fc808005",
          2900 => x"70902c5a",
          2901 => x"40547380",
          2902 => x"24e53874",
          2903 => x"81065372",
          2904 => x"802eb238",
          2905 => x"78798180",
          2906 => x"0a2981ff",
          2907 => x"0a057098",
          2908 => x"2c5b5555",
          2909 => x"8075259d",
          2910 => x"387c52b0",
          2911 => x"5187ef3f",
          2912 => x"78798180",
          2913 => x"0a2981ff",
          2914 => x"0a057098",
          2915 => x"2c5b5555",
          2916 => x"748024e5",
          2917 => x"387a872a",
          2918 => x"7081065c",
          2919 => x"557a802e",
          2920 => x"81b93876",
          2921 => x"80e32e84",
          2922 => x"d8387680",
          2923 => x"f32e81ca",
          2924 => x"387680d3",
          2925 => x"2e81e238",
          2926 => x"7d84b9d8",
          2927 => x"2e96387c",
          2928 => x"52ff1e70",
          2929 => x"33525e87",
          2930 => x"a53f7d84",
          2931 => x"b9d82e09",
          2932 => x"8106ec38",
          2933 => x"7481065b",
          2934 => x"7a802efc",
          2935 => x"a7387778",
          2936 => x"84808029",
          2937 => x"fc808005",
          2938 => x"70902c5a",
          2939 => x"40558075",
          2940 => x"25fc9138",
          2941 => x"7c52a051",
          2942 => x"86f43fe2",
          2943 => x"397a9007",
          2944 => x"5b7aa007",
          2945 => x"7c33585b",
          2946 => x"76fa8738",
          2947 => x"fac8397a",
          2948 => x"80c0075b",
          2949 => x"80f85790",
          2950 => x"60618405",
          2951 => x"71087e83",
          2952 => x"ffcf065f",
          2953 => x"5942555a",
          2954 => x"fbfd397f",
          2955 => x"60840577",
          2956 => x"fe800a06",
          2957 => x"83133370",
          2958 => x"982b7207",
          2959 => x"7c848080",
          2960 => x"29fc8080",
          2961 => x"0570902c",
          2962 => x"5e525a56",
          2963 => x"57415f7a",
          2964 => x"872a7081",
          2965 => x"065c557a",
          2966 => x"fec93877",
          2967 => x"78848080",
          2968 => x"29fc8080",
          2969 => x"0570902c",
          2970 => x"5a545f80",
          2971 => x"7f25feb3",
          2972 => x"387c52a0",
          2973 => x"5185f73f",
          2974 => x"e239ff1a",
          2975 => x"7083ffff",
          2976 => x"065b5779",
          2977 => x"83ffff2e",
          2978 => x"feca387c",
          2979 => x"52757081",
          2980 => x"05573351",
          2981 => x"85d83fe2",
          2982 => x"39ff1a70",
          2983 => x"83ffff06",
          2984 => x"5b547983",
          2985 => x"ffff2efe",
          2986 => x"ab387c52",
          2987 => x"75708105",
          2988 => x"57335185",
          2989 => x"b93fe239",
          2990 => x"75fc0a06",
          2991 => x"81fc0a07",
          2992 => x"78848080",
          2993 => x"29fc8080",
          2994 => x"0570902c",
          2995 => x"5a585680",
          2996 => x"e37b872a",
          2997 => x"7081065d",
          2998 => x"56577afd",
          2999 => x"c638fefb",
          3000 => x"397f6084",
          3001 => x"05710870",
          3002 => x"53404156",
          3003 => x"807e2482",
          3004 => x"df387a83",
          3005 => x"ffbf065b",
          3006 => x"84b9d85e",
          3007 => x"faad397a",
          3008 => x"84077c33",
          3009 => x"585b76f8",
          3010 => x"8938f8ca",
          3011 => x"397a8807",
          3012 => x"5b807c33",
          3013 => x"585976f7",
          3014 => x"f938f8ba",
          3015 => x"397f6084",
          3016 => x"05710877",
          3017 => x"81065658",
          3018 => x"415f7282",
          3019 => x"8a387551",
          3020 => x"87f63f84",
          3021 => x"b9c80883",
          3022 => x"ffff0678",
          3023 => x"7131902b",
          3024 => x"545a7290",
          3025 => x"2c58fe87",
          3026 => x"397a80c0",
          3027 => x"077c3358",
          3028 => x"5b76f7be",
          3029 => x"38f7ff39",
          3030 => x"7f608405",
          3031 => x"71087781",
          3032 => x"065d5841",
          3033 => x"547981cf",
          3034 => x"38755187",
          3035 => x"bb3f84b9",
          3036 => x"c80883ff",
          3037 => x"ff067871",
          3038 => x"31902b54",
          3039 => x"5ac4397a",
          3040 => x"8180077c",
          3041 => x"33585b76",
          3042 => x"f78838f7",
          3043 => x"c9397778",
          3044 => x"84808029",
          3045 => x"fc808005",
          3046 => x"70902c5a",
          3047 => x"54548074",
          3048 => x"25fad638",
          3049 => x"7c52a051",
          3050 => x"83c43fe2",
          3051 => x"397c52b0",
          3052 => x"5183bb3f",
          3053 => x"79902e09",
          3054 => x"8106fae3",
          3055 => x"387c5276",
          3056 => x"5183ab3f",
          3057 => x"7a882a81",
          3058 => x"065f7e80",
          3059 => x"2efb8c38",
          3060 => x"fad83975",
          3061 => x"982c7871",
          3062 => x"31902b70",
          3063 => x"902c7d83",
          3064 => x"8006575a",
          3065 => x"515373fa",
          3066 => x"9038ffa2",
          3067 => x"397c52ad",
          3068 => x"5182fb3f",
          3069 => x"7e810654",
          3070 => x"73802efa",
          3071 => x"a238ffad",
          3072 => x"397c5275",
          3073 => x"982a5182",
          3074 => x"e53f7481",
          3075 => x"065b7a80",
          3076 => x"2ef7f138",
          3077 => x"fbc83978",
          3078 => x"7431982b",
          3079 => x"70982c5a",
          3080 => x"53f9b739",
          3081 => x"7c52ab51",
          3082 => x"82c43fc8",
          3083 => x"397c52a0",
          3084 => x"5182bb3f",
          3085 => x"ffbe3978",
          3086 => x"52755188",
          3087 => x"8b3f84b9",
          3088 => x"c80883ff",
          3089 => x"ff067871",
          3090 => x"31902b54",
          3091 => x"5afdf339",
          3092 => x"7a82077e",
          3093 => x"307183ff",
          3094 => x"bf065257",
          3095 => x"5bfd9939",
          3096 => x"fe3d0d84",
          3097 => x"d5a80853",
          3098 => x"75527451",
          3099 => x"f3b53f84",
          3100 => x"3d0d04fa",
          3101 => x"3d0d7855",
          3102 => x"800b84d5",
          3103 => x"ac088511",
          3104 => x"3370812a",
          3105 => x"81327081",
          3106 => x"06515658",
          3107 => x"5557ff56",
          3108 => x"72772e09",
          3109 => x"810680d5",
          3110 => x"38747081",
          3111 => x"05563353",
          3112 => x"72772eb0",
          3113 => x"3884d5ac",
          3114 => x"08527251",
          3115 => x"90140853",
          3116 => x"722d84b9",
          3117 => x"c808802e",
          3118 => x"8338ff57",
          3119 => x"74708105",
          3120 => x"56335372",
          3121 => x"802e8838",
          3122 => x"84d5ac08",
          3123 => x"54d73984",
          3124 => x"d5ac0854",
          3125 => x"84d5ac08",
          3126 => x"528a5190",
          3127 => x"14085574",
          3128 => x"2d84b9c8",
          3129 => x"08802e83",
          3130 => x"38ff5776",
          3131 => x"567584b9",
          3132 => x"c80c883d",
          3133 => x"0d04fa3d",
          3134 => x"0d787a56",
          3135 => x"54800b85",
          3136 => x"16337081",
          3137 => x"2a813270",
          3138 => x"81065155",
          3139 => x"5757ff56",
          3140 => x"72772e09",
          3141 => x"81069238",
          3142 => x"73708105",
          3143 => x"55335372",
          3144 => x"772e0981",
          3145 => x"06983876",
          3146 => x"567584b9",
          3147 => x"c80c883d",
          3148 => x"0d047370",
          3149 => x"81055533",
          3150 => x"5372802e",
          3151 => x"ea387452",
          3152 => x"72519015",
          3153 => x"0853722d",
          3154 => x"84b9c808",
          3155 => x"802ee338",
          3156 => x"ff747081",
          3157 => x"05563354",
          3158 => x"5772e338",
          3159 => x"ca39ff3d",
          3160 => x"0d84d5ac",
          3161 => x"08527351",
          3162 => x"853f833d",
          3163 => x"0d04fa3d",
          3164 => x"0d787a85",
          3165 => x"11337081",
          3166 => x"2a813281",
          3167 => x"06565656",
          3168 => x"57ff5672",
          3169 => x"ae387382",
          3170 => x"2a810654",
          3171 => x"73802eac",
          3172 => x"388c1508",
          3173 => x"53728816",
          3174 => x"08259138",
          3175 => x"74085676",
          3176 => x"76347408",
          3177 => x"8105750c",
          3178 => x"8c150853",
          3179 => x"81138c16",
          3180 => x"0c765675",
          3181 => x"84b9c80c",
          3182 => x"883d0d04",
          3183 => x"74527681",
          3184 => x"ff065190",
          3185 => x"15085473",
          3186 => x"2dff5684",
          3187 => x"b9c808e3",
          3188 => x"388c1508",
          3189 => x"81058c16",
          3190 => x"0c7656d7",
          3191 => x"39fb3d0d",
          3192 => x"77851133",
          3193 => x"7081ff06",
          3194 => x"70813281",
          3195 => x"06555556",
          3196 => x"56ff5471",
          3197 => x"b3387286",
          3198 => x"2a810652",
          3199 => x"71b33872",
          3200 => x"822a8106",
          3201 => x"5271802e",
          3202 => x"80c33875",
          3203 => x"08703353",
          3204 => x"5371802e",
          3205 => x"80f03881",
          3206 => x"13760c8c",
          3207 => x"16088105",
          3208 => x"8c170c71",
          3209 => x"81ff0654",
          3210 => x"7384b9c8",
          3211 => x"0c873d0d",
          3212 => x"0474ffbf",
          3213 => x"06537285",
          3214 => x"17348c16",
          3215 => x"0881058c",
          3216 => x"170c8416",
          3217 => x"3384b9c8",
          3218 => x"0c873d0d",
          3219 => x"04755194",
          3220 => x"16085574",
          3221 => x"2d84b9c8",
          3222 => x"085284b9",
          3223 => x"c8088025",
          3224 => x"ffb93885",
          3225 => x"16337090",
          3226 => x"07545284",
          3227 => x"b9c808ff",
          3228 => x"2e853871",
          3229 => x"a0075372",
          3230 => x"851734ff",
          3231 => x"547384b9",
          3232 => x"c80c873d",
          3233 => x"0d0474a0",
          3234 => x"07537285",
          3235 => x"1734ff54",
          3236 => x"ec39fd3d",
          3237 => x"0d757771",
          3238 => x"54545471",
          3239 => x"70810553",
          3240 => x"335170f7",
          3241 => x"38ff1252",
          3242 => x"72708105",
          3243 => x"54335170",
          3244 => x"72708105",
          3245 => x"543470f0",
          3246 => x"387384b9",
          3247 => x"c80c853d",
          3248 => x"0d04fc3d",
          3249 => x"0d767971",
          3250 => x"7a555552",
          3251 => x"5470802e",
          3252 => x"9d387372",
          3253 => x"27a13870",
          3254 => x"802e9338",
          3255 => x"71708105",
          3256 => x"53337370",
          3257 => x"81055534",
          3258 => x"ff115170",
          3259 => x"ef387384",
          3260 => x"b9c80c86",
          3261 => x"3d0d0470",
          3262 => x"12557375",
          3263 => x"27d93870",
          3264 => x"14755353",
          3265 => x"ff13ff13",
          3266 => x"53537133",
          3267 => x"7334ff11",
          3268 => x"5170802e",
          3269 => x"d938ff13",
          3270 => x"ff135353",
          3271 => x"71337334",
          3272 => x"ff115170",
          3273 => x"df38c739",
          3274 => x"fe3d0d74",
          3275 => x"70535371",
          3276 => x"70810553",
          3277 => x"335170f7",
          3278 => x"38ff1270",
          3279 => x"743184b9",
          3280 => x"c80c5184",
          3281 => x"3d0d04fd",
          3282 => x"3d0d7577",
          3283 => x"71545454",
          3284 => x"72708105",
          3285 => x"54335170",
          3286 => x"72708105",
          3287 => x"543470f0",
          3288 => x"387384b9",
          3289 => x"c80c853d",
          3290 => x"0d04fd3d",
          3291 => x"0d757871",
          3292 => x"79555552",
          3293 => x"5470802e",
          3294 => x"93387170",
          3295 => x"81055333",
          3296 => x"73708105",
          3297 => x"5534ff11",
          3298 => x"5170ef38",
          3299 => x"7384b9c8",
          3300 => x"0c853d0d",
          3301 => x"04fc3d0d",
          3302 => x"76787a55",
          3303 => x"56547280",
          3304 => x"2ea13873",
          3305 => x"33757081",
          3306 => x"05573352",
          3307 => x"5271712e",
          3308 => x"0981069a",
          3309 => x"38811454",
          3310 => x"71802eb7",
          3311 => x"38ff1353",
          3312 => x"72e13880",
          3313 => x"517084b9",
          3314 => x"c80c863d",
          3315 => x"0d047280",
          3316 => x"2ef13873",
          3317 => x"3353ff51",
          3318 => x"72802ee9",
          3319 => x"38ff1533",
          3320 => x"52815171",
          3321 => x"802ede38",
          3322 => x"72723184",
          3323 => x"b9c80c86",
          3324 => x"3d0d0471",
          3325 => x"84b9c80c",
          3326 => x"863d0d04",
          3327 => x"fb3d0d77",
          3328 => x"79537052",
          3329 => x"5680c13f",
          3330 => x"84b9c808",
          3331 => x"84b9c808",
          3332 => x"81055255",
          3333 => x"81b2ea3f",
          3334 => x"84b9c808",
          3335 => x"5484b9c8",
          3336 => x"08802e9b",
          3337 => x"3884b9c8",
          3338 => x"08155480",
          3339 => x"74347453",
          3340 => x"755284b9",
          3341 => x"c80851fe",
          3342 => x"b13f84b9",
          3343 => x"c8085473",
          3344 => x"84b9c80c",
          3345 => x"873d0d04",
          3346 => x"fd3d0d75",
          3347 => x"77717154",
          3348 => x"55535471",
          3349 => x"802e9f38",
          3350 => x"72708105",
          3351 => x"54335170",
          3352 => x"802e8c38",
          3353 => x"ff125271",
          3354 => x"ff2e0981",
          3355 => x"06ea38ff",
          3356 => x"13707531",
          3357 => x"52527084",
          3358 => x"b9c80c85",
          3359 => x"3d0d04fd",
          3360 => x"3d0d7577",
          3361 => x"79725553",
          3362 => x"54547080",
          3363 => x"2e8e3872",
          3364 => x"72708105",
          3365 => x"5434ff11",
          3366 => x"5170f438",
          3367 => x"7384b9c8",
          3368 => x"0c853d0d",
          3369 => x"04fa3d0d",
          3370 => x"787a5854",
          3371 => x"a0527680",
          3372 => x"2e8b3876",
          3373 => x"5180f53f",
          3374 => x"84b9c808",
          3375 => x"52e01253",
          3376 => x"73802e8d",
          3377 => x"38735180",
          3378 => x"e33f7184",
          3379 => x"b9c80831",
          3380 => x"53805272",
          3381 => x"9f2680cb",
          3382 => x"38735272",
          3383 => x"9f2e80c3",
          3384 => x"38811374",
          3385 => x"712aa072",
          3386 => x"3176712b",
          3387 => x"57545455",
          3388 => x"80567476",
          3389 => x"2ea83872",
          3390 => x"10749f2a",
          3391 => x"07741077",
          3392 => x"07787231",
          3393 => x"ff119f2c",
          3394 => x"7081067b",
          3395 => x"72067571",
          3396 => x"31ff1c5c",
          3397 => x"56525255",
          3398 => x"58555374",
          3399 => x"da387310",
          3400 => x"76075271",
          3401 => x"84b9c80c",
          3402 => x"883d0d04",
          3403 => x"fc3d0d76",
          3404 => x"70fc8080",
          3405 => x"06703070",
          3406 => x"72078025",
          3407 => x"70842b90",
          3408 => x"71317571",
          3409 => x"2a7083fe",
          3410 => x"80067030",
          3411 => x"70802583",
          3412 => x"2b887131",
          3413 => x"74712a70",
          3414 => x"81f00670",
          3415 => x"30708025",
          3416 => x"822b8471",
          3417 => x"3174712a",
          3418 => x"5553751b",
          3419 => x"05738c06",
          3420 => x"70307080",
          3421 => x"25108271",
          3422 => x"3177712a",
          3423 => x"70812a81",
          3424 => x"32708106",
          3425 => x"70308274",
          3426 => x"31067519",
          3427 => x"0584b9c8",
          3428 => x"0c515254",
          3429 => x"55515456",
          3430 => x"5a535555",
          3431 => x"55515656",
          3432 => x"56565158",
          3433 => x"56545286",
          3434 => x"3d0d04fd",
          3435 => x"3d0d7577",
          3436 => x"70547153",
          3437 => x"54548194",
          3438 => x"3f84b9c8",
          3439 => x"08732974",
          3440 => x"713184b9",
          3441 => x"c80c5385",
          3442 => x"3d0d04fa",
          3443 => x"3d0d787a",
          3444 => x"5854a053",
          3445 => x"76802e8b",
          3446 => x"387651fe",
          3447 => x"cf3f84b9",
          3448 => x"c80853e0",
          3449 => x"13527380",
          3450 => x"2e8d3873",
          3451 => x"51febd3f",
          3452 => x"7284b9c8",
          3453 => x"08315273",
          3454 => x"53719f26",
          3455 => x"80c53880",
          3456 => x"53719f2e",
          3457 => x"be388112",
          3458 => x"74712aa0",
          3459 => x"72317671",
          3460 => x"2b575454",
          3461 => x"55805674",
          3462 => x"762ea838",
          3463 => x"7210749f",
          3464 => x"2a077410",
          3465 => x"77077872",
          3466 => x"31ff119f",
          3467 => x"2c708106",
          3468 => x"7b720675",
          3469 => x"7131ff1c",
          3470 => x"5c565252",
          3471 => x"55585553",
          3472 => x"74da3872",
          3473 => x"84b9c80c",
          3474 => x"883d0d04",
          3475 => x"fa3d0d78",
          3476 => x"9f2c7a9f",
          3477 => x"2c7a9f2c",
          3478 => x"7b327c9f",
          3479 => x"2c7d3273",
          3480 => x"73327174",
          3481 => x"31577275",
          3482 => x"31565956",
          3483 => x"595556fc",
          3484 => x"b43f84b9",
          3485 => x"c8087532",
          3486 => x"753184b9",
          3487 => x"c80c883d",
          3488 => x"0d04f73d",
          3489 => x"0d7b7d5b",
          3490 => x"5780707b",
          3491 => x"0c770870",
          3492 => x"33565659",
          3493 => x"73a02e09",
          3494 => x"81068f38",
          3495 => x"81157078",
          3496 => x"0c703355",
          3497 => x"5573a02e",
          3498 => x"f33873ad",
          3499 => x"2e80f538",
          3500 => x"73b02e81",
          3501 => x"8338d014",
          3502 => x"58805677",
          3503 => x"892680db",
          3504 => x"388a5880",
          3505 => x"56a07427",
          3506 => x"80c43880",
          3507 => x"e0742789",
          3508 => x"38e01470",
          3509 => x"81ff0655",
          3510 => x"53d01470",
          3511 => x"81ff0651",
          3512 => x"53907327",
          3513 => x"8f38f913",
          3514 => x"7081ff06",
          3515 => x"54548973",
          3516 => x"27818938",
          3517 => x"72782781",
          3518 => x"83387776",
          3519 => x"29138116",
          3520 => x"70790c70",
          3521 => x"33565656",
          3522 => x"73a026ff",
          3523 => x"be387880",
          3524 => x"2e843875",
          3525 => x"3056757a",
          3526 => x"0c815675",
          3527 => x"84b9c80c",
          3528 => x"8b3d0d04",
          3529 => x"81701670",
          3530 => x"790c7033",
          3531 => x"56565973",
          3532 => x"b02e0981",
          3533 => x"06feff38",
          3534 => x"81157078",
          3535 => x"0c703355",
          3536 => x"557380e2",
          3537 => x"2ea63890",
          3538 => x"587380f8",
          3539 => x"2ea03881",
          3540 => x"56a07427",
          3541 => x"c638d014",
          3542 => x"53805688",
          3543 => x"58897327",
          3544 => x"fee13875",
          3545 => x"84b9c80c",
          3546 => x"8b3d0d04",
          3547 => x"82588115",
          3548 => x"70780c70",
          3549 => x"33555580",
          3550 => x"56feca39",
          3551 => x"800b84b9",
          3552 => x"c80c8b3d",
          3553 => x"0d04f73d",
          3554 => x"0d7b7d5b",
          3555 => x"5780707b",
          3556 => x"0c770870",
          3557 => x"33565659",
          3558 => x"73a02e09",
          3559 => x"81068f38",
          3560 => x"81157078",
          3561 => x"0c703355",
          3562 => x"5573a02e",
          3563 => x"f33873ad",
          3564 => x"2e80f538",
          3565 => x"73b02e81",
          3566 => x"8338d014",
          3567 => x"58805677",
          3568 => x"892680db",
          3569 => x"388a5880",
          3570 => x"56a07427",
          3571 => x"80c43880",
          3572 => x"e0742789",
          3573 => x"38e01470",
          3574 => x"81ff0655",
          3575 => x"53d01470",
          3576 => x"81ff0651",
          3577 => x"53907327",
          3578 => x"8f38f913",
          3579 => x"7081ff06",
          3580 => x"54548973",
          3581 => x"27818938",
          3582 => x"72782781",
          3583 => x"83387776",
          3584 => x"29138116",
          3585 => x"70790c70",
          3586 => x"33565656",
          3587 => x"73a026ff",
          3588 => x"be387880",
          3589 => x"2e843875",
          3590 => x"3056757a",
          3591 => x"0c815675",
          3592 => x"84b9c80c",
          3593 => x"8b3d0d04",
          3594 => x"81701670",
          3595 => x"790c7033",
          3596 => x"56565973",
          3597 => x"b02e0981",
          3598 => x"06feff38",
          3599 => x"81157078",
          3600 => x"0c703355",
          3601 => x"557380e2",
          3602 => x"2ea63890",
          3603 => x"587380f8",
          3604 => x"2ea03881",
          3605 => x"56a07427",
          3606 => x"c638d014",
          3607 => x"53805688",
          3608 => x"58897327",
          3609 => x"fee13875",
          3610 => x"84b9c80c",
          3611 => x"8b3d0d04",
          3612 => x"82588115",
          3613 => x"70780c70",
          3614 => x"33555580",
          3615 => x"56feca39",
          3616 => x"800b84b9",
          3617 => x"c80c8b3d",
          3618 => x"0d0480d6",
          3619 => x"e23f84b9",
          3620 => x"c80881ff",
          3621 => x"0684b9c8",
          3622 => x"0c04ff3d",
          3623 => x"0d735271",
          3624 => x"93268c38",
          3625 => x"71101083",
          3626 => x"be840552",
          3627 => x"71080483",
          3628 => x"ce9c51ef",
          3629 => x"be3f833d",
          3630 => x"0d0483ce",
          3631 => x"ac51efb3",
          3632 => x"3f833d0d",
          3633 => x"0483cec4",
          3634 => x"51efa83f",
          3635 => x"833d0d04",
          3636 => x"83cedc51",
          3637 => x"ef9d3f83",
          3638 => x"3d0d0483",
          3639 => x"cef451ef",
          3640 => x"923f833d",
          3641 => x"0d0483cf",
          3642 => x"8451ef87",
          3643 => x"3f833d0d",
          3644 => x"0483cfa4",
          3645 => x"51eefc3f",
          3646 => x"833d0d04",
          3647 => x"83cfb451",
          3648 => x"eef13f83",
          3649 => x"3d0d0483",
          3650 => x"cfdc51ee",
          3651 => x"e63f833d",
          3652 => x"0d0483cf",
          3653 => x"f051eedb",
          3654 => x"3f833d0d",
          3655 => x"0483d08c",
          3656 => x"51eed03f",
          3657 => x"833d0d04",
          3658 => x"83d0a451",
          3659 => x"eec53f83",
          3660 => x"3d0d0483",
          3661 => x"d0bc51ee",
          3662 => x"ba3f833d",
          3663 => x"0d0483d0",
          3664 => x"d451eeaf",
          3665 => x"3f833d0d",
          3666 => x"0483d0e4",
          3667 => x"51eea43f",
          3668 => x"833d0d04",
          3669 => x"83d0f851",
          3670 => x"ee993f83",
          3671 => x"3d0d0483",
          3672 => x"d18851ee",
          3673 => x"8e3f833d",
          3674 => x"0d0483d1",
          3675 => x"9851ee83",
          3676 => x"3f833d0d",
          3677 => x"0483d1a8",
          3678 => x"51edf83f",
          3679 => x"833d0d04",
          3680 => x"83d1b851",
          3681 => x"eded3f83",
          3682 => x"3d0d0483",
          3683 => x"d1c451ed",
          3684 => x"e23f833d",
          3685 => x"0d04ec3d",
          3686 => x"0d660284",
          3687 => x"0580e305",
          3688 => x"335b5880",
          3689 => x"68793070",
          3690 => x"7b077325",
          3691 => x"51575759",
          3692 => x"78577587",
          3693 => x"ff268338",
          3694 => x"81577477",
          3695 => x"077081ff",
          3696 => x"06515593",
          3697 => x"577480e2",
          3698 => x"38815377",
          3699 => x"528c3d70",
          3700 => x"52588295",
          3701 => x"d93f84b9",
          3702 => x"c8085784",
          3703 => x"b9c80880",
          3704 => x"2e80d038",
          3705 => x"775182af",
          3706 => x"973f7630",
          3707 => x"70780780",
          3708 => x"257b3070",
          3709 => x"9f2a7206",
          3710 => x"53575758",
          3711 => x"77802eaa",
          3712 => x"3887c098",
          3713 => x"88085574",
          3714 => x"87e72680",
          3715 => x"e0387452",
          3716 => x"7887e829",
          3717 => x"51f58e3f",
          3718 => x"84b9c808",
          3719 => x"5483d1f4",
          3720 => x"53785283",
          3721 => x"d1d051df",
          3722 => x"df3f7684",
          3723 => x"b9c80c96",
          3724 => x"3d0d0484",
          3725 => x"b9c80887",
          3726 => x"c098880c",
          3727 => x"84b9c808",
          3728 => x"59963dd4",
          3729 => x"05548480",
          3730 => x"53755277",
          3731 => x"51829dce",
          3732 => x"3f84b9c8",
          3733 => x"085784b9",
          3734 => x"c808ff88",
          3735 => x"387a5574",
          3736 => x"802eff80",
          3737 => x"38741975",
          3738 => x"175759d5",
          3739 => x"3987e852",
          3740 => x"7451f4b1",
          3741 => x"3f84b9c8",
          3742 => x"08527851",
          3743 => x"f4a73f84",
          3744 => x"b9c80854",
          3745 => x"83d1f453",
          3746 => x"785283d1",
          3747 => x"d051def8",
          3748 => x"3fff9739",
          3749 => x"f83d0d7c",
          3750 => x"028405b7",
          3751 => x"05335859",
          3752 => x"ff588053",
          3753 => x"7b527a51",
          3754 => x"fdec3f84",
          3755 => x"b9c8088b",
          3756 => x"3876802e",
          3757 => x"91387681",
          3758 => x"2e8a3877",
          3759 => x"84b9c80c",
          3760 => x"8a3d0d04",
          3761 => x"780484d5",
          3762 => x"a8566155",
          3763 => x"605484b9",
          3764 => x"c8537f52",
          3765 => x"7e51782d",
          3766 => x"84b9c808",
          3767 => x"84b9c80c",
          3768 => x"8a3d0d04",
          3769 => x"f33d0d7f",
          3770 => x"6163028c",
          3771 => x"0580cf05",
          3772 => x"33737315",
          3773 => x"68415f5c",
          3774 => x"5c5f5d5e",
          3775 => x"78802e83",
          3776 => x"82387a52",
          3777 => x"83d1fc51",
          3778 => x"ddfe3f83",
          3779 => x"d28451dd",
          3780 => x"f73f8054",
          3781 => x"737927b2",
          3782 => x"387c902e",
          3783 => x"81ed387c",
          3784 => x"a02e82a8",
          3785 => x"38731853",
          3786 => x"727a2781",
          3787 => x"a7387233",
          3788 => x"5283d288",
          3789 => x"51ddd13f",
          3790 => x"811484d5",
          3791 => x"ac085354",
          3792 => x"a051ecaa",
          3793 => x"3f787426",
          3794 => x"dc3883d2",
          3795 => x"9051ddb8",
          3796 => x"3f805675",
          3797 => x"792780c0",
          3798 => x"38751870",
          3799 => x"33555380",
          3800 => x"55727a27",
          3801 => x"83388155",
          3802 => x"80539f74",
          3803 => x"27833881",
          3804 => x"53747306",
          3805 => x"7081ff06",
          3806 => x"56577480",
          3807 => x"2e883880",
          3808 => x"fe742781",
          3809 => x"ee3884d5",
          3810 => x"ac0852a0",
          3811 => x"51ebdf3f",
          3812 => x"81165678",
          3813 => x"7626c238",
          3814 => x"83d29451",
          3815 => x"e9d53f78",
          3816 => x"18791c5c",
          3817 => x"5880519d",
          3818 => x"c33f84b9",
          3819 => x"c808982b",
          3820 => x"70982c58",
          3821 => x"5476a02e",
          3822 => x"81ee3876",
          3823 => x"9b2e82c3",
          3824 => x"387b1e57",
          3825 => x"767826fe",
          3826 => x"b938ff0b",
          3827 => x"84b9c80c",
          3828 => x"8f3d0d04",
          3829 => x"83d29851",
          3830 => x"dcae3f81",
          3831 => x"1484d5ac",
          3832 => x"085354a0",
          3833 => x"51eb873f",
          3834 => x"787426fe",
          3835 => x"b838feda",
          3836 => x"3983d2a8",
          3837 => x"51dc913f",
          3838 => x"821484d5",
          3839 => x"ac085354",
          3840 => x"a051eaea",
          3841 => x"3f737927",
          3842 => x"fec03873",
          3843 => x"1853727a",
          3844 => x"27df3872",
          3845 => x"225283d2",
          3846 => x"9c51dbec",
          3847 => x"3f821484",
          3848 => x"d5ac0853",
          3849 => x"54a051ea",
          3850 => x"c53f7874",
          3851 => x"26dd38fe",
          3852 => x"993983d2",
          3853 => x"a451dbd0",
          3854 => x"3f841484",
          3855 => x"d5ac0853",
          3856 => x"54a051ea",
          3857 => x"a93f7379",
          3858 => x"27fdff38",
          3859 => x"73185372",
          3860 => x"7a27df38",
          3861 => x"72085283",
          3862 => x"d1fc51db",
          3863 => x"ab3f8414",
          3864 => x"84d5ac08",
          3865 => x"5354a051",
          3866 => x"ea843f78",
          3867 => x"7426dd38",
          3868 => x"fdd83984",
          3869 => x"d5ac0852",
          3870 => x"7351e9f2",
          3871 => x"3f811656",
          3872 => x"fe913980",
          3873 => x"cee93f84",
          3874 => x"b9c80881",
          3875 => x"ff065388",
          3876 => x"5972a82e",
          3877 => x"fcec38a0",
          3878 => x"597280d0",
          3879 => x"2e098106",
          3880 => x"fce03890",
          3881 => x"59fcdb39",
          3882 => x"80519bc0",
          3883 => x"3f84b9c8",
          3884 => x"08982b70",
          3885 => x"982c70a0",
          3886 => x"32703072",
          3887 => x"9b327030",
          3888 => x"70720773",
          3889 => x"75070651",
          3890 => x"55585957",
          3891 => x"58537280",
          3892 => x"25fde838",
          3893 => x"80519b94",
          3894 => x"3f84b9c8",
          3895 => x"08982b70",
          3896 => x"982c70a0",
          3897 => x"32703072",
          3898 => x"9b327030",
          3899 => x"70720773",
          3900 => x"75070651",
          3901 => x"55585957",
          3902 => x"58538073",
          3903 => x"24ffa938",
          3904 => x"fdb93980",
          3905 => x"0b84b9c8",
          3906 => x"0c8f3d0d",
          3907 => x"04fe3d0d",
          3908 => x"87c09680",
          3909 => x"0853aad7",
          3910 => x"3f81519d",
          3911 => x"883f83d3",
          3912 => x"c0519d99",
          3913 => x"3f80519c",
          3914 => x"fc3f7281",
          3915 => x"2a708106",
          3916 => x"51527182",
          3917 => x"b7387282",
          3918 => x"2a708106",
          3919 => x"51527182",
          3920 => x"89387283",
          3921 => x"2a708106",
          3922 => x"51527181",
          3923 => x"db387284",
          3924 => x"2a708106",
          3925 => x"51527181",
          3926 => x"ad387285",
          3927 => x"2a708106",
          3928 => x"51527180",
          3929 => x"ff387286",
          3930 => x"2a708106",
          3931 => x"51527180",
          3932 => x"d2387287",
          3933 => x"2a708106",
          3934 => x"515271a9",
          3935 => x"3872882a",
          3936 => x"81065372",
          3937 => x"8838a9ef",
          3938 => x"3f843d0d",
          3939 => x"0481519c",
          3940 => x"943f83d3",
          3941 => x"d8519ca5",
          3942 => x"3f80519c",
          3943 => x"883fa9d7",
          3944 => x"3f843d0d",
          3945 => x"0481519b",
          3946 => x"fc3f83d3",
          3947 => x"ec519c8d",
          3948 => x"3f80519b",
          3949 => x"f03f7288",
          3950 => x"2a810653",
          3951 => x"72802ec6",
          3952 => x"38cb3981",
          3953 => x"519bde3f",
          3954 => x"83d48051",
          3955 => x"9bef3f80",
          3956 => x"519bd23f",
          3957 => x"72872a70",
          3958 => x"81065152",
          3959 => x"71802eff",
          3960 => x"9c38c239",
          3961 => x"81519bbd",
          3962 => x"3f83d494",
          3963 => x"519bce3f",
          3964 => x"80519bb1",
          3965 => x"3f72862a",
          3966 => x"70810651",
          3967 => x"5271802e",
          3968 => x"fef038ff",
          3969 => x"be398151",
          3970 => x"9b9b3f83",
          3971 => x"d4a8519b",
          3972 => x"ac3f8051",
          3973 => x"9b8f3f72",
          3974 => x"852a7081",
          3975 => x"06515271",
          3976 => x"802efec2",
          3977 => x"38ffbd39",
          3978 => x"81519af9",
          3979 => x"3f83d4bc",
          3980 => x"519b8a3f",
          3981 => x"80519aed",
          3982 => x"3f72842a",
          3983 => x"70810651",
          3984 => x"5271802e",
          3985 => x"fe9438ff",
          3986 => x"bd398151",
          3987 => x"9ad73f83",
          3988 => x"d4d0519a",
          3989 => x"e83f8051",
          3990 => x"9acb3f72",
          3991 => x"832a7081",
          3992 => x"06515271",
          3993 => x"802efde6",
          3994 => x"38ffbd39",
          3995 => x"81519ab5",
          3996 => x"3f83d4e0",
          3997 => x"519ac63f",
          3998 => x"80519aa9",
          3999 => x"3f72822a",
          4000 => x"70810651",
          4001 => x"5271802e",
          4002 => x"fdb838ff",
          4003 => x"bd39ca3d",
          4004 => x"0d807041",
          4005 => x"41ff6184",
          4006 => x"d0d40c42",
          4007 => x"81526051",
          4008 => x"81b68c3f",
          4009 => x"84b9c808",
          4010 => x"81ff069b",
          4011 => x"3d405978",
          4012 => x"612e84b1",
          4013 => x"3883d5b4",
          4014 => x"51e3b83f",
          4015 => x"983d4383",
          4016 => x"d5ec51d6",
          4017 => x"c33f7e48",
          4018 => x"80f85380",
          4019 => x"527e51eb",
          4020 => x"ae3f0b0b",
          4021 => x"83eebc33",
          4022 => x"7081ff06",
          4023 => x"5b597980",
          4024 => x"2e82f138",
          4025 => x"79812e83",
          4026 => x"88387881",
          4027 => x"ff065e7d",
          4028 => x"822e83c1",
          4029 => x"3867705a",
          4030 => x"5a79802e",
          4031 => x"83dc3879",
          4032 => x"335c7ba0",
          4033 => x"2e098106",
          4034 => x"8c38811a",
          4035 => x"70335d5a",
          4036 => x"7ba02ef6",
          4037 => x"38805c7b",
          4038 => x"9b26be38",
          4039 => x"7b902983",
          4040 => x"eec00570",
          4041 => x"08525be7",
          4042 => x"ff3f84b9",
          4043 => x"c80884b9",
          4044 => x"c808547a",
          4045 => x"537b0852",
          4046 => x"5de8da3f",
          4047 => x"84b9c808",
          4048 => x"8b38841b",
          4049 => x"335e7d81",
          4050 => x"2e838038",
          4051 => x"811c7081",
          4052 => x"ff065d5b",
          4053 => x"9b7c27c4",
          4054 => x"389a3d33",
          4055 => x"5c7b802e",
          4056 => x"fedd3880",
          4057 => x"f8527e51",
          4058 => x"e9923f84",
          4059 => x"b9c8085e",
          4060 => x"84b9c808",
          4061 => x"802e8dc9",
          4062 => x"3884b9c8",
          4063 => x"0848b83d",
          4064 => x"ff800551",
          4065 => x"91a43f84",
          4066 => x"b9c80860",
          4067 => x"62065c5c",
          4068 => x"7a802e81",
          4069 => x"843884b9",
          4070 => x"c80851e7",
          4071 => x"8b3f84b9",
          4072 => x"c8088f26",
          4073 => x"80f33881",
          4074 => x"0ba53d5e",
          4075 => x"5b7a822e",
          4076 => x"8d85387a",
          4077 => x"82248ce2",
          4078 => x"387a812e",
          4079 => x"82e4387b",
          4080 => x"54805383",
          4081 => x"d5f0527c",
          4082 => x"51d5dd3f",
          4083 => x"83f28458",
          4084 => x"84b9f857",
          4085 => x"7d566755",
          4086 => x"80549080",
          4087 => x"0a539080",
          4088 => x"0a527c51",
          4089 => x"f5ae3f84",
          4090 => x"b9c80884",
          4091 => x"b9c80809",
          4092 => x"70307072",
          4093 => x"07802551",
          4094 => x"5b5b4280",
          4095 => x"5a7a8326",
          4096 => x"8338815a",
          4097 => x"787a0659",
          4098 => x"78802e8d",
          4099 => x"38811b70",
          4100 => x"81ff065c",
          4101 => x"5a7aff95",
          4102 => x"387f8132",
          4103 => x"61813207",
          4104 => x"5d7c81ee",
          4105 => x"3861ff2e",
          4106 => x"81e8387d",
          4107 => x"518194e1",
          4108 => x"3f83d5ec",
          4109 => x"51d3d13f",
          4110 => x"7e4880f8",
          4111 => x"5380527e",
          4112 => x"51e8bc3f",
          4113 => x"0b0b83ee",
          4114 => x"bc337081",
          4115 => x"ff065b59",
          4116 => x"79fd9138",
          4117 => x"815383d5",
          4118 => x"985284d0",
          4119 => x"d8518288",
          4120 => x"cd3f84b9",
          4121 => x"c80880c5",
          4122 => x"38810b0b",
          4123 => x"0b83eebc",
          4124 => x"3484d0d8",
          4125 => x"5380f852",
          4126 => x"7e5182f6",
          4127 => x"c83f84b9",
          4128 => x"c808802e",
          4129 => x"a03884b9",
          4130 => x"c80851df",
          4131 => x"e63f0b0b",
          4132 => x"83eebc33",
          4133 => x"7081ff06",
          4134 => x"5f597d82",
          4135 => x"2e098106",
          4136 => x"fcd33891",
          4137 => x"3984d0d8",
          4138 => x"5182a1d4",
          4139 => x"3f820b0b",
          4140 => x"0b83eebc",
          4141 => x"3483d5a8",
          4142 => x"5380f852",
          4143 => x"7e51a7d4",
          4144 => x"3f67705a",
          4145 => x"5a79fcb7",
          4146 => x"3890397c",
          4147 => x"1a630c85",
          4148 => x"1b335978",
          4149 => x"818926fd",
          4150 => x"80387810",
          4151 => x"1083bed4",
          4152 => x"055a7908",
          4153 => x"04835383",
          4154 => x"d5f8527e",
          4155 => x"51e4fb3f",
          4156 => x"60537e52",
          4157 => x"84baf451",
          4158 => x"8285843f",
          4159 => x"84b9c808",
          4160 => x"612e0981",
          4161 => x"06fbae38",
          4162 => x"81709a3d",
          4163 => x"454141fb",
          4164 => x"ae3983d5",
          4165 => x"fc51dedb",
          4166 => x"3f7d5181",
          4167 => x"92f33ffe",
          4168 => x"903983d6",
          4169 => x"8c567b55",
          4170 => x"83d69054",
          4171 => x"805383d6",
          4172 => x"94527c51",
          4173 => x"d2f23ffd",
          4174 => x"9339818c",
          4175 => x"ab3ffaff",
          4176 => x"399af83f",
          4177 => x"faf93981",
          4178 => x"528351bf",
          4179 => x"a43ffaef",
          4180 => x"39818dd6",
          4181 => x"3ffae839",
          4182 => x"83d6a451",
          4183 => x"de953f80",
          4184 => x"59780483",
          4185 => x"d6b851de",
          4186 => x"8a3fd0fd",
          4187 => x"3ffad039",
          4188 => x"b83dff84",
          4189 => x"1153ff80",
          4190 => x"0551ec8a",
          4191 => x"3f84b9c8",
          4192 => x"08802efa",
          4193 => x"ba386852",
          4194 => x"83d6d451",
          4195 => x"d0fa3f68",
          4196 => x"5a792d84",
          4197 => x"b9c80880",
          4198 => x"2efaa438",
          4199 => x"84b9c808",
          4200 => x"5283d6f0",
          4201 => x"51d0e13f",
          4202 => x"fa9539b8",
          4203 => x"3dff8411",
          4204 => x"53ff8005",
          4205 => x"51ebcf3f",
          4206 => x"84b9c808",
          4207 => x"802ef9ff",
          4208 => x"38685283",
          4209 => x"d78c51d0",
          4210 => x"bf3f6859",
          4211 => x"7804b83d",
          4212 => x"fef41153",
          4213 => x"ff800551",
          4214 => x"e9a83f84",
          4215 => x"b9c80880",
          4216 => x"2ef9dc38",
          4217 => x"b83dfef0",
          4218 => x"1153ff80",
          4219 => x"0551e992",
          4220 => x"3f84b9c8",
          4221 => x"0886d038",
          4222 => x"64597808",
          4223 => x"53785283",
          4224 => x"d7a851d0",
          4225 => x"833f84d5",
          4226 => x"a8085380",
          4227 => x"f8527e51",
          4228 => x"d0913f7e",
          4229 => x"487e3359",
          4230 => x"78ae2ef9",
          4231 => x"a238789f",
          4232 => x"2687d338",
          4233 => x"64840570",
          4234 => x"4659cf39",
          4235 => x"b83dfef4",
          4236 => x"1153ff80",
          4237 => x"0551e8ca",
          4238 => x"3f84b9c8",
          4239 => x"08802ef8",
          4240 => x"fe38b83d",
          4241 => x"fef01153",
          4242 => x"ff800551",
          4243 => x"e8b43f84",
          4244 => x"b9c80886",
          4245 => x"b0386459",
          4246 => x"78225378",
          4247 => x"5283d7b8",
          4248 => x"51cfa53f",
          4249 => x"84d5a808",
          4250 => x"5380f852",
          4251 => x"7e51cfb3",
          4252 => x"3f7e487e",
          4253 => x"335978ae",
          4254 => x"2ef8c438",
          4255 => x"789f2687",
          4256 => x"ca386482",
          4257 => x"05704659",
          4258 => x"cf39b83d",
          4259 => x"ff841153",
          4260 => x"ff800551",
          4261 => x"e9f03f84",
          4262 => x"b9c80880",
          4263 => x"2ef8a038",
          4264 => x"b83dfefc",
          4265 => x"1153ff80",
          4266 => x"0551e9da",
          4267 => x"3f84b9c8",
          4268 => x"08802ef8",
          4269 => x"8a38b83d",
          4270 => x"fef81153",
          4271 => x"ff800551",
          4272 => x"e9c43f84",
          4273 => x"b9c80880",
          4274 => x"2ef7f438",
          4275 => x"83d7c451",
          4276 => x"ceb63f68",
          4277 => x"675d5978",
          4278 => x"7c27838d",
          4279 => x"38657033",
          4280 => x"7a335f5c",
          4281 => x"5a7a7d2e",
          4282 => x"95387a55",
          4283 => x"79547833",
          4284 => x"53785283",
          4285 => x"d7d451ce",
          4286 => x"8f3f6666",
          4287 => x"5b5c8119",
          4288 => x"811b4759",
          4289 => x"d239b83d",
          4290 => x"ff841153",
          4291 => x"ff800551",
          4292 => x"e8f43f84",
          4293 => x"b9c80880",
          4294 => x"2ef7a438",
          4295 => x"b83dfefc",
          4296 => x"1153ff80",
          4297 => x"0551e8de",
          4298 => x"3f84b9c8",
          4299 => x"08802ef7",
          4300 => x"8e38b83d",
          4301 => x"fef81153",
          4302 => x"ff800551",
          4303 => x"e8c83f84",
          4304 => x"b9c80880",
          4305 => x"2ef6f838",
          4306 => x"83d7f051",
          4307 => x"cdba3f68",
          4308 => x"5a796727",
          4309 => x"82933865",
          4310 => x"5c797081",
          4311 => x"055b337c",
          4312 => x"34658105",
          4313 => x"46eb39b8",
          4314 => x"3dff8411",
          4315 => x"53ff8005",
          4316 => x"51e8933f",
          4317 => x"84b9c808",
          4318 => x"802ef6c3",
          4319 => x"38b83dfe",
          4320 => x"fc1153ff",
          4321 => x"800551e7",
          4322 => x"fd3f84b9",
          4323 => x"c808b138",
          4324 => x"68703354",
          4325 => x"5283d7fc",
          4326 => x"51cced3f",
          4327 => x"84d5a808",
          4328 => x"5380f852",
          4329 => x"7e51ccfb",
          4330 => x"3f7e487e",
          4331 => x"335978ae",
          4332 => x"2ef68c38",
          4333 => x"789f2684",
          4334 => x"97386881",
          4335 => x"0549d139",
          4336 => x"68590280",
          4337 => x"db053379",
          4338 => x"34688105",
          4339 => x"49b83dfe",
          4340 => x"fc1153ff",
          4341 => x"800551e7",
          4342 => x"ad3f84b9",
          4343 => x"c808802e",
          4344 => x"f5dd3868",
          4345 => x"590280db",
          4346 => x"05337934",
          4347 => x"68810549",
          4348 => x"b83dfefc",
          4349 => x"1153ff80",
          4350 => x"0551e78a",
          4351 => x"3f84b9c8",
          4352 => x"08ffbd38",
          4353 => x"f5b939b8",
          4354 => x"3dff8411",
          4355 => x"53ff8005",
          4356 => x"51e6f33f",
          4357 => x"84b9c808",
          4358 => x"802ef5a3",
          4359 => x"38b83dfe",
          4360 => x"fc1153ff",
          4361 => x"800551e6",
          4362 => x"dd3f84b9",
          4363 => x"c808802e",
          4364 => x"f58d38b8",
          4365 => x"3dfef811",
          4366 => x"53ff8005",
          4367 => x"51e6c73f",
          4368 => x"84b9c808",
          4369 => x"863884b9",
          4370 => x"c8084683",
          4371 => x"d88851cb",
          4372 => x"b73f6867",
          4373 => x"5b59787a",
          4374 => x"278f3865",
          4375 => x"5b7a7970",
          4376 => x"84055b0c",
          4377 => x"797926f5",
          4378 => x"388a51d9",
          4379 => x"f13ff4cf",
          4380 => x"39b83dff",
          4381 => x"80055187",
          4382 => x"b13f84b9",
          4383 => x"c808b93d",
          4384 => x"ff800552",
          4385 => x"5988f33f",
          4386 => x"815384b9",
          4387 => x"c8085278",
          4388 => x"51ea833f",
          4389 => x"84b9c808",
          4390 => x"802ef4a3",
          4391 => x"3884b9c8",
          4392 => x"0851e7f6",
          4393 => x"3ff49839",
          4394 => x"b83dff84",
          4395 => x"1153ff80",
          4396 => x"0551e5d2",
          4397 => x"3f84b9c8",
          4398 => x"08913883",
          4399 => x"f2cc335a",
          4400 => x"79802e83",
          4401 => x"c03883f2",
          4402 => x"840849b8",
          4403 => x"3dfefc11",
          4404 => x"53ff8005",
          4405 => x"51e5af3f",
          4406 => x"84b9c808",
          4407 => x"913883f2",
          4408 => x"cc335a79",
          4409 => x"802e838a",
          4410 => x"3883f288",
          4411 => x"0847b83d",
          4412 => x"fef81153",
          4413 => x"ff800551",
          4414 => x"e58c3f84",
          4415 => x"b9c80880",
          4416 => x"2ea53880",
          4417 => x"665c5c7a",
          4418 => x"882e8338",
          4419 => x"815c7a90",
          4420 => x"32703070",
          4421 => x"72079f2a",
          4422 => x"7e065c5f",
          4423 => x"5d79802e",
          4424 => x"88387aa0",
          4425 => x"2e833888",
          4426 => x"4683d898",
          4427 => x"51d6c43f",
          4428 => x"80556854",
          4429 => x"65536652",
          4430 => x"6851eba8",
          4431 => x"3f83d8a4",
          4432 => x"51d6b03f",
          4433 => x"f2f93964",
          4434 => x"64710c59",
          4435 => x"64840545",
          4436 => x"b83dfef0",
          4437 => x"1153ff80",
          4438 => x"0551e2a6",
          4439 => x"3f84b9c8",
          4440 => x"08802ef2",
          4441 => x"da386464",
          4442 => x"710c5964",
          4443 => x"840545b8",
          4444 => x"3dfef011",
          4445 => x"53ff8005",
          4446 => x"51e2873f",
          4447 => x"84b9c808",
          4448 => x"c638f2bb",
          4449 => x"39645e02",
          4450 => x"80ce0522",
          4451 => x"7e708205",
          4452 => x"40237d45",
          4453 => x"b83dfef0",
          4454 => x"1153ff80",
          4455 => x"0551e1e2",
          4456 => x"3f84b9c8",
          4457 => x"08802ef2",
          4458 => x"9638645e",
          4459 => x"0280ce05",
          4460 => x"227e7082",
          4461 => x"0540237d",
          4462 => x"45b83dfe",
          4463 => x"f01153ff",
          4464 => x"800551e1",
          4465 => x"bd3f84b9",
          4466 => x"c808ffb9",
          4467 => x"38f1f039",
          4468 => x"b83dfefc",
          4469 => x"1153ff80",
          4470 => x"0551e3aa",
          4471 => x"3f84b9c8",
          4472 => x"08802e81",
          4473 => x"dc38685c",
          4474 => x"0280db05",
          4475 => x"337c3468",
          4476 => x"810549fb",
          4477 => x"9b39b83d",
          4478 => x"fef01153",
          4479 => x"ff800551",
          4480 => x"e1803f84",
          4481 => x"b9c80880",
          4482 => x"2e819838",
          4483 => x"6464710c",
          4484 => x"5d648405",
          4485 => x"704659f7",
          4486 => x"e1397a83",
          4487 => x"2e098106",
          4488 => x"f39d387b",
          4489 => x"5583d690",
          4490 => x"54805383",
          4491 => x"d8b0527c",
          4492 => x"51c8f53f",
          4493 => x"f396397b",
          4494 => x"527c51da",
          4495 => x"8a3ff38c",
          4496 => x"3983d8bc",
          4497 => x"51d4ac3f",
          4498 => x"f0f539b8",
          4499 => x"3dfef011",
          4500 => x"53ff8005",
          4501 => x"51e0ab3f",
          4502 => x"84b9c808",
          4503 => x"802eb838",
          4504 => x"64590280",
          4505 => x"ce052279",
          4506 => x"7082055b",
          4507 => x"237845f7",
          4508 => x"e73983f2",
          4509 => x"cd335c7b",
          4510 => x"802e80cf",
          4511 => x"3883f290",
          4512 => x"0847fcea",
          4513 => x"3983f2cd",
          4514 => x"335c7b80",
          4515 => x"2ea13883",
          4516 => x"f28c0849",
          4517 => x"fcb53983",
          4518 => x"d8e851d3",
          4519 => x"d63f6459",
          4520 => x"f7b63983",
          4521 => x"d8e851d3",
          4522 => x"ca3f6459",
          4523 => x"f6cc3983",
          4524 => x"f2ce3359",
          4525 => x"78802ea5",
          4526 => x"3883f294",
          4527 => x"0849fc8b",
          4528 => x"3983d8e8",
          4529 => x"51d3ac3f",
          4530 => x"f9c63983",
          4531 => x"f2ce3359",
          4532 => x"78802e9b",
          4533 => x"3883f298",
          4534 => x"0847fc92",
          4535 => x"3983f2cf",
          4536 => x"335e7d80",
          4537 => x"2e9b3883",
          4538 => x"f29c0849",
          4539 => x"fbdd3983",
          4540 => x"f2cf335e",
          4541 => x"7d802e9b",
          4542 => x"3883f2a0",
          4543 => x"0847fbee",
          4544 => x"3983f2ca",
          4545 => x"335d7c80",
          4546 => x"2e9b3883",
          4547 => x"f2a40849",
          4548 => x"fbb93983",
          4549 => x"f2ca335d",
          4550 => x"7c802e94",
          4551 => x"3883f2a8",
          4552 => x"0847fbca",
          4553 => x"3983f2b4",
          4554 => x"08fc8005",
          4555 => x"49fb9c39",
          4556 => x"83f2b408",
          4557 => x"880547fb",
          4558 => x"b539f33d",
          4559 => x"0d800b84",
          4560 => x"b9f83487",
          4561 => x"c0948c70",
          4562 => x"08565787",
          4563 => x"84805274",
          4564 => x"51dad23f",
          4565 => x"84b9c808",
          4566 => x"902b7708",
          4567 => x"57558784",
          4568 => x"80527551",
          4569 => x"dabf3f74",
          4570 => x"84b9c808",
          4571 => x"07770c87",
          4572 => x"c0949c70",
          4573 => x"08565787",
          4574 => x"84805274",
          4575 => x"51daa63f",
          4576 => x"84b9c808",
          4577 => x"902b7708",
          4578 => x"57558784",
          4579 => x"80527551",
          4580 => x"da933f74",
          4581 => x"84b9c808",
          4582 => x"07770c8c",
          4583 => x"80830b87",
          4584 => x"c094840c",
          4585 => x"8c80830b",
          4586 => x"87c09494",
          4587 => x"0c81bcf2",
          4588 => x"5c81c7f1",
          4589 => x"5d830284",
          4590 => x"05a10534",
          4591 => x"805e84d5",
          4592 => x"a80b893d",
          4593 => x"7088130c",
          4594 => x"70720c84",
          4595 => x"d5ac0c56",
          4596 => x"b7853f89",
          4597 => x"9e3f9597",
          4598 => x"3fba8d51",
          4599 => x"958c3f83",
          4600 => x"d2b05283",
          4601 => x"d2b451c4",
          4602 => x"9f3f83f2",
          4603 => x"b8702252",
          4604 => x"5594973f",
          4605 => x"83d2bc54",
          4606 => x"83d2c853",
          4607 => x"81153352",
          4608 => x"83d2d051",
          4609 => x"c4823f8d",
          4610 => x"b23f83d2",
          4611 => x"ec51d0e3",
          4612 => x"3f805283",
          4613 => x"d2f051c3",
          4614 => x"ef3f9080",
          4615 => x"0a5283d3",
          4616 => x"9851c3e4",
          4617 => x"3fece73f",
          4618 => x"8004fb3d",
          4619 => x"0d777008",
          4620 => x"56568075",
          4621 => x"52537473",
          4622 => x"2e818338",
          4623 => x"74337081",
          4624 => x"ff065252",
          4625 => x"70a02e09",
          4626 => x"81069138",
          4627 => x"81157033",
          4628 => x"7081ff06",
          4629 => x"53535570",
          4630 => x"a02ef138",
          4631 => x"7181ff06",
          4632 => x"5473a22e",
          4633 => x"81823874",
          4634 => x"5272812e",
          4635 => x"80e73880",
          4636 => x"72337081",
          4637 => x"ff065354",
          4638 => x"5470a02e",
          4639 => x"83388154",
          4640 => x"70802e8b",
          4641 => x"3873802e",
          4642 => x"86388112",
          4643 => x"52e13980",
          4644 => x"7381ff06",
          4645 => x"525470a0",
          4646 => x"2e098106",
          4647 => x"83388154",
          4648 => x"70a23270",
          4649 => x"30708025",
          4650 => x"76075252",
          4651 => x"5372802e",
          4652 => x"88388072",
          4653 => x"70810554",
          4654 => x"3471760c",
          4655 => x"74517084",
          4656 => x"b9c80c87",
          4657 => x"3d0d0470",
          4658 => x"802ec438",
          4659 => x"73802eff",
          4660 => x"be388112",
          4661 => x"52807233",
          4662 => x"7081ff06",
          4663 => x"53545470",
          4664 => x"a22ee438",
          4665 => x"8154e039",
          4666 => x"81155581",
          4667 => x"75535372",
          4668 => x"812e0981",
          4669 => x"06fef838",
          4670 => x"dc39fc3d",
          4671 => x"0d765372",
          4672 => x"088b3880",
          4673 => x"0b84b9c8",
          4674 => x"0c863d0d",
          4675 => x"04863dfc",
          4676 => x"05527251",
          4677 => x"daec3f84",
          4678 => x"b9c80880",
          4679 => x"2ee53874",
          4680 => x"84b9c80c",
          4681 => x"863d0d04",
          4682 => x"fc3d0d76",
          4683 => x"821133ff",
          4684 => x"05525381",
          4685 => x"52708b26",
          4686 => x"81983883",
          4687 => x"1333ff05",
          4688 => x"54825273",
          4689 => x"9e26818a",
          4690 => x"38841333",
          4691 => x"51835270",
          4692 => x"972680fe",
          4693 => x"38851333",
          4694 => x"54845273",
          4695 => x"bb2680f2",
          4696 => x"38861333",
          4697 => x"55855274",
          4698 => x"bb2680e6",
          4699 => x"38881322",
          4700 => x"55865274",
          4701 => x"87e72680",
          4702 => x"d9388a13",
          4703 => x"22548752",
          4704 => x"7387e726",
          4705 => x"80cc3881",
          4706 => x"0b87c098",
          4707 => x"9c0c7222",
          4708 => x"87c098bc",
          4709 => x"0c821333",
          4710 => x"87c098b8",
          4711 => x"0c831333",
          4712 => x"87c098b4",
          4713 => x"0c841333",
          4714 => x"87c098b0",
          4715 => x"0c851333",
          4716 => x"87c098ac",
          4717 => x"0c861333",
          4718 => x"87c098a8",
          4719 => x"0c7487c0",
          4720 => x"98a40c73",
          4721 => x"87c098a0",
          4722 => x"0c800b87",
          4723 => x"c0989c0c",
          4724 => x"80527184",
          4725 => x"b9c80c86",
          4726 => x"3d0d04f3",
          4727 => x"3d0d7f5b",
          4728 => x"87c0989c",
          4729 => x"5d817d0c",
          4730 => x"87c098bc",
          4731 => x"085e7d7b",
          4732 => x"2387c098",
          4733 => x"b8085c7b",
          4734 => x"821c3487",
          4735 => x"c098b408",
          4736 => x"5a79831c",
          4737 => x"3487c098",
          4738 => x"b0085c7b",
          4739 => x"841c3487",
          4740 => x"c098ac08",
          4741 => x"5a79851c",
          4742 => x"3487c098",
          4743 => x"a8085c7b",
          4744 => x"861c3487",
          4745 => x"c098a408",
          4746 => x"5c7b881c",
          4747 => x"2387c098",
          4748 => x"a0085a79",
          4749 => x"8a1c2380",
          4750 => x"7d0c7983",
          4751 => x"ffff0659",
          4752 => x"7b83ffff",
          4753 => x"0658861b",
          4754 => x"3357851b",
          4755 => x"3356841b",
          4756 => x"3355831b",
          4757 => x"3354821b",
          4758 => x"33537d83",
          4759 => x"ffff0652",
          4760 => x"83d8ec51",
          4761 => x"ffbfa13f",
          4762 => x"8f3d0d04",
          4763 => x"fe3d0d02",
          4764 => x"93053353",
          4765 => x"72812ea8",
          4766 => x"38725180",
          4767 => x"e8a63f84",
          4768 => x"b9c80898",
          4769 => x"2b70982c",
          4770 => x"515271ff",
          4771 => x"2e098106",
          4772 => x"86387283",
          4773 => x"2ee33871",
          4774 => x"84b9c80c",
          4775 => x"843d0d04",
          4776 => x"725180e7",
          4777 => x"ff3f84b9",
          4778 => x"c808982b",
          4779 => x"70982c51",
          4780 => x"5271ff2e",
          4781 => x"098106df",
          4782 => x"38725180",
          4783 => x"e7e63f84",
          4784 => x"b9c80898",
          4785 => x"2b70982c",
          4786 => x"515271ff",
          4787 => x"2ed238c7",
          4788 => x"39fd3d0d",
          4789 => x"80705452",
          4790 => x"71882b54",
          4791 => x"815180e7",
          4792 => x"c33f84b9",
          4793 => x"c808982b",
          4794 => x"70982c51",
          4795 => x"5271ff2e",
          4796 => x"eb387372",
          4797 => x"07811454",
          4798 => x"52837325",
          4799 => x"db387184",
          4800 => x"b9c80c85",
          4801 => x"3d0d04fc",
          4802 => x"3d0d029b",
          4803 => x"053383f2",
          4804 => x"80337081",
          4805 => x"ff065355",
          4806 => x"5570802e",
          4807 => x"80f43887",
          4808 => x"c0949408",
          4809 => x"70962a70",
          4810 => x"81065354",
          4811 => x"5270802e",
          4812 => x"8c387191",
          4813 => x"2a708106",
          4814 => x"515170e3",
          4815 => x"38728132",
          4816 => x"81065372",
          4817 => x"802e8a38",
          4818 => x"71932a81",
          4819 => x"065271cf",
          4820 => x"387381ff",
          4821 => x"065187c0",
          4822 => x"94805270",
          4823 => x"802e8638",
          4824 => x"87c09490",
          4825 => x"5274720c",
          4826 => x"7484b9c8",
          4827 => x"0c863d0d",
          4828 => x"0471912a",
          4829 => x"70810651",
          4830 => x"51709738",
          4831 => x"72813281",
          4832 => x"06537280",
          4833 => x"2ecb3871",
          4834 => x"932a8106",
          4835 => x"5271802e",
          4836 => x"c03887c0",
          4837 => x"94840870",
          4838 => x"962a7081",
          4839 => x"06535452",
          4840 => x"70cf38d8",
          4841 => x"39ff3d0d",
          4842 => x"028f0533",
          4843 => x"7030709f",
          4844 => x"2a515252",
          4845 => x"7083f280",
          4846 => x"34833d0d",
          4847 => x"04fa3d0d",
          4848 => x"78558075",
          4849 => x"33705652",
          4850 => x"5770772e",
          4851 => x"80e73881",
          4852 => x"1583f280",
          4853 => x"337081ff",
          4854 => x"06545755",
          4855 => x"71802e80",
          4856 => x"ff3887c0",
          4857 => x"94940870",
          4858 => x"962a7081",
          4859 => x"06535452",
          4860 => x"70802e8c",
          4861 => x"3871912a",
          4862 => x"70810651",
          4863 => x"5170e338",
          4864 => x"72813281",
          4865 => x"06537280",
          4866 => x"2e8a3871",
          4867 => x"932a8106",
          4868 => x"5271cf38",
          4869 => x"7581ff06",
          4870 => x"5187c094",
          4871 => x"80527080",
          4872 => x"2e863887",
          4873 => x"c0949052",
          4874 => x"73720c81",
          4875 => x"17753355",
          4876 => x"5773ff9b",
          4877 => x"387684b9",
          4878 => x"c80c883d",
          4879 => x"0d047191",
          4880 => x"2a708106",
          4881 => x"51517098",
          4882 => x"38728132",
          4883 => x"81065372",
          4884 => x"802ec138",
          4885 => x"71932a81",
          4886 => x"06527180",
          4887 => x"2effb538",
          4888 => x"87c09484",
          4889 => x"0870962a",
          4890 => x"70810653",
          4891 => x"545270ce",
          4892 => x"38d739ff",
          4893 => x"3d0d87c0",
          4894 => x"9e800870",
          4895 => x"9c2a8a06",
          4896 => x"52527080",
          4897 => x"2e84ab38",
          4898 => x"87c09ea4",
          4899 => x"0883f284",
          4900 => x"0c87c09e",
          4901 => x"a80883f2",
          4902 => x"880c87c0",
          4903 => x"9e940883",
          4904 => x"f28c0c87",
          4905 => x"c09e9808",
          4906 => x"83f2900c",
          4907 => x"87c09e9c",
          4908 => x"0883f294",
          4909 => x"0c87c09e",
          4910 => x"a00883f2",
          4911 => x"980c87c0",
          4912 => x"9eac0883",
          4913 => x"f29c0c87",
          4914 => x"c09eb008",
          4915 => x"83f2a00c",
          4916 => x"87c09eb4",
          4917 => x"0883f2a4",
          4918 => x"0c87c09e",
          4919 => x"b80883f2",
          4920 => x"a80c87c0",
          4921 => x"9ebc0883",
          4922 => x"f2ac0c87",
          4923 => x"c09ec008",
          4924 => x"83f2b00c",
          4925 => x"87c09ec4",
          4926 => x"0883f2b4",
          4927 => x"0c87c09e",
          4928 => x"80085271",
          4929 => x"83f2b823",
          4930 => x"87c09e84",
          4931 => x"0883f2bc",
          4932 => x"0c87c09e",
          4933 => x"880883f2",
          4934 => x"c00c87c0",
          4935 => x"9e8c0883",
          4936 => x"f2c40c81",
          4937 => x"0b83f2c8",
          4938 => x"34800b87",
          4939 => x"c09e9008",
          4940 => x"7084800a",
          4941 => x"06515252",
          4942 => x"7082fb38",
          4943 => x"7183f2c9",
          4944 => x"34800b87",
          4945 => x"c09e9008",
          4946 => x"7088800a",
          4947 => x"06515252",
          4948 => x"70802e83",
          4949 => x"38815271",
          4950 => x"83f2ca34",
          4951 => x"800b87c0",
          4952 => x"9e900870",
          4953 => x"90800a06",
          4954 => x"51525270",
          4955 => x"802e8338",
          4956 => x"81527183",
          4957 => x"f2cb3480",
          4958 => x"0b87c09e",
          4959 => x"90087088",
          4960 => x"80800651",
          4961 => x"52527080",
          4962 => x"2e833881",
          4963 => x"527183f2",
          4964 => x"cc34800b",
          4965 => x"87c09e90",
          4966 => x"0870a080",
          4967 => x"80065152",
          4968 => x"5270802e",
          4969 => x"83388152",
          4970 => x"7183f2cd",
          4971 => x"34800b87",
          4972 => x"c09e9008",
          4973 => x"70908080",
          4974 => x"06515252",
          4975 => x"70802e83",
          4976 => x"38815271",
          4977 => x"83f2ce34",
          4978 => x"800b87c0",
          4979 => x"9e900870",
          4980 => x"84808006",
          4981 => x"51525270",
          4982 => x"802e8338",
          4983 => x"81527183",
          4984 => x"f2cf3480",
          4985 => x"0b87c09e",
          4986 => x"90087082",
          4987 => x"80800651",
          4988 => x"52527080",
          4989 => x"2e833881",
          4990 => x"527183f2",
          4991 => x"d034800b",
          4992 => x"87c09e90",
          4993 => x"08708180",
          4994 => x"80065152",
          4995 => x"5270802e",
          4996 => x"83388152",
          4997 => x"7183f2d1",
          4998 => x"34800b87",
          4999 => x"c09e9008",
          5000 => x"7080c080",
          5001 => x"06515252",
          5002 => x"70802e83",
          5003 => x"38815271",
          5004 => x"83f2d234",
          5005 => x"800b87c0",
          5006 => x"9e900870",
          5007 => x"a0800651",
          5008 => x"52527080",
          5009 => x"2e833881",
          5010 => x"527183f2",
          5011 => x"d33487c0",
          5012 => x"9e900898",
          5013 => x"8006708a",
          5014 => x"2a535171",
          5015 => x"83f2d434",
          5016 => x"800b87c0",
          5017 => x"9e900870",
          5018 => x"84800651",
          5019 => x"52527080",
          5020 => x"2e833881",
          5021 => x"527183f2",
          5022 => x"d53487c0",
          5023 => x"9e900883",
          5024 => x"f0067084",
          5025 => x"2a535171",
          5026 => x"83f2d634",
          5027 => x"800b87c0",
          5028 => x"9e900870",
          5029 => x"88065152",
          5030 => x"5270802e",
          5031 => x"83388152",
          5032 => x"7183f2d7",
          5033 => x"3487c09e",
          5034 => x"90088706",
          5035 => x"517083f2",
          5036 => x"d834833d",
          5037 => x"0d048152",
          5038 => x"fd8239fb",
          5039 => x"3d0d83d9",
          5040 => x"8451ffb6",
          5041 => x"c33f83f2",
          5042 => x"c8335473",
          5043 => x"869f3883",
          5044 => x"d99851c3",
          5045 => x"9e3f83f2",
          5046 => x"ca335574",
          5047 => x"85ef3883",
          5048 => x"f2cf3354",
          5049 => x"7385c638",
          5050 => x"83f2cc33",
          5051 => x"5675859d",
          5052 => x"3883f2cd",
          5053 => x"33557484",
          5054 => x"f43883f2",
          5055 => x"ce335473",
          5056 => x"84cb3883",
          5057 => x"f2d33356",
          5058 => x"7584a838",
          5059 => x"83f2d733",
          5060 => x"54738485",
          5061 => x"3883f2d5",
          5062 => x"33557483",
          5063 => x"e23883f2",
          5064 => x"c9335675",
          5065 => x"83c43883",
          5066 => x"f2cb3354",
          5067 => x"7383a638",
          5068 => x"83f2d033",
          5069 => x"55748388",
          5070 => x"3883f2d1",
          5071 => x"33567582",
          5072 => x"e93883f2",
          5073 => x"d2335473",
          5074 => x"81e13883",
          5075 => x"d9b051c2",
          5076 => x"a23f83f2",
          5077 => x"ac085283",
          5078 => x"d9bc51ff",
          5079 => x"b5aa3f83",
          5080 => x"f2b00852",
          5081 => x"83d9e451",
          5082 => x"ffb59d3f",
          5083 => x"83f2b408",
          5084 => x"5283da8c",
          5085 => x"51ffb590",
          5086 => x"3f83dab4",
          5087 => x"51c1f43f",
          5088 => x"83f2b822",
          5089 => x"5283dabc",
          5090 => x"51ffb4fc",
          5091 => x"3f83f2bc",
          5092 => x"0856bd84",
          5093 => x"c0527551",
          5094 => x"ca8b3f84",
          5095 => x"b9c808bd",
          5096 => x"84c02976",
          5097 => x"71315454",
          5098 => x"84b9c808",
          5099 => x"5283dae4",
          5100 => x"51ffb4d4",
          5101 => x"3f83f2cf",
          5102 => x"335574b9",
          5103 => x"3883f2ca",
          5104 => x"33557485",
          5105 => x"38873d0d",
          5106 => x"0483f2c4",
          5107 => x"0856bd84",
          5108 => x"c0527551",
          5109 => x"c9cf3f84",
          5110 => x"b9c808bd",
          5111 => x"84c02976",
          5112 => x"71315454",
          5113 => x"84b9c808",
          5114 => x"5283db90",
          5115 => x"51ffb498",
          5116 => x"3f873d0d",
          5117 => x"0483f2c0",
          5118 => x"0856bd84",
          5119 => x"c0527551",
          5120 => x"c9a33f84",
          5121 => x"b9c808bd",
          5122 => x"84c02976",
          5123 => x"71315454",
          5124 => x"84b9c808",
          5125 => x"5283dbbc",
          5126 => x"51ffb3ec",
          5127 => x"3f83f2ca",
          5128 => x"33557480",
          5129 => x"2eff9e38",
          5130 => x"ff9f3983",
          5131 => x"dbe851c0",
          5132 => x"c23f83d9",
          5133 => x"b051c0bb",
          5134 => x"3f83f2ac",
          5135 => x"085283d9",
          5136 => x"bc51ffb3",
          5137 => x"c33f83f2",
          5138 => x"b0085283",
          5139 => x"d9e451ff",
          5140 => x"b3b63f83",
          5141 => x"f2b40852",
          5142 => x"83da8c51",
          5143 => x"ffb3a93f",
          5144 => x"83dab451",
          5145 => x"c08d3f83",
          5146 => x"f2b82252",
          5147 => x"83dabc51",
          5148 => x"ffb3953f",
          5149 => x"83f2bc08",
          5150 => x"56bd84c0",
          5151 => x"527551c8",
          5152 => x"a43f84b9",
          5153 => x"c808bd84",
          5154 => x"c0297671",
          5155 => x"31545484",
          5156 => x"b9c80852",
          5157 => x"83dae451",
          5158 => x"ffb2ed3f",
          5159 => x"83f2cf33",
          5160 => x"5574802e",
          5161 => x"fe9738fe",
          5162 => x"cc3983db",
          5163 => x"f051ffbf",
          5164 => x"c23f83f2",
          5165 => x"d2335473",
          5166 => x"802efd8f",
          5167 => x"38feec39",
          5168 => x"83dbf851",
          5169 => x"ffbfac3f",
          5170 => x"83f2d133",
          5171 => x"5675802e",
          5172 => x"fcf038d6",
          5173 => x"3983dc84",
          5174 => x"51ffbf97",
          5175 => x"3f83f2d0",
          5176 => x"33557480",
          5177 => x"2efcd238",
          5178 => x"d73983dc",
          5179 => x"9051ffbf",
          5180 => x"823f83f2",
          5181 => x"cb335473",
          5182 => x"802efcb4",
          5183 => x"38d73983",
          5184 => x"f2d63352",
          5185 => x"83dca451",
          5186 => x"ffb1fd3f",
          5187 => x"83f2c933",
          5188 => x"5675802e",
          5189 => x"fc9138d2",
          5190 => x"3983f2d8",
          5191 => x"335283dc",
          5192 => x"c451ffb1",
          5193 => x"e33f83f2",
          5194 => x"d5335574",
          5195 => x"802efbee",
          5196 => x"38cd3983",
          5197 => x"f2d43352",
          5198 => x"83dce451",
          5199 => x"ffb1c93f",
          5200 => x"83f2d733",
          5201 => x"5473802e",
          5202 => x"fbcb38cd",
          5203 => x"3983f294",
          5204 => x"0883f298",
          5205 => x"08115452",
          5206 => x"83dd8451",
          5207 => x"ffb1a93f",
          5208 => x"83f2d333",
          5209 => x"5675802e",
          5210 => x"fba238c7",
          5211 => x"3983f28c",
          5212 => x"0883f290",
          5213 => x"08115452",
          5214 => x"83dda051",
          5215 => x"ffb1893f",
          5216 => x"83f2ce33",
          5217 => x"5473802e",
          5218 => x"faf938c1",
          5219 => x"3983f284",
          5220 => x"0883f288",
          5221 => x"08115452",
          5222 => x"83ddbc51",
          5223 => x"ffb0e93f",
          5224 => x"83f2cd33",
          5225 => x"5574802e",
          5226 => x"fad038c1",
          5227 => x"3983f29c",
          5228 => x"0883f2a0",
          5229 => x"08115452",
          5230 => x"83ddd851",
          5231 => x"ffb0c93f",
          5232 => x"83f2cc33",
          5233 => x"5675802e",
          5234 => x"faa738c1",
          5235 => x"3983f2a4",
          5236 => x"0883f2a8",
          5237 => x"08115452",
          5238 => x"83ddf451",
          5239 => x"ffb0a93f",
          5240 => x"83f2cf33",
          5241 => x"5473802e",
          5242 => x"f9fe38c1",
          5243 => x"3983de90",
          5244 => x"51ffb094",
          5245 => x"3f83d998",
          5246 => x"51ffbcf7",
          5247 => x"3f83f2ca",
          5248 => x"33557480",
          5249 => x"2ef9d838",
          5250 => x"c439ff3d",
          5251 => x"0d028e05",
          5252 => x"33527185",
          5253 => x"268c3871",
          5254 => x"101083c2",
          5255 => x"fc055271",
          5256 => x"080483de",
          5257 => x"a451ffaf",
          5258 => x"df3f833d",
          5259 => x"0d0483de",
          5260 => x"ac51ffaf",
          5261 => x"d33f833d",
          5262 => x"0d0483de",
          5263 => x"b451ffaf",
          5264 => x"c73f833d",
          5265 => x"0d0483de",
          5266 => x"bc51ffaf",
          5267 => x"bb3f833d",
          5268 => x"0d0483de",
          5269 => x"c451ffaf",
          5270 => x"af3f833d",
          5271 => x"0d0483de",
          5272 => x"cc51ffaf",
          5273 => x"a33f833d",
          5274 => x"0d047188",
          5275 => x"800c0480",
          5276 => x"0b87c096",
          5277 => x"840c0483",
          5278 => x"f2dc0887",
          5279 => x"c096840c",
          5280 => x"04d93d0d",
          5281 => x"aa3d08ad",
          5282 => x"3d085a5a",
          5283 => x"81705758",
          5284 => x"805283f3",
          5285 => x"b4085182",
          5286 => x"88833f84",
          5287 => x"b9c80880",
          5288 => x"ed388b3d",
          5289 => x"57ff0b83",
          5290 => x"f3b40854",
          5291 => x"5580f852",
          5292 => x"765182d2",
          5293 => x"903f84b9",
          5294 => x"c808802e",
          5295 => x"a4387651",
          5296 => x"c0e63f84",
          5297 => x"b9c80881",
          5298 => x"17575580",
          5299 => x"0b84b9c8",
          5300 => x"08258e38",
          5301 => x"84b9c808",
          5302 => x"ff057018",
          5303 => x"55558074",
          5304 => x"34740970",
          5305 => x"30707207",
          5306 => x"9f2a5155",
          5307 => x"5578762e",
          5308 => x"853873ff",
          5309 => x"b03883f3",
          5310 => x"b4088c11",
          5311 => x"08535182",
          5312 => x"879b3f84",
          5313 => x"b9c8088f",
          5314 => x"3878762e",
          5315 => x"9a387784",
          5316 => x"b9c80ca9",
          5317 => x"3d0d0483",
          5318 => x"e1fc51ff",
          5319 => x"adea3f78",
          5320 => x"762e0981",
          5321 => x"06e83876",
          5322 => x"527951c0",
          5323 => x"9a3f7951",
          5324 => x"ffbff53f",
          5325 => x"ab3d0856",
          5326 => x"84b9c808",
          5327 => x"76347652",
          5328 => x"83e2a851",
          5329 => x"ffadc13f",
          5330 => x"800b84b9",
          5331 => x"c80ca93d",
          5332 => x"0d04d83d",
          5333 => x"0dab3d08",
          5334 => x"ad3d0871",
          5335 => x"725d7233",
          5336 => x"57575a57",
          5337 => x"73a02e81",
          5338 => x"9138800b",
          5339 => x"8d3d5956",
          5340 => x"75101010",
          5341 => x"83f3bc05",
          5342 => x"70085254",
          5343 => x"ffbfa93f",
          5344 => x"84b9c808",
          5345 => x"53795273",
          5346 => x"0851c089",
          5347 => x"3f84b9c8",
          5348 => x"08903884",
          5349 => x"14335473",
          5350 => x"812e8188",
          5351 => x"3873822e",
          5352 => x"99388116",
          5353 => x"7081ff06",
          5354 => x"57548276",
          5355 => x"27c23880",
          5356 => x"547384b9",
          5357 => x"c80caa3d",
          5358 => x"0d04811a",
          5359 => x"5aaa3dff",
          5360 => x"841153ff",
          5361 => x"800551c7",
          5362 => x"bd3f84b9",
          5363 => x"c808802e",
          5364 => x"d138ff1b",
          5365 => x"53785276",
          5366 => x"51fda63f",
          5367 => x"84b9c808",
          5368 => x"81ff0654",
          5369 => x"73802ec9",
          5370 => x"38811670",
          5371 => x"81ff0657",
          5372 => x"54827627",
          5373 => x"fefa38ff",
          5374 => x"b6397833",
          5375 => x"77055676",
          5376 => x"7627fee6",
          5377 => x"38811570",
          5378 => x"5b703355",
          5379 => x"5573a02e",
          5380 => x"098106fe",
          5381 => x"d5387575",
          5382 => x"26eb3880",
          5383 => x"0b8d3d59",
          5384 => x"56fecd39",
          5385 => x"7384b9c8",
          5386 => x"085383f3",
          5387 => x"b4085256",
          5388 => x"8284ea3f",
          5389 => x"84b9c808",
          5390 => x"80d03883",
          5391 => x"f3b40853",
          5392 => x"80f85277",
          5393 => x"5182cefd",
          5394 => x"3f84b9c8",
          5395 => x"08802eba",
          5396 => x"387751ff",
          5397 => x"bdd23f84",
          5398 => x"b9c80855",
          5399 => x"800b84b9",
          5400 => x"c808259d",
          5401 => x"3884b9c8",
          5402 => x"08ff0570",
          5403 => x"19585580",
          5404 => x"77347753",
          5405 => x"75528116",
          5406 => x"83e1f052",
          5407 => x"56ffab88",
          5408 => x"3f74ff2e",
          5409 => x"098106ff",
          5410 => x"b238810b",
          5411 => x"84b9c80c",
          5412 => x"aa3d0d04",
          5413 => x"ce3d0db5",
          5414 => x"3d08b73d",
          5415 => x"08b93d08",
          5416 => x"5a415c80",
          5417 => x"0bb43d34",
          5418 => x"83f3b833",
          5419 => x"83f3b408",
          5420 => x"565d749e",
          5421 => x"387483f3",
          5422 => x"b0335656",
          5423 => x"74802e82",
          5424 => x"cb387780",
          5425 => x"2e918d38",
          5426 => x"81707706",
          5427 => x"5a577890",
          5428 => x"a0387780",
          5429 => x"2e90fd38",
          5430 => x"933db43d",
          5431 => x"5f5f8051",
          5432 => x"eb8a3f84",
          5433 => x"b9c80898",
          5434 => x"2b70982c",
          5435 => x"5b5679ff",
          5436 => x"2eec3879",
          5437 => x"81ff0684",
          5438 => x"d1843370",
          5439 => x"982b7098",
          5440 => x"2c84d180",
          5441 => x"3370982b",
          5442 => x"70972c71",
          5443 => x"982c0570",
          5444 => x"101083de",
          5445 => x"d0057008",
          5446 => x"15703352",
          5447 => x"535c5d46",
          5448 => x"525b585c",
          5449 => x"59815774",
          5450 => x"792e80cd",
          5451 => x"38787527",
          5452 => x"81873875",
          5453 => x"81800a29",
          5454 => x"81ff0a05",
          5455 => x"70982c57",
          5456 => x"55807624",
          5457 => x"81cb3875",
          5458 => x"10167082",
          5459 => x"2b565780",
          5460 => x"0b83ded4",
          5461 => x"16334257",
          5462 => x"77612591",
          5463 => x"3883ded0",
          5464 => x"15081870",
          5465 => x"33564178",
          5466 => x"752e8195",
          5467 => x"3876802e",
          5468 => x"c2387584",
          5469 => x"d1803481",
          5470 => x"5776802e",
          5471 => x"81993881",
          5472 => x"1b70982b",
          5473 => x"70982c84",
          5474 => x"d1803370",
          5475 => x"982b7097",
          5476 => x"2c71982c",
          5477 => x"0570822b",
          5478 => x"83ded411",
          5479 => x"335f535f",
          5480 => x"5d585d57",
          5481 => x"577a782e",
          5482 => x"81903876",
          5483 => x"84d18434",
          5484 => x"feac3981",
          5485 => x"5776ffba",
          5486 => x"38758180",
          5487 => x"0a298180",
          5488 => x"0a057098",
          5489 => x"2c7081ff",
          5490 => x"06595741",
          5491 => x"76952680",
          5492 => x"c0387510",
          5493 => x"1670822b",
          5494 => x"5155800b",
          5495 => x"83ded416",
          5496 => x"33425777",
          5497 => x"6125ce38",
          5498 => x"83ded015",
          5499 => x"08187033",
          5500 => x"42557861",
          5501 => x"2effbc38",
          5502 => x"76802eff",
          5503 => x"bc38fef2",
          5504 => x"39815776",
          5505 => x"802efeab",
          5506 => x"38fee739",
          5507 => x"8156fdb2",
          5508 => x"39805776",
          5509 => x"fee93876",
          5510 => x"84d18434",
          5511 => x"7684d180",
          5512 => x"34797e34",
          5513 => x"767f0c62",
          5514 => x"55749526",
          5515 => x"fdb03874",
          5516 => x"101083c3",
          5517 => x"94055776",
          5518 => x"080483de",
          5519 => x"d815087f",
          5520 => x"0c800b84",
          5521 => x"d1843480",
          5522 => x"0b84d180",
          5523 => x"34d93984",
          5524 => x"d18c3356",
          5525 => x"75802efd",
          5526 => x"853884d5",
          5527 => x"ac085288",
          5528 => x"51ffb68a",
          5529 => x"3f84d18c",
          5530 => x"33ff0557",
          5531 => x"7684d18c",
          5532 => x"34fceb39",
          5533 => x"84d18c33",
          5534 => x"7081ff06",
          5535 => x"84d18833",
          5536 => x"5b575575",
          5537 => x"7927fcd6",
          5538 => x"3884d5ac",
          5539 => x"08528115",
          5540 => x"587784d1",
          5541 => x"8c347b16",
          5542 => x"70335255",
          5543 => x"ffb5cf3f",
          5544 => x"fcbc397c",
          5545 => x"932e8bda",
          5546 => x"387c1010",
          5547 => x"83f2e405",
          5548 => x"70085759",
          5549 => x"758f8338",
          5550 => x"7584d188",
          5551 => x"34757c34",
          5552 => x"84d18833",
          5553 => x"84d18c33",
          5554 => x"56567480",
          5555 => x"2eb63884",
          5556 => x"d5ac0852",
          5557 => x"8851ffb5",
          5558 => x"953f84d5",
          5559 => x"ac0852a0",
          5560 => x"51ffb58a",
          5561 => x"3f84d5ac",
          5562 => x"08528851",
          5563 => x"ffb4ff3f",
          5564 => x"84d18c33",
          5565 => x"ff055b7a",
          5566 => x"84d18c34",
          5567 => x"7a81ff06",
          5568 => x"5574cc38",
          5569 => x"7b51ffa5",
          5570 => x"ff3f7584",
          5571 => x"d18c34fb",
          5572 => x"cd397c8a",
          5573 => x"3883f3ac",
          5574 => x"0856758d",
          5575 => x"9e387c10",
          5576 => x"1083f2e0",
          5577 => x"05fc1108",
          5578 => x"5755758e",
          5579 => x"f9387408",
          5580 => x"5675802e",
          5581 => x"fba83875",
          5582 => x"51ffb7ec",
          5583 => x"3f84b9c8",
          5584 => x"0884d188",
          5585 => x"3484b9c8",
          5586 => x"0881ff06",
          5587 => x"81055375",
          5588 => x"527b51ff",
          5589 => x"b8943f84",
          5590 => x"d1883384",
          5591 => x"d18c3356",
          5592 => x"5674802e",
          5593 => x"ff9e3884",
          5594 => x"d5ac0852",
          5595 => x"8851ffb3",
          5596 => x"fd3f84d5",
          5597 => x"ac0852a0",
          5598 => x"51ffb3f2",
          5599 => x"3f84d5ac",
          5600 => x"08528851",
          5601 => x"ffb3e73f",
          5602 => x"84d18c33",
          5603 => x"ff055574",
          5604 => x"84d18c34",
          5605 => x"7481ff06",
          5606 => x"55c73984",
          5607 => x"d18c3370",
          5608 => x"81ff0684",
          5609 => x"d188335b",
          5610 => x"57557579",
          5611 => x"27faaf38",
          5612 => x"84d5ac08",
          5613 => x"52811557",
          5614 => x"7684d18c",
          5615 => x"347b1670",
          5616 => x"335255ff",
          5617 => x"b3a83f84",
          5618 => x"d18c3370",
          5619 => x"81ff0684",
          5620 => x"d188335a",
          5621 => x"57557578",
          5622 => x"27fa8338",
          5623 => x"84d5ac08",
          5624 => x"52811557",
          5625 => x"7684d18c",
          5626 => x"347b1670",
          5627 => x"335255ff",
          5628 => x"b2fc3f84",
          5629 => x"d18c3370",
          5630 => x"81ff0684",
          5631 => x"d188335a",
          5632 => x"57557776",
          5633 => x"26ffa938",
          5634 => x"f9d43984",
          5635 => x"d18c3384",
          5636 => x"d1883356",
          5637 => x"5674762e",
          5638 => x"f9c438ff",
          5639 => x"155b7a84",
          5640 => x"d1883475",
          5641 => x"982b7098",
          5642 => x"2c7c81ff",
          5643 => x"0643575a",
          5644 => x"60762480",
          5645 => x"ef3884d5",
          5646 => x"ac0852a0",
          5647 => x"51ffb2ae",
          5648 => x"3f84d18c",
          5649 => x"3370982b",
          5650 => x"70982c84",
          5651 => x"d188335a",
          5652 => x"57574174",
          5653 => x"7724f986",
          5654 => x"3884d5ac",
          5655 => x"08528851",
          5656 => x"ffb28b3f",
          5657 => x"7481800a",
          5658 => x"2981800a",
          5659 => x"0570982c",
          5660 => x"84d18833",
          5661 => x"5d565a74",
          5662 => x"7b24f8e2",
          5663 => x"3884d5ac",
          5664 => x"08528851",
          5665 => x"ffb1e73f",
          5666 => x"7481800a",
          5667 => x"2981800a",
          5668 => x"0570982c",
          5669 => x"84d18833",
          5670 => x"5d565a7a",
          5671 => x"7525ffb9",
          5672 => x"38f8bb39",
          5673 => x"7b165881",
          5674 => x"18337834",
          5675 => x"84d5ac08",
          5676 => x"52773351",
          5677 => x"ffb1b73f",
          5678 => x"7581800a",
          5679 => x"2981800a",
          5680 => x"0570982c",
          5681 => x"84d18833",
          5682 => x"5b575575",
          5683 => x"7925fee6",
          5684 => x"387b1658",
          5685 => x"81183378",
          5686 => x"3484d5ac",
          5687 => x"08527733",
          5688 => x"51ffb18a",
          5689 => x"3f758180",
          5690 => x"0a298180",
          5691 => x"0a057098",
          5692 => x"2c84d188",
          5693 => x"335b5755",
          5694 => x"787624ff",
          5695 => x"a738feb6",
          5696 => x"3984d18c",
          5697 => x"33557480",
          5698 => x"2ef7d338",
          5699 => x"84d5ac08",
          5700 => x"528851ff",
          5701 => x"b0d83f84",
          5702 => x"d18c33ff",
          5703 => x"05577684",
          5704 => x"d18c3476",
          5705 => x"81ff0655",
          5706 => x"dd3984d1",
          5707 => x"88337c05",
          5708 => x"5f807f34",
          5709 => x"84d5ac08",
          5710 => x"528a51ff",
          5711 => x"b0b03f84",
          5712 => x"d188527b",
          5713 => x"51f48b3f",
          5714 => x"84b9c808",
          5715 => x"81ff0658",
          5716 => x"7789cf38",
          5717 => x"84d18833",
          5718 => x"5776802e",
          5719 => x"80d83883",
          5720 => x"f3b83370",
          5721 => x"101083f2",
          5722 => x"e0057008",
          5723 => x"575e5674",
          5724 => x"8ba03875",
          5725 => x"822b87fc",
          5726 => x"0683f2e0",
          5727 => x"05811870",
          5728 => x"53575b80",
          5729 => x"e7fb3f84",
          5730 => x"b9c8087b",
          5731 => x"0c83f3b8",
          5732 => x"33701010",
          5733 => x"83f2e005",
          5734 => x"70085741",
          5735 => x"41748bad",
          5736 => x"3883f3b4",
          5737 => x"08567580",
          5738 => x"2e8c3883",
          5739 => x"f3b03358",
          5740 => x"77802e8b",
          5741 => x"bc38800b",
          5742 => x"84d18c34",
          5743 => x"800b84d1",
          5744 => x"88347b84",
          5745 => x"b9c80cb4",
          5746 => x"3d0d0484",
          5747 => x"d18c3355",
          5748 => x"74802eb6",
          5749 => x"3884d5ac",
          5750 => x"08528851",
          5751 => x"ffaf8f3f",
          5752 => x"84d5ac08",
          5753 => x"52a051ff",
          5754 => x"af843f84",
          5755 => x"d5ac0852",
          5756 => x"8851ffae",
          5757 => x"f93f84d1",
          5758 => x"8c33ff05",
          5759 => x"567584d1",
          5760 => x"8c347581",
          5761 => x"ff065574",
          5762 => x"cc3883d1",
          5763 => x"f051ff9f",
          5764 => x"f73f800b",
          5765 => x"84d18c34",
          5766 => x"800b84d1",
          5767 => x"8834f5be",
          5768 => x"39837c34",
          5769 => x"800b811d",
          5770 => x"3484d18c",
          5771 => x"33557480",
          5772 => x"2eb63884",
          5773 => x"d5ac0852",
          5774 => x"8851ffae",
          5775 => x"b13f84d5",
          5776 => x"ac0852a0",
          5777 => x"51ffaea6",
          5778 => x"3f84d5ac",
          5779 => x"08528851",
          5780 => x"ffae9b3f",
          5781 => x"84d18c33",
          5782 => x"ff055d7c",
          5783 => x"84d18c34",
          5784 => x"7c81ff06",
          5785 => x"5574cc38",
          5786 => x"83d1f051",
          5787 => x"ff9f993f",
          5788 => x"800b84d1",
          5789 => x"8c34800b",
          5790 => x"84d18834",
          5791 => x"7b84b9c8",
          5792 => x"0cb43d0d",
          5793 => x"0484d18c",
          5794 => x"337081ff",
          5795 => x"065c567a",
          5796 => x"802ef4ca",
          5797 => x"3884d188",
          5798 => x"33ff0559",
          5799 => x"7884d188",
          5800 => x"34ff1658",
          5801 => x"7784d18c",
          5802 => x"3484d5ac",
          5803 => x"08528851",
          5804 => x"ffadbb3f",
          5805 => x"84d18c33",
          5806 => x"70982b70",
          5807 => x"982c84d1",
          5808 => x"88335a52",
          5809 => x"5b567676",
          5810 => x"2480ef38",
          5811 => x"84d5ac08",
          5812 => x"52a051ff",
          5813 => x"ad983f84",
          5814 => x"d18c3370",
          5815 => x"982b7098",
          5816 => x"2c84d188",
          5817 => x"335d5759",
          5818 => x"56747a24",
          5819 => x"f3f03884",
          5820 => x"d5ac0852",
          5821 => x"8851ffac",
          5822 => x"f53f7481",
          5823 => x"800a2981",
          5824 => x"800a0570",
          5825 => x"982c84d1",
          5826 => x"88335b51",
          5827 => x"55747924",
          5828 => x"f3cc3884",
          5829 => x"d5ac0852",
          5830 => x"8851ffac",
          5831 => x"d13f7481",
          5832 => x"800a2981",
          5833 => x"800a0570",
          5834 => x"982c84d1",
          5835 => x"88335b51",
          5836 => x"55787525",
          5837 => x"ffb938f3",
          5838 => x"a5397b16",
          5839 => x"57811733",
          5840 => x"773484d5",
          5841 => x"ac085276",
          5842 => x"3351ffac",
          5843 => x"a13f7581",
          5844 => x"800a2981",
          5845 => x"800a0570",
          5846 => x"982c84d1",
          5847 => x"88334357",
          5848 => x"5b756125",
          5849 => x"fee6387b",
          5850 => x"16578117",
          5851 => x"33773484",
          5852 => x"d5ac0852",
          5853 => x"763351ff",
          5854 => x"abf43f75",
          5855 => x"81800a29",
          5856 => x"81800a05",
          5857 => x"70982c84",
          5858 => x"d1883343",
          5859 => x"575b6076",
          5860 => x"24ffa738",
          5861 => x"feb63984",
          5862 => x"d18c3370",
          5863 => x"81ff0658",
          5864 => x"5876602e",
          5865 => x"f2b83884",
          5866 => x"d1883355",
          5867 => x"767527ae",
          5868 => x"3874982b",
          5869 => x"70982c57",
          5870 => x"41767624",
          5871 => x"a1387b16",
          5872 => x"5b7a3381",
          5873 => x"1c347581",
          5874 => x"800a2981",
          5875 => x"ff0a0570",
          5876 => x"982c84d1",
          5877 => x"8c335257",
          5878 => x"58757825",
          5879 => x"e1388118",
          5880 => x"557484d1",
          5881 => x"8c347781",
          5882 => x"ff067c05",
          5883 => x"5ab33d33",
          5884 => x"7a3484d1",
          5885 => x"88335776",
          5886 => x"60258b38",
          5887 => x"81175675",
          5888 => x"84d18834",
          5889 => x"755784d1",
          5890 => x"8c337081",
          5891 => x"800a2981",
          5892 => x"ff0a0570",
          5893 => x"982c7981",
          5894 => x"ff064458",
          5895 => x"5c586076",
          5896 => x"2481ef38",
          5897 => x"77982b70",
          5898 => x"982c7881",
          5899 => x"ff065c57",
          5900 => x"59757a25",
          5901 => x"f1a83884",
          5902 => x"d5ac0852",
          5903 => x"8851ffaa",
          5904 => x"ad3f7581",
          5905 => x"800a2981",
          5906 => x"800a0570",
          5907 => x"982c84d1",
          5908 => x"88335757",
          5909 => x"41757525",
          5910 => x"f1843884",
          5911 => x"d5ac0852",
          5912 => x"8851ffaa",
          5913 => x"893f7581",
          5914 => x"800a2981",
          5915 => x"800a0570",
          5916 => x"982c84d1",
          5917 => x"88335757",
          5918 => x"41747624",
          5919 => x"ffb938f0",
          5920 => x"dd3983f2",
          5921 => x"e0085675",
          5922 => x"802ef49d",
          5923 => x"387551ff",
          5924 => x"ad963f84",
          5925 => x"b9c80884",
          5926 => x"d1883484",
          5927 => x"b9c80881",
          5928 => x"ff068105",
          5929 => x"5375527b",
          5930 => x"51ffadbe",
          5931 => x"3f84d188",
          5932 => x"3384d18c",
          5933 => x"33565674",
          5934 => x"802ef4c8",
          5935 => x"3884d5ac",
          5936 => x"08528851",
          5937 => x"ffa9a73f",
          5938 => x"84d5ac08",
          5939 => x"52a051ff",
          5940 => x"a99c3f84",
          5941 => x"d5ac0852",
          5942 => x"8851ffa9",
          5943 => x"913f84d1",
          5944 => x"8c33ff05",
          5945 => x"5b7a84d1",
          5946 => x"8c347a81",
          5947 => x"ff0655c7",
          5948 => x"39a85180",
          5949 => x"e18b3f84",
          5950 => x"b9c80883",
          5951 => x"f3b40c84",
          5952 => x"b9c80885",
          5953 => x"a5387683",
          5954 => x"f3b03477",
          5955 => x"efca3880",
          5956 => x"c33984d5",
          5957 => x"ac08527b",
          5958 => x"16703352",
          5959 => x"58ffa8ce",
          5960 => x"3f758180",
          5961 => x"0a298180",
          5962 => x"0a057098",
          5963 => x"2c84d188",
          5964 => x"33525757",
          5965 => x"767624da",
          5966 => x"3884d18c",
          5967 => x"3370982b",
          5968 => x"70982c79",
          5969 => x"81ff065d",
          5970 => x"585a5875",
          5971 => x"7a25ef8e",
          5972 => x"38fde439",
          5973 => x"83f3b408",
          5974 => x"802eeefc",
          5975 => x"3883f2e0",
          5976 => x"57935676",
          5977 => x"085574bb",
          5978 => x"38ff1684",
          5979 => x"18585675",
          5980 => x"8025f038",
          5981 => x"800b83f3",
          5982 => x"b83483f3",
          5983 => x"b4085574",
          5984 => x"802eeed4",
          5985 => x"38745181",
          5986 => x"e7f63f83",
          5987 => x"f3b40851",
          5988 => x"80d9fe3f",
          5989 => x"800b83f3",
          5990 => x"b40c933d",
          5991 => x"b43d5f5f",
          5992 => x"eebc3974",
          5993 => x"5180d9e9",
          5994 => x"3f80770c",
          5995 => x"ff168418",
          5996 => x"58567580",
          5997 => x"25ffac38",
          5998 => x"ffba3975",
          5999 => x"51ffaae8",
          6000 => x"3f84b9c8",
          6001 => x"0884d188",
          6002 => x"3484b9c8",
          6003 => x"0881ff06",
          6004 => x"81055375",
          6005 => x"527b51ff",
          6006 => x"ab903f93",
          6007 => x"0b84d188",
          6008 => x"3384d18c",
          6009 => x"3357575d",
          6010 => x"74802ef2",
          6011 => x"973884d5",
          6012 => x"ac085288",
          6013 => x"51ffa6f6",
          6014 => x"3f84d5ac",
          6015 => x"0852a051",
          6016 => x"ffa6eb3f",
          6017 => x"84d5ac08",
          6018 => x"528851ff",
          6019 => x"a6e03f84",
          6020 => x"d18c33ff",
          6021 => x"055a7984",
          6022 => x"d18c3479",
          6023 => x"81ff0655",
          6024 => x"c739807c",
          6025 => x"34800b84",
          6026 => x"d18c3480",
          6027 => x"0b84d188",
          6028 => x"347b84b9",
          6029 => x"c80cb43d",
          6030 => x"0d047551",
          6031 => x"ffa9e93f",
          6032 => x"84b9c808",
          6033 => x"84d18834",
          6034 => x"84b9c808",
          6035 => x"81ff0681",
          6036 => x"05537552",
          6037 => x"7b51ffaa",
          6038 => x"913f811d",
          6039 => x"7081ff06",
          6040 => x"84d18833",
          6041 => x"84d18c33",
          6042 => x"58525e56",
          6043 => x"74802ef1",
          6044 => x"933884d5",
          6045 => x"ac085288",
          6046 => x"51ffa5f2",
          6047 => x"3f84d5ac",
          6048 => x"0852a051",
          6049 => x"ffa5e73f",
          6050 => x"84d5ac08",
          6051 => x"528851ff",
          6052 => x"a5dc3f84",
          6053 => x"d18c33ff",
          6054 => x"05577684",
          6055 => x"d18c3476",
          6056 => x"81ff0655",
          6057 => x"c7397551",
          6058 => x"ffa8fd3f",
          6059 => x"84b9c808",
          6060 => x"84d18834",
          6061 => x"84b9c808",
          6062 => x"81ff0681",
          6063 => x"05537552",
          6064 => x"7b51ffa9",
          6065 => x"a53fff1d",
          6066 => x"7081ff06",
          6067 => x"84d18833",
          6068 => x"84d18c33",
          6069 => x"58585e58",
          6070 => x"74802ef0",
          6071 => x"a73884d5",
          6072 => x"ac085288",
          6073 => x"51ffa586",
          6074 => x"3f84d5ac",
          6075 => x"0852a051",
          6076 => x"ffa4fb3f",
          6077 => x"84d5ac08",
          6078 => x"528851ff",
          6079 => x"a4f03f84",
          6080 => x"d18c33ff",
          6081 => x"05416084",
          6082 => x"d18c3460",
          6083 => x"81ff0655",
          6084 => x"c7397451",
          6085 => x"80d6fa3f",
          6086 => x"83f3b833",
          6087 => x"70822b87",
          6088 => x"fc0683f2",
          6089 => x"e0058119",
          6090 => x"7054525c",
          6091 => x"5680dcd1",
          6092 => x"3f84b9c8",
          6093 => x"087b0c83",
          6094 => x"f3b83370",
          6095 => x"101083f2",
          6096 => x"e0057008",
          6097 => x"57414174",
          6098 => x"802ef4d5",
          6099 => x"3875537b",
          6100 => x"527451ff",
          6101 => x"a8943f83",
          6102 => x"f3b83381",
          6103 => x"057081ff",
          6104 => x"065a5693",
          6105 => x"792782f2",
          6106 => x"387783f3",
          6107 => x"b834f4b1",
          6108 => x"39b43dfe",
          6109 => x"f8055476",
          6110 => x"537b5275",
          6111 => x"5181d8c0",
          6112 => x"3f83f3b4",
          6113 => x"08528a51",
          6114 => x"82ba883f",
          6115 => x"83f3b408",
          6116 => x"5181dff3",
          6117 => x"3f800b84",
          6118 => x"d18c3480",
          6119 => x"0b84d188",
          6120 => x"347b84b9",
          6121 => x"c80cb43d",
          6122 => x"0d049353",
          6123 => x"775284b9",
          6124 => x"c8085181",
          6125 => x"c9f83f84",
          6126 => x"b9c80882",
          6127 => x"a53884b9",
          6128 => x"c808963d",
          6129 => x"5c5d83f3",
          6130 => x"b4085380",
          6131 => x"f8527a51",
          6132 => x"82b7f23f",
          6133 => x"84b9c808",
          6134 => x"5a84b9c8",
          6135 => x"087b2e09",
          6136 => x"8106e9ee",
          6137 => x"3884b9c8",
          6138 => x"0851ffa6",
          6139 => x"bb3f84b9",
          6140 => x"c8085680",
          6141 => x"0b84b9c8",
          6142 => x"082580e3",
          6143 => x"3884b9c8",
          6144 => x"08ff0570",
          6145 => x"1b585680",
          6146 => x"77347581",
          6147 => x"ff0683f3",
          6148 => x"b8337010",
          6149 => x"1083f2e0",
          6150 => x"05700858",
          6151 => x"40585974",
          6152 => x"80f23876",
          6153 => x"822b87fc",
          6154 => x"0683f2e0",
          6155 => x"05811a70",
          6156 => x"53585580",
          6157 => x"dacb3f84",
          6158 => x"b9c80875",
          6159 => x"0c83f3b8",
          6160 => x"33701010",
          6161 => x"83f2e005",
          6162 => x"70085740",
          6163 => x"4174a038",
          6164 => x"811d7081",
          6165 => x"ff065e57",
          6166 => x"937d2783",
          6167 => x"38805d75",
          6168 => x"ff2e0981",
          6169 => x"06fedf38",
          6170 => x"77e8ed38",
          6171 => x"f9e63976",
          6172 => x"53795274",
          6173 => x"51ffa5f2",
          6174 => x"3f83f3b8",
          6175 => x"33810570",
          6176 => x"81ff065b",
          6177 => x"57937a27",
          6178 => x"80c83880",
          6179 => x"0b83f3b8",
          6180 => x"34ffbd39",
          6181 => x"745180d3",
          6182 => x"f83f83f3",
          6183 => x"b8337082",
          6184 => x"2b87fc06",
          6185 => x"83f2e005",
          6186 => x"811b7054",
          6187 => x"52565780",
          6188 => x"d9cf3f84",
          6189 => x"b9c80875",
          6190 => x"0c83f3b8",
          6191 => x"33701010",
          6192 => x"83f2e005",
          6193 => x"70085740",
          6194 => x"4174802e",
          6195 => x"ff8238ff",
          6196 => x"9e397683",
          6197 => x"f3b834fe",
          6198 => x"f7397583",
          6199 => x"f3b834f1",
          6200 => x"c03983e1",
          6201 => x"b051ff9f",
          6202 => x"8a3f77e7",
          6203 => x"eb38f8e4",
          6204 => x"39f23d0d",
          6205 => x"0280c305",
          6206 => x"33028405",
          6207 => x"80c70533",
          6208 => x"5b537283",
          6209 => x"26818d38",
          6210 => x"72812e81",
          6211 => x"8b388173",
          6212 => x"25839e38",
          6213 => x"72822e82",
          6214 => x"a83886a7",
          6215 => x"a0805986",
          6216 => x"a7b08070",
          6217 => x"5e578056",
          6218 => x"9fa05879",
          6219 => x"762e9038",
          6220 => x"7583f8f8",
          6221 => x"347583f8",
          6222 => x"f9347583",
          6223 => x"f8f62383",
          6224 => x"f8f43370",
          6225 => x"982b7190",
          6226 => x"2b077188",
          6227 => x"2b077107",
          6228 => x"7a7f5656",
          6229 => x"565b7877",
          6230 => x"27943880",
          6231 => x"74708405",
          6232 => x"560c7473",
          6233 => x"70840555",
          6234 => x"0c767426",
          6235 => x"ee387578",
          6236 => x"27a23883",
          6237 => x"f8f43384",
          6238 => x"989a1779",
          6239 => x"78315555",
          6240 => x"55a00be0",
          6241 => x"e0153474",
          6242 => x"74708105",
          6243 => x"5634ff13",
          6244 => x"5372ee38",
          6245 => x"903d0d04",
          6246 => x"86a7a080",
          6247 => x"0b83f8f8",
          6248 => x"33701010",
          6249 => x"1183f8f9",
          6250 => x"33719029",
          6251 => x"1174055b",
          6252 => x"41584059",
          6253 => x"86a7b080",
          6254 => x"0b84b7bc",
          6255 => x"337081ff",
          6256 => x"0684b7bb",
          6257 => x"337081ff",
          6258 => x"0683f8f6",
          6259 => x"227083ff",
          6260 => x"ff067075",
          6261 => x"295d595d",
          6262 => x"585e575b",
          6263 => x"5d737326",
          6264 => x"87387274",
          6265 => x"31752956",
          6266 => x"7981ff06",
          6267 => x"7e81ff06",
          6268 => x"7c81ff06",
          6269 => x"7a83ffff",
          6270 => x"066281ff",
          6271 => x"06707529",
          6272 => x"145d4257",
          6273 => x"575b5c74",
          6274 => x"74268f38",
          6275 => x"83f8f833",
          6276 => x"74763105",
          6277 => x"707d291b",
          6278 => x"595f7683",
          6279 => x"065c7b80",
          6280 => x"2efe9c38",
          6281 => x"787d5553",
          6282 => x"727726fe",
          6283 => x"c1388073",
          6284 => x"70810555",
          6285 => x"3483f8f4",
          6286 => x"33747081",
          6287 => x"055634e8",
          6288 => x"3986a7a0",
          6289 => x"805986a7",
          6290 => x"b0807084",
          6291 => x"b7bc3370",
          6292 => x"81ff0684",
          6293 => x"b7bb3370",
          6294 => x"81ff0683",
          6295 => x"f8f62270",
          6296 => x"74295d5b",
          6297 => x"5d575e56",
          6298 => x"5e577478",
          6299 => x"2781df38",
          6300 => x"7381ff06",
          6301 => x"7381ff06",
          6302 => x"71712918",
          6303 => x"5a545479",
          6304 => x"802efdbb",
          6305 => x"38800b83",
          6306 => x"f8f83480",
          6307 => x"0b83f8f9",
          6308 => x"3483f8f4",
          6309 => x"3370982b",
          6310 => x"71902b07",
          6311 => x"71882b07",
          6312 => x"71077a7f",
          6313 => x"5656565b",
          6314 => x"767926fd",
          6315 => x"ae38fdbe",
          6316 => x"3972fce6",
          6317 => x"3883f8f8",
          6318 => x"337081ff",
          6319 => x"06701010",
          6320 => x"1183f8f9",
          6321 => x"33719029",
          6322 => x"1186a7a0",
          6323 => x"80115e57",
          6324 => x"5b56565f",
          6325 => x"86a7b080",
          6326 => x"701484b7",
          6327 => x"bc337081",
          6328 => x"ff0684b7",
          6329 => x"bb337081",
          6330 => x"ff0683f8",
          6331 => x"f6227083",
          6332 => x"ffff067c",
          6333 => x"75296005",
          6334 => x"5e5a415f",
          6335 => x"585f405e",
          6336 => x"57797326",
          6337 => x"8b38727a",
          6338 => x"3115707d",
          6339 => x"29195753",
          6340 => x"7d81ff06",
          6341 => x"7481ff06",
          6342 => x"7171297d",
          6343 => x"83ffff06",
          6344 => x"6281ff06",
          6345 => x"70752958",
          6346 => x"5f5b5c5d",
          6347 => x"557b7826",
          6348 => x"85387775",
          6349 => x"29537973",
          6350 => x"31167983",
          6351 => x"065b5879",
          6352 => x"fde23876",
          6353 => x"83065c7b",
          6354 => x"fdda38fb",
          6355 => x"f2397478",
          6356 => x"317b2956",
          6357 => x"fe9a39fb",
          6358 => x"3d0d86ee",
          6359 => x"808c53ff",
          6360 => x"8a733487",
          6361 => x"73348573",
          6362 => x"34817334",
          6363 => x"86ee809c",
          6364 => x"5580f475",
          6365 => x"34ffb075",
          6366 => x"3486ee80",
          6367 => x"98568076",
          6368 => x"34807634",
          6369 => x"86ee8094",
          6370 => x"548a7434",
          6371 => x"807434ff",
          6372 => x"80753481",
          6373 => x"528351fa",
          6374 => x"d83f86a0",
          6375 => x"87e07008",
          6376 => x"545481f8",
          6377 => x"5686a081",
          6378 => x"f8737706",
          6379 => x"84075455",
          6380 => x"72753473",
          6381 => x"087080ff",
          6382 => x"0680c007",
          6383 => x"51537275",
          6384 => x"3486a087",
          6385 => x"cc087077",
          6386 => x"06810751",
          6387 => x"537286a0",
          6388 => x"81f33473",
          6389 => x"0881f706",
          6390 => x"88075372",
          6391 => x"753480d0",
          6392 => x"0b84b7bc",
          6393 => x"34800b84",
          6394 => x"b9c80c87",
          6395 => x"3d0d0484",
          6396 => x"b7bc3384",
          6397 => x"b9c80c04",
          6398 => x"f73d0d02",
          6399 => x"af053302",
          6400 => x"8405b305",
          6401 => x"3384b7bb",
          6402 => x"335b5956",
          6403 => x"81537579",
          6404 => x"2682da38",
          6405 => x"84b7bc33",
          6406 => x"83f8f933",
          6407 => x"83f8f833",
          6408 => x"72712912",
          6409 => x"86a7a080",
          6410 => x"1183f8f6",
          6411 => x"225f5157",
          6412 => x"59717c29",
          6413 => x"057083ff",
          6414 => x"ff0683f7",
          6415 => x"ce335357",
          6416 => x"58537281",
          6417 => x"2e83c438",
          6418 => x"83f8f622",
          6419 => x"76055574",
          6420 => x"83f8f623",
          6421 => x"83f8f833",
          6422 => x"76057081",
          6423 => x"ff067a81",
          6424 => x"ff06555b",
          6425 => x"55727a26",
          6426 => x"828c38ff",
          6427 => x"19537283",
          6428 => x"f8f83483",
          6429 => x"f8f62270",
          6430 => x"83ffff06",
          6431 => x"84b7ba33",
          6432 => x"5c555779",
          6433 => x"74268289",
          6434 => x"3884b7bc",
          6435 => x"33767129",
          6436 => x"54588054",
          6437 => x"729f9f26",
          6438 => x"ac388498",
          6439 => x"9a701454",
          6440 => x"55e0e013",
          6441 => x"33e0e016",
          6442 => x"34727081",
          6443 => x"05543375",
          6444 => x"70810557",
          6445 => x"34811454",
          6446 => x"84b7b973",
          6447 => x"27e33873",
          6448 => x"9f9f26a1",
          6449 => x"3883f8f4",
          6450 => x"3384989a",
          6451 => x"155455a0",
          6452 => x"0be0e014",
          6453 => x"34747370",
          6454 => x"81055534",
          6455 => x"8114549f",
          6456 => x"9f7427eb",
          6457 => x"3884b7ba",
          6458 => x"33ff0556",
          6459 => x"7583f8f6",
          6460 => x"23755778",
          6461 => x"81ff0677",
          6462 => x"83ffff06",
          6463 => x"54547373",
          6464 => x"2681fd38",
          6465 => x"72743181",
          6466 => x"0584b7bc",
          6467 => x"33717129",
          6468 => x"58555775",
          6469 => x"5586a7a0",
          6470 => x"805886a7",
          6471 => x"b0807981",
          6472 => x"ff067581",
          6473 => x"ff067171",
          6474 => x"29195c5c",
          6475 => x"54577579",
          6476 => x"27b93884",
          6477 => x"989a1654",
          6478 => x"e0e01433",
          6479 => x"5384b7c4",
          6480 => x"13337870",
          6481 => x"81055a34",
          6482 => x"73708105",
          6483 => x"55337770",
          6484 => x"81055934",
          6485 => x"811584b7",
          6486 => x"bc3384b7",
          6487 => x"bb337171",
          6488 => x"2919565c",
          6489 => x"5a557275",
          6490 => x"26ce3880",
          6491 => x"537284b9",
          6492 => x"c80c8b3d",
          6493 => x"0d047483",
          6494 => x"f8f83483",
          6495 => x"f8f62270",
          6496 => x"83ffff06",
          6497 => x"84b7ba33",
          6498 => x"5c555773",
          6499 => x"7a27fdf9",
          6500 => x"3877802e",
          6501 => x"fedd3878",
          6502 => x"81ff06ff",
          6503 => x"0583f8f8",
          6504 => x"33565372",
          6505 => x"752e0981",
          6506 => x"06fec838",
          6507 => x"73763181",
          6508 => x"0584b7bc",
          6509 => x"33717129",
          6510 => x"78722911",
          6511 => x"56525954",
          6512 => x"737327fe",
          6513 => x"ae3883f8",
          6514 => x"f4338498",
          6515 => x"9a157476",
          6516 => x"31555656",
          6517 => x"a00be0e0",
          6518 => x"16347575",
          6519 => x"70810557",
          6520 => x"34ff1353",
          6521 => x"72802efe",
          6522 => x"8a38a00b",
          6523 => x"e0e01634",
          6524 => x"75757081",
          6525 => x"055734ff",
          6526 => x"135372d8",
          6527 => x"38fdf439",
          6528 => x"800b84b7",
          6529 => x"bc335556",
          6530 => x"fe893983",
          6531 => x"f8fa1533",
          6532 => x"5984b7c4",
          6533 => x"19337434",
          6534 => x"84b7bb33",
          6535 => x"59fca939",
          6536 => x"fc3d0d76",
          6537 => x"0284059f",
          6538 => x"05335351",
          6539 => x"7086269b",
          6540 => x"38701010",
          6541 => x"83c3ec05",
          6542 => x"51700804",
          6543 => x"84b7bc33",
          6544 => x"51717127",
          6545 => x"86387183",
          6546 => x"f8f93480",
          6547 => x"0b84b9c8",
          6548 => x"0c863d0d",
          6549 => x"04800b83",
          6550 => x"f8f93483",
          6551 => x"f8f83370",
          6552 => x"81ff0654",
          6553 => x"5272802e",
          6554 => x"e238ff12",
          6555 => x"517083f8",
          6556 => x"f834800b",
          6557 => x"84b9c80c",
          6558 => x"863d0d04",
          6559 => x"83f8f833",
          6560 => x"70733170",
          6561 => x"09709f2c",
          6562 => x"72065455",
          6563 => x"53547083",
          6564 => x"f8f834de",
          6565 => x"3983f8f8",
          6566 => x"33720584",
          6567 => x"b7bb33ff",
          6568 => x"11555651",
          6569 => x"70752583",
          6570 => x"38705372",
          6571 => x"83f8f834",
          6572 => x"800b84b9",
          6573 => x"c80c863d",
          6574 => x"0d0483f8",
          6575 => x"f9337073",
          6576 => x"31700970",
          6577 => x"9f2c7206",
          6578 => x"54565355",
          6579 => x"7083f8f9",
          6580 => x"34800b84",
          6581 => x"b9c80c86",
          6582 => x"3d0d0483",
          6583 => x"f8f93372",
          6584 => x"0584b7bc",
          6585 => x"33ff1155",
          6586 => x"55517074",
          6587 => x"25833870",
          6588 => x"537283f8",
          6589 => x"f934800b",
          6590 => x"84b9c80c",
          6591 => x"863d0d04",
          6592 => x"800b83f8",
          6593 => x"f93483f8",
          6594 => x"f83384b7",
          6595 => x"bb33ff05",
          6596 => x"56527175",
          6597 => x"25feb438",
          6598 => x"81125170",
          6599 => x"83f8f834",
          6600 => x"fed039ff",
          6601 => x"3d0d028f",
          6602 => x"05335170",
          6603 => x"b126b338",
          6604 => x"70101083",
          6605 => x"c4880551",
          6606 => x"70080483",
          6607 => x"f8f43370",
          6608 => x"80f00671",
          6609 => x"842b80f0",
          6610 => x"06707284",
          6611 => x"2a075152",
          6612 => x"53517180",
          6613 => x"f02e0981",
          6614 => x"069c3880",
          6615 => x"f20b83f8",
          6616 => x"f434800b",
          6617 => x"84b9c80c",
          6618 => x"833d0d04",
          6619 => x"83f8f433",
          6620 => x"819f0690",
          6621 => x"07517083",
          6622 => x"f8f43480",
          6623 => x"0b84b9c8",
          6624 => x"0c833d0d",
          6625 => x"0483f8f4",
          6626 => x"3380f007",
          6627 => x"517083f8",
          6628 => x"f434e839",
          6629 => x"83f8f433",
          6630 => x"81fe0686",
          6631 => x"07517083",
          6632 => x"f8f434d7",
          6633 => x"3980f10b",
          6634 => x"83f8f434",
          6635 => x"800b84b9",
          6636 => x"c80c833d",
          6637 => x"0d0483f8",
          6638 => x"f43381fc",
          6639 => x"06840751",
          6640 => x"7083f8f4",
          6641 => x"34ffb439",
          6642 => x"83f8f433",
          6643 => x"87075170",
          6644 => x"83f8f434",
          6645 => x"ffa53983",
          6646 => x"f8f43381",
          6647 => x"fd068507",
          6648 => x"517083f8",
          6649 => x"f434ff93",
          6650 => x"3983f8f4",
          6651 => x"3381fb06",
          6652 => x"83075170",
          6653 => x"83f8f434",
          6654 => x"ff813983",
          6655 => x"f8f43381",
          6656 => x"f9068107",
          6657 => x"517083f8",
          6658 => x"f434feef",
          6659 => x"3983f8f4",
          6660 => x"3381f806",
          6661 => x"517083f8",
          6662 => x"f434fedf",
          6663 => x"3983f8f4",
          6664 => x"3381df06",
          6665 => x"80d00751",
          6666 => x"7083f8f4",
          6667 => x"34fecc39",
          6668 => x"83f8f433",
          6669 => x"81bf06b0",
          6670 => x"07517083",
          6671 => x"f8f434fe",
          6672 => x"ba3983f8",
          6673 => x"f43381ef",
          6674 => x"0680e007",
          6675 => x"517083f8",
          6676 => x"f434fea7",
          6677 => x"3983f8f4",
          6678 => x"3381cf06",
          6679 => x"80c00751",
          6680 => x"7083f8f4",
          6681 => x"34fe9439",
          6682 => x"83f8f433",
          6683 => x"81af06a0",
          6684 => x"07517083",
          6685 => x"f8f434fe",
          6686 => x"823983f8",
          6687 => x"f433818f",
          6688 => x"06517083",
          6689 => x"f8f434fd",
          6690 => x"f23983f8",
          6691 => x"f43381fa",
          6692 => x"06820751",
          6693 => x"7083f8f4",
          6694 => x"34fde039",
          6695 => x"f33d0d02",
          6696 => x"bf053302",
          6697 => x"840580c3",
          6698 => x"053383f8",
          6699 => x"f83383f8",
          6700 => x"f73383f8",
          6701 => x"f93384b7",
          6702 => x"be334341",
          6703 => x"5f5d5b59",
          6704 => x"78822e82",
          6705 => x"a1387882",
          6706 => x"24a53878",
          6707 => x"812e8182",
          6708 => x"387d84b7",
          6709 => x"be34800b",
          6710 => x"84b7c034",
          6711 => x"7a83f8f8",
          6712 => x"347b83f8",
          6713 => x"f6237c83",
          6714 => x"f8f9348f",
          6715 => x"3d0d0478",
          6716 => x"832e0981",
          6717 => x"06db3880",
          6718 => x"0b84b7be",
          6719 => x"34810b84",
          6720 => x"b7c03482",
          6721 => x"0b83f8f8",
          6722 => x"34a80b83",
          6723 => x"f8f93482",
          6724 => x"0b83f8f6",
          6725 => x"23795884",
          6726 => x"b7bc3357",
          6727 => x"84b7bb33",
          6728 => x"5684b7ba",
          6729 => x"33557b54",
          6730 => x"7c537a52",
          6731 => x"83e3bc51",
          6732 => x"ff81d53f",
          6733 => x"7d84b7be",
          6734 => x"34800b84",
          6735 => x"b7c0347a",
          6736 => x"83f8f834",
          6737 => x"7b83f8f6",
          6738 => x"237c83f8",
          6739 => x"f9348f3d",
          6740 => x"0d04800b",
          6741 => x"84b7be34",
          6742 => x"810b84b7",
          6743 => x"c034800b",
          6744 => x"83f8f834",
          6745 => x"a80b83f8",
          6746 => x"f934800b",
          6747 => x"83f8f623",
          6748 => x"84b8cb33",
          6749 => x"5884b8ca",
          6750 => x"335784b8",
          6751 => x"c9335679",
          6752 => x"557b547c",
          6753 => x"537a5283",
          6754 => x"e3d851ff",
          6755 => x"80fa3f80",
          6756 => x"0b84b8c9",
          6757 => x"335a5a79",
          6758 => x"7927a538",
          6759 => x"791084b9",
          6760 => x"9c057022",
          6761 => x"535983e3",
          6762 => x"f051ff80",
          6763 => x"db3f811a",
          6764 => x"7081ff06",
          6765 => x"84b8c933",
          6766 => x"525b5978",
          6767 => x"7a26dd38",
          6768 => x"83d2a451",
          6769 => x"ff80c13f",
          6770 => x"7d84b7be",
          6771 => x"34800b84",
          6772 => x"b7c0347a",
          6773 => x"83f8f834",
          6774 => x"7b83f8f6",
          6775 => x"237c83f8",
          6776 => x"f9348f3d",
          6777 => x"0d04800b",
          6778 => x"84b7be34",
          6779 => x"810b84b7",
          6780 => x"c034810b",
          6781 => x"83f8f834",
          6782 => x"a80b83f8",
          6783 => x"f934810b",
          6784 => x"83f8f623",
          6785 => x"83f7ac51",
          6786 => x"ff929d3f",
          6787 => x"84b9c808",
          6788 => x"5283e3f4",
          6789 => x"51fefff0",
          6790 => x"3f805983",
          6791 => x"f7ac51ff",
          6792 => x"92863f78",
          6793 => x"84b9c808",
          6794 => x"27fda638",
          6795 => x"83f7ac19",
          6796 => x"335283e3",
          6797 => x"fc51feff",
          6798 => x"cf3f8119",
          6799 => x"7081ff06",
          6800 => x"5a5ad839",
          6801 => x"f93d0d7a",
          6802 => x"028405a7",
          6803 => x"053384b7",
          6804 => x"bc3383f8",
          6805 => x"f93383f8",
          6806 => x"f8337271",
          6807 => x"291286a7",
          6808 => x"a0801183",
          6809 => x"f8f62253",
          6810 => x"51595c71",
          6811 => x"7c290570",
          6812 => x"83ffff06",
          6813 => x"83f7ce33",
          6814 => x"52595155",
          6815 => x"57577281",
          6816 => x"2e81e938",
          6817 => x"75892e81",
          6818 => x"f9387589",
          6819 => x"2481b938",
          6820 => x"75812e83",
          6821 => x"85387588",
          6822 => x"2e82d538",
          6823 => x"84b7bc33",
          6824 => x"83f8f833",
          6825 => x"83f8f933",
          6826 => x"72722905",
          6827 => x"55565484",
          6828 => x"b7c41633",
          6829 => x"86a7a080",
          6830 => x"143484b7",
          6831 => x"bc3383f8",
          6832 => x"f93383f8",
          6833 => x"f6227271",
          6834 => x"29125a5a",
          6835 => x"56537583",
          6836 => x"f8fa1834",
          6837 => x"83f8f833",
          6838 => x"73712916",
          6839 => x"585483f8",
          6840 => x"f43386a7",
          6841 => x"b0801834",
          6842 => x"84b7bc33",
          6843 => x"7081ff06",
          6844 => x"83f8f622",
          6845 => x"83f8f933",
          6846 => x"72722911",
          6847 => x"575b5755",
          6848 => x"5783f8f4",
          6849 => x"3384989a",
          6850 => x"14348118",
          6851 => x"7081ff06",
          6852 => x"59557378",
          6853 => x"26819938",
          6854 => x"84b7bd33",
          6855 => x"587781ea",
          6856 => x"38ff1753",
          6857 => x"7283f8f9",
          6858 => x"3484b7bf",
          6859 => x"33537280",
          6860 => x"2e8c3884",
          6861 => x"b7c03357",
          6862 => x"76802e80",
          6863 => x"fb38800b",
          6864 => x"84b9c80c",
          6865 => x"893d0d04",
          6866 => x"758d2e97",
          6867 => x"38758d24",
          6868 => x"80f73875",
          6869 => x"8a2e0981",
          6870 => x"06fec138",
          6871 => x"81528151",
          6872 => x"f1963f80",
          6873 => x"0b83f8f9",
          6874 => x"34ffbe39",
          6875 => x"83f8fa15",
          6876 => x"335384b7",
          6877 => x"c4133374",
          6878 => x"3475892e",
          6879 => x"098106fe",
          6880 => x"89388053",
          6881 => x"7652a051",
          6882 => x"fdba3f81",
          6883 => x"137081ff",
          6884 => x"06545472",
          6885 => x"8326ff91",
          6886 => x"387652a0",
          6887 => x"51fda53f",
          6888 => x"81137081",
          6889 => x"ff065454",
          6890 => x"837327d8",
          6891 => x"38fefa39",
          6892 => x"7483f8f9",
          6893 => x"34fef239",
          6894 => x"75528351",
          6895 => x"f9de3f80",
          6896 => x"0b84b9c8",
          6897 => x"0c893d0d",
          6898 => x"047580ff",
          6899 => x"2e098106",
          6900 => x"fdca3883",
          6901 => x"f8f93370",
          6902 => x"81ff0655",
          6903 => x"ff055373",
          6904 => x"83387353",
          6905 => x"7283f8f9",
          6906 => x"347652a0",
          6907 => x"51fcd53f",
          6908 => x"83f8f933",
          6909 => x"7081ff06",
          6910 => x"55ff0553",
          6911 => x"73fea538",
          6912 => x"73537283",
          6913 => x"f8f934fe",
          6914 => x"a039800b",
          6915 => x"83f8f934",
          6916 => x"81528151",
          6917 => x"efe23ffe",
          6918 => x"90398052",
          6919 => x"7551efd8",
          6920 => x"3ffe8639",
          6921 => x"e63d0d02",
          6922 => x"80f30533",
          6923 => x"84b8c408",
          6924 => x"57597581",
          6925 => x"2e81b838",
          6926 => x"75822e83",
          6927 => x"8238788a",
          6928 => x"2e84b538",
          6929 => x"788a2482",
          6930 => x"d1387888",
          6931 => x"2e84b938",
          6932 => x"78892e88",
          6933 => x"8f3884b7",
          6934 => x"bc3383f8",
          6935 => x"f83383f8",
          6936 => x"f9337272",
          6937 => x"2905585e",
          6938 => x"5c84b7c4",
          6939 => x"193386a7",
          6940 => x"a0801734",
          6941 => x"84b7bc33",
          6942 => x"83f8f933",
          6943 => x"83f8f622",
          6944 => x"72712912",
          6945 => x"5a5a4240",
          6946 => x"7883f8fa",
          6947 => x"183483f8",
          6948 => x"f8336071",
          6949 => x"29620540",
          6950 => x"5a83f8f4",
          6951 => x"337f86a7",
          6952 => x"b0800534",
          6953 => x"84b7bc33",
          6954 => x"7081ff06",
          6955 => x"83f8f622",
          6956 => x"83f8f933",
          6957 => x"72722911",
          6958 => x"42405d58",
          6959 => x"5983f8f4",
          6960 => x"3384989a",
          6961 => x"1f34811d",
          6962 => x"7081ff06",
          6963 => x"42587661",
          6964 => x"2681b838",
          6965 => x"84b7bd33",
          6966 => x"5a7986f1",
          6967 => x"38ff1956",
          6968 => x"7583f8f9",
          6969 => x"34800b84",
          6970 => x"b9c80c9c",
          6971 => x"3d0d0478",
          6972 => x"b72e848a",
          6973 => x"38b77925",
          6974 => x"81fd3878",
          6975 => x"b82e9bb3",
          6976 => x"387880db",
          6977 => x"2e89cc38",
          6978 => x"800b84b8",
          6979 => x"c40c84b7",
          6980 => x"bc3383f8",
          6981 => x"f83383f8",
          6982 => x"f9337272",
          6983 => x"29055e40",
          6984 => x"4084b7c4",
          6985 => x"193386a7",
          6986 => x"a0801d34",
          6987 => x"84b7bc33",
          6988 => x"83f8f933",
          6989 => x"83f8f622",
          6990 => x"72712912",
          6991 => x"415f5956",
          6992 => x"7883f8fa",
          6993 => x"1f3483f8",
          6994 => x"f8337671",
          6995 => x"29195b57",
          6996 => x"83f8f433",
          6997 => x"86a7b080",
          6998 => x"1b3484b7",
          6999 => x"bc337081",
          7000 => x"ff0683f8",
          7001 => x"f62283f8",
          7002 => x"f9337272",
          7003 => x"29114442",
          7004 => x"43585983",
          7005 => x"f8f43360",
          7006 => x"84989a05",
          7007 => x"34811f58",
          7008 => x"7781ff06",
          7009 => x"41607727",
          7010 => x"feca3877",
          7011 => x"83f8f934",
          7012 => x"800b84b9",
          7013 => x"c80c9c3d",
          7014 => x"0d04789b",
          7015 => x"2e82b738",
          7016 => x"789b2483",
          7017 => x"8138788d",
          7018 => x"2e098106",
          7019 => x"fda83880",
          7020 => x"0b83f8f9",
          7021 => x"34800b84",
          7022 => x"b9c80c9c",
          7023 => x"3d0d0478",
          7024 => x"9b2e82aa",
          7025 => x"38d01956",
          7026 => x"75892684",
          7027 => x"d03884b8",
          7028 => x"c8338111",
          7029 => x"59577784",
          7030 => x"b8c83478",
          7031 => x"84b8cc18",
          7032 => x"347781ff",
          7033 => x"0659800b",
          7034 => x"84b8cc1a",
          7035 => x"34800b84",
          7036 => x"b9c80c9c",
          7037 => x"3d0d0478",
          7038 => x"9b2efde9",
          7039 => x"38800b84",
          7040 => x"b8c40c84",
          7041 => x"b7bc3383",
          7042 => x"f8f83383",
          7043 => x"f8f93372",
          7044 => x"7229055e",
          7045 => x"404084b7",
          7046 => x"c4193386",
          7047 => x"a7a0801d",
          7048 => x"3484b7bc",
          7049 => x"3383f8f9",
          7050 => x"3383f8f6",
          7051 => x"22727129",
          7052 => x"12415f59",
          7053 => x"567883f8",
          7054 => x"fa1f3483",
          7055 => x"f8f83376",
          7056 => x"7129195b",
          7057 => x"5783f8f4",
          7058 => x"3386a7b0",
          7059 => x"801b3484",
          7060 => x"b7bc3370",
          7061 => x"81ff0683",
          7062 => x"f8f62283",
          7063 => x"f8f93372",
          7064 => x"72291144",
          7065 => x"42435859",
          7066 => x"83f8f433",
          7067 => x"6084989a",
          7068 => x"0534811f",
          7069 => x"58fe8939",
          7070 => x"81528151",
          7071 => x"eafa3f80",
          7072 => x"0b83f8f9",
          7073 => x"34feae39",
          7074 => x"84b7bc33",
          7075 => x"83f8f933",
          7076 => x"7081ff06",
          7077 => x"83f8f833",
          7078 => x"73712912",
          7079 => x"86a7a080",
          7080 => x"0583f8f6",
          7081 => x"2240515d",
          7082 => x"727e2905",
          7083 => x"7083ffff",
          7084 => x"0683f7ce",
          7085 => x"335a5159",
          7086 => x"5a5c7581",
          7087 => x"2e86a438",
          7088 => x"7881ff06",
          7089 => x"ff1a5757",
          7090 => x"76fc9538",
          7091 => x"76567583",
          7092 => x"f8f934fc",
          7093 => x"9039800b",
          7094 => x"84b8c834",
          7095 => x"800b84b8",
          7096 => x"c934800b",
          7097 => x"84b8ca34",
          7098 => x"800b84b8",
          7099 => x"cb34810b",
          7100 => x"84b8c40c",
          7101 => x"800b84b9",
          7102 => x"c80c9c3d",
          7103 => x"0d0483f8",
          7104 => x"f83384b9",
          7105 => x"b03483f8",
          7106 => x"f93384b9",
          7107 => x"b13483f8",
          7108 => x"f73384b9",
          7109 => x"b234800b",
          7110 => x"84b8c40c",
          7111 => x"800b84b9",
          7112 => x"c80c9c3d",
          7113 => x"0d047880",
          7114 => x"ff2e0981",
          7115 => x"06faa738",
          7116 => x"83f8f833",
          7117 => x"84b7bc33",
          7118 => x"7081ff06",
          7119 => x"83f8f933",
          7120 => x"7081ff06",
          7121 => x"72752911",
          7122 => x"86a7a080",
          7123 => x"0583f8f6",
          7124 => x"225c4072",
          7125 => x"7b290570",
          7126 => x"83ffff06",
          7127 => x"83f7ce33",
          7128 => x"445c435c",
          7129 => x"425b5c7d",
          7130 => x"812e85fe",
          7131 => x"387881ff",
          7132 => x"06ff1a58",
          7133 => x"56758338",
          7134 => x"75577683",
          7135 => x"f8f9347b",
          7136 => x"81ff067a",
          7137 => x"81ff0678",
          7138 => x"81ff0672",
          7139 => x"7229055f",
          7140 => x"405b84b7",
          7141 => x"e43386a7",
          7142 => x"a0801e34",
          7143 => x"84b7bc33",
          7144 => x"83f8f933",
          7145 => x"83f8f622",
          7146 => x"72712912",
          7147 => x"5a5e4240",
          7148 => x"a00b83f8",
          7149 => x"fa183483",
          7150 => x"f8f83360",
          7151 => x"71296205",
          7152 => x"5a5683f8",
          7153 => x"f43386a7",
          7154 => x"b0801a34",
          7155 => x"84b7bc33",
          7156 => x"7081ff06",
          7157 => x"83f8f622",
          7158 => x"83f8f933",
          7159 => x"72722911",
          7160 => x"435d5a5e",
          7161 => x"5983f8f4",
          7162 => x"337f8498",
          7163 => x"9a053481",
          7164 => x"1a7081ff",
          7165 => x"065c587c",
          7166 => x"7b2695ea",
          7167 => x"3884b7bd",
          7168 => x"335a7996",
          7169 => x"d038ff19",
          7170 => x"587783f8",
          7171 => x"f93483f8",
          7172 => x"f9337081",
          7173 => x"ff0658ff",
          7174 => x"0556fdac",
          7175 => x"3978bb2e",
          7176 => x"95d83878",
          7177 => x"bd2e83d7",
          7178 => x"3878bf2e",
          7179 => x"95a83884",
          7180 => x"b8c8335f",
          7181 => x"7e83f938",
          7182 => x"ffbf1956",
          7183 => x"75b42684",
          7184 => x"c8387510",
          7185 => x"1083c5d0",
          7186 => x"05587708",
          7187 => x"04800b83",
          7188 => x"f8f93480",
          7189 => x"528151e7",
          7190 => x"9f3f800b",
          7191 => x"84b9c80c",
          7192 => x"9c3d0d04",
          7193 => x"83f8f833",
          7194 => x"84b7bc33",
          7195 => x"7081ff06",
          7196 => x"83f8f933",
          7197 => x"7081ff06",
          7198 => x"72752911",
          7199 => x"86a7a080",
          7200 => x"0583f8f6",
          7201 => x"225c4172",
          7202 => x"7b290570",
          7203 => x"83ffff06",
          7204 => x"83f7ce33",
          7205 => x"4653455c",
          7206 => x"595b5b7f",
          7207 => x"812e82ef",
          7208 => x"38805c7a",
          7209 => x"81ff067a",
          7210 => x"81ff067a",
          7211 => x"81ff0672",
          7212 => x"7229055c",
          7213 => x"584084b7",
          7214 => x"e43386a7",
          7215 => x"a0801b34",
          7216 => x"84b7bc33",
          7217 => x"83f8f933",
          7218 => x"83f8f622",
          7219 => x"72712912",
          7220 => x"5e415e56",
          7221 => x"a00b83f8",
          7222 => x"fa1c3483",
          7223 => x"f8f83376",
          7224 => x"71291e5a",
          7225 => x"5e83f8f4",
          7226 => x"3386a7b0",
          7227 => x"801a3484",
          7228 => x"b7bc3370",
          7229 => x"81ff0683",
          7230 => x"f8f62283",
          7231 => x"f8f93372",
          7232 => x"7229115b",
          7233 => x"445a4059",
          7234 => x"83f8f433",
          7235 => x"84989a18",
          7236 => x"34608105",
          7237 => x"7081ff06",
          7238 => x"5b587e7a",
          7239 => x"2681ac38",
          7240 => x"84b7bd33",
          7241 => x"587792fb",
          7242 => x"38ff1956",
          7243 => x"7583f8f9",
          7244 => x"34811c70",
          7245 => x"81ff065d",
          7246 => x"597b8326",
          7247 => x"f7a73883",
          7248 => x"f8f83384",
          7249 => x"b7bc3383",
          7250 => x"f8f93372",
          7251 => x"81ff0672",
          7252 => x"81ff0672",
          7253 => x"81ff0672",
          7254 => x"72290554",
          7255 => x"5b435b5b",
          7256 => x"5b84b7e4",
          7257 => x"3386a7a0",
          7258 => x"801b3484",
          7259 => x"b7bc3383",
          7260 => x"f8f93383",
          7261 => x"f8f62272",
          7262 => x"7129125e",
          7263 => x"415e56a0",
          7264 => x"0b83f8fa",
          7265 => x"1c3483f8",
          7266 => x"f8337671",
          7267 => x"291e5a5e",
          7268 => x"83f8f433",
          7269 => x"86a7b080",
          7270 => x"1a3484b7",
          7271 => x"bc337081",
          7272 => x"ff0683f8",
          7273 => x"f62283f8",
          7274 => x"f9337272",
          7275 => x"29115b44",
          7276 => x"5a405983",
          7277 => x"f8f43384",
          7278 => x"989a1834",
          7279 => x"60810570",
          7280 => x"81ff065b",
          7281 => x"58797f27",
          7282 => x"fed63877",
          7283 => x"83f8f934",
          7284 => x"fedf3982",
          7285 => x"0b84b8c4",
          7286 => x"0c800b84",
          7287 => x"b9c80c9c",
          7288 => x"3d0d0483",
          7289 => x"f8fa1733",
          7290 => x"5984b7c4",
          7291 => x"19337a34",
          7292 => x"83f8f933",
          7293 => x"7081ff06",
          7294 => x"58ff0556",
          7295 => x"f9ca3981",
          7296 => x"0b84b8ca",
          7297 => x"34800b84",
          7298 => x"b9c80c9c",
          7299 => x"3d0d0483",
          7300 => x"f8fa1733",
          7301 => x"5b84b7c4",
          7302 => x"1b337c34",
          7303 => x"83f8f833",
          7304 => x"84b7bc33",
          7305 => x"83f8f933",
          7306 => x"5b5b5b80",
          7307 => x"5cfcf439",
          7308 => x"84b8cc42",
          7309 => x"9c3ddc11",
          7310 => x"53d80551",
          7311 => x"ff8ac73f",
          7312 => x"84b9c808",
          7313 => x"802efbf0",
          7314 => x"3884b8c9",
          7315 => x"33811157",
          7316 => x"5a7584b8",
          7317 => x"c9347910",
          7318 => x"83fe0641",
          7319 => x"0280ca05",
          7320 => x"226184b9",
          7321 => x"9c0523fb",
          7322 => x"cf3983f8",
          7323 => x"fa17335c",
          7324 => x"84b7c41c",
          7325 => x"337b3483",
          7326 => x"f8f83384",
          7327 => x"b7bc3383",
          7328 => x"f8f9335b",
          7329 => x"5b5cf9e5",
          7330 => x"3984b7bc",
          7331 => x"3383f8f8",
          7332 => x"3383f8f9",
          7333 => x"33727229",
          7334 => x"05415d5b",
          7335 => x"84b7c419",
          7336 => x"337f86a7",
          7337 => x"a0800534",
          7338 => x"84b7bc33",
          7339 => x"83f8f933",
          7340 => x"83f8f622",
          7341 => x"72712912",
          7342 => x"5a435b56",
          7343 => x"7883f8fa",
          7344 => x"183483f8",
          7345 => x"f8337671",
          7346 => x"291b415e",
          7347 => x"83f8f433",
          7348 => x"6086a7b0",
          7349 => x"80053484",
          7350 => x"b7bc3370",
          7351 => x"81ff0683",
          7352 => x"f8f62283",
          7353 => x"f8f93372",
          7354 => x"72291141",
          7355 => x"5f5a425a",
          7356 => x"83f8f433",
          7357 => x"84989a1e",
          7358 => x"34811c70",
          7359 => x"81ff065c",
          7360 => x"58607b26",
          7361 => x"90a23884",
          7362 => x"b7bd3358",
          7363 => x"7790e238",
          7364 => x"ff1a5675",
          7365 => x"83f8f934",
          7366 => x"800b84b8",
          7367 => x"c40c84b7",
          7368 => x"bf33407f",
          7369 => x"802ef3bd",
          7370 => x"3884b7c0",
          7371 => x"335675f3",
          7372 => x"b4387852",
          7373 => x"8151eae4",
          7374 => x"3f800b84",
          7375 => x"b9c80c9c",
          7376 => x"3d0d0484",
          7377 => x"b9b03383",
          7378 => x"f8f83484",
          7379 => x"b9b13383",
          7380 => x"f8f93484",
          7381 => x"b9b23357",
          7382 => x"7683f8f6",
          7383 => x"23ffb939",
          7384 => x"83f8f833",
          7385 => x"84b9b034",
          7386 => x"83f8f933",
          7387 => x"84b9b134",
          7388 => x"83f8f733",
          7389 => x"84b9b234",
          7390 => x"ff9e3984",
          7391 => x"b8c9335b",
          7392 => x"7a802eff",
          7393 => x"933884b9",
          7394 => x"9c225d7c",
          7395 => x"862e0981",
          7396 => x"06ff8538",
          7397 => x"83f8f933",
          7398 => x"81055583",
          7399 => x"f8f83381",
          7400 => x"05549b53",
          7401 => x"83e48452",
          7402 => x"943d7052",
          7403 => x"57feedf8",
          7404 => x"3f7651fe",
          7405 => x"fef23f84",
          7406 => x"b9c80881",
          7407 => x"ff0683f7",
          7408 => x"cc335776",
          7409 => x"054160a0",
          7410 => x"24fecd38",
          7411 => x"765283f7",
          7412 => x"ac51fefd",
          7413 => x"bd3ffec0",
          7414 => x"39800b84",
          7415 => x"b8c9335b",
          7416 => x"587981ff",
          7417 => x"065b777b",
          7418 => x"27fead38",
          7419 => x"771084b9",
          7420 => x"9c058111",
          7421 => x"33574175",
          7422 => x"b1268aa5",
          7423 => x"38751010",
          7424 => x"83c7a405",
          7425 => x"5f7e0804",
          7426 => x"84b8c933",
          7427 => x"5e7d802e",
          7428 => x"8fa43883",
          7429 => x"f8f83384",
          7430 => x"b99d3371",
          7431 => x"71317009",
          7432 => x"709f2c72",
          7433 => x"065a4259",
          7434 => x"5e5c7583",
          7435 => x"f8f834fd",
          7436 => x"e73984b8",
          7437 => x"c9335675",
          7438 => x"802e8ee7",
          7439 => x"3884b99d",
          7440 => x"33ff0570",
          7441 => x"81ff0684",
          7442 => x"b7bc335d",
          7443 => x"575f757b",
          7444 => x"27fdc538",
          7445 => x"7583f8f9",
          7446 => x"34fdbd39",
          7447 => x"800b83f8",
          7448 => x"f93483f8",
          7449 => x"f8337081",
          7450 => x"ff065d57",
          7451 => x"7b802efd",
          7452 => x"a738ff17",
          7453 => x"567583f8",
          7454 => x"f834fd9c",
          7455 => x"39800b83",
          7456 => x"f8f93483",
          7457 => x"f8f83384",
          7458 => x"b7bb33ff",
          7459 => x"05575776",
          7460 => x"7625fd84",
          7461 => x"38811756",
          7462 => x"7583f8f8",
          7463 => x"34fcf939",
          7464 => x"84b8c933",
          7465 => x"407f802e",
          7466 => x"8de03883",
          7467 => x"f8f93384",
          7468 => x"b99d3371",
          7469 => x"71317009",
          7470 => x"709f2c72",
          7471 => x"065a4159",
          7472 => x"425a7583",
          7473 => x"f8f934fc",
          7474 => x"cf3984b8",
          7475 => x"c9335b7a",
          7476 => x"802efcc4",
          7477 => x"3884b99c",
          7478 => x"22416099",
          7479 => x"2e098106",
          7480 => x"fcb63884",
          7481 => x"b7bc3383",
          7482 => x"f8f93383",
          7483 => x"f8f83372",
          7484 => x"71291286",
          7485 => x"a7a08011",
          7486 => x"83f8f622",
          7487 => x"43515a58",
          7488 => x"71602905",
          7489 => x"7083ffff",
          7490 => x"0683f7cc",
          7491 => x"0887fffe",
          7492 => x"8006425a",
          7493 => x"5d5d7e84",
          7494 => x"82802e92",
          7495 => x"bf38800b",
          7496 => x"83f7cd34",
          7497 => x"fbf23984",
          7498 => x"b8c9335a",
          7499 => x"79802efb",
          7500 => x"e73884b9",
          7501 => x"9c225877",
          7502 => x"992e0981",
          7503 => x"06fbd938",
          7504 => x"810b83f7",
          7505 => x"cd34fbd0",
          7506 => x"3984b8c9",
          7507 => x"33567580",
          7508 => x"2e90be38",
          7509 => x"84b99d33",
          7510 => x"83f8f933",
          7511 => x"5d7c0584",
          7512 => x"b7bc33ff",
          7513 => x"11595e56",
          7514 => x"757d2583",
          7515 => x"38755776",
          7516 => x"83f8f934",
          7517 => x"fba23984",
          7518 => x"b8c93357",
          7519 => x"76802e8c",
          7520 => x"c83884b9",
          7521 => x"9d3383f8",
          7522 => x"f8334261",
          7523 => x"0584b7bb",
          7524 => x"33ff1159",
          7525 => x"41567560",
          7526 => x"25833875",
          7527 => x"577683f8",
          7528 => x"f834faf4",
          7529 => x"3983e490",
          7530 => x"51fee8dc",
          7531 => x"3f800b84",
          7532 => x"b8c93357",
          7533 => x"57767627",
          7534 => x"8bc73876",
          7535 => x"1084b99c",
          7536 => x"05702253",
          7537 => x"5a83e3f0",
          7538 => x"51fee8bc",
          7539 => x"3f811770",
          7540 => x"81ff0684",
          7541 => x"b8c93358",
          7542 => x"5858da39",
          7543 => x"820b84b8",
          7544 => x"c9335f57",
          7545 => x"7d802e8d",
          7546 => x"3884b99c",
          7547 => x"22567583",
          7548 => x"26833875",
          7549 => x"57815276",
          7550 => x"81ff0651",
          7551 => x"d5f33ffa",
          7552 => x"973984b8",
          7553 => x"c9335781",
          7554 => x"77278eb7",
          7555 => x"3884b99f",
          7556 => x"33ff0570",
          7557 => x"81ff0684",
          7558 => x"b99d33ff",
          7559 => x"057081ff",
          7560 => x"0684b7bb",
          7561 => x"337081ff",
          7562 => x"06ff1140",
          7563 => x"43525b59",
          7564 => x"5c5c777e",
          7565 => x"27833877",
          7566 => x"5a7983f8",
          7567 => x"f6237681",
          7568 => x"ff06ff18",
          7569 => x"585f777f",
          7570 => x"27833877",
          7571 => x"577683f8",
          7572 => x"f83484b7",
          7573 => x"bc33ff11",
          7574 => x"57407a60",
          7575 => x"27f9b438",
          7576 => x"7a567583",
          7577 => x"f8f934f9",
          7578 => x"af3984b8",
          7579 => x"c9335f7e",
          7580 => x"802e8aef",
          7581 => x"3884b99d",
          7582 => x"3384b7bb",
          7583 => x"33405b7a",
          7584 => x"7f26f994",
          7585 => x"3883f8f8",
          7586 => x"3384b7bc",
          7587 => x"337081ff",
          7588 => x"0683f8f9",
          7589 => x"33717429",
          7590 => x"1186a7a0",
          7591 => x"800583f8",
          7592 => x"f6225f40",
          7593 => x"717e2905",
          7594 => x"7083ffff",
          7595 => x"0683f7ce",
          7596 => x"33465259",
          7597 => x"595f5d60",
          7598 => x"812e84f0",
          7599 => x"387983ff",
          7600 => x"ff06707c",
          7601 => x"315d5780",
          7602 => x"7c248efe",
          7603 => x"3884b7bb",
          7604 => x"33567676",
          7605 => x"278ed638",
          7606 => x"ff165675",
          7607 => x"83f8f623",
          7608 => x"7c81ff06",
          7609 => x"707c3141",
          7610 => x"57806024",
          7611 => x"8ee53884",
          7612 => x"b7bb3356",
          7613 => x"7676278d",
          7614 => x"ee38ff16",
          7615 => x"567583f8",
          7616 => x"f8347e81",
          7617 => x"ff0683f8",
          7618 => x"f6225757",
          7619 => x"805a7676",
          7620 => x"26903875",
          7621 => x"77318105",
          7622 => x"7e81ff06",
          7623 => x"7171295c",
          7624 => x"5e5b7958",
          7625 => x"86a7a080",
          7626 => x"5b86a7b0",
          7627 => x"807f81ff",
          7628 => x"067f81ff",
          7629 => x"06717129",
          7630 => x"1d425842",
          7631 => x"5c797f27",
          7632 => x"f7d63884",
          7633 => x"989a1a57",
          7634 => x"e0e01733",
          7635 => x"5f84b7c4",
          7636 => x"1f337b70",
          7637 => x"81055d34",
          7638 => x"76708105",
          7639 => x"58337c70",
          7640 => x"81055e34",
          7641 => x"811884b7",
          7642 => x"bc3384b7",
          7643 => x"bb337171",
          7644 => x"291d4340",
          7645 => x"5e587760",
          7646 => x"27f79d38",
          7647 => x"e0e01733",
          7648 => x"5f84b7c4",
          7649 => x"1f337b70",
          7650 => x"81055d34",
          7651 => x"76708105",
          7652 => x"58337c70",
          7653 => x"81055e34",
          7654 => x"811884b7",
          7655 => x"bc3384b7",
          7656 => x"bb337171",
          7657 => x"291d4340",
          7658 => x"5e587f78",
          7659 => x"26ff9938",
          7660 => x"f6e63984",
          7661 => x"b8c93356",
          7662 => x"75802e87",
          7663 => x"e0388052",
          7664 => x"84b99d33",
          7665 => x"51d8b13f",
          7666 => x"f6ce3980",
          7667 => x"0b84b7bc",
          7668 => x"33ff1184",
          7669 => x"b8c9335d",
          7670 => x"59405879",
          7671 => x"782e9438",
          7672 => x"84b99c22",
          7673 => x"5675782e",
          7674 => x"0981068b",
          7675 => x"be3883f8",
          7676 => x"f9335876",
          7677 => x"81ff0683",
          7678 => x"f8f83379",
          7679 => x"435c5c76",
          7680 => x"ff2e81ed",
          7681 => x"3884b7bb",
          7682 => x"33407a60",
          7683 => x"26f68938",
          7684 => x"7e81ff06",
          7685 => x"56607626",
          7686 => x"f5fe387b",
          7687 => x"7626617d",
          7688 => x"27075776",
          7689 => x"f5f2387a",
          7690 => x"10101b70",
          7691 => x"90296205",
          7692 => x"86a7a080",
          7693 => x"11701f5d",
          7694 => x"5a86a7b0",
          7695 => x"80057983",
          7696 => x"0658515d",
          7697 => x"758bac38",
          7698 => x"79830657",
          7699 => x"768ba438",
          7700 => x"83f8f433",
          7701 => x"70982b71",
          7702 => x"902b0771",
          7703 => x"882b0771",
          7704 => x"07797f59",
          7705 => x"525f5777",
          7706 => x"7a279e38",
          7707 => x"80777084",
          7708 => x"05590c7d",
          7709 => x"76708405",
          7710 => x"580c7977",
          7711 => x"26ee3884",
          7712 => x"b7bc3384",
          7713 => x"b7bb3341",
          7714 => x"5f7e81ff",
          7715 => x"066081ff",
          7716 => x"0683f8f6",
          7717 => x"227d7329",
          7718 => x"64055959",
          7719 => x"595a7777",
          7720 => x"268c3876",
          7721 => x"78311b70",
          7722 => x"7b296205",
          7723 => x"57407576",
          7724 => x"1d575776",
          7725 => x"7626f4e0",
          7726 => x"3883f8f4",
          7727 => x"3384989a",
          7728 => x"18595aa0",
          7729 => x"0be0e019",
          7730 => x"34797870",
          7731 => x"81055a34",
          7732 => x"81175776",
          7733 => x"7626f4c0",
          7734 => x"38a00be0",
          7735 => x"e0193479",
          7736 => x"78708105",
          7737 => x"5a348117",
          7738 => x"57757727",
          7739 => x"d638f4a8",
          7740 => x"39ff1f70",
          7741 => x"81ff065d",
          7742 => x"58fe8a39",
          7743 => x"83f8f433",
          7744 => x"7080f006",
          7745 => x"71842b80",
          7746 => x"f0067184",
          7747 => x"2a07585d",
          7748 => x"577b80f0",
          7749 => x"2e098106",
          7750 => x"be3880f2",
          7751 => x"0b83f8f4",
          7752 => x"34811870",
          7753 => x"81ff0659",
          7754 => x"56f5b639",
          7755 => x"83f8fa17",
          7756 => x"335e84b7",
          7757 => x"c41e337c",
          7758 => x"3483f8f8",
          7759 => x"3384b7bc",
          7760 => x"3383f8f6",
          7761 => x"2284b7bb",
          7762 => x"33425c5f",
          7763 => x"5dfaee39",
          7764 => x"83f8f433",
          7765 => x"87075675",
          7766 => x"83f8f434",
          7767 => x"81187081",
          7768 => x"ff065956",
          7769 => x"f4fb3983",
          7770 => x"f8f43381",
          7771 => x"fd068507",
          7772 => x"567583f8",
          7773 => x"f434e539",
          7774 => x"83f8f433",
          7775 => x"81fb0683",
          7776 => x"07567583",
          7777 => x"f8f434d4",
          7778 => x"3983f8f4",
          7779 => x"3381f906",
          7780 => x"81075675",
          7781 => x"83f8f434",
          7782 => x"c33983f8",
          7783 => x"f433819f",
          7784 => x"06900756",
          7785 => x"7583f8f4",
          7786 => x"34ffb139",
          7787 => x"80f10b83",
          7788 => x"f8f43481",
          7789 => x"187081ff",
          7790 => x"065956f4",
          7791 => x"a43983f8",
          7792 => x"f433818f",
          7793 => x"06567583",
          7794 => x"f8f434ff",
          7795 => x"8f3983f8",
          7796 => x"f433819f",
          7797 => x"06900756",
          7798 => x"7583f8f4",
          7799 => x"34fefd39",
          7800 => x"83f8f433",
          7801 => x"81ef0680",
          7802 => x"e0075675",
          7803 => x"83f8f434",
          7804 => x"feea3983",
          7805 => x"f8f43381",
          7806 => x"cf0680c0",
          7807 => x"07567583",
          7808 => x"f8f434fe",
          7809 => x"d73983f8",
          7810 => x"f43381af",
          7811 => x"06a00756",
          7812 => x"7583f8f4",
          7813 => x"34fec539",
          7814 => x"83f8f433",
          7815 => x"81fe0686",
          7816 => x"07567583",
          7817 => x"f8f434fe",
          7818 => x"b33983f8",
          7819 => x"f43381fc",
          7820 => x"06840756",
          7821 => x"7583f8f4",
          7822 => x"34fea139",
          7823 => x"83f8f433",
          7824 => x"81fa0682",
          7825 => x"07567583",
          7826 => x"f8f434fe",
          7827 => x"8f3983f8",
          7828 => x"f43381f8",
          7829 => x"06567583",
          7830 => x"f8f434fd",
          7831 => x"ff3983f8",
          7832 => x"f43380f0",
          7833 => x"07567583",
          7834 => x"f8f434fd",
          7835 => x"ef3983f8",
          7836 => x"f43380f0",
          7837 => x"07567583",
          7838 => x"f8f434fd",
          7839 => x"df3983f8",
          7840 => x"f43381df",
          7841 => x"0680d007",
          7842 => x"567583f8",
          7843 => x"f434fdcc",
          7844 => x"3983f8f4",
          7845 => x"3381bf06",
          7846 => x"b0075675",
          7847 => x"83f8f434",
          7848 => x"fdba3980",
          7849 => x"0b83f8f9",
          7850 => x"34805281",
          7851 => x"51d2c93f",
          7852 => x"ecff3984",
          7853 => x"b9b03383",
          7854 => x"f8f83484",
          7855 => x"b9b13383",
          7856 => x"f8f93484",
          7857 => x"b9b23359",
          7858 => x"7883f8f6",
          7859 => x"23800b84",
          7860 => x"b8c40ce8",
          7861 => x"c739810b",
          7862 => x"84b8cb34",
          7863 => x"800b84b9",
          7864 => x"c80c9c3d",
          7865 => x"0d047783",
          7866 => x"f8f93483",
          7867 => x"f8f93370",
          7868 => x"81ff0658",
          7869 => x"ff0556e7",
          7870 => x"cf3984b8",
          7871 => x"cc429c3d",
          7872 => x"dc1153d8",
          7873 => x"0551fef8",
          7874 => x"fd3f84b9",
          7875 => x"c808a138",
          7876 => x"84b9c808",
          7877 => x"84b8c40c",
          7878 => x"800b84b8",
          7879 => x"c834800b",
          7880 => x"84b9c80c",
          7881 => x"9c3d0d04",
          7882 => x"7783f8f9",
          7883 => x"34efe939",
          7884 => x"84b8c933",
          7885 => x"81115c5c",
          7886 => x"7a84b8c9",
          7887 => x"347b1083",
          7888 => x"fe065d02",
          7889 => x"80ca0522",
          7890 => x"84b99c1e",
          7891 => x"23800b84",
          7892 => x"b8c834ca",
          7893 => x"39800b83",
          7894 => x"f8f93480",
          7895 => x"528151d1",
          7896 => x"973f83f8",
          7897 => x"f9337081",
          7898 => x"ff0658ff",
          7899 => x"0556e6d8",
          7900 => x"39800b83",
          7901 => x"f8f93480",
          7902 => x"528151d0",
          7903 => x"fb3fef98",
          7904 => x"398a51fe",
          7905 => x"ebd83fef",
          7906 => x"8f3983f8",
          7907 => x"f933ff05",
          7908 => x"7009709f",
          7909 => x"2c720658",
          7910 => x"5f57f2a6",
          7911 => x"39755281",
          7912 => x"51d93984",
          7913 => x"b7bc3340",
          7914 => x"756027ee",
          7915 => x"eb387583",
          7916 => x"f8f934ee",
          7917 => x"e33983f8",
          7918 => x"f833ff05",
          7919 => x"7009709f",
          7920 => x"2c720658",
          7921 => x"4057f0e2",
          7922 => x"3983f8f8",
          7923 => x"33810584",
          7924 => x"b7bb33ff",
          7925 => x"11595956",
          7926 => x"757825f3",
          7927 => x"c0387557",
          7928 => x"f3bb3984",
          7929 => x"b7bb3370",
          7930 => x"81ff0658",
          7931 => x"5c817726",
          7932 => x"eea63883",
          7933 => x"f8f83384",
          7934 => x"b7bc3370",
          7935 => x"81ff0683",
          7936 => x"f8f93371",
          7937 => x"74291186",
          7938 => x"a7a08005",
          7939 => x"83f8f622",
          7940 => x"5f5f717e",
          7941 => x"29057083",
          7942 => x"ffff0683",
          7943 => x"f7ce335d",
          7944 => x"5b44425f",
          7945 => x"5d77812e",
          7946 => x"81f53879",
          7947 => x"83ffff06",
          7948 => x"ff115c57",
          7949 => x"807b2484",
          7950 => x"893884b7",
          7951 => x"bb335676",
          7952 => x"76278398",
          7953 => x"38ff1656",
          7954 => x"7583f8f6",
          7955 => x"237c81ff",
          7956 => x"06ff1157",
          7957 => x"57807624",
          7958 => x"83df3884",
          7959 => x"b7bb3356",
          7960 => x"76762782",
          7961 => x"ec38ff16",
          7962 => x"567583f8",
          7963 => x"f8347b81",
          7964 => x"ff0683f8",
          7965 => x"f6225757",
          7966 => x"805a7676",
          7967 => x"26903875",
          7968 => x"77318105",
          7969 => x"7e81ff06",
          7970 => x"7171295c",
          7971 => x"5e5f7958",
          7972 => x"86a7a080",
          7973 => x"5b86a7b0",
          7974 => x"807c81ff",
          7975 => x"067f81ff",
          7976 => x"06717129",
          7977 => x"1d414242",
          7978 => x"5d797e27",
          7979 => x"ecea3884",
          7980 => x"989a1a57",
          7981 => x"e0e01733",
          7982 => x"5e84b7c4",
          7983 => x"1e337b70",
          7984 => x"81055d34",
          7985 => x"76708105",
          7986 => x"58337d70",
          7987 => x"81055f34",
          7988 => x"811884b7",
          7989 => x"bc3384b7",
          7990 => x"bb337171",
          7991 => x"291d5941",
          7992 => x"5d587776",
          7993 => x"27ecb138",
          7994 => x"e0e01733",
          7995 => x"5e84b7c4",
          7996 => x"1e337b70",
          7997 => x"81055d34",
          7998 => x"76708105",
          7999 => x"58337d70",
          8000 => x"81055f34",
          8001 => x"811884b7",
          8002 => x"bc3384b7",
          8003 => x"bb337171",
          8004 => x"291d5941",
          8005 => x"5d587578",
          8006 => x"26ff9938",
          8007 => x"ebfa3983",
          8008 => x"f8fa1733",
          8009 => x"5c84b7c4",
          8010 => x"1c337b34",
          8011 => x"83f8f833",
          8012 => x"84b7bc33",
          8013 => x"83f8f622",
          8014 => x"84b7bb33",
          8015 => x"5f5c5f5d",
          8016 => x"fde93976",
          8017 => x"ebd23884",
          8018 => x"b7bb3370",
          8019 => x"81ff06ff",
          8020 => x"115c4258",
          8021 => x"76612783",
          8022 => x"38765a79",
          8023 => x"83f8f623",
          8024 => x"7781ff06",
          8025 => x"ff19585a",
          8026 => x"807a2783",
          8027 => x"38805776",
          8028 => x"83f8f834",
          8029 => x"84b7bc33",
          8030 => x"7081ff06",
          8031 => x"ff125259",
          8032 => x"56807827",
          8033 => x"eb8d3880",
          8034 => x"567583f8",
          8035 => x"f934eb88",
          8036 => x"3983f8f9",
          8037 => x"33810584",
          8038 => x"b7bc33ff",
          8039 => x"11594056",
          8040 => x"757f25ef",
          8041 => x"ca387557",
          8042 => x"efc53975",
          8043 => x"812e0981",
          8044 => x"06f4c038",
          8045 => x"83f8f933",
          8046 => x"7081ff06",
          8047 => x"83f8f833",
          8048 => x"7a445d5d",
          8049 => x"5776ff2e",
          8050 => x"098106f4",
          8051 => x"b838f6a1",
          8052 => x"39ff1d56",
          8053 => x"7583f8f8",
          8054 => x"34fd9339",
          8055 => x"ff1a5675",
          8056 => x"83f8f623",
          8057 => x"fce7397c",
          8058 => x"7b315675",
          8059 => x"83f8f834",
          8060 => x"f2903977",
          8061 => x"7d585677",
          8062 => x"7a26f58d",
          8063 => x"38807670",
          8064 => x"81055834",
          8065 => x"83f8f433",
          8066 => x"77708105",
          8067 => x"5934757a",
          8068 => x"26f4ec38",
          8069 => x"80767081",
          8070 => x"05583483",
          8071 => x"f8f43377",
          8072 => x"70810559",
          8073 => x"34797627",
          8074 => x"d438f4d3",
          8075 => x"39797b31",
          8076 => x"567583f8",
          8077 => x"f623f1a8",
          8078 => x"39800b83",
          8079 => x"f8f834fc",
          8080 => x"ad397e83",
          8081 => x"f8f623fc",
          8082 => x"8439800b",
          8083 => x"83f8f623",
          8084 => x"f18e3980",
          8085 => x"0b83f8f8",
          8086 => x"34f1a739",
          8087 => x"83f8fa18",
          8088 => x"335a84b7",
          8089 => x"c41a3377",
          8090 => x"34800b83",
          8091 => x"f7cd34e9",
          8092 => x"a739fd3d",
          8093 => x"0d029705",
          8094 => x"3384b7be",
          8095 => x"33545472",
          8096 => x"802e9038",
          8097 => x"7351db9c",
          8098 => x"3f800b84",
          8099 => x"b9c80c85",
          8100 => x"3d0d0476",
          8101 => x"527351d7",
          8102 => x"ab3f800b",
          8103 => x"84b9c80c",
          8104 => x"853d0d04",
          8105 => x"f33d0d02",
          8106 => x"bf05335c",
          8107 => x"ff0b83f7",
          8108 => x"cc337081",
          8109 => x"ff0683f7",
          8110 => x"ac113358",
          8111 => x"55555974",
          8112 => x"802e80d6",
          8113 => x"38811456",
          8114 => x"7583f7cc",
          8115 => x"34745978",
          8116 => x"84b9c80c",
          8117 => x"8f3d0d04",
          8118 => x"83f7a808",
          8119 => x"54825373",
          8120 => x"802e9138",
          8121 => x"73733270",
          8122 => x"30710770",
          8123 => x"09709f2a",
          8124 => x"565d5e58",
          8125 => x"7283f7a8",
          8126 => x"0cff5980",
          8127 => x"547b812e",
          8128 => x"09810683",
          8129 => x"387b547b",
          8130 => x"83327030",
          8131 => x"70802576",
          8132 => x"075c5c5d",
          8133 => x"79802e85",
          8134 => x"c43884b7",
          8135 => x"bc3383f8",
          8136 => x"f93383f8",
          8137 => x"f8337271",
          8138 => x"291286a7",
          8139 => x"a0800583",
          8140 => x"f8f6225b",
          8141 => x"595d7179",
          8142 => x"29057083",
          8143 => x"ffff0683",
          8144 => x"f7cd3358",
          8145 => x"59555874",
          8146 => x"812e838c",
          8147 => x"3881f054",
          8148 => x"7386ee80",
          8149 => x"8034800b",
          8150 => x"87c09888",
          8151 => x"0c87c098",
          8152 => x"88085675",
          8153 => x"802ef638",
          8154 => x"86ee8084",
          8155 => x"08577683",
          8156 => x"f4f81534",
          8157 => x"81147081",
          8158 => x"ff065555",
          8159 => x"81f97427",
          8160 => x"cf388054",
          8161 => x"83f6e814",
          8162 => x"337081ff",
          8163 => x"0683f6f2",
          8164 => x"16335854",
          8165 => x"5572762e",
          8166 => x"85c13872",
          8167 => x"81ff2e86",
          8168 => x"b4387483",
          8169 => x"f6fc1534",
          8170 => x"7581ff06",
          8171 => x"5a7981ff",
          8172 => x"2e85cd38",
          8173 => x"7583f786",
          8174 => x"153483f6",
          8175 => x"e8143383",
          8176 => x"f6f21534",
          8177 => x"81147081",
          8178 => x"ff06555e",
          8179 => x"897427ff",
          8180 => x"b33883f6",
          8181 => x"f0337098",
          8182 => x"2b708025",
          8183 => x"58565475",
          8184 => x"83f7a034",
          8185 => x"7381ff06",
          8186 => x"70862a81",
          8187 => x"32708106",
          8188 => x"51545872",
          8189 => x"802e85e7",
          8190 => x"38810b83",
          8191 => x"f7a13473",
          8192 => x"09810653",
          8193 => x"72802e85",
          8194 => x"e438810b",
          8195 => x"83f7a234",
          8196 => x"800b83f7",
          8197 => x"a13383f7",
          8198 => x"a80883f7",
          8199 => x"a2337083",
          8200 => x"f7a43383",
          8201 => x"f7a3335d",
          8202 => x"5d425e5c",
          8203 => x"5e5683f6",
          8204 => x"fc163355",
          8205 => x"7481ff2e",
          8206 => x"8d3883f7",
          8207 => x"90163354",
          8208 => x"73802e82",
          8209 => x"823883f7",
          8210 => x"86163353",
          8211 => x"7281ff2e",
          8212 => x"8b3883f7",
          8213 => x"90163354",
          8214 => x"7381ec38",
          8215 => x"7481ff06",
          8216 => x"547381ff",
          8217 => x"2e8d3883",
          8218 => x"f7901633",
          8219 => x"5372812e",
          8220 => x"81da3874",
          8221 => x"81ff0653",
          8222 => x"7281ff2e",
          8223 => x"848c3883",
          8224 => x"f7901633",
          8225 => x"54817427",
          8226 => x"84803883",
          8227 => x"f79c0887",
          8228 => x"e80587c0",
          8229 => x"989c0854",
          8230 => x"54737327",
          8231 => x"83ec3881",
          8232 => x"0b87c098",
          8233 => x"9c0883f7",
          8234 => x"9c0c5881",
          8235 => x"167081ff",
          8236 => x"06575489",
          8237 => x"7627fef6",
          8238 => x"387683f7",
          8239 => x"a3347783",
          8240 => x"f7a434fe",
          8241 => x"9e195372",
          8242 => x"9c26828b",
          8243 => x"38721010",
          8244 => x"83c8ec05",
          8245 => x"5a790804",
          8246 => x"83f7d008",
          8247 => x"5473802e",
          8248 => x"913883f4",
          8249 => x"1487c098",
          8250 => x"9c085e5e",
          8251 => x"7d7d27fc",
          8252 => x"dc38800b",
          8253 => x"83f7ce33",
          8254 => x"54547281",
          8255 => x"2e833874",
          8256 => x"547383f7",
          8257 => x"ce3487c0",
          8258 => x"989c0883",
          8259 => x"f7d00c73",
          8260 => x"81ff0658",
          8261 => x"77812e94",
          8262 => x"3883f8fa",
          8263 => x"17335484",
          8264 => x"b7c41433",
          8265 => x"763481f0",
          8266 => x"54fca539",
          8267 => x"83f7a808",
          8268 => x"5372802e",
          8269 => x"829c3872",
          8270 => x"812e83f4",
          8271 => x"3880c376",
          8272 => x"3481f054",
          8273 => x"fc8a3980",
          8274 => x"58fee039",
          8275 => x"80745657",
          8276 => x"83597c81",
          8277 => x"2e9b3879",
          8278 => x"772e0981",
          8279 => x"0683b438",
          8280 => x"7d812e80",
          8281 => x"ed387981",
          8282 => x"2e80d738",
          8283 => x"7981ff06",
          8284 => x"59877727",
          8285 => x"75982b54",
          8286 => x"54728025",
          8287 => x"a1387380",
          8288 => x"2e9c3881",
          8289 => x"177081ff",
          8290 => x"06761081",
          8291 => x"fe068772",
          8292 => x"2771982b",
          8293 => x"57535758",
          8294 => x"54807324",
          8295 => x"e1387810",
          8296 => x"10107910",
          8297 => x"05761183",
          8298 => x"2b780583",
          8299 => x"f3d80570",
          8300 => x"335b5654",
          8301 => x"7887c098",
          8302 => x"9c0883f7",
          8303 => x"9c0c57fd",
          8304 => x"ea398059",
          8305 => x"7d812eff",
          8306 => x"a8387981",
          8307 => x"ff0659ff",
          8308 => x"a0398259",
          8309 => x"ff9b3978",
          8310 => x"ff2efa9f",
          8311 => x"38800b84",
          8312 => x"b7be3354",
          8313 => x"5472812e",
          8314 => x"83e8387b",
          8315 => x"82327030",
          8316 => x"70802576",
          8317 => x"07405956",
          8318 => x"7d8a387b",
          8319 => x"832e0981",
          8320 => x"06f9cc38",
          8321 => x"78ff2ef9",
          8322 => x"c6388053",
          8323 => x"72101010",
          8324 => x"83f7d405",
          8325 => x"70335d54",
          8326 => x"787c2e83",
          8327 => x"ba388113",
          8328 => x"7081ff06",
          8329 => x"54579373",
          8330 => x"27e23884",
          8331 => x"b7bf3353",
          8332 => x"72802ef9",
          8333 => x"9a3884b7",
          8334 => x"c0335574",
          8335 => x"f9913878",
          8336 => x"81ff0652",
          8337 => x"8251ccd4",
          8338 => x"3f7884b9",
          8339 => x"c80c8f3d",
          8340 => x"0d04be76",
          8341 => x"3481f054",
          8342 => x"f9f63972",
          8343 => x"81ff2e92",
          8344 => x"3883f790",
          8345 => x"14338105",
          8346 => x"5b7a83f7",
          8347 => x"901534fa",
          8348 => x"c939800b",
          8349 => x"83f79015",
          8350 => x"34ff0b83",
          8351 => x"f6fc1534",
          8352 => x"ff0b83f7",
          8353 => x"861534fa",
          8354 => x"b1397481",
          8355 => x"ff065372",
          8356 => x"81ff2efc",
          8357 => x"963883f7",
          8358 => x"90163355",
          8359 => x"817527fc",
          8360 => x"8a387781",
          8361 => x"ff065473",
          8362 => x"812e0981",
          8363 => x"06fbfc38",
          8364 => x"83f79c08",
          8365 => x"81fa0587",
          8366 => x"c0989c08",
          8367 => x"54557473",
          8368 => x"27fbe838",
          8369 => x"87c0989c",
          8370 => x"0883f79c",
          8371 => x"0c7681ff",
          8372 => x"0659fbd7",
          8373 => x"39ff0b83",
          8374 => x"f6fc1534",
          8375 => x"f9ca3972",
          8376 => x"83f7a134",
          8377 => x"73098106",
          8378 => x"5372fa9e",
          8379 => x"387283f7",
          8380 => x"a234800b",
          8381 => x"83f7a133",
          8382 => x"83f7a808",
          8383 => x"83f7a233",
          8384 => x"7083f7a4",
          8385 => x"3383f7a3",
          8386 => x"335d5d42",
          8387 => x"5e5c5e56",
          8388 => x"fa9c3979",
          8389 => x"822e0981",
          8390 => x"06fccb38",
          8391 => x"7a597a81",
          8392 => x"2efcce38",
          8393 => x"79812e09",
          8394 => x"8106fcc0",
          8395 => x"38fd9339",
          8396 => x"ef763481",
          8397 => x"f054f898",
          8398 => x"39800b84",
          8399 => x"b7bf3357",
          8400 => x"54758338",
          8401 => x"81547384",
          8402 => x"b7bf34ff",
          8403 => x"59f7ac39",
          8404 => x"800b84b7",
          8405 => x"be335854",
          8406 => x"76833881",
          8407 => x"547384b7",
          8408 => x"be34ff59",
          8409 => x"f7953981",
          8410 => x"5383f7a8",
          8411 => x"08842ef7",
          8412 => x"8338840b",
          8413 => x"83f7a80c",
          8414 => x"f6ff3984",
          8415 => x"b7bb3370",
          8416 => x"81ff06ff",
          8417 => x"11575a54",
          8418 => x"80792783",
          8419 => x"38805574",
          8420 => x"83f8f623",
          8421 => x"7381ff06",
          8422 => x"ff155553",
          8423 => x"80732783",
          8424 => x"38805473",
          8425 => x"83f8f834",
          8426 => x"84b7bc33",
          8427 => x"7081ff06",
          8428 => x"56ff0553",
          8429 => x"80752783",
          8430 => x"38805372",
          8431 => x"83f8f934",
          8432 => x"ff59f6b7",
          8433 => x"39815283",
          8434 => x"51ffbaa5",
          8435 => x"3fff59f6",
          8436 => x"aa397254",
          8437 => x"fc953984",
          8438 => x"14085283",
          8439 => x"f7ac51fe",
          8440 => x"dee53f81",
          8441 => x"0b83f7cc",
          8442 => x"3483f7ac",
          8443 => x"3359fcbb",
          8444 => x"39803d0d",
          8445 => x"8151f5ac",
          8446 => x"3f823d0d",
          8447 => x"04fa3d0d",
          8448 => x"800b83f3",
          8449 => x"d4085357",
          8450 => x"02a30533",
          8451 => x"82133483",
          8452 => x"f3d40851",
          8453 => x"80e07134",
          8454 => x"850b83f3",
          8455 => x"d4085556",
          8456 => x"fe0b8115",
          8457 => x"34800b86",
          8458 => x"f080e834",
          8459 => x"87c0989c",
          8460 => x"0883f3d4",
          8461 => x"085580ce",
          8462 => x"90055387",
          8463 => x"c0989c08",
          8464 => x"5287c098",
          8465 => x"9c085170",
          8466 => x"722ef638",
          8467 => x"81143387",
          8468 => x"c0989c08",
          8469 => x"56527473",
          8470 => x"27873871",
          8471 => x"81fe2edb",
          8472 => x"3887c098",
          8473 => x"a40851ff",
          8474 => x"55707327",
          8475 => x"80c83871",
          8476 => x"5571ff2e",
          8477 => x"80c03887",
          8478 => x"c0989c08",
          8479 => x"80ce9005",
          8480 => x"5387c098",
          8481 => x"9c085287",
          8482 => x"c0989c08",
          8483 => x"5574722e",
          8484 => x"f6388114",
          8485 => x"3387c098",
          8486 => x"9c085252",
          8487 => x"70732787",
          8488 => x"387181ff",
          8489 => x"2edb3887",
          8490 => x"c098a408",
          8491 => x"55727526",
          8492 => x"8338ff52",
          8493 => x"7155ff16",
          8494 => x"7081ff06",
          8495 => x"57537580",
          8496 => x"2e983874",
          8497 => x"81ff0652",
          8498 => x"71fed538",
          8499 => x"74ff2e8a",
          8500 => x"387684b9",
          8501 => x"c80c883d",
          8502 => x"0d04810b",
          8503 => x"84b9c80c",
          8504 => x"883d0d04",
          8505 => x"fa3d0d79",
          8506 => x"028405a3",
          8507 => x"05335652",
          8508 => x"800b83f3",
          8509 => x"d4087388",
          8510 => x"2b87fc80",
          8511 => x"80067075",
          8512 => x"982a0751",
          8513 => x"55555771",
          8514 => x"83153472",
          8515 => x"902a5170",
          8516 => x"84153471",
          8517 => x"902a5675",
          8518 => x"85153472",
          8519 => x"86153483",
          8520 => x"f3d40852",
          8521 => x"74821334",
          8522 => x"83f3d408",
          8523 => x"5180e171",
          8524 => x"34850b83",
          8525 => x"f3d40855",
          8526 => x"56fe0b81",
          8527 => x"1534800b",
          8528 => x"86f080e8",
          8529 => x"3487c098",
          8530 => x"9c0883f3",
          8531 => x"d4085580",
          8532 => x"ce900553",
          8533 => x"87c0989c",
          8534 => x"085287c0",
          8535 => x"989c0851",
          8536 => x"70722ef6",
          8537 => x"38811433",
          8538 => x"87c0989c",
          8539 => x"08565274",
          8540 => x"73278738",
          8541 => x"7181fe2e",
          8542 => x"db3887c0",
          8543 => x"98a40851",
          8544 => x"ff557073",
          8545 => x"2780c838",
          8546 => x"715571ff",
          8547 => x"2e80c038",
          8548 => x"87c0989c",
          8549 => x"0880ce90",
          8550 => x"055387c0",
          8551 => x"989c0852",
          8552 => x"87c0989c",
          8553 => x"08557472",
          8554 => x"2ef63881",
          8555 => x"143387c0",
          8556 => x"989c0852",
          8557 => x"52707327",
          8558 => x"87387181",
          8559 => x"ff2edb38",
          8560 => x"87c098a4",
          8561 => x"08557275",
          8562 => x"268338ff",
          8563 => x"527155ff",
          8564 => x"167081ff",
          8565 => x"06575375",
          8566 => x"802e80c7",
          8567 => x"387481ff",
          8568 => x"065271fe",
          8569 => x"d4387451",
          8570 => x"7081ff06",
          8571 => x"5675aa38",
          8572 => x"80c6147b",
          8573 => x"84801155",
          8574 => x"52527073",
          8575 => x"27923871",
          8576 => x"70810553",
          8577 => x"33717081",
          8578 => x"05533472",
          8579 => x"7126f038",
          8580 => x"7684b9c8",
          8581 => x"0c883d0d",
          8582 => x"04810b84",
          8583 => x"b9c80c88",
          8584 => x"3d0d04ff",
          8585 => x"51c239fa",
          8586 => x"3d0d7902",
          8587 => x"8405a305",
          8588 => x"33565680",
          8589 => x"0b83f3d4",
          8590 => x"0877882b",
          8591 => x"87fc8080",
          8592 => x"06707998",
          8593 => x"2a075155",
          8594 => x"55577583",
          8595 => x"15347290",
          8596 => x"2a517084",
          8597 => x"15347590",
          8598 => x"2a527185",
          8599 => x"15347286",
          8600 => x"15347a83",
          8601 => x"f3d40880",
          8602 => x"c6118480",
          8603 => x"13565455",
          8604 => x"51707327",
          8605 => x"97387070",
          8606 => x"81055233",
          8607 => x"72708105",
          8608 => x"54347271",
          8609 => x"26f03883",
          8610 => x"f3d40854",
          8611 => x"74821534",
          8612 => x"83f3d408",
          8613 => x"5580e275",
          8614 => x"34850b83",
          8615 => x"f3d40855",
          8616 => x"56fe0b81",
          8617 => x"1534800b",
          8618 => x"86f080e8",
          8619 => x"3487c098",
          8620 => x"9c0883f3",
          8621 => x"d4085580",
          8622 => x"ce900553",
          8623 => x"87c0989c",
          8624 => x"085287c0",
          8625 => x"989c0851",
          8626 => x"70722ef6",
          8627 => x"38811433",
          8628 => x"87c0989c",
          8629 => x"08565274",
          8630 => x"73278738",
          8631 => x"7181fe2e",
          8632 => x"db3887c0",
          8633 => x"98a40851",
          8634 => x"ff557073",
          8635 => x"2780c838",
          8636 => x"715571ff",
          8637 => x"2e80c038",
          8638 => x"87c0989c",
          8639 => x"0880ce90",
          8640 => x"055387c0",
          8641 => x"989c0852",
          8642 => x"87c0989c",
          8643 => x"08557472",
          8644 => x"2ef63881",
          8645 => x"143387c0",
          8646 => x"989c0852",
          8647 => x"52707327",
          8648 => x"87387181",
          8649 => x"ff2edb38",
          8650 => x"87c098a4",
          8651 => x"08557275",
          8652 => x"268338ff",
          8653 => x"527155ff",
          8654 => x"167081ff",
          8655 => x"06575375",
          8656 => x"802ea138",
          8657 => x"7481ff06",
          8658 => x"5271fed5",
          8659 => x"38745170",
          8660 => x"81ff0654",
          8661 => x"73802e83",
          8662 => x"38815776",
          8663 => x"84b9c80c",
          8664 => x"883d0d04",
          8665 => x"ff51e839",
          8666 => x"fb3d0d83",
          8667 => x"f3d40851",
          8668 => x"80d07134",
          8669 => x"850b83f3",
          8670 => x"d4085656",
          8671 => x"fe0b8116",
          8672 => x"34800b86",
          8673 => x"f080e834",
          8674 => x"87c0989c",
          8675 => x"0883f3d4",
          8676 => x"085680ce",
          8677 => x"90055487",
          8678 => x"c0989c08",
          8679 => x"5287c098",
          8680 => x"9c085372",
          8681 => x"722ef638",
          8682 => x"81153387",
          8683 => x"c0989c08",
          8684 => x"52527074",
          8685 => x"27873871",
          8686 => x"81fe2edb",
          8687 => x"3887c098",
          8688 => x"a40851ff",
          8689 => x"53707427",
          8690 => x"80c83871",
          8691 => x"5371ff2e",
          8692 => x"80c03887",
          8693 => x"c0989c08",
          8694 => x"80ce9005",
          8695 => x"5387c098",
          8696 => x"9c085287",
          8697 => x"c0989c08",
          8698 => x"5170722e",
          8699 => x"f6388115",
          8700 => x"3387c098",
          8701 => x"9c085552",
          8702 => x"73732787",
          8703 => x"387181ff",
          8704 => x"2edb3887",
          8705 => x"c098a408",
          8706 => x"51727126",
          8707 => x"8338ff52",
          8708 => x"7153ff16",
          8709 => x"7081ff06",
          8710 => x"57527580",
          8711 => x"2e8a3872",
          8712 => x"81ff0654",
          8713 => x"73fed538",
          8714 => x"ff39803d",
          8715 => x"0d83e4cc",
          8716 => x"51fed0bf",
          8717 => x"3f823d0d",
          8718 => x"04f93d0d",
          8719 => x"84b9b808",
          8720 => x"7a713183",
          8721 => x"2a7083ff",
          8722 => x"ff067083",
          8723 => x"2b731170",
          8724 => x"33811233",
          8725 => x"718b2b71",
          8726 => x"832b0777",
          8727 => x"11703381",
          8728 => x"12337198",
          8729 => x"2b71902b",
          8730 => x"075c5441",
          8731 => x"53535d57",
          8732 => x"59525657",
          8733 => x"53807124",
          8734 => x"81af3872",
          8735 => x"16821133",
          8736 => x"83123371",
          8737 => x"8b2b7183",
          8738 => x"2b077605",
          8739 => x"70338112",
          8740 => x"3371982b",
          8741 => x"71902b07",
          8742 => x"57535c52",
          8743 => x"59565280",
          8744 => x"7124839e",
          8745 => x"38841333",
          8746 => x"85143371",
          8747 => x"8b2b7183",
          8748 => x"2b077505",
          8749 => x"76882a52",
          8750 => x"54565774",
          8751 => x"86133473",
          8752 => x"81ff0654",
          8753 => x"73871334",
          8754 => x"84b9b808",
          8755 => x"70178412",
          8756 => x"33851333",
          8757 => x"71882b07",
          8758 => x"70882a5c",
          8759 => x"55595451",
          8760 => x"77841434",
          8761 => x"71851434",
          8762 => x"84b9b808",
          8763 => x"1652800b",
          8764 => x"86133480",
          8765 => x"0b871334",
          8766 => x"84b9b808",
          8767 => x"53748414",
          8768 => x"34738514",
          8769 => x"3484b9b8",
          8770 => x"08167033",
          8771 => x"81123371",
          8772 => x"882b0782",
          8773 => x"80800770",
          8774 => x"882a5858",
          8775 => x"52527472",
          8776 => x"34758113",
          8777 => x"34893d0d",
          8778 => x"04861233",
          8779 => x"87133371",
          8780 => x"8b2b7183",
          8781 => x"2b077511",
          8782 => x"84163385",
          8783 => x"17337188",
          8784 => x"2b077088",
          8785 => x"2a585854",
          8786 => x"51535858",
          8787 => x"71841234",
          8788 => x"72851234",
          8789 => x"84b9b808",
          8790 => x"70168411",
          8791 => x"33851233",
          8792 => x"718b2b71",
          8793 => x"832b0756",
          8794 => x"5a5a5272",
          8795 => x"05861233",
          8796 => x"87133371",
          8797 => x"882b0770",
          8798 => x"882a5255",
          8799 => x"59527786",
          8800 => x"13347287",
          8801 => x"133484b9",
          8802 => x"b8081570",
          8803 => x"33811233",
          8804 => x"71882b07",
          8805 => x"81ffff06",
          8806 => x"70882a5a",
          8807 => x"5a545276",
          8808 => x"72347781",
          8809 => x"133484b9",
          8810 => x"b8087017",
          8811 => x"70338112",
          8812 => x"33718b2b",
          8813 => x"71832b07",
          8814 => x"74057033",
          8815 => x"81123371",
          8816 => x"882b0770",
          8817 => x"832b8fff",
          8818 => x"f8067705",
          8819 => x"7b882a54",
          8820 => x"5253545c",
          8821 => x"5a575452",
          8822 => x"77821434",
          8823 => x"73831434",
          8824 => x"84b9b808",
          8825 => x"70177033",
          8826 => x"81123371",
          8827 => x"8b2b7183",
          8828 => x"2b077405",
          8829 => x"70338112",
          8830 => x"3371882b",
          8831 => x"0781ffff",
          8832 => x"0670882a",
          8833 => x"5f525355",
          8834 => x"5a575452",
          8835 => x"77733470",
          8836 => x"81143484",
          8837 => x"b9b80870",
          8838 => x"17821133",
          8839 => x"83123371",
          8840 => x"8b2b7183",
          8841 => x"2b077405",
          8842 => x"70338112",
          8843 => x"3371982b",
          8844 => x"71902b07",
          8845 => x"58535d52",
          8846 => x"5a575353",
          8847 => x"708025fc",
          8848 => x"e4387133",
          8849 => x"81133371",
          8850 => x"882b0782",
          8851 => x"80800770",
          8852 => x"882a5959",
          8853 => x"54767534",
          8854 => x"77811634",
          8855 => x"84b9b808",
          8856 => x"70177033",
          8857 => x"81123371",
          8858 => x"8b2b7183",
          8859 => x"2b077405",
          8860 => x"82143383",
          8861 => x"15337188",
          8862 => x"2b077088",
          8863 => x"2a575c5c",
          8864 => x"52585652",
          8865 => x"53728215",
          8866 => x"34758315",
          8867 => x"34893d0d",
          8868 => x"04f93d0d",
          8869 => x"7984b9b8",
          8870 => x"08585876",
          8871 => x"802e8f38",
          8872 => x"77802e86",
          8873 => x"387751fb",
          8874 => x"903f893d",
          8875 => x"0d0484ff",
          8876 => x"f40b84b9",
          8877 => x"b80ca080",
          8878 => x"0b84b9b4",
          8879 => x"23828080",
          8880 => x"53765284",
          8881 => x"fff451fe",
          8882 => x"d3b53f84",
          8883 => x"b9b80855",
          8884 => x"76753481",
          8885 => x"0b811634",
          8886 => x"84b9b808",
          8887 => x"54768415",
          8888 => x"34810b85",
          8889 => x"153484b9",
          8890 => x"b8085676",
          8891 => x"86173481",
          8892 => x"0b871734",
          8893 => x"84b9b808",
          8894 => x"84b9b422",
          8895 => x"ff05fe80",
          8896 => x"80077083",
          8897 => x"ffff0670",
          8898 => x"882a5851",
          8899 => x"55567488",
          8900 => x"17347389",
          8901 => x"173484b9",
          8902 => x"b4227010",
          8903 => x"101084b9",
          8904 => x"b80805f8",
          8905 => x"05555576",
          8906 => x"82153481",
          8907 => x"0b831534",
          8908 => x"feee39f7",
          8909 => x"3d0d7b52",
          8910 => x"80538151",
          8911 => x"8472278e",
          8912 => x"38fb1283",
          8913 => x"2a820570",
          8914 => x"83ffff06",
          8915 => x"51517083",
          8916 => x"ffff0684",
          8917 => x"b9b80884",
          8918 => x"11338512",
          8919 => x"3371882b",
          8920 => x"07705259",
          8921 => x"5a585581",
          8922 => x"ffff5475",
          8923 => x"802e80cc",
          8924 => x"38751010",
          8925 => x"10177033",
          8926 => x"81123371",
          8927 => x"882b0770",
          8928 => x"81ffff06",
          8929 => x"79317083",
          8930 => x"ffff0670",
          8931 => x"7a275653",
          8932 => x"5c5c5452",
          8933 => x"7274278a",
          8934 => x"3870802e",
          8935 => x"85387573",
          8936 => x"55588412",
          8937 => x"33851333",
          8938 => x"71882b07",
          8939 => x"575a75c1",
          8940 => x"387381ff",
          8941 => x"ff2e8538",
          8942 => x"77745456",
          8943 => x"8076832b",
          8944 => x"78117033",
          8945 => x"81123371",
          8946 => x"882b0770",
          8947 => x"81ffff06",
          8948 => x"56565d56",
          8949 => x"59597079",
          8950 => x"2e833881",
          8951 => x"59805174",
          8952 => x"7326828d",
          8953 => x"38785178",
          8954 => x"802e8285",
          8955 => x"3872752e",
          8956 => x"82883874",
          8957 => x"1670832b",
          8958 => x"78117482",
          8959 => x"80800770",
          8960 => x"882a5b5c",
          8961 => x"56565a76",
          8962 => x"74347881",
          8963 => x"153484b9",
          8964 => x"b8081576",
          8965 => x"882a5353",
          8966 => x"71821434",
          8967 => x"75831434",
          8968 => x"84b9b808",
          8969 => x"70197033",
          8970 => x"81123371",
          8971 => x"882b0770",
          8972 => x"832b8fff",
          8973 => x"f8067405",
          8974 => x"7e83ffff",
          8975 => x"0670882a",
          8976 => x"5c585357",
          8977 => x"59525275",
          8978 => x"82123472",
          8979 => x"81ff0653",
          8980 => x"72831234",
          8981 => x"84b9b808",
          8982 => x"18547574",
          8983 => x"34728115",
          8984 => x"3484b9b8",
          8985 => x"08701986",
          8986 => x"11338712",
          8987 => x"33718b2b",
          8988 => x"71832b07",
          8989 => x"7405585c",
          8990 => x"5c535775",
          8991 => x"84153472",
          8992 => x"85153484",
          8993 => x"b9b80870",
          8994 => x"16557805",
          8995 => x"86113387",
          8996 => x"12337188",
          8997 => x"2b077088",
          8998 => x"2a545458",
          8999 => x"59708615",
          9000 => x"34718715",
          9001 => x"3484b9b8",
          9002 => x"08701984",
          9003 => x"11338512",
          9004 => x"33718b2b",
          9005 => x"71832b07",
          9006 => x"7405585a",
          9007 => x"5c5a5275",
          9008 => x"86153472",
          9009 => x"87153484",
          9010 => x"b9b80870",
          9011 => x"16557805",
          9012 => x"84113385",
          9013 => x"12337188",
          9014 => x"2b077088",
          9015 => x"2a545c57",
          9016 => x"59708415",
          9017 => x"34798515",
          9018 => x"3484b9b8",
          9019 => x"08188405",
          9020 => x"517084b9",
          9021 => x"c80c8b3d",
          9022 => x"0d048614",
          9023 => x"33871533",
          9024 => x"718b2b71",
          9025 => x"832b0779",
          9026 => x"05841733",
          9027 => x"85183371",
          9028 => x"882b0770",
          9029 => x"882a5a5b",
          9030 => x"59535452",
          9031 => x"74841234",
          9032 => x"76851234",
          9033 => x"84b9b808",
          9034 => x"70198411",
          9035 => x"33851233",
          9036 => x"718b2b71",
          9037 => x"832b0774",
          9038 => x"05861433",
          9039 => x"87153371",
          9040 => x"882b0770",
          9041 => x"882a585d",
          9042 => x"5f52565b",
          9043 => x"57527086",
          9044 => x"1a347687",
          9045 => x"1a3484b9",
          9046 => x"b8081870",
          9047 => x"33811233",
          9048 => x"71882b07",
          9049 => x"81ffff06",
          9050 => x"70882a59",
          9051 => x"57545775",
          9052 => x"77347481",
          9053 => x"183484b9",
          9054 => x"b8081884",
          9055 => x"0551fef1",
          9056 => x"39f93d0d",
          9057 => x"7984b9b8",
          9058 => x"08585876",
          9059 => x"802ea038",
          9060 => x"7754778a",
          9061 => x"387384b9",
          9062 => x"c80c893d",
          9063 => x"0d047751",
          9064 => x"fb913f84",
          9065 => x"b9c80884",
          9066 => x"b9c80c89",
          9067 => x"3d0d0484",
          9068 => x"fff40b84",
          9069 => x"b9b80ca0",
          9070 => x"800b84b9",
          9071 => x"b4238280",
          9072 => x"80537652",
          9073 => x"84fff451",
          9074 => x"fecdb43f",
          9075 => x"84b9b808",
          9076 => x"55767534",
          9077 => x"810b8116",
          9078 => x"3484b9b8",
          9079 => x"08547684",
          9080 => x"1534810b",
          9081 => x"85153484",
          9082 => x"b9b80856",
          9083 => x"76861734",
          9084 => x"810b8717",
          9085 => x"3484b9b8",
          9086 => x"0884b9b4",
          9087 => x"22ff05fe",
          9088 => x"80800770",
          9089 => x"83ffff06",
          9090 => x"70882a58",
          9091 => x"51555674",
          9092 => x"88173473",
          9093 => x"89173484",
          9094 => x"b9b42270",
          9095 => x"10101084",
          9096 => x"b9b80805",
          9097 => x"f8055555",
          9098 => x"76821534",
          9099 => x"810b8315",
          9100 => x"34775477",
          9101 => x"802efedd",
          9102 => x"38fee339",
          9103 => x"ed3d0d65",
          9104 => x"67415f80",
          9105 => x"7084b9b8",
          9106 => x"08594541",
          9107 => x"76612e84",
          9108 => x"aa387e80",
          9109 => x"2e85af38",
          9110 => x"7f802e88",
          9111 => x"d7388154",
          9112 => x"8460278f",
          9113 => x"387ffb05",
          9114 => x"832a8205",
          9115 => x"7083ffff",
          9116 => x"06555873",
          9117 => x"83ffff06",
          9118 => x"7f783183",
          9119 => x"2a7083ff",
          9120 => x"ff067083",
          9121 => x"2b7a1170",
          9122 => x"33811233",
          9123 => x"71882b07",
          9124 => x"70753170",
          9125 => x"83ffff06",
          9126 => x"70101010",
          9127 => x"fc057383",
          9128 => x"2b611170",
          9129 => x"33811233",
          9130 => x"71882b07",
          9131 => x"70902b70",
          9132 => x"902c5342",
          9133 => x"45464453",
          9134 => x"5443445c",
          9135 => x"4859525e",
          9136 => x"5f42807a",
          9137 => x"2485fd38",
          9138 => x"82153383",
          9139 => x"16337188",
          9140 => x"2b077010",
          9141 => x"10101970",
          9142 => x"33811233",
          9143 => x"71982b71",
          9144 => x"902b0753",
          9145 => x"5c535656",
          9146 => x"56807424",
          9147 => x"85c9387a",
          9148 => x"622782f6",
          9149 => x"38631b58",
          9150 => x"77622e87",
          9151 => x"a2386080",
          9152 => x"2e85f938",
          9153 => x"601b5877",
          9154 => x"622587be",
          9155 => x"38631859",
          9156 => x"61792492",
          9157 => x"f738761e",
          9158 => x"70338112",
          9159 => x"33718b2b",
          9160 => x"71832b07",
          9161 => x"7a117033",
          9162 => x"81123371",
          9163 => x"982b7190",
          9164 => x"2b074743",
          9165 => x"59525357",
          9166 => x"5b588060",
          9167 => x"248cba38",
          9168 => x"761e8211",
          9169 => x"33831233",
          9170 => x"718b2b71",
          9171 => x"832b077a",
          9172 => x"11861133",
          9173 => x"87123371",
          9174 => x"8b2b7183",
          9175 => x"2b077e05",
          9176 => x"84143385",
          9177 => x"15337188",
          9178 => x"2b077088",
          9179 => x"2a595748",
          9180 => x"525b4158",
          9181 => x"535c5956",
          9182 => x"77841d34",
          9183 => x"79851d34",
          9184 => x"84b9b808",
          9185 => x"70178411",
          9186 => x"33851233",
          9187 => x"718b2b71",
          9188 => x"832b0774",
          9189 => x"05861433",
          9190 => x"87153371",
          9191 => x"882b0770",
          9192 => x"882a5f42",
          9193 => x"5e524057",
          9194 => x"41577786",
          9195 => x"16347b87",
          9196 => x"163484b9",
          9197 => x"b8081670",
          9198 => x"33811233",
          9199 => x"71882b07",
          9200 => x"81ffff06",
          9201 => x"70882a5a",
          9202 => x"5c5e5976",
          9203 => x"79347981",
          9204 => x"1a3484b9",
          9205 => x"b808701f",
          9206 => x"82113383",
          9207 => x"1233718b",
          9208 => x"2b71832b",
          9209 => x"07740573",
          9210 => x"33811533",
          9211 => x"71882b07",
          9212 => x"70882a41",
          9213 => x"5c455d5f",
          9214 => x"5a555579",
          9215 => x"79347581",
          9216 => x"1a3484b9",
          9217 => x"b808701f",
          9218 => x"70338112",
          9219 => x"33718b2b",
          9220 => x"71832b07",
          9221 => x"74058214",
          9222 => x"33831533",
          9223 => x"71882b07",
          9224 => x"70882a41",
          9225 => x"5c455d5f",
          9226 => x"5a555579",
          9227 => x"821a3475",
          9228 => x"831a3484",
          9229 => x"b9b80870",
          9230 => x"1f821133",
          9231 => x"83123371",
          9232 => x"882b0766",
          9233 => x"57625670",
          9234 => x"832b4252",
          9235 => x"5a5d7e05",
          9236 => x"840551fe",
          9237 => x"c4ec3f84",
          9238 => x"b9b8081e",
          9239 => x"84056165",
          9240 => x"051c7083",
          9241 => x"ffff065d",
          9242 => x"445f7a62",
          9243 => x"2681b638",
          9244 => x"7e547384",
          9245 => x"b9c80c95",
          9246 => x"3d0d0484",
          9247 => x"fff40b84",
          9248 => x"b9b80ca0",
          9249 => x"800b84b9",
          9250 => x"b4238280",
          9251 => x"80536052",
          9252 => x"84fff451",
          9253 => x"fec7e83f",
          9254 => x"84b9b808",
          9255 => x"5e607e34",
          9256 => x"810b811f",
          9257 => x"3484b9b8",
          9258 => x"085d6084",
          9259 => x"1e34810b",
          9260 => x"851e3484",
          9261 => x"b9b8085c",
          9262 => x"60861d34",
          9263 => x"810b871d",
          9264 => x"3484b9b8",
          9265 => x"0884b9b4",
          9266 => x"22ff05fe",
          9267 => x"80800770",
          9268 => x"83ffff06",
          9269 => x"70882a5c",
          9270 => x"5a5b5778",
          9271 => x"88183477",
          9272 => x"89183484",
          9273 => x"b9b42270",
          9274 => x"10101084",
          9275 => x"b9b80805",
          9276 => x"f8055556",
          9277 => x"60821534",
          9278 => x"810b8315",
          9279 => x"3484b9b8",
          9280 => x"08577efa",
          9281 => x"d3387680",
          9282 => x"2e828c38",
          9283 => x"7e547f80",
          9284 => x"2efedf38",
          9285 => x"7f51f49b",
          9286 => x"3f84b9c8",
          9287 => x"0884b9c8",
          9288 => x"0c953d0d",
          9289 => x"04611c84",
          9290 => x"b9b80871",
          9291 => x"832b7111",
          9292 => x"5e447f05",
          9293 => x"70338112",
          9294 => x"3371882b",
          9295 => x"0781ffff",
          9296 => x"0670882a",
          9297 => x"48445b5e",
          9298 => x"40637b34",
          9299 => x"60811c34",
          9300 => x"6184b9b8",
          9301 => x"08057c88",
          9302 => x"2a575875",
          9303 => x"8219347b",
          9304 => x"83193484",
          9305 => x"b9b80870",
          9306 => x"1f703381",
          9307 => x"12337188",
          9308 => x"2b077083",
          9309 => x"2b8ffff8",
          9310 => x"06740564",
          9311 => x"83ffff06",
          9312 => x"70882a4a",
          9313 => x"5c47575e",
          9314 => x"5b5d6363",
          9315 => x"82053476",
          9316 => x"81ff0641",
          9317 => x"60638305",
          9318 => x"3484b9b8",
          9319 => x"081e5b63",
          9320 => x"7b346081",
          9321 => x"1c346184",
          9322 => x"b9b80805",
          9323 => x"840551ed",
          9324 => x"883f7e54",
          9325 => x"fdbc397b",
          9326 => x"75317083",
          9327 => x"ffff0642",
          9328 => x"54faac39",
          9329 => x"7781ffff",
          9330 => x"06763170",
          9331 => x"83ffff06",
          9332 => x"82173383",
          9333 => x"18337188",
          9334 => x"2b077010",
          9335 => x"10101b70",
          9336 => x"33811233",
          9337 => x"71982b71",
          9338 => x"902b0753",
          9339 => x"5e535458",
          9340 => x"58455473",
          9341 => x"8025f9f7",
          9342 => x"38ffbc39",
          9343 => x"617824fa",
          9344 => x"8338807a",
          9345 => x"248b8f38",
          9346 => x"7783ffff",
          9347 => x"065b617b",
          9348 => x"27fcdd38",
          9349 => x"fe8f3984",
          9350 => x"fff40b84",
          9351 => x"b9b80ca0",
          9352 => x"800b84b9",
          9353 => x"b4238280",
          9354 => x"80537e52",
          9355 => x"84fff451",
          9356 => x"fec4cc3f",
          9357 => x"84b9b808",
          9358 => x"5a7e7a34",
          9359 => x"810b811b",
          9360 => x"3484b9b8",
          9361 => x"08597e84",
          9362 => x"1a34810b",
          9363 => x"851a3484",
          9364 => x"b9b80858",
          9365 => x"7e861934",
          9366 => x"810b8719",
          9367 => x"3484b9b8",
          9368 => x"0884b9b4",
          9369 => x"22ff05fe",
          9370 => x"80800770",
          9371 => x"83ffff06",
          9372 => x"70882a58",
          9373 => x"56574474",
          9374 => x"64880534",
          9375 => x"73648905",
          9376 => x"3484b9b4",
          9377 => x"22701010",
          9378 => x"1084b9b8",
          9379 => x"0805f805",
          9380 => x"42437e61",
          9381 => x"82053481",
          9382 => x"61830534",
          9383 => x"fcee3980",
          9384 => x"7a2483de",
          9385 => x"386183ff",
          9386 => x"ff065b61",
          9387 => x"7b27fbc0",
          9388 => x"38fcf239",
          9389 => x"76802e82",
          9390 => x"bd387e51",
          9391 => x"eafb3f7f",
          9392 => x"547384b9",
          9393 => x"c80c953d",
          9394 => x"0d04761e",
          9395 => x"82113383",
          9396 => x"1233718b",
          9397 => x"2b71832b",
          9398 => x"077a1186",
          9399 => x"11338712",
          9400 => x"33718b2b",
          9401 => x"71832b07",
          9402 => x"7e058414",
          9403 => x"33851533",
          9404 => x"71882b07",
          9405 => x"70882a43",
          9406 => x"4445565b",
          9407 => x"4658535c",
          9408 => x"45567864",
          9409 => x"8405347a",
          9410 => x"64850534",
          9411 => x"84b9b808",
          9412 => x"70178411",
          9413 => x"33851233",
          9414 => x"718b2b71",
          9415 => x"832b0774",
          9416 => x"05861433",
          9417 => x"87153371",
          9418 => x"882b0770",
          9419 => x"882a5b41",
          9420 => x"42485d59",
          9421 => x"5d417364",
          9422 => x"8605347a",
          9423 => x"64870534",
          9424 => x"84b9b808",
          9425 => x"16703381",
          9426 => x"12337188",
          9427 => x"2b0781ff",
          9428 => x"ff067088",
          9429 => x"2a5f5c5a",
          9430 => x"5d7b7d34",
          9431 => x"79811e34",
          9432 => x"84b9b808",
          9433 => x"701f8211",
          9434 => x"33831233",
          9435 => x"718b2b71",
          9436 => x"832b0774",
          9437 => x"05733381",
          9438 => x"15337188",
          9439 => x"2b077088",
          9440 => x"2a5e5c5e",
          9441 => x"40435745",
          9442 => x"54767c34",
          9443 => x"75811d34",
          9444 => x"84b9b808",
          9445 => x"701f7033",
          9446 => x"81123371",
          9447 => x"8b2b7183",
          9448 => x"2b077405",
          9449 => x"82143383",
          9450 => x"15337188",
          9451 => x"2b077088",
          9452 => x"2a404740",
          9453 => x"5b405c55",
          9454 => x"55788218",
          9455 => x"34608318",
          9456 => x"3484b9b8",
          9457 => x"08701f82",
          9458 => x"11338312",
          9459 => x"3371882b",
          9460 => x"07665762",
          9461 => x"5670832b",
          9462 => x"4252585d",
          9463 => x"7e058405",
          9464 => x"51febdde",
          9465 => x"3f84b9b8",
          9466 => x"081e8405",
          9467 => x"7883ffff",
          9468 => x"065c5ffc",
          9469 => x"993984ff",
          9470 => x"f40b84b9",
          9471 => x"b80ca080",
          9472 => x"0b84b9b4",
          9473 => x"23828080",
          9474 => x"537f5284",
          9475 => x"fff451fe",
          9476 => x"c0ed3f84",
          9477 => x"b9b80856",
          9478 => x"7f763481",
          9479 => x"0b811734",
          9480 => x"84b9b808",
          9481 => x"557f8416",
          9482 => x"34810b85",
          9483 => x"163484b9",
          9484 => x"b808547f",
          9485 => x"86153481",
          9486 => x"0b871534",
          9487 => x"84b9b808",
          9488 => x"84b9b422",
          9489 => x"ff05fe80",
          9490 => x"80077083",
          9491 => x"ffff0670",
          9492 => x"882a4543",
          9493 => x"445e6188",
          9494 => x"1f346089",
          9495 => x"1f3484b9",
          9496 => x"b4227010",
          9497 => x"101084b9",
          9498 => x"b80805f8",
          9499 => x"055c5d7f",
          9500 => x"821c3481",
          9501 => x"0b831c34",
          9502 => x"7e51e7bd",
          9503 => x"3f7f54fc",
          9504 => x"c0398619",
          9505 => x"33871a33",
          9506 => x"718b2b71",
          9507 => x"832b0779",
          9508 => x"05841c33",
          9509 => x"851d3371",
          9510 => x"882b0770",
          9511 => x"882a5c48",
          9512 => x"5e435955",
          9513 => x"76618405",
          9514 => x"34636185",
          9515 => x"053484b9",
          9516 => x"b808701e",
          9517 => x"84113385",
          9518 => x"1233718b",
          9519 => x"2b71832b",
          9520 => x"07740586",
          9521 => x"14338715",
          9522 => x"3371882b",
          9523 => x"0770882a",
          9524 => x"415f4848",
          9525 => x"59565940",
          9526 => x"79648605",
          9527 => x"34786487",
          9528 => x"053484b9",
          9529 => x"b8081d70",
          9530 => x"33811233",
          9531 => x"71882b07",
          9532 => x"81ffff06",
          9533 => x"70882a59",
          9534 => x"42585875",
          9535 => x"78347f81",
          9536 => x"193484b9",
          9537 => x"b808701f",
          9538 => x"70338112",
          9539 => x"33718b2b",
          9540 => x"71832b07",
          9541 => x"74057033",
          9542 => x"81123371",
          9543 => x"882b0770",
          9544 => x"832b8fff",
          9545 => x"f8067705",
          9546 => x"63882a48",
          9547 => x"5d5d5a5d",
          9548 => x"405d4441",
          9549 => x"7f821734",
          9550 => x"7b831734",
          9551 => x"84b9b808",
          9552 => x"701f7033",
          9553 => x"81123371",
          9554 => x"8b2b7183",
          9555 => x"2b077405",
          9556 => x"70338112",
          9557 => x"3371882b",
          9558 => x"0781ffff",
          9559 => x"0670882a",
          9560 => x"485d5e5e",
          9561 => x"465a415b",
          9562 => x"60603476",
          9563 => x"60810534",
          9564 => x"6183ffff",
          9565 => x"065bfab3",
          9566 => x"39861533",
          9567 => x"87163371",
          9568 => x"8b2b7183",
          9569 => x"2b077905",
          9570 => x"84183385",
          9571 => x"19337188",
          9572 => x"2b077088",
          9573 => x"2a5e5e5a",
          9574 => x"52415d78",
          9575 => x"841e3479",
          9576 => x"851e3484",
          9577 => x"b9b80870",
          9578 => x"19841133",
          9579 => x"85123371",
          9580 => x"8b2b7183",
          9581 => x"2b077405",
          9582 => x"86143387",
          9583 => x"15337188",
          9584 => x"2b077088",
          9585 => x"2a44565e",
          9586 => x"525a4255",
          9587 => x"567c6086",
          9588 => x"05347560",
          9589 => x"87053484",
          9590 => x"b9b80818",
          9591 => x"70338112",
          9592 => x"3371882b",
          9593 => x"0781ffff",
          9594 => x"0670882a",
          9595 => x"5b5b5855",
          9596 => x"77753478",
          9597 => x"81163484",
          9598 => x"b9b80870",
          9599 => x"1f703381",
          9600 => x"1233718b",
          9601 => x"2b71832b",
          9602 => x"07740570",
          9603 => x"33811233",
          9604 => x"71882b07",
          9605 => x"70832b8f",
          9606 => x"fff80677",
          9607 => x"0563882a",
          9608 => x"56545f5f",
          9609 => x"5859425e",
          9610 => x"557f8217",
          9611 => x"347b8317",
          9612 => x"3484b9b8",
          9613 => x"08701f70",
          9614 => x"33811233",
          9615 => x"718b2b71",
          9616 => x"832b0774",
          9617 => x"05703381",
          9618 => x"12337188",
          9619 => x"2b0781ff",
          9620 => x"ff067088",
          9621 => x"2a5d545e",
          9622 => x"585b595d",
          9623 => x"55757c34",
          9624 => x"76811d34",
          9625 => x"84b9b808",
          9626 => x"701f8211",
          9627 => x"33831233",
          9628 => x"718b2b71",
          9629 => x"832b0774",
          9630 => x"11861133",
          9631 => x"87123371",
          9632 => x"8b2b7183",
          9633 => x"2b077805",
          9634 => x"84143385",
          9635 => x"15337188",
          9636 => x"2b077088",
          9637 => x"2a595749",
          9638 => x"525c4259",
          9639 => x"535d5a57",
          9640 => x"5777841d",
          9641 => x"3479851d",
          9642 => x"3484b9b8",
          9643 => x"08701784",
          9644 => x"11338512",
          9645 => x"33718b2b",
          9646 => x"71832b07",
          9647 => x"74058614",
          9648 => x"33871533",
          9649 => x"71882b07",
          9650 => x"70882a5f",
          9651 => x"425e5240",
          9652 => x"57415777",
          9653 => x"8616347b",
          9654 => x"87163484",
          9655 => x"b9b80816",
          9656 => x"70338112",
          9657 => x"3371882b",
          9658 => x"0781ffff",
          9659 => x"0670882a",
          9660 => x"5a5c5e59",
          9661 => x"76793479",
          9662 => x"811a3484",
          9663 => x"b9b80870",
          9664 => x"1f821133",
          9665 => x"83123371",
          9666 => x"8b2b7183",
          9667 => x"2b077405",
          9668 => x"73338115",
          9669 => x"3371882b",
          9670 => x"0770882a",
          9671 => x"415c455d",
          9672 => x"5f5a5555",
          9673 => x"79793475",
          9674 => x"811a3484",
          9675 => x"b9b80870",
          9676 => x"1f703381",
          9677 => x"1233718b",
          9678 => x"2b71832b",
          9679 => x"07740582",
          9680 => x"14338315",
          9681 => x"3371882b",
          9682 => x"0770882a",
          9683 => x"415c455d",
          9684 => x"5f5a5555",
          9685 => x"79821a34",
          9686 => x"75831a34",
          9687 => x"84b9b808",
          9688 => x"701f8211",
          9689 => x"33831233",
          9690 => x"71882b07",
          9691 => x"66576256",
          9692 => x"70832b42",
          9693 => x"525a5d7e",
          9694 => x"05840551",
          9695 => x"feb6c33f",
          9696 => x"84b9b808",
          9697 => x"1e840561",
          9698 => x"65051c70",
          9699 => x"83ffff06",
          9700 => x"5d445ff1",
          9701 => x"d5398619",
          9702 => x"33871a33",
          9703 => x"718b2b71",
          9704 => x"832b0779",
          9705 => x"05841c33",
          9706 => x"851d3371",
          9707 => x"882b0770",
          9708 => x"882a4048",
          9709 => x"5d434155",
          9710 => x"7a618405",
          9711 => x"34636185",
          9712 => x"053484b9",
          9713 => x"b808701e",
          9714 => x"84113385",
          9715 => x"1233718b",
          9716 => x"2b71832b",
          9717 => x"07740586",
          9718 => x"14338715",
          9719 => x"3371882b",
          9720 => x"0770882a",
          9721 => x"5b415f48",
          9722 => x"5c594156",
          9723 => x"73648605",
          9724 => x"347a6487",
          9725 => x"053484b9",
          9726 => x"b8081d70",
          9727 => x"33811233",
          9728 => x"71882b07",
          9729 => x"81ffff06",
          9730 => x"70882a5c",
          9731 => x"5f425578",
          9732 => x"75347c81",
          9733 => x"163484b9",
          9734 => x"b808701f",
          9735 => x"70338112",
          9736 => x"33718b2b",
          9737 => x"71832b07",
          9738 => x"74057033",
          9739 => x"81123371",
          9740 => x"882b0770",
          9741 => x"832b8fff",
          9742 => x"f8067705",
          9743 => x"63882a5d",
          9744 => x"445c4958",
          9745 => x"5e455840",
          9746 => x"74821e34",
          9747 => x"7b831e34",
          9748 => x"84b9b808",
          9749 => x"701f7033",
          9750 => x"81123371",
          9751 => x"8b2b7183",
          9752 => x"2b077405",
          9753 => x"70338112",
          9754 => x"3371882b",
          9755 => x"0781ffff",
          9756 => x"0670882a",
          9757 => x"475f4958",
          9758 => x"46595e5b",
          9759 => x"7f7d3478",
          9760 => x"811e3477",
          9761 => x"83ffff06",
          9762 => x"5bf38339",
          9763 => x"7e605254",
          9764 => x"e5a13f84",
          9765 => x"b9c8085f",
          9766 => x"84b9c808",
          9767 => x"802e9338",
          9768 => x"62537352",
          9769 => x"84b9c808",
          9770 => x"51feb5be",
          9771 => x"3f7351df",
          9772 => x"883f615b",
          9773 => x"617b27ef",
          9774 => x"b738f0e9",
          9775 => x"39f93d0d",
          9776 => x"7a7a2984",
          9777 => x"b9b80858",
          9778 => x"5876802e",
          9779 => x"b7387754",
          9780 => x"778a3873",
          9781 => x"84b9c80c",
          9782 => x"893d0d04",
          9783 => x"7751e4d3",
          9784 => x"3f84b9c8",
          9785 => x"085484b9",
          9786 => x"c808802e",
          9787 => x"e6387753",
          9788 => x"805284b9",
          9789 => x"c80851fe",
          9790 => x"b7853f73",
          9791 => x"84b9c80c",
          9792 => x"893d0d04",
          9793 => x"84fff40b",
          9794 => x"84b9b80c",
          9795 => x"a0800b84",
          9796 => x"b9b42382",
          9797 => x"80805376",
          9798 => x"5284fff4",
          9799 => x"51feb6df",
          9800 => x"3f84b9b8",
          9801 => x"08557675",
          9802 => x"34810b81",
          9803 => x"163484b9",
          9804 => x"b8085476",
          9805 => x"84153481",
          9806 => x"0b851534",
          9807 => x"84b9b808",
          9808 => x"56768617",
          9809 => x"34810b87",
          9810 => x"173484b9",
          9811 => x"b80884b9",
          9812 => x"b422ff05",
          9813 => x"fe808007",
          9814 => x"7083ffff",
          9815 => x"0670882a",
          9816 => x"58515556",
          9817 => x"74881734",
          9818 => x"73891734",
          9819 => x"84b9b422",
          9820 => x"70101010",
          9821 => x"84b9b808",
          9822 => x"05f80555",
          9823 => x"55768215",
          9824 => x"34810b83",
          9825 => x"15347754",
          9826 => x"77802efe",
          9827 => x"c638fecc",
          9828 => x"39ff3d0d",
          9829 => x"028f0533",
          9830 => x"51815270",
          9831 => x"72268738",
          9832 => x"84b9c411",
          9833 => x"33527184",
          9834 => x"b9c80c83",
          9835 => x"3d0d04fe",
          9836 => x"3d0d0293",
          9837 => x"05335283",
          9838 => x"53718126",
          9839 => x"9d387151",
          9840 => x"d4bb3f84",
          9841 => x"b9c80881",
          9842 => x"ff065372",
          9843 => x"87387284",
          9844 => x"b9c41334",
          9845 => x"84b9c412",
          9846 => x"33537284",
          9847 => x"b9c80c84",
          9848 => x"3d0d04f7",
          9849 => x"3d0d7c7e",
          9850 => x"60028c05",
          9851 => x"af05335a",
          9852 => x"5c575981",
          9853 => x"54767426",
          9854 => x"873884b9",
          9855 => x"c4173354",
          9856 => x"73810654",
          9857 => x"835573bd",
          9858 => x"38735885",
          9859 => x"0b87c098",
          9860 => x"8c0c7853",
          9861 => x"75527651",
          9862 => x"d5ca3f84",
          9863 => x"b9c80881",
          9864 => x"ff065574",
          9865 => x"802ea738",
          9866 => x"87c0988c",
          9867 => x"085473e2",
          9868 => x"38797826",
          9869 => x"d63874fc",
          9870 => x"80800654",
          9871 => x"73802e83",
          9872 => x"38815473",
          9873 => x"557484b9",
          9874 => x"c80c8b3d",
          9875 => x"0d048480",
          9876 => x"16811970",
          9877 => x"81ff065a",
          9878 => x"55567978",
          9879 => x"26ffac38",
          9880 => x"d539f73d",
          9881 => x"0d7c7e60",
          9882 => x"028c05af",
          9883 => x"05335a5c",
          9884 => x"57598154",
          9885 => x"76742687",
          9886 => x"3884b9c4",
          9887 => x"17335473",
          9888 => x"81065483",
          9889 => x"5573bd38",
          9890 => x"7358850b",
          9891 => x"87c0988c",
          9892 => x"0c785375",
          9893 => x"527651d7",
          9894 => x"8e3f84b9",
          9895 => x"c80881ff",
          9896 => x"06557480",
          9897 => x"2ea73887",
          9898 => x"c0988c08",
          9899 => x"5473e238",
          9900 => x"797826d6",
          9901 => x"3874fc80",
          9902 => x"80065473",
          9903 => x"802e8338",
          9904 => x"81547355",
          9905 => x"7484b9c8",
          9906 => x"0c8b3d0d",
          9907 => x"04848016",
          9908 => x"81197081",
          9909 => x"ff065a55",
          9910 => x"56797826",
          9911 => x"ffac38d5",
          9912 => x"39fc3d0d",
          9913 => x"78028405",
          9914 => x"9b053302",
          9915 => x"88059f05",
          9916 => x"33535355",
          9917 => x"81537173",
          9918 => x"26873884",
          9919 => x"b9c41233",
          9920 => x"53728106",
          9921 => x"54835373",
          9922 => x"9b38850b",
          9923 => x"87c0988c",
          9924 => x"0c815370",
          9925 => x"732e9638",
          9926 => x"727125ad",
          9927 => x"3870832e",
          9928 => x"9a388453",
          9929 => x"7284b9c8",
          9930 => x"0c863d0d",
          9931 => x"0488800a",
          9932 => x"750c7384",
          9933 => x"b9c80c86",
          9934 => x"3d0d0481",
          9935 => x"80750c80",
          9936 => x"0b84b9c8",
          9937 => x"0c863d0d",
          9938 => x"0471842b",
          9939 => x"87c0928c",
          9940 => x"11535470",
          9941 => x"cd387108",
          9942 => x"70812a81",
          9943 => x"06515170",
          9944 => x"802e8a38",
          9945 => x"87c0988c",
          9946 => x"085574ea",
          9947 => x"3887c098",
          9948 => x"8c085170",
          9949 => x"ca388172",
          9950 => x"0c87c092",
          9951 => x"8c145271",
          9952 => x"08820654",
          9953 => x"73802eff",
          9954 => x"9b387108",
          9955 => x"82065473",
          9956 => x"ee38ff90",
          9957 => x"39f63d0d",
          9958 => x"7c58800b",
          9959 => x"83193371",
          9960 => x"5b565774",
          9961 => x"772e0981",
          9962 => x"06a83877",
          9963 => x"33567583",
          9964 => x"2e818738",
          9965 => x"80538052",
          9966 => x"81183351",
          9967 => x"fea33f84",
          9968 => x"b9c80880",
          9969 => x"2e833881",
          9970 => x"597884b9",
          9971 => x"c80c8c3d",
          9972 => x"0d048154",
          9973 => x"b4180853",
          9974 => x"b8187053",
          9975 => x"81193352",
          9976 => x"5afcff3f",
          9977 => x"815984b9",
          9978 => x"c808772e",
          9979 => x"098106d9",
          9980 => x"3884b9c8",
          9981 => x"08831934",
          9982 => x"b4180870",
          9983 => x"a81a0831",
          9984 => x"a01a0884",
          9985 => x"b9c8085c",
          9986 => x"58565b74",
          9987 => x"7627ff9b",
          9988 => x"38821833",
          9989 => x"5574822e",
          9990 => x"098106ff",
          9991 => x"8e388154",
          9992 => x"751b5379",
          9993 => x"52811833",
          9994 => x"51fcb73f",
          9995 => x"76783357",
          9996 => x"5975832e",
          9997 => x"098106fe",
          9998 => x"fb388418",
          9999 => x"33577681",
         10000 => x"2e098106",
         10001 => x"feee38b8",
         10002 => x"185a8480",
         10003 => x"7a565780",
         10004 => x"75708105",
         10005 => x"5734ff17",
         10006 => x"5776f438",
         10007 => x"80d50b84",
         10008 => x"b61934ff",
         10009 => x"aa0b84b7",
         10010 => x"193480d2",
         10011 => x"7a3480d2",
         10012 => x"0bb91934",
         10013 => x"80e10bba",
         10014 => x"193480c1",
         10015 => x"0bbb1934",
         10016 => x"80f20b84",
         10017 => x"9c193480",
         10018 => x"f20b849d",
         10019 => x"193480c1",
         10020 => x"0b849e19",
         10021 => x"3480e10b",
         10022 => x"849f1934",
         10023 => x"94180855",
         10024 => x"7484a019",
         10025 => x"3474882a",
         10026 => x"5b7a84a1",
         10027 => x"19347490",
         10028 => x"2a567584",
         10029 => x"a2193474",
         10030 => x"982a5b7a",
         10031 => x"84a31934",
         10032 => x"9018085b",
         10033 => x"7a84a419",
         10034 => x"347a882a",
         10035 => x"557484a5",
         10036 => x"19347a90",
         10037 => x"2a567584",
         10038 => x"a619347a",
         10039 => x"982a5574",
         10040 => x"84a71934",
         10041 => x"a4180881",
         10042 => x"0570b41a",
         10043 => x"0c5b8154",
         10044 => x"7a537952",
         10045 => x"81183351",
         10046 => x"fae83f76",
         10047 => x"84193480",
         10048 => x"53805281",
         10049 => x"183351fb",
         10050 => x"d83f84b9",
         10051 => x"c808802e",
         10052 => x"fdb738fd",
         10053 => x"b239f33d",
         10054 => x"0d606070",
         10055 => x"08595656",
         10056 => x"81762788",
         10057 => x"389c1708",
         10058 => x"76268c38",
         10059 => x"81587784",
         10060 => x"b9c80c8f",
         10061 => x"3d0d04ff",
         10062 => x"77335658",
         10063 => x"74822e81",
         10064 => x"cc387482",
         10065 => x"2482a538",
         10066 => x"74812e09",
         10067 => x"8106dd38",
         10068 => x"75812a16",
         10069 => x"70892aa8",
         10070 => x"1908055a",
         10071 => x"5a805bb4",
         10072 => x"1708792e",
         10073 => x"b0388317",
         10074 => x"335c7b7b",
         10075 => x"2e098106",
         10076 => x"83de3881",
         10077 => x"547853b8",
         10078 => x"17528117",
         10079 => x"3351f8e3",
         10080 => x"3f84b9c8",
         10081 => x"08802e85",
         10082 => x"38ff5981",
         10083 => x"5b78b418",
         10084 => x"0c7aff9a",
         10085 => x"387983ff",
         10086 => x"0617b811",
         10087 => x"33811c70",
         10088 => x"892aa81b",
         10089 => x"0805535d",
         10090 => x"5d59b417",
         10091 => x"08792eb5",
         10092 => x"38800b83",
         10093 => x"1833715c",
         10094 => x"565d747d",
         10095 => x"2e098106",
         10096 => x"84b53881",
         10097 => x"547853b8",
         10098 => x"17528117",
         10099 => x"3351f893",
         10100 => x"3f84b9c8",
         10101 => x"08802e85",
         10102 => x"38ff5981",
         10103 => x"5a78b418",
         10104 => x"0c79feca",
         10105 => x"387a83ff",
         10106 => x"0617b811",
         10107 => x"3370882b",
         10108 => x"7e077881",
         10109 => x"0671842a",
         10110 => x"535d5959",
         10111 => x"5d79feae",
         10112 => x"38769fff",
         10113 => x"0684b9c8",
         10114 => x"0c8f3d0d",
         10115 => x"0475882a",
         10116 => x"a8180805",
         10117 => x"59b41708",
         10118 => x"792eb538",
         10119 => x"800b8318",
         10120 => x"33715c5d",
         10121 => x"5b7b7b2e",
         10122 => x"09810681",
         10123 => x"c2388154",
         10124 => x"7853b817",
         10125 => x"52811733",
         10126 => x"51f7a83f",
         10127 => x"84b9c808",
         10128 => x"802e8538",
         10129 => x"ff59815a",
         10130 => x"78b4180c",
         10131 => x"79fddf38",
         10132 => x"751083fe",
         10133 => x"067705b8",
         10134 => x"05811133",
         10135 => x"71337188",
         10136 => x"2b0784b9",
         10137 => x"c80c575b",
         10138 => x"8f3d0d04",
         10139 => x"74832e09",
         10140 => x"8106fdb8",
         10141 => x"3875872a",
         10142 => x"a8180805",
         10143 => x"59b41708",
         10144 => x"792eb538",
         10145 => x"800b8318",
         10146 => x"33715c5e",
         10147 => x"5b7c7b2e",
         10148 => x"09810682",
         10149 => x"81388154",
         10150 => x"7853b817",
         10151 => x"52811733",
         10152 => x"51f6c03f",
         10153 => x"84b9c808",
         10154 => x"802e8538",
         10155 => x"ff59815a",
         10156 => x"78b4180c",
         10157 => x"79fcf738",
         10158 => x"75822b83",
         10159 => x"fc067705",
         10160 => x"b8058311",
         10161 => x"33821233",
         10162 => x"71902b71",
         10163 => x"882b0781",
         10164 => x"14337072",
         10165 => x"07882b75",
         10166 => x"337180ff",
         10167 => x"fffe8006",
         10168 => x"0784b9c8",
         10169 => x"0c415c5e",
         10170 => x"595a568f",
         10171 => x"3d0d0481",
         10172 => x"54b41708",
         10173 => x"53b81770",
         10174 => x"53811833",
         10175 => x"525cf6e2",
         10176 => x"3f815a84",
         10177 => x"b9c8087b",
         10178 => x"2e098106",
         10179 => x"febe3884",
         10180 => x"b9c80883",
         10181 => x"1834b417",
         10182 => x"08a81808",
         10183 => x"3184b9c8",
         10184 => x"085b5e7d",
         10185 => x"a0180827",
         10186 => x"fe843882",
         10187 => x"17335574",
         10188 => x"822e0981",
         10189 => x"06fdf738",
         10190 => x"8154b417",
         10191 => x"08a01808",
         10192 => x"05537b52",
         10193 => x"81173351",
         10194 => x"f6983f7a",
         10195 => x"5afddf39",
         10196 => x"8154b417",
         10197 => x"0853b817",
         10198 => x"70538118",
         10199 => x"33525cf6",
         10200 => x"813f84b9",
         10201 => x"c8087b2e",
         10202 => x"09810682",
         10203 => x"813884b9",
         10204 => x"c8088318",
         10205 => x"34b41708",
         10206 => x"a8180831",
         10207 => x"5d7ca018",
         10208 => x"08278b38",
         10209 => x"8217335e",
         10210 => x"7d822e81",
         10211 => x"cb3884b9",
         10212 => x"c8085bfb",
         10213 => x"de398154",
         10214 => x"b4170853",
         10215 => x"b8177053",
         10216 => x"81183352",
         10217 => x"5cf5bb3f",
         10218 => x"815a84b9",
         10219 => x"c8087b2e",
         10220 => x"098106fd",
         10221 => x"ff3884b9",
         10222 => x"c8088318",
         10223 => x"34b41708",
         10224 => x"a8180831",
         10225 => x"84b9c808",
         10226 => x"5b5e7da0",
         10227 => x"180827fd",
         10228 => x"c5388217",
         10229 => x"33557482",
         10230 => x"2e098106",
         10231 => x"fdb83881",
         10232 => x"54b41708",
         10233 => x"a0180805",
         10234 => x"537b5281",
         10235 => x"173351f4",
         10236 => x"f13f7a5a",
         10237 => x"fda03981",
         10238 => x"54b41708",
         10239 => x"53b81770",
         10240 => x"53811833",
         10241 => x"525ef4da",
         10242 => x"3f815a84",
         10243 => x"b9c8087d",
         10244 => x"2e098106",
         10245 => x"fbcb3884",
         10246 => x"b9c80883",
         10247 => x"1834b417",
         10248 => x"08a81808",
         10249 => x"3184b9c8",
         10250 => x"085b5574",
         10251 => x"a0180827",
         10252 => x"fb913882",
         10253 => x"17335574",
         10254 => x"822e0981",
         10255 => x"06fb8438",
         10256 => x"8154b417",
         10257 => x"08a01808",
         10258 => x"05537d52",
         10259 => x"81173351",
         10260 => x"f4903f7c",
         10261 => x"5afaec39",
         10262 => x"8154b417",
         10263 => x"08a01808",
         10264 => x"05537b52",
         10265 => x"81173351",
         10266 => x"f3f83ffa",
         10267 => x"8639815b",
         10268 => x"7af9bb38",
         10269 => x"fa9f39f2",
         10270 => x"3d0d6062",
         10271 => x"645d5759",
         10272 => x"82588176",
         10273 => x"279c3875",
         10274 => x"9c1a0827",
         10275 => x"95387833",
         10276 => x"5574782e",
         10277 => x"96387478",
         10278 => x"24818038",
         10279 => x"74812e82",
         10280 => x"8a387784",
         10281 => x"b9c80c90",
         10282 => x"3d0d0475",
         10283 => x"882aa81a",
         10284 => x"08055880",
         10285 => x"0bb41a08",
         10286 => x"585c7678",
         10287 => x"2e86b638",
         10288 => x"8319337c",
         10289 => x"5b5d7c7c",
         10290 => x"2e098106",
         10291 => x"83fa3881",
         10292 => x"547753b8",
         10293 => x"19528119",
         10294 => x"3351f287",
         10295 => x"3f84b9c8",
         10296 => x"08802e85",
         10297 => x"38ff5881",
         10298 => x"5a77b41a",
         10299 => x"0c795879",
         10300 => x"ffb03875",
         10301 => x"1083fe06",
         10302 => x"79057b83",
         10303 => x"ffff0658",
         10304 => x"5e76b81f",
         10305 => x"3476882a",
         10306 => x"5a79b91f",
         10307 => x"34810b83",
         10308 => x"1a347784",
         10309 => x"b9c80c90",
         10310 => x"3d0d0474",
         10311 => x"832e0981",
         10312 => x"06feff38",
         10313 => x"75872aa8",
         10314 => x"1a080558",
         10315 => x"800bb41a",
         10316 => x"08585c76",
         10317 => x"782e85e1",
         10318 => x"38831933",
         10319 => x"7c5b5d7c",
         10320 => x"7c2e0981",
         10321 => x"0684bd38",
         10322 => x"81547753",
         10323 => x"b8195281",
         10324 => x"193351f1",
         10325 => x"8e3f84b9",
         10326 => x"c808802e",
         10327 => x"8538ff58",
         10328 => x"815a77b4",
         10329 => x"1a0c7958",
         10330 => x"79feb738",
         10331 => x"75822b83",
         10332 => x"fc067905",
         10333 => x"b8118311",
         10334 => x"3370982b",
         10335 => x"8f0a067e",
         10336 => x"f00a0607",
         10337 => x"41575e5c",
         10338 => x"7d7d347d",
         10339 => x"882a5675",
         10340 => x"b91d347d",
         10341 => x"902a5a79",
         10342 => x"ba1d347d",
         10343 => x"982a5b7a",
         10344 => x"bb1d3481",
         10345 => x"0b831a34",
         10346 => x"fee83975",
         10347 => x"812a1670",
         10348 => x"892aa81b",
         10349 => x"0805b41b",
         10350 => x"0859595a",
         10351 => x"76782eb7",
         10352 => x"38800b83",
         10353 => x"1a33715e",
         10354 => x"565d747d",
         10355 => x"2e098106",
         10356 => x"82d43881",
         10357 => x"547753b8",
         10358 => x"19528119",
         10359 => x"3351f083",
         10360 => x"3f84b9c8",
         10361 => x"08802e85",
         10362 => x"38ff5881",
         10363 => x"5c77b41a",
         10364 => x"0c7b587b",
         10365 => x"fdac3879",
         10366 => x"83ff0619",
         10367 => x"b805811b",
         10368 => x"7781065f",
         10369 => x"5f577a55",
         10370 => x"7c802e8f",
         10371 => x"387a842b",
         10372 => x"9ff00677",
         10373 => x"338f0671",
         10374 => x"07565a74",
         10375 => x"7734810b",
         10376 => x"831a347d",
         10377 => x"892aa81a",
         10378 => x"08055680",
         10379 => x"0bb41a08",
         10380 => x"565f7476",
         10381 => x"2e83dd38",
         10382 => x"81547453",
         10383 => x"b8197053",
         10384 => x"811a3352",
         10385 => x"57f09b3f",
         10386 => x"815884b9",
         10387 => x"c8087f2e",
         10388 => x"09810680",
         10389 => x"c73884b9",
         10390 => x"c808831a",
         10391 => x"34b41908",
         10392 => x"70a81b08",
         10393 => x"31a01b08",
         10394 => x"84b9c808",
         10395 => x"5b5c565c",
         10396 => x"747a278b",
         10397 => x"38821933",
         10398 => x"5574822e",
         10399 => x"82e43881",
         10400 => x"54755376",
         10401 => x"52811933",
         10402 => x"51eed83f",
         10403 => x"84b9c808",
         10404 => x"802e8538",
         10405 => x"ff568158",
         10406 => x"75b41a0c",
         10407 => x"77fc8338",
         10408 => x"7d83ff06",
         10409 => x"19b8057b",
         10410 => x"842a5656",
         10411 => x"7c8f387a",
         10412 => x"882a7633",
         10413 => x"81f00671",
         10414 => x"8f060756",
         10415 => x"5c747634",
         10416 => x"810b831a",
         10417 => x"34fccb39",
         10418 => x"81547653",
         10419 => x"b8197053",
         10420 => x"811a3352",
         10421 => x"5def8b3f",
         10422 => x"815a84b9",
         10423 => x"c8087c2e",
         10424 => x"098106fc",
         10425 => x"883884b9",
         10426 => x"c808831a",
         10427 => x"34b41908",
         10428 => x"70a81b08",
         10429 => x"31a01b08",
         10430 => x"84b9c808",
         10431 => x"5d59405e",
         10432 => x"7e7727fb",
         10433 => x"ca388219",
         10434 => x"33557482",
         10435 => x"2e098106",
         10436 => x"fbbd3881",
         10437 => x"54761e53",
         10438 => x"7c528119",
         10439 => x"3351eec2",
         10440 => x"3f7b5afb",
         10441 => x"aa398154",
         10442 => x"7653b819",
         10443 => x"7053811a",
         10444 => x"335257ee",
         10445 => x"ad3f815c",
         10446 => x"84b9c808",
         10447 => x"7d2e0981",
         10448 => x"06fdae38",
         10449 => x"84b9c808",
         10450 => x"831a34b4",
         10451 => x"190870a8",
         10452 => x"1b0831a0",
         10453 => x"1b0884b9",
         10454 => x"c8085f40",
         10455 => x"565f747e",
         10456 => x"27fcf038",
         10457 => x"82193355",
         10458 => x"74822e09",
         10459 => x"8106fce3",
         10460 => x"3881547d",
         10461 => x"1f537652",
         10462 => x"81193351",
         10463 => x"ede43f7c",
         10464 => x"5cfcd039",
         10465 => x"81547653",
         10466 => x"b8197053",
         10467 => x"811a3352",
         10468 => x"57edcf3f",
         10469 => x"815a84b9",
         10470 => x"c8087c2e",
         10471 => x"098106fb",
         10472 => x"c53884b9",
         10473 => x"c808831a",
         10474 => x"34b41908",
         10475 => x"70a81b08",
         10476 => x"31a01b08",
         10477 => x"84b9c808",
         10478 => x"5d5f405e",
         10479 => x"7e7d27fb",
         10480 => x"87388219",
         10481 => x"33557482",
         10482 => x"2e098106",
         10483 => x"fafa3881",
         10484 => x"547c1e53",
         10485 => x"76528119",
         10486 => x"3351ed86",
         10487 => x"3f7b5afa",
         10488 => x"e7398154",
         10489 => x"791c5376",
         10490 => x"52811933",
         10491 => x"51ecf33f",
         10492 => x"7e58fd8b",
         10493 => x"397b7610",
         10494 => x"83fe067a",
         10495 => x"057c83ff",
         10496 => x"ff06595f",
         10497 => x"5876b81f",
         10498 => x"3476882a",
         10499 => x"5a79b91f",
         10500 => x"34f9fa39",
         10501 => x"7e58fd88",
         10502 => x"397b7682",
         10503 => x"2b83fc06",
         10504 => x"7a05b811",
         10505 => x"83113370",
         10506 => x"982b8f0a",
         10507 => x"067ff00a",
         10508 => x"06074258",
         10509 => x"5f5d587d",
         10510 => x"7d347d88",
         10511 => x"2a5675b9",
         10512 => x"1d347d90",
         10513 => x"2a5a79ba",
         10514 => x"1d347d98",
         10515 => x"2a5b7abb",
         10516 => x"1d34facf",
         10517 => x"39f63d0d",
         10518 => x"7c7e7108",
         10519 => x"5b5c5a7a",
         10520 => x"818a3890",
         10521 => x"19085776",
         10522 => x"802e80f4",
         10523 => x"38769c1a",
         10524 => x"082780ec",
         10525 => x"38941908",
         10526 => x"70565473",
         10527 => x"802e80d7",
         10528 => x"38767b2e",
         10529 => x"81933876",
         10530 => x"56811656",
         10531 => x"9c190876",
         10532 => x"26893882",
         10533 => x"56757726",
         10534 => x"82b23875",
         10535 => x"527951f0",
         10536 => x"f53f84b9",
         10537 => x"c808802e",
         10538 => x"81d03880",
         10539 => x"5884b9c8",
         10540 => x"08812eb1",
         10541 => x"3884b9c8",
         10542 => x"08097030",
         10543 => x"70720780",
         10544 => x"25707b07",
         10545 => x"51515555",
         10546 => x"7382aa38",
         10547 => x"75772e09",
         10548 => x"8106ffb5",
         10549 => x"38735574",
         10550 => x"84b9c80c",
         10551 => x"8c3d0d04",
         10552 => x"8157ff91",
         10553 => x"3984b9c8",
         10554 => x"0858ca39",
         10555 => x"7a527951",
         10556 => x"f0a43f81",
         10557 => x"557484b9",
         10558 => x"c80827db",
         10559 => x"3884b9c8",
         10560 => x"085584b9",
         10561 => x"c808ff2e",
         10562 => x"ce389c19",
         10563 => x"0884b9c8",
         10564 => x"0826c438",
         10565 => x"7a57fedd",
         10566 => x"39811b56",
         10567 => x"9c190876",
         10568 => x"26833882",
         10569 => x"56755279",
         10570 => x"51efeb3f",
         10571 => x"805884b9",
         10572 => x"c808812e",
         10573 => x"81a03884",
         10574 => x"b9c80809",
         10575 => x"70307072",
         10576 => x"07802570",
         10577 => x"7b0784b9",
         10578 => x"c8085451",
         10579 => x"51555573",
         10580 => x"ff853884",
         10581 => x"b9c80880",
         10582 => x"2e9a3890",
         10583 => x"19085481",
         10584 => x"7427fea3",
         10585 => x"38739c1a",
         10586 => x"0827fe9b",
         10587 => x"38737057",
         10588 => x"57fe9639",
         10589 => x"75802efe",
         10590 => x"8e38ff53",
         10591 => x"75527851",
         10592 => x"f5f53f84",
         10593 => x"b9c80884",
         10594 => x"b9c80830",
         10595 => x"7084b9c8",
         10596 => x"08078025",
         10597 => x"5658557a",
         10598 => x"80c43874",
         10599 => x"80e33875",
         10600 => x"901a0c9c",
         10601 => x"1908fe05",
         10602 => x"941a0856",
         10603 => x"58747826",
         10604 => x"8638ff15",
         10605 => x"941a0c84",
         10606 => x"19338107",
         10607 => x"5a79841a",
         10608 => x"34755574",
         10609 => x"84b9c80c",
         10610 => x"8c3d0d04",
         10611 => x"800b84b9",
         10612 => x"c80c8c3d",
         10613 => x"0d0484b9",
         10614 => x"c80858fe",
         10615 => x"da397380",
         10616 => x"2effb838",
         10617 => x"75537a52",
         10618 => x"7851f58b",
         10619 => x"3f84b9c8",
         10620 => x"0855ffa7",
         10621 => x"3984b9c8",
         10622 => x"0884b9c8",
         10623 => x"0c8c3d0d",
         10624 => x"04ff5674",
         10625 => x"812effb9",
         10626 => x"388155ff",
         10627 => x"b639f83d",
         10628 => x"0d7a7c71",
         10629 => x"08595558",
         10630 => x"73f0800a",
         10631 => x"2680df38",
         10632 => x"739f0653",
         10633 => x"7280d738",
         10634 => x"7390190c",
         10635 => x"88180855",
         10636 => x"7480df38",
         10637 => x"76335675",
         10638 => x"822680cc",
         10639 => x"3873852a",
         10640 => x"53820b88",
         10641 => x"18225a56",
         10642 => x"727927a9",
         10643 => x"38ac1708",
         10644 => x"98190c74",
         10645 => x"94190c98",
         10646 => x"18085382",
         10647 => x"5672802e",
         10648 => x"94387389",
         10649 => x"2a139819",
         10650 => x"0c7383ff",
         10651 => x"0617b805",
         10652 => x"9c190c80",
         10653 => x"567584b9",
         10654 => x"c80c8a3d",
         10655 => x"0d04820b",
         10656 => x"84b9c80c",
         10657 => x"8a3d0d04",
         10658 => x"ac170855",
         10659 => x"74802eff",
         10660 => x"ac388a17",
         10661 => x"2270892b",
         10662 => x"57597376",
         10663 => x"27a5389c",
         10664 => x"170853fe",
         10665 => x"15fe1454",
         10666 => x"56805975",
         10667 => x"73278d38",
         10668 => x"8a172276",
         10669 => x"7129b019",
         10670 => x"08055a53",
         10671 => x"7898190c",
         10672 => x"ff913974",
         10673 => x"527751ec",
         10674 => x"cd3f84b9",
         10675 => x"c8085584",
         10676 => x"b9c808ff",
         10677 => x"2ea43881",
         10678 => x"0b84b9c8",
         10679 => x"0827ff9e",
         10680 => x"389c1708",
         10681 => x"5384b9c8",
         10682 => x"087327ff",
         10683 => x"91387376",
         10684 => x"31547376",
         10685 => x"27cd38ff",
         10686 => x"aa39810b",
         10687 => x"84b9c80c",
         10688 => x"8a3d0d04",
         10689 => x"f33d0d7f",
         10690 => x"70089012",
         10691 => x"08a0055c",
         10692 => x"5a57f080",
         10693 => x"0a7a2786",
         10694 => x"38800b98",
         10695 => x"180c9817",
         10696 => x"08558456",
         10697 => x"74802eb2",
         10698 => x"387983ff",
         10699 => x"065b7a9d",
         10700 => x"38811594",
         10701 => x"18085758",
         10702 => x"75a93879",
         10703 => x"852a881a",
         10704 => x"22575574",
         10705 => x"762781f5",
         10706 => x"38779818",
         10707 => x"0c799018",
         10708 => x"0c781bb8",
         10709 => x"059c180c",
         10710 => x"80567584",
         10711 => x"b9c80c8f",
         10712 => x"3d0d0477",
         10713 => x"98180c8a",
         10714 => x"1922ff05",
         10715 => x"7a892a06",
         10716 => x"5c7bda38",
         10717 => x"75527651",
         10718 => x"eb9c3f84",
         10719 => x"b9c8085d",
         10720 => x"8256810b",
         10721 => x"84b9c808",
         10722 => x"27d03881",
         10723 => x"5684b9c8",
         10724 => x"08ff2ec6",
         10725 => x"389c1908",
         10726 => x"84b9c808",
         10727 => x"26829138",
         10728 => x"60802e81",
         10729 => x"98389417",
         10730 => x"08527651",
         10731 => x"f9a73f84",
         10732 => x"b9c8085d",
         10733 => x"875684b9",
         10734 => x"c808802e",
         10735 => x"ff9c3882",
         10736 => x"5684b9c8",
         10737 => x"08812eff",
         10738 => x"91388156",
         10739 => x"84b9c808",
         10740 => x"ff2eff86",
         10741 => x"3884b9c8",
         10742 => x"08831a33",
         10743 => x"5f587d80",
         10744 => x"ea38fe18",
         10745 => x"9c1a08fe",
         10746 => x"05595680",
         10747 => x"5c757827",
         10748 => x"8d388a19",
         10749 => x"22767129",
         10750 => x"b01b0805",
         10751 => x"5d5e7bb4",
         10752 => x"1a0cb819",
         10753 => x"58848078",
         10754 => x"57558076",
         10755 => x"70810558",
         10756 => x"34ff1555",
         10757 => x"74f43874",
         10758 => x"568a1922",
         10759 => x"55757527",
         10760 => x"81803881",
         10761 => x"54751c53",
         10762 => x"77528119",
         10763 => x"3351e4b2",
         10764 => x"3f84b9c8",
         10765 => x"0880e738",
         10766 => x"811656dd",
         10767 => x"397a9818",
         10768 => x"0c840b84",
         10769 => x"b9c80c8f",
         10770 => x"3d0d0475",
         10771 => x"54b41908",
         10772 => x"53b81970",
         10773 => x"53811a33",
         10774 => x"5256e486",
         10775 => x"3f84b9c8",
         10776 => x"0880f338",
         10777 => x"84b9c808",
         10778 => x"831a34b4",
         10779 => x"1908a81a",
         10780 => x"08315574",
         10781 => x"a01a0827",
         10782 => x"fee83882",
         10783 => x"19335c7b",
         10784 => x"822e0981",
         10785 => x"06fedb38",
         10786 => x"8154b419",
         10787 => x"08a01a08",
         10788 => x"05537552",
         10789 => x"81193351",
         10790 => x"e3c83ffe",
         10791 => x"c5398a19",
         10792 => x"22557483",
         10793 => x"ffff0655",
         10794 => x"74762e09",
         10795 => x"8106a738",
         10796 => x"7c94180c",
         10797 => x"fe1d9c1a",
         10798 => x"08fe055e",
         10799 => x"56805875",
         10800 => x"7d27fd85",
         10801 => x"388a1922",
         10802 => x"767129b0",
         10803 => x"1b080598",
         10804 => x"190c5cfc",
         10805 => x"f839810b",
         10806 => x"84b9c80c",
         10807 => x"8f3d0d04",
         10808 => x"ee3d0d64",
         10809 => x"66415c84",
         10810 => x"7c085a5b",
         10811 => x"81ff7098",
         10812 => x"1e08585e",
         10813 => x"5e75802e",
         10814 => x"82d238b8",
         10815 => x"195f755a",
         10816 => x"8058b419",
         10817 => x"08762e82",
         10818 => x"d1388319",
         10819 => x"33785855",
         10820 => x"74782e09",
         10821 => x"81068194",
         10822 => x"38815475",
         10823 => x"53b81952",
         10824 => x"81193351",
         10825 => x"e1bd3f84",
         10826 => x"b9c80880",
         10827 => x"2e8538ff",
         10828 => x"5a815779",
         10829 => x"b41a0c76",
         10830 => x"5b768290",
         10831 => x"389c1c08",
         10832 => x"70335858",
         10833 => x"76802e82",
         10834 => x"81388b18",
         10835 => x"33bf0670",
         10836 => x"81ff065b",
         10837 => x"4160861d",
         10838 => x"347681e5",
         10839 => x"32703078",
         10840 => x"ae327030",
         10841 => x"72802571",
         10842 => x"80250754",
         10843 => x"45455755",
         10844 => x"74933874",
         10845 => x"7adf0643",
         10846 => x"5661882e",
         10847 => x"81bf3875",
         10848 => x"602e8186",
         10849 => x"3881ff5d",
         10850 => x"80527b51",
         10851 => x"faf63f84",
         10852 => x"b9c8085b",
         10853 => x"84b9c808",
         10854 => x"81b23898",
         10855 => x"1c085675",
         10856 => x"fedc387a",
         10857 => x"84b9c80c",
         10858 => x"943d0d04",
         10859 => x"8154b419",
         10860 => x"08537e52",
         10861 => x"81193351",
         10862 => x"e1a83f81",
         10863 => x"5784b9c8",
         10864 => x"08782e09",
         10865 => x"8106feef",
         10866 => x"3884b9c8",
         10867 => x"08831a34",
         10868 => x"b41908a8",
         10869 => x"1a083184",
         10870 => x"b9c80858",
         10871 => x"5b7aa01a",
         10872 => x"0827feb5",
         10873 => x"38821933",
         10874 => x"4160822e",
         10875 => x"098106fe",
         10876 => x"a8388154",
         10877 => x"b41908a0",
         10878 => x"1a080553",
         10879 => x"7e528119",
         10880 => x"3351e0de",
         10881 => x"3f7757fe",
         10882 => x"9039798f",
         10883 => x"2e098106",
         10884 => x"81e73876",
         10885 => x"862a8106",
         10886 => x"5b7a802e",
         10887 => x"93388d18",
         10888 => x"337781bf",
         10889 => x"0670901f",
         10890 => x"087fac05",
         10891 => x"0c595e5e",
         10892 => x"767d2eab",
         10893 => x"3881ff55",
         10894 => x"745dfecc",
         10895 => x"39815675",
         10896 => x"602e0981",
         10897 => x"06febe38",
         10898 => x"c139845b",
         10899 => x"800b981d",
         10900 => x"0c7a84b9",
         10901 => x"c80c943d",
         10902 => x"0d04775b",
         10903 => x"fddf398d",
         10904 => x"1833577d",
         10905 => x"772e0981",
         10906 => x"06cb388c",
         10907 => x"19089b19",
         10908 => x"339a1a33",
         10909 => x"71882b07",
         10910 => x"58564175",
         10911 => x"ffb73877",
         10912 => x"337081bf",
         10913 => x"068d29f3",
         10914 => x"05515a81",
         10915 => x"76585b83",
         10916 => x"e5c81733",
         10917 => x"78058111",
         10918 => x"33713371",
         10919 => x"882b0752",
         10920 => x"44567a80",
         10921 => x"2e80c538",
         10922 => x"7981fe26",
         10923 => x"ff873879",
         10924 => x"10610576",
         10925 => x"5c427562",
         10926 => x"23811a5a",
         10927 => x"8117578c",
         10928 => x"7727cc38",
         10929 => x"77337086",
         10930 => x"2a810659",
         10931 => x"5777802e",
         10932 => x"90387981",
         10933 => x"fe26fedd",
         10934 => x"38791061",
         10935 => x"05438063",
         10936 => x"23ff1d70",
         10937 => x"81ff065e",
         10938 => x"41fd9d39",
         10939 => x"7583ffff",
         10940 => x"2eca3881",
         10941 => x"ff55fec0",
         10942 => x"397ca838",
         10943 => x"7c558b57",
         10944 => x"74812a75",
         10945 => x"81802905",
         10946 => x"78708105",
         10947 => x"5a33407f",
         10948 => x"057081ff",
         10949 => x"06ff1959",
         10950 => x"565976e4",
         10951 => x"38747e2e",
         10952 => x"fd8138ff",
         10953 => x"0bac1d0c",
         10954 => x"7a84b9c8",
         10955 => x"0c943d0d",
         10956 => x"04ef3d0d",
         10957 => x"6370085c",
         10958 => x"5c80527b",
         10959 => x"51f5cf3f",
         10960 => x"84b9c808",
         10961 => x"5a84b9c8",
         10962 => x"08828038",
         10963 => x"81ff7040",
         10964 => x"5dff0bac",
         10965 => x"1d0cb81b",
         10966 => x"5e981c08",
         10967 => x"568058b4",
         10968 => x"1b08762e",
         10969 => x"82cc3883",
         10970 => x"1b337858",
         10971 => x"5574782e",
         10972 => x"09810681",
         10973 => x"df388154",
         10974 => x"7553b81b",
         10975 => x"52811b33",
         10976 => x"51dce03f",
         10977 => x"84b9c808",
         10978 => x"802e8538",
         10979 => x"ff568157",
         10980 => x"75b41c0c",
         10981 => x"765a7681",
         10982 => x"b2389c1c",
         10983 => x"08703358",
         10984 => x"5976802e",
         10985 => x"8499388b",
         10986 => x"1933bf06",
         10987 => x"7081ff06",
         10988 => x"57587786",
         10989 => x"1d347681",
         10990 => x"e52e80f2",
         10991 => x"3875832a",
         10992 => x"81065575",
         10993 => x"8f2e81ef",
         10994 => x"387480e2",
         10995 => x"38758f2e",
         10996 => x"81e5387c",
         10997 => x"aa38787d",
         10998 => x"56588b57",
         10999 => x"74812a75",
         11000 => x"81802905",
         11001 => x"78708105",
         11002 => x"5a335776",
         11003 => x"057081ff",
         11004 => x"06ff1959",
         11005 => x"565d76e4",
         11006 => x"38747f2e",
         11007 => x"80cd38ab",
         11008 => x"1c338106",
         11009 => x"5776a738",
         11010 => x"8b0ba01d",
         11011 => x"59577870",
         11012 => x"81055a33",
         11013 => x"78708105",
         11014 => x"5a337171",
         11015 => x"31ff1a5a",
         11016 => x"58424076",
         11017 => x"802e81dc",
         11018 => x"3875802e",
         11019 => x"e13881ff",
         11020 => x"5dff0bac",
         11021 => x"1d0c8052",
         11022 => x"7b51f5c8",
         11023 => x"3f84b9c8",
         11024 => x"085a84b9",
         11025 => x"c808802e",
         11026 => x"fe8f3879",
         11027 => x"84b9c80c",
         11028 => x"933d0d04",
         11029 => x"8154b41b",
         11030 => x"08537d52",
         11031 => x"811b3351",
         11032 => x"dc803f81",
         11033 => x"5784b9c8",
         11034 => x"08782e09",
         11035 => x"8106fea4",
         11036 => x"3884b9c8",
         11037 => x"08831c34",
         11038 => x"b41b08a8",
         11039 => x"1c083184",
         11040 => x"b9c80858",
         11041 => x"5978a01c",
         11042 => x"0827fdea",
         11043 => x"38821b33",
         11044 => x"5a79822e",
         11045 => x"098106fd",
         11046 => x"dd388154",
         11047 => x"b41b08a0",
         11048 => x"1c080553",
         11049 => x"7d52811b",
         11050 => x"3351dbb6",
         11051 => x"3f7757fd",
         11052 => x"c539775a",
         11053 => x"fde439ab",
         11054 => x"1c337086",
         11055 => x"2a810642",
         11056 => x"5560fef2",
         11057 => x"3876862a",
         11058 => x"81065a79",
         11059 => x"802e9338",
         11060 => x"8d193377",
         11061 => x"81bf0670",
         11062 => x"901f087f",
         11063 => x"ac050c59",
         11064 => x"5e5f767d",
         11065 => x"2eaf3881",
         11066 => x"ff55745d",
         11067 => x"80527b51",
         11068 => x"f4923f84",
         11069 => x"b9c8085a",
         11070 => x"84b9c808",
         11071 => x"802efcd9",
         11072 => x"38fec839",
         11073 => x"75802efe",
         11074 => x"c23881ff",
         11075 => x"5dff0bac",
         11076 => x"1d0cfea2",
         11077 => x"398d1933",
         11078 => x"577e772e",
         11079 => x"098106c7",
         11080 => x"388c1b08",
         11081 => x"9b1a339a",
         11082 => x"1b337188",
         11083 => x"2b075942",
         11084 => x"4076ffb3",
         11085 => x"38783370",
         11086 => x"bf068d29",
         11087 => x"f3055b55",
         11088 => x"81775956",
         11089 => x"83e5c818",
         11090 => x"33790581",
         11091 => x"11337133",
         11092 => x"71882b07",
         11093 => x"52425775",
         11094 => x"802e80ed",
         11095 => x"387981fe",
         11096 => x"26ff8438",
         11097 => x"765181a1",
         11098 => x"8a3f84b9",
         11099 => x"c8087a10",
         11100 => x"61057022",
         11101 => x"5343811b",
         11102 => x"5b5681a0",
         11103 => x"f63f7584",
         11104 => x"b9c8082e",
         11105 => x"098106fe",
         11106 => x"de387656",
         11107 => x"8118588c",
         11108 => x"7827ffb0",
         11109 => x"38783370",
         11110 => x"862a8106",
         11111 => x"56597580",
         11112 => x"2e923874",
         11113 => x"802e8d38",
         11114 => x"79106005",
         11115 => x"70224141",
         11116 => x"7ffeb438",
         11117 => x"ff1d7081",
         11118 => x"ff065e5a",
         11119 => x"feae3984",
         11120 => x"0b84b9c8",
         11121 => x"0c933d0d",
         11122 => x"047683ff",
         11123 => x"ff2effbc",
         11124 => x"3881ff55",
         11125 => x"fe9439ea",
         11126 => x"3d0d6870",
         11127 => x"0870ab13",
         11128 => x"3381a006",
         11129 => x"585a5d5e",
         11130 => x"86567485",
         11131 => x"b538748c",
         11132 => x"1d087022",
         11133 => x"57575d74",
         11134 => x"802e8e38",
         11135 => x"811d7010",
         11136 => x"17702251",
         11137 => x"565d74f4",
         11138 => x"38953da0",
         11139 => x"1f5b408c",
         11140 => x"607b5858",
         11141 => x"55757081",
         11142 => x"05573377",
         11143 => x"70810559",
         11144 => x"34ff1555",
         11145 => x"74ef3802",
         11146 => x"80db0533",
         11147 => x"70810658",
         11148 => x"5676802e",
         11149 => x"82aa3880",
         11150 => x"c00bab1f",
         11151 => x"34810b94",
         11152 => x"3d405b8c",
         11153 => x"1c087b58",
         11154 => x"598b7a61",
         11155 => x"5a575577",
         11156 => x"70810559",
         11157 => x"33767081",
         11158 => x"055834ff",
         11159 => x"155574ef",
         11160 => x"38857b27",
         11161 => x"80c2387a",
         11162 => x"79225657",
         11163 => x"74802eb8",
         11164 => x"3874821a",
         11165 => x"5a568f58",
         11166 => x"75810677",
         11167 => x"10077681",
         11168 => x"2a7083ff",
         11169 => x"ff067290",
         11170 => x"2a810644",
         11171 => x"58565760",
         11172 => x"802e8738",
         11173 => x"7684a0a1",
         11174 => x"3257ff18",
         11175 => x"58778025",
         11176 => x"d7387822",
         11177 => x"5574ca38",
         11178 => x"87028405",
         11179 => x"80cf0557",
         11180 => x"5876b007",
         11181 => x"bf0655b9",
         11182 => x"75278438",
         11183 => x"87155574",
         11184 => x"7634ff16",
         11185 => x"ff197884",
         11186 => x"2a595956",
         11187 => x"76e33877",
         11188 => x"1f5980fe",
         11189 => x"7934767a",
         11190 => x"58568078",
         11191 => x"27a03879",
         11192 => x"335574a0",
         11193 => x"2e983881",
         11194 => x"16567578",
         11195 => x"2788a238",
         11196 => x"751a7033",
         11197 => x"565774a0",
         11198 => x"2e098106",
         11199 => x"ea388116",
         11200 => x"56a05577",
         11201 => x"87268e38",
         11202 => x"983d7805",
         11203 => x"ec058119",
         11204 => x"71335759",
         11205 => x"41747734",
         11206 => x"87762787",
         11207 => x"f4387d51",
         11208 => x"f88f3f84",
         11209 => x"b9c8088b",
         11210 => x"38811b5b",
         11211 => x"80e37b27",
         11212 => x"fe913887",
         11213 => x"567a80e4",
         11214 => x"2e82e738",
         11215 => x"84b9c808",
         11216 => x"5684b9c8",
         11217 => x"08842e09",
         11218 => x"810682d6",
         11219 => x"380280db",
         11220 => x"0533ab1f",
         11221 => x"347d0802",
         11222 => x"840580db",
         11223 => x"05335758",
         11224 => x"75812a81",
         11225 => x"065f815b",
         11226 => x"7e802e90",
         11227 => x"388d528c",
         11228 => x"1d51fe8a",
         11229 => x"b03f84b9",
         11230 => x"c8081b5b",
         11231 => x"80527d51",
         11232 => x"ed8c3f84",
         11233 => x"b9c80856",
         11234 => x"84b9c808",
         11235 => x"81823884",
         11236 => x"b9c808b8",
         11237 => x"195e5998",
         11238 => x"1e085680",
         11239 => x"57b41808",
         11240 => x"762e85f3",
         11241 => x"38831833",
         11242 => x"407f772e",
         11243 => x"09810682",
         11244 => x"a3388154",
         11245 => x"7553b818",
         11246 => x"52811833",
         11247 => x"51d4a43f",
         11248 => x"84b9c808",
         11249 => x"802e8538",
         11250 => x"ff568157",
         11251 => x"75b4190c",
         11252 => x"765676bc",
         11253 => x"389c1e08",
         11254 => x"70335642",
         11255 => x"7481e52e",
         11256 => x"81c93874",
         11257 => x"30708025",
         11258 => x"7807565f",
         11259 => x"74802e81",
         11260 => x"c9388119",
         11261 => x"59787b2e",
         11262 => x"86893881",
         11263 => x"527d51ee",
         11264 => x"833f84b9",
         11265 => x"c8085684",
         11266 => x"b9c80880",
         11267 => x"2eff8838",
         11268 => x"87587584",
         11269 => x"2e818938",
         11270 => x"75587581",
         11271 => x"8338ff1b",
         11272 => x"407f81f3",
         11273 => x"38981e08",
         11274 => x"57b41c08",
         11275 => x"772eaf38",
         11276 => x"831c3378",
         11277 => x"57407f84",
         11278 => x"82388154",
         11279 => x"7653b81c",
         11280 => x"52811c33",
         11281 => x"51d39c3f",
         11282 => x"84b9c808",
         11283 => x"802e8538",
         11284 => x"ff578156",
         11285 => x"76b41d0c",
         11286 => x"75587580",
         11287 => x"c338a00b",
         11288 => x"9c1f0857",
         11289 => x"55807670",
         11290 => x"81055834",
         11291 => x"ff155574",
         11292 => x"f4388b0b",
         11293 => x"9c1f087b",
         11294 => x"58585575",
         11295 => x"70810557",
         11296 => x"33777081",
         11297 => x"055934ff",
         11298 => x"155574ef",
         11299 => x"389c1e08",
         11300 => x"ab1f3398",
         11301 => x"065e5a7c",
         11302 => x"8c1b3481",
         11303 => x"0b831d34",
         11304 => x"77567584",
         11305 => x"b9c80c98",
         11306 => x"3d0d0481",
         11307 => x"75307080",
         11308 => x"25720757",
         11309 => x"405774fe",
         11310 => x"b9387459",
         11311 => x"81527d51",
         11312 => x"ecc23f84",
         11313 => x"b9c80856",
         11314 => x"84b9c808",
         11315 => x"802efdc7",
         11316 => x"38febd39",
         11317 => x"8154b418",
         11318 => x"08537c52",
         11319 => x"81183351",
         11320 => x"d3803f84",
         11321 => x"b9c80877",
         11322 => x"2e098106",
         11323 => x"83bf3884",
         11324 => x"b9c80883",
         11325 => x"1934b418",
         11326 => x"08a81908",
         11327 => x"315574a0",
         11328 => x"1908278b",
         11329 => x"38821833",
         11330 => x"4160822e",
         11331 => x"84ac3884",
         11332 => x"b9c80857",
         11333 => x"fd9c397f",
         11334 => x"852b901f",
         11335 => x"08713153",
         11336 => x"587d51e9",
         11337 => x"e93f84b9",
         11338 => x"c8085884",
         11339 => x"b9c808fe",
         11340 => x"ef387984",
         11341 => x"b9c80856",
         11342 => x"588b5774",
         11343 => x"812a7581",
         11344 => x"80290578",
         11345 => x"7081055a",
         11346 => x"33577605",
         11347 => x"7081ff06",
         11348 => x"ff195956",
         11349 => x"5d76e438",
         11350 => x"7481ff06",
         11351 => x"b81d4341",
         11352 => x"981e0857",
         11353 => x"8056b41c",
         11354 => x"08772eb2",
         11355 => x"38831c33",
         11356 => x"5b7a762e",
         11357 => x"09810682",
         11358 => x"c9388154",
         11359 => x"7653b81c",
         11360 => x"52811c33",
         11361 => x"51d0dc3f",
         11362 => x"84b9c808",
         11363 => x"802e8538",
         11364 => x"ff578156",
         11365 => x"76b41d0c",
         11366 => x"755875fe",
         11367 => x"83388c1c",
         11368 => x"089c1f08",
         11369 => x"6181ff06",
         11370 => x"5f5c5f60",
         11371 => x"8d1c348f",
         11372 => x"0b8b1c34",
         11373 => x"758c1c34",
         11374 => x"759a1c34",
         11375 => x"759b1c34",
         11376 => x"7c8d29f3",
         11377 => x"0576775a",
         11378 => x"58597683",
         11379 => x"ffff2e8b",
         11380 => x"3878101f",
         11381 => x"7022811b",
         11382 => x"5b585683",
         11383 => x"e5c81833",
         11384 => x"7b055576",
         11385 => x"75708105",
         11386 => x"57347688",
         11387 => x"2a567575",
         11388 => x"34768538",
         11389 => x"83ffff57",
         11390 => x"8118588c",
         11391 => x"7827cb38",
         11392 => x"7683ffff",
         11393 => x"2e81b338",
         11394 => x"78101f70",
         11395 => x"22585876",
         11396 => x"802e81a6",
         11397 => x"387c7b34",
         11398 => x"810b831d",
         11399 => x"3480527d",
         11400 => x"51e9e13f",
         11401 => x"84b9c808",
         11402 => x"5884b9c8",
         11403 => x"08fcf138",
         11404 => x"7fff0540",
         11405 => x"7ffea938",
         11406 => x"fbeb3981",
         11407 => x"54b41c08",
         11408 => x"53b81c70",
         11409 => x"53811d33",
         11410 => x"5259d096",
         11411 => x"3f815684",
         11412 => x"b9c808fc",
         11413 => x"833884b9",
         11414 => x"c808831d",
         11415 => x"34b41c08",
         11416 => x"a81d0831",
         11417 => x"84b9c808",
         11418 => x"574160a0",
         11419 => x"1d0827fb",
         11420 => x"c938821c",
         11421 => x"33426182",
         11422 => x"2e098106",
         11423 => x"fbbc3881",
         11424 => x"54b41c08",
         11425 => x"a01d0805",
         11426 => x"53785281",
         11427 => x"1c3351cf",
         11428 => x"d13f7756",
         11429 => x"fba43976",
         11430 => x"9c1f0870",
         11431 => x"33574356",
         11432 => x"7481e52e",
         11433 => x"098106fa",
         11434 => x"ba38fbff",
         11435 => x"39817057",
         11436 => x"5776802e",
         11437 => x"fa9f38fa",
         11438 => x"d7397c80",
         11439 => x"c0075dfe",
         11440 => x"d4398154",
         11441 => x"b41c0853",
         11442 => x"6152811c",
         11443 => x"3351cf92",
         11444 => x"3f84b9c8",
         11445 => x"08762e09",
         11446 => x"8106bc38",
         11447 => x"84b9c808",
         11448 => x"831d34b4",
         11449 => x"1c08a81d",
         11450 => x"08315574",
         11451 => x"a01d0827",
         11452 => x"8a38821c",
         11453 => x"335f7e82",
         11454 => x"2eaa3884",
         11455 => x"b9c80856",
         11456 => x"fcf83975",
         11457 => x"ff1c4158",
         11458 => x"7f802efa",
         11459 => x"9838fc87",
         11460 => x"39751a57",
         11461 => x"f7e83981",
         11462 => x"70595675",
         11463 => x"802efcfe",
         11464 => x"38fafd39",
         11465 => x"8154b41c",
         11466 => x"08a01d08",
         11467 => x"05536152",
         11468 => x"811c3351",
         11469 => x"ceac3ffc",
         11470 => x"c1398154",
         11471 => x"b41808a0",
         11472 => x"19080553",
         11473 => x"7c528118",
         11474 => x"3351ce96",
         11475 => x"3ff8e339",
         11476 => x"f33d0d7f",
         11477 => x"61710840",
         11478 => x"5e5c800b",
         11479 => x"961e3498",
         11480 => x"1c08802e",
         11481 => x"82b538ac",
         11482 => x"1c08ff2e",
         11483 => x"80d93880",
         11484 => x"7071608c",
         11485 => x"05087022",
         11486 => x"57585b5c",
         11487 => x"5872782e",
         11488 => x"bc387754",
         11489 => x"74147022",
         11490 => x"811b5b55",
         11491 => x"567a8295",
         11492 => x"3880d080",
         11493 => x"147083ff",
         11494 => x"ff06585a",
         11495 => x"768fff26",
         11496 => x"82833873",
         11497 => x"791a7611",
         11498 => x"70225d58",
         11499 => x"555b79d4",
         11500 => x"387a3070",
         11501 => x"80257030",
         11502 => x"7a065a5c",
         11503 => x"5e7c1894",
         11504 => x"0557800b",
         11505 => x"82183480",
         11506 => x"70891f59",
         11507 => x"57589c1c",
         11508 => x"08167033",
         11509 => x"81185856",
         11510 => x"5374a02e",
         11511 => x"b2387485",
         11512 => x"2e81bc38",
         11513 => x"75893270",
         11514 => x"30707207",
         11515 => x"8025555b",
         11516 => x"54778b26",
         11517 => x"90387280",
         11518 => x"2e8b38ae",
         11519 => x"77708105",
         11520 => x"59348118",
         11521 => x"58747770",
         11522 => x"81055934",
         11523 => x"8118588a",
         11524 => x"7627ffba",
         11525 => x"387c1888",
         11526 => x"0555800b",
         11527 => x"81163496",
         11528 => x"1d335372",
         11529 => x"a5387781",
         11530 => x"f338bf0b",
         11531 => x"961e3481",
         11532 => x"577c1794",
         11533 => x"0556800b",
         11534 => x"8217349c",
         11535 => x"1c088c11",
         11536 => x"33555373",
         11537 => x"89387389",
         11538 => x"1e349c1c",
         11539 => x"08538b13",
         11540 => x"33881e34",
         11541 => x"9c1c089c",
         11542 => x"11831133",
         11543 => x"82123371",
         11544 => x"902b7188",
         11545 => x"2b078114",
         11546 => x"33707207",
         11547 => x"882b7533",
         11548 => x"7107640c",
         11549 => x"59971633",
         11550 => x"96173371",
         11551 => x"882b075f",
         11552 => x"415b405a",
         11553 => x"565b5577",
         11554 => x"861e2399",
         11555 => x"15339816",
         11556 => x"3371882b",
         11557 => x"075d547b",
         11558 => x"841e238f",
         11559 => x"3d0d0481",
         11560 => x"e555fec0",
         11561 => x"39771d96",
         11562 => x"1181ff7a",
         11563 => x"31585b57",
         11564 => x"83b5527a",
         11565 => x"902b7407",
         11566 => x"51819189",
         11567 => x"3f84b9c8",
         11568 => x"0883ffff",
         11569 => x"065581ff",
         11570 => x"7527ad38",
         11571 => x"81762781",
         11572 => x"b3387488",
         11573 => x"2a54737a",
         11574 => x"34749718",
         11575 => x"34827805",
         11576 => x"58800b8c",
         11577 => x"1f08565b",
         11578 => x"78197511",
         11579 => x"70225c57",
         11580 => x"5479fd90",
         11581 => x"38fdba39",
         11582 => x"74307630",
         11583 => x"70780780",
         11584 => x"25728025",
         11585 => x"07585557",
         11586 => x"7580f938",
         11587 => x"747a3481",
         11588 => x"78055880",
         11589 => x"0b8c1f08",
         11590 => x"565bcd39",
         11591 => x"7273891f",
         11592 => x"335a5757",
         11593 => x"77802efe",
         11594 => x"88387c96",
         11595 => x"1e7e5759",
         11596 => x"54891433",
         11597 => x"ffbf115a",
         11598 => x"54789926",
         11599 => x"a4389c1c",
         11600 => x"088c1133",
         11601 => x"545b8876",
         11602 => x"27b43872",
         11603 => x"842a5372",
         11604 => x"81065e7d",
         11605 => x"802e8a38",
         11606 => x"a0147083",
         11607 => x"ffff0655",
         11608 => x"53737870",
         11609 => x"81055a34",
         11610 => x"81168116",
         11611 => x"81197189",
         11612 => x"13335e57",
         11613 => x"59565679",
         11614 => x"ffb738fd",
         11615 => x"b4397283",
         11616 => x"2a53cc39",
         11617 => x"807b3070",
         11618 => x"80257030",
         11619 => x"7306535d",
         11620 => x"5f58fca9",
         11621 => x"39ef3d0d",
         11622 => x"63700870",
         11623 => x"42575c80",
         11624 => x"65703357",
         11625 => x"555374af",
         11626 => x"2e833881",
         11627 => x"537480dc",
         11628 => x"2e81df38",
         11629 => x"72802e81",
         11630 => x"d9389816",
         11631 => x"08881d0c",
         11632 => x"7333963d",
         11633 => x"943d4142",
         11634 => x"559f7527",
         11635 => x"82a73873",
         11636 => x"428c1608",
         11637 => x"58805761",
         11638 => x"70708105",
         11639 => x"52335553",
         11640 => x"7381df38",
         11641 => x"727f0c73",
         11642 => x"ff2e81ec",
         11643 => x"3883ffff",
         11644 => x"74278b38",
         11645 => x"76101856",
         11646 => x"80762381",
         11647 => x"17577383",
         11648 => x"ffff0670",
         11649 => x"af327030",
         11650 => x"9f732771",
         11651 => x"80250757",
         11652 => x"5b5b5573",
         11653 => x"82903874",
         11654 => x"80dc2e82",
         11655 => x"89387480",
         11656 => x"ff26b238",
         11657 => x"83e4e40b",
         11658 => x"83e4e433",
         11659 => x"7081ff06",
         11660 => x"56545673",
         11661 => x"802e81ab",
         11662 => x"3873752e",
         11663 => x"8f388116",
         11664 => x"70337081",
         11665 => x"ff065654",
         11666 => x"5673ee38",
         11667 => x"7281ff06",
         11668 => x"5b7a8184",
         11669 => x"387681fe",
         11670 => x"2680fd38",
         11671 => x"7610185d",
         11672 => x"747d2381",
         11673 => x"17627070",
         11674 => x"81055233",
         11675 => x"56545773",
         11676 => x"802efef0",
         11677 => x"3880cb39",
         11678 => x"817380dc",
         11679 => x"32703070",
         11680 => x"80257307",
         11681 => x"51555855",
         11682 => x"72802ea1",
         11683 => x"38811470",
         11684 => x"46548074",
         11685 => x"33545572",
         11686 => x"af2edd38",
         11687 => x"7280dc32",
         11688 => x"70307080",
         11689 => x"25770751",
         11690 => x"545772e1",
         11691 => x"3872881d",
         11692 => x"0c733396",
         11693 => x"3d943d41",
         11694 => x"4255749f",
         11695 => x"26fe9038",
         11696 => x"b43983b5",
         11697 => x"52735181",
         11698 => x"8de73f84",
         11699 => x"b9c80883",
         11700 => x"ffff0654",
         11701 => x"73fe8d38",
         11702 => x"86547384",
         11703 => x"b9c80c93",
         11704 => x"3d0d0483",
         11705 => x"e4e43370",
         11706 => x"81ff065c",
         11707 => x"537a802e",
         11708 => x"fee338e4",
         11709 => x"39ff800b",
         11710 => x"ab1d3480",
         11711 => x"527b51de",
         11712 => x"8d3f84b9",
         11713 => x"c80884b9",
         11714 => x"c80c933d",
         11715 => x"0d048173",
         11716 => x"80dc3270",
         11717 => x"30708025",
         11718 => x"73074155",
         11719 => x"5a567d80",
         11720 => x"2ea13881",
         11721 => x"14428062",
         11722 => x"70335555",
         11723 => x"5672af2e",
         11724 => x"dd387280",
         11725 => x"dc327030",
         11726 => x"70802578",
         11727 => x"07405459",
         11728 => x"7de13873",
         11729 => x"610c9f75",
         11730 => x"27822b5a",
         11731 => x"76812e84",
         11732 => x"f8387682",
         11733 => x"2e83d138",
         11734 => x"76175976",
         11735 => x"802ea738",
         11736 => x"76177811",
         11737 => x"fe057022",
         11738 => x"70a03270",
         11739 => x"30709f2a",
         11740 => x"5242565f",
         11741 => x"56597cae",
         11742 => x"2e843872",
         11743 => x"8938ff17",
         11744 => x"5776dd38",
         11745 => x"76597719",
         11746 => x"56807623",
         11747 => x"76802efe",
         11748 => x"c7388078",
         11749 => x"227083ff",
         11750 => x"ff067258",
         11751 => x"5d55567a",
         11752 => x"a02e82e6",
         11753 => x"387383ff",
         11754 => x"ff065372",
         11755 => x"ae2e82f1",
         11756 => x"3876802e",
         11757 => x"aa387719",
         11758 => x"fe057022",
         11759 => x"5a5478ae",
         11760 => x"2e9d3876",
         11761 => x"1018fe05",
         11762 => x"54ff1757",
         11763 => x"76802e8f",
         11764 => x"38fe1470",
         11765 => x"225e547c",
         11766 => x"ae2e0981",
         11767 => x"06eb388b",
         11768 => x"0ba01d55",
         11769 => x"53a07470",
         11770 => x"81055634",
         11771 => x"ff135372",
         11772 => x"f4387273",
         11773 => x"5c5e8878",
         11774 => x"16702281",
         11775 => x"19595754",
         11776 => x"5d74802e",
         11777 => x"80ed3874",
         11778 => x"a02e83d0",
         11779 => x"3874ae32",
         11780 => x"70307080",
         11781 => x"25555a54",
         11782 => x"75772e85",
         11783 => x"ce387283",
         11784 => x"bb387259",
         11785 => x"7c7b2683",
         11786 => x"38815975",
         11787 => x"77327030",
         11788 => x"70720780",
         11789 => x"25707c07",
         11790 => x"51515454",
         11791 => x"72802e83",
         11792 => x"e0387c8b",
         11793 => x"2e868338",
         11794 => x"75772e8a",
         11795 => x"38798307",
         11796 => x"5a757726",
         11797 => x"9e387656",
         11798 => x"885b8b7e",
         11799 => x"822b81fc",
         11800 => x"06771857",
         11801 => x"5f5d7715",
         11802 => x"70228118",
         11803 => x"58565374",
         11804 => x"ff9538a0",
         11805 => x"1c335776",
         11806 => x"81e52e83",
         11807 => x"84387c88",
         11808 => x"2e82e338",
         11809 => x"7d8c0658",
         11810 => x"778c2e82",
         11811 => x"ed387d83",
         11812 => x"06557483",
         11813 => x"2e82e338",
         11814 => x"79812a81",
         11815 => x"0656759d",
         11816 => x"387d8106",
         11817 => x"5d7c802e",
         11818 => x"85387990",
         11819 => x"075a7d82",
         11820 => x"2a81065e",
         11821 => x"7d802e85",
         11822 => x"38798807",
         11823 => x"5a79ab1d",
         11824 => x"347b51e4",
         11825 => x"ec3f84b9",
         11826 => x"c808ab1d",
         11827 => x"33565484",
         11828 => x"b9c80880",
         11829 => x"2e81ac38",
         11830 => x"84b9c808",
         11831 => x"842e0981",
         11832 => x"06fbf738",
         11833 => x"74852a81",
         11834 => x"065a7980",
         11835 => x"2e84f038",
         11836 => x"74822a81",
         11837 => x"06597882",
         11838 => x"98387b08",
         11839 => x"65555673",
         11840 => x"428c1608",
         11841 => x"588057f9",
         11842 => x"ce398116",
         11843 => x"70117911",
         11844 => x"70224040",
         11845 => x"56567ca0",
         11846 => x"2ef03875",
         11847 => x"802efd85",
         11848 => x"38798307",
         11849 => x"5afd8a39",
         11850 => x"82182256",
         11851 => x"75ae2e09",
         11852 => x"8106fcac",
         11853 => x"38772254",
         11854 => x"73ae2e09",
         11855 => x"8106fca0",
         11856 => x"38761018",
         11857 => x"5b807b23",
         11858 => x"800ba01d",
         11859 => x"5653ae54",
         11860 => x"76732683",
         11861 => x"38a05473",
         11862 => x"75708105",
         11863 => x"57348113",
         11864 => x"538a7327",
         11865 => x"e93879a0",
         11866 => x"075877ab",
         11867 => x"1d347b51",
         11868 => x"e3bf3f84",
         11869 => x"b9c808ab",
         11870 => x"1d335654",
         11871 => x"84b9c808",
         11872 => x"fed63874",
         11873 => x"822a8106",
         11874 => x"5877face",
         11875 => x"38861c33",
         11876 => x"70842a81",
         11877 => x"06565d74",
         11878 => x"802e83cd",
         11879 => x"38901c08",
         11880 => x"83ff0660",
         11881 => x"0580d311",
         11882 => x"3380d212",
         11883 => x"3371882b",
         11884 => x"07623341",
         11885 => x"5754547d",
         11886 => x"832e82d8",
         11887 => x"3874881d",
         11888 => x"0c7b0865",
         11889 => x"5556feb7",
         11890 => x"39772255",
         11891 => x"74ae2efe",
         11892 => x"f0387617",
         11893 => x"5976fb88",
         11894 => x"38fbab39",
         11895 => x"79830776",
         11896 => x"17565afd",
         11897 => x"81397d82",
         11898 => x"2b81fc06",
         11899 => x"708c0659",
         11900 => x"5e778c2e",
         11901 => x"098106fd",
         11902 => x"95387982",
         11903 => x"075afd98",
         11904 => x"39850ba0",
         11905 => x"1d347c88",
         11906 => x"2e098106",
         11907 => x"fcf638d6",
         11908 => x"39ff800b",
         11909 => x"ab1d3480",
         11910 => x"0b84b9c8",
         11911 => x"0c933d0d",
         11912 => x"047480ff",
         11913 => x"269d3881",
         11914 => x"ff752780",
         11915 => x"c938ff1d",
         11916 => x"59787b26",
         11917 => x"81f73879",
         11918 => x"83077d77",
         11919 => x"18575c5a",
         11920 => x"fca43979",
         11921 => x"82075a83",
         11922 => x"b5527451",
         11923 => x"8185f63f",
         11924 => x"84b9c808",
         11925 => x"83ffff06",
         11926 => x"70872a81",
         11927 => x"065a5578",
         11928 => x"802ec438",
         11929 => x"7480ff06",
         11930 => x"83e5d811",
         11931 => x"33565474",
         11932 => x"81ff26ff",
         11933 => x"b9387480",
         11934 => x"2e818538",
         11935 => x"83e4f00b",
         11936 => x"83e4f033",
         11937 => x"7081ff06",
         11938 => x"56545973",
         11939 => x"802e80e0",
         11940 => x"3873752e",
         11941 => x"8f388119",
         11942 => x"70337081",
         11943 => x"ff065654",
         11944 => x"5973ee38",
         11945 => x"7281ff06",
         11946 => x"597880d4",
         11947 => x"38ffbf15",
         11948 => x"54739926",
         11949 => x"8a387d82",
         11950 => x"077081ff",
         11951 => x"065f53ff",
         11952 => x"9f155978",
         11953 => x"99269338",
         11954 => x"7d810770",
         11955 => x"81ff06e0",
         11956 => x"177083ff",
         11957 => x"ff065856",
         11958 => x"5f537b1b",
         11959 => x"a0055974",
         11960 => x"7934811b",
         11961 => x"5b751655",
         11962 => x"fafc3980",
         11963 => x"53fab339",
         11964 => x"83e4f033",
         11965 => x"7081ff06",
         11966 => x"5a537880",
         11967 => x"2effae38",
         11968 => x"80df7a83",
         11969 => x"077d1da0",
         11970 => x"055b5b55",
         11971 => x"74793481",
         11972 => x"1b5bd239",
         11973 => x"80cd1433",
         11974 => x"80cc1533",
         11975 => x"71982b71",
         11976 => x"902b0777",
         11977 => x"07881f0c",
         11978 => x"5a57fd95",
         11979 => x"397b1ba0",
         11980 => x"0575882a",
         11981 => x"54547274",
         11982 => x"34811b7c",
         11983 => x"11a0055a",
         11984 => x"5b747934",
         11985 => x"811b5bff",
         11986 => x"9c397983",
         11987 => x"07a01d33",
         11988 => x"585a7681",
         11989 => x"e52e0981",
         11990 => x"06faa338",
         11991 => x"fda33974",
         11992 => x"822a8106",
         11993 => x"5c7bf6f2",
         11994 => x"38850b84",
         11995 => x"b9c80c93",
         11996 => x"3d0d04eb",
         11997 => x"3d0d6769",
         11998 => x"02880580",
         11999 => x"e7053342",
         12000 => x"425e8061",
         12001 => x"0cff7e08",
         12002 => x"70595b42",
         12003 => x"79802e85",
         12004 => x"d7387970",
         12005 => x"81055b33",
         12006 => x"709f2656",
         12007 => x"5675ba2e",
         12008 => x"85d03874",
         12009 => x"ed3875ba",
         12010 => x"2e85c738",
         12011 => x"84d1a433",
         12012 => x"56807624",
         12013 => x"85b23875",
         12014 => x"101084d1",
         12015 => x"90057008",
         12016 => x"585a8c58",
         12017 => x"76802e85",
         12018 => x"96387661",
         12019 => x"0c7f81fe",
         12020 => x"0677335d",
         12021 => x"597b802e",
         12022 => x"9b388117",
         12023 => x"3351ffbb",
         12024 => x"b03f84b9",
         12025 => x"c80881ff",
         12026 => x"06708106",
         12027 => x"5e587c80",
         12028 => x"2e869638",
         12029 => x"80773475",
         12030 => x"165d84b9",
         12031 => x"bc1d3381",
         12032 => x"18348152",
         12033 => x"81173351",
         12034 => x"ffbba43f",
         12035 => x"84b9c808",
         12036 => x"81ff0670",
         12037 => x"81064156",
         12038 => x"83587f84",
         12039 => x"c2387880",
         12040 => x"2e8d3875",
         12041 => x"822a8106",
         12042 => x"418a5860",
         12043 => x"84b13880",
         12044 => x"5b7a8318",
         12045 => x"34ff0bb4",
         12046 => x"180c7a7b",
         12047 => x"5a558154",
         12048 => x"7a53b817",
         12049 => x"70538118",
         12050 => x"335258ff",
         12051 => x"bb953f84",
         12052 => x"b9c8087b",
         12053 => x"2e8538ff",
         12054 => x"55815974",
         12055 => x"b4180c84",
         12056 => x"56789938",
         12057 => x"84b71733",
         12058 => x"84b61833",
         12059 => x"71882b07",
         12060 => x"56568356",
         12061 => x"7482d4d5",
         12062 => x"2e85a538",
         12063 => x"7581268b",
         12064 => x"3884b9bd",
         12065 => x"1d334261",
         12066 => x"85bf3881",
         12067 => x"5875842e",
         12068 => x"83cd388d",
         12069 => x"58758126",
         12070 => x"83c53880",
         12071 => x"c4173380",
         12072 => x"c3183371",
         12073 => x"882b075e",
         12074 => x"597c8480",
         12075 => x"2e098106",
         12076 => x"83ad3880",
         12077 => x"cf173380",
         12078 => x"ce183371",
         12079 => x"882b0757",
         12080 => x"5a75a438",
         12081 => x"80dc1783",
         12082 => x"11338212",
         12083 => x"3371902b",
         12084 => x"71882b07",
         12085 => x"81143370",
         12086 => x"7207882b",
         12087 => x"75337107",
         12088 => x"565a4543",
         12089 => x"5e5f5675",
         12090 => x"a0180c80",
         12091 => x"c8173382",
         12092 => x"183480c8",
         12093 => x"1733ff11",
         12094 => x"7081ff06",
         12095 => x"5f40598d",
         12096 => x"587c8126",
         12097 => x"82d93878",
         12098 => x"81ff0676",
         12099 => x"712980c5",
         12100 => x"19335a5f",
         12101 => x"5a778a18",
         12102 => x"23775977",
         12103 => x"802e87c4",
         12104 => x"38ff1878",
         12105 => x"06426187",
         12106 => x"bb3880ca",
         12107 => x"173380c9",
         12108 => x"18337188",
         12109 => x"2b075640",
         12110 => x"74881823",
         12111 => x"74758f06",
         12112 => x"5e5a8d58",
         12113 => x"7c829838",
         12114 => x"80cc1733",
         12115 => x"80cb1833",
         12116 => x"71882b07",
         12117 => x"565c74a4",
         12118 => x"3880d817",
         12119 => x"83113382",
         12120 => x"12337190",
         12121 => x"2b71882b",
         12122 => x"07811433",
         12123 => x"70720788",
         12124 => x"2b753371",
         12125 => x"0753445a",
         12126 => x"58424242",
         12127 => x"80c71733",
         12128 => x"80c61833",
         12129 => x"71882b07",
         12130 => x"5d588d58",
         12131 => x"7b802e81",
         12132 => x"ce387d1c",
         12133 => x"7a842a05",
         12134 => x"5a797526",
         12135 => x"81c13878",
         12136 => x"52747a31",
         12137 => x"51fdedfd",
         12138 => x"3f84b9c8",
         12139 => x"085684b9",
         12140 => x"c808802e",
         12141 => x"81a93884",
         12142 => x"b9c80880",
         12143 => x"fffffff5",
         12144 => x"26833883",
         12145 => x"5d7583ff",
         12146 => x"f5268338",
         12147 => x"825d759f",
         12148 => x"f52685eb",
         12149 => x"38815d82",
         12150 => x"16709c19",
         12151 => x"0c7ba419",
         12152 => x"0c7b1d70",
         12153 => x"a81a0c7b",
         12154 => x"1db01a0c",
         12155 => x"57597c83",
         12156 => x"2e8a8738",
         12157 => x"8817225c",
         12158 => x"8d587b80",
         12159 => x"2e80e038",
         12160 => x"7d16ac18",
         12161 => x"0c781955",
         12162 => x"7c822e8d",
         12163 => x"38781019",
         12164 => x"70812a7a",
         12165 => x"81060556",
         12166 => x"5a83ff15",
         12167 => x"892a598d",
         12168 => x"5878a018",
         12169 => x"0826b838",
         12170 => x"ff0b9418",
         12171 => x"0cff0b90",
         12172 => x"180cff80",
         12173 => x"0b841834",
         12174 => x"7c832e86",
         12175 => x"96387c77",
         12176 => x"3484d1a0",
         12177 => x"2281055d",
         12178 => x"7c84d1a0",
         12179 => x"237c8618",
         12180 => x"2384d1a8",
         12181 => x"0b8c180c",
         12182 => x"800b9818",
         12183 => x"0c805877",
         12184 => x"84b9c80c",
         12185 => x"973d0d04",
         12186 => x"8b0b84b9",
         12187 => x"c80c973d",
         12188 => x"0d047633",
         12189 => x"d0117081",
         12190 => x"ff065757",
         12191 => x"58748926",
         12192 => x"91388217",
         12193 => x"7881ff06",
         12194 => x"d0055d59",
         12195 => x"787a2e87",
         12196 => x"fe38807e",
         12197 => x"0883e5b8",
         12198 => x"5f405c7c",
         12199 => x"087f5a5b",
         12200 => x"7a708105",
         12201 => x"5c337970",
         12202 => x"81055b33",
         12203 => x"ff9f125a",
         12204 => x"58567799",
         12205 => x"268938e0",
         12206 => x"167081ff",
         12207 => x"065755ff",
         12208 => x"9f175877",
         12209 => x"99268938",
         12210 => x"e0177081",
         12211 => x"ff065855",
         12212 => x"7530709f",
         12213 => x"2a595575",
         12214 => x"772e0981",
         12215 => x"06853877",
         12216 => x"ffbe3878",
         12217 => x"7a327030",
         12218 => x"7072079f",
         12219 => x"2a7a075d",
         12220 => x"58557a80",
         12221 => x"2e879838",
         12222 => x"811c841e",
         12223 => x"5e5c837c",
         12224 => x"25ff9838",
         12225 => x"6156f9a9",
         12226 => x"3978802e",
         12227 => x"fecf3877",
         12228 => x"822a8106",
         12229 => x"5e8a587d",
         12230 => x"fec53880",
         12231 => x"58fec039",
         12232 => x"7a783357",
         12233 => x"597581e9",
         12234 => x"2e098106",
         12235 => x"83388159",
         12236 => x"7581eb32",
         12237 => x"70307080",
         12238 => x"257b075a",
         12239 => x"5b5c7783",
         12240 => x"ad387581",
         12241 => x"e82e83a6",
         12242 => x"38933d77",
         12243 => x"575a8359",
         12244 => x"83fa1633",
         12245 => x"70595b7a",
         12246 => x"802ea538",
         12247 => x"84811633",
         12248 => x"84801733",
         12249 => x"71902b71",
         12250 => x"882b0783",
         12251 => x"ff193370",
         12252 => x"7207882b",
         12253 => x"83fe1b33",
         12254 => x"71075259",
         12255 => x"5b404040",
         12256 => x"777a7084",
         12257 => x"055c0cff",
         12258 => x"19901757",
         12259 => x"59788025",
         12260 => x"ffbe3884",
         12261 => x"b9bd1d33",
         12262 => x"7030709f",
         12263 => x"2a727131",
         12264 => x"9b3d7110",
         12265 => x"1005f005",
         12266 => x"84b61c44",
         12267 => x"5d52435b",
         12268 => x"4278085b",
         12269 => x"83567a80",
         12270 => x"2e80fb38",
         12271 => x"800b8318",
         12272 => x"34ff0bb4",
         12273 => x"180c7a55",
         12274 => x"80567aff",
         12275 => x"2ea53881",
         12276 => x"547a53b8",
         12277 => x"17528117",
         12278 => x"3351ffb4",
         12279 => x"863f84b9",
         12280 => x"c808762e",
         12281 => x"8538ff55",
         12282 => x"815674b4",
         12283 => x"180c8458",
         12284 => x"75bf3881",
         12285 => x"1f337f33",
         12286 => x"71882b07",
         12287 => x"5d5e8358",
         12288 => x"7b82d4d5",
         12289 => x"2e098106",
         12290 => x"a838800b",
         12291 => x"b8183357",
         12292 => x"587581e9",
         12293 => x"2e82b738",
         12294 => x"7581eb32",
         12295 => x"70307080",
         12296 => x"257a0742",
         12297 => x"42427fbc",
         12298 => x"387581e8",
         12299 => x"2eb63882",
         12300 => x"587781ff",
         12301 => x"0656800b",
         12302 => x"84b9bd1e",
         12303 => x"335d587b",
         12304 => x"782e0981",
         12305 => x"06833881",
         12306 => x"58817627",
         12307 => x"f8bd3877",
         12308 => x"802ef8b7",
         12309 => x"38811a84",
         12310 => x"1a5a5a83",
         12311 => x"7a27fed1",
         12312 => x"38f8a839",
         12313 => x"830b80ee",
         12314 => x"1883e4f8",
         12315 => x"405d587b",
         12316 => x"7081055d",
         12317 => x"337e7081",
         12318 => x"05403371",
         12319 => x"7131ff1b",
         12320 => x"5b525656",
         12321 => x"77802e80",
         12322 => x"c5387580",
         12323 => x"2ee13885",
         12324 => x"0b818a18",
         12325 => x"83e4fc40",
         12326 => x"5d587b70",
         12327 => x"81055d33",
         12328 => x"7e708105",
         12329 => x"40337171",
         12330 => x"31ff1b5b",
         12331 => x"58424077",
         12332 => x"802e858e",
         12333 => x"3875802e",
         12334 => x"e1388258",
         12335 => x"fef3398d",
         12336 => x"587cfa93",
         12337 => x"387784b9",
         12338 => x"c80c973d",
         12339 => x"0d047558",
         12340 => x"75802efe",
         12341 => x"dc38850b",
         12342 => x"818a1883",
         12343 => x"e4fc405d",
         12344 => x"58ffb739",
         12345 => x"8d0b84b9",
         12346 => x"c80c973d",
         12347 => x"0d04830b",
         12348 => x"80ee1883",
         12349 => x"e4f85c5a",
         12350 => x"58787081",
         12351 => x"055a337a",
         12352 => x"7081055c",
         12353 => x"33717131",
         12354 => x"ff1b5b57",
         12355 => x"5f5f7780",
         12356 => x"2e83d138",
         12357 => x"74802ee1",
         12358 => x"38850b81",
         12359 => x"8a1883e4",
         12360 => x"fc5c5a58",
         12361 => x"78708105",
         12362 => x"5a337a70",
         12363 => x"81055c33",
         12364 => x"717131ff",
         12365 => x"1b5b5842",
         12366 => x"4077802e",
         12367 => x"84913875",
         12368 => x"802ee138",
         12369 => x"933d7757",
         12370 => x"5a8359fc",
         12371 => x"83398158",
         12372 => x"fdc63980",
         12373 => x"e9173380",
         12374 => x"e8183371",
         12375 => x"882b0757",
         12376 => x"5575812e",
         12377 => x"098106f9",
         12378 => x"d538811b",
         12379 => x"58805ab4",
         12380 => x"1708782e",
         12381 => x"b1388317",
         12382 => x"335b7a7a",
         12383 => x"2e098106",
         12384 => x"829b3881",
         12385 => x"547753b8",
         12386 => x"17528117",
         12387 => x"3351ffb0",
         12388 => x"d23f84b9",
         12389 => x"c808802e",
         12390 => x"8538ff58",
         12391 => x"815a77b4",
         12392 => x"180c79f9",
         12393 => x"99387984",
         12394 => x"183484b7",
         12395 => x"173384b6",
         12396 => x"18337188",
         12397 => x"2b07575e",
         12398 => x"7582d4d5",
         12399 => x"2e098106",
         12400 => x"f8fc38b8",
         12401 => x"17831133",
         12402 => x"82123371",
         12403 => x"902b7188",
         12404 => x"2b078114",
         12405 => x"33707207",
         12406 => x"882b7533",
         12407 => x"71075e41",
         12408 => x"5945425c",
         12409 => x"5977848b",
         12410 => x"85a4d22e",
         12411 => x"098106f8",
         12412 => x"cd38849c",
         12413 => x"17831133",
         12414 => x"82123371",
         12415 => x"902b7188",
         12416 => x"2b078114",
         12417 => x"33707207",
         12418 => x"882b7533",
         12419 => x"71074744",
         12420 => x"405b5c5a",
         12421 => x"5e60868a",
         12422 => x"85e4f22e",
         12423 => x"098106f8",
         12424 => x"9d3884a0",
         12425 => x"17831133",
         12426 => x"82123371",
         12427 => x"902b7188",
         12428 => x"2b078114",
         12429 => x"33707207",
         12430 => x"882b7533",
         12431 => x"7107941e",
         12432 => x"0c5d84a4",
         12433 => x"1c831133",
         12434 => x"82123371",
         12435 => x"902b7188",
         12436 => x"2b078114",
         12437 => x"33707207",
         12438 => x"882b7533",
         12439 => x"71076290",
         12440 => x"050c5944",
         12441 => x"49465c45",
         12442 => x"40455b56",
         12443 => x"5a7c7734",
         12444 => x"84d1a022",
         12445 => x"81055d7c",
         12446 => x"84d1a023",
         12447 => x"7c861823",
         12448 => x"84d1a80b",
         12449 => x"8c180c80",
         12450 => x"0b98180c",
         12451 => x"f7cf397b",
         12452 => x"8324f8f0",
         12453 => x"387b7a7f",
         12454 => x"0c56f295",
         12455 => x"397554b4",
         12456 => x"170853b8",
         12457 => x"17705381",
         12458 => x"18335259",
         12459 => x"ffafb33f",
         12460 => x"84b9c808",
         12461 => x"7a2e0981",
         12462 => x"0681a438",
         12463 => x"84b9c808",
         12464 => x"831834b4",
         12465 => x"1708a818",
         12466 => x"0831407f",
         12467 => x"a0180827",
         12468 => x"8b388217",
         12469 => x"33416082",
         12470 => x"2e818d38",
         12471 => x"84b9c808",
         12472 => x"5afda039",
         12473 => x"74567480",
         12474 => x"2ef39138",
         12475 => x"850b818a",
         12476 => x"1883e4fc",
         12477 => x"5c5a58fc",
         12478 => x"ab3980e3",
         12479 => x"173380e2",
         12480 => x"18337188",
         12481 => x"2b075f5a",
         12482 => x"8d587df6",
         12483 => x"d2388817",
         12484 => x"224261f6",
         12485 => x"ca3880e4",
         12486 => x"17831133",
         12487 => x"82123371",
         12488 => x"902b7188",
         12489 => x"2b078114",
         12490 => x"33707207",
         12491 => x"882b7533",
         12492 => x"7107ac1e",
         12493 => x"0c5a7d82",
         12494 => x"2b5a4344",
         12495 => x"405940f5",
         12496 => x"d8397558",
         12497 => x"75802ef9",
         12498 => x"e8388258",
         12499 => x"f9e33975",
         12500 => x"802ef2a8",
         12501 => x"38933d77",
         12502 => x"575a8359",
         12503 => x"f7f23975",
         12504 => x"5a79f5da",
         12505 => x"38fcbf39",
         12506 => x"7554b417",
         12507 => x"08a01808",
         12508 => x"05537852",
         12509 => x"81173351",
         12510 => x"ffade73f",
         12511 => x"fc8539f0",
         12512 => x"3d0d0280",
         12513 => x"d3053364",
         12514 => x"7043933d",
         12515 => x"41575dff",
         12516 => x"765a4075",
         12517 => x"802e80e9",
         12518 => x"38787081",
         12519 => x"055a3370",
         12520 => x"9f265555",
         12521 => x"74ba2e80",
         12522 => x"e23873ed",
         12523 => x"3874ba2e",
         12524 => x"80d93884",
         12525 => x"d1a43354",
         12526 => x"80742480",
         12527 => x"c4387310",
         12528 => x"1084d190",
         12529 => x"05700855",
         12530 => x"5573802e",
         12531 => x"84388074",
         12532 => x"34625473",
         12533 => x"802e8638",
         12534 => x"80743462",
         12535 => x"5473750c",
         12536 => x"7c547c80",
         12537 => x"2e923880",
         12538 => x"53933d70",
         12539 => x"53840551",
         12540 => x"ef813f84",
         12541 => x"b9c80854",
         12542 => x"7384b9c8",
         12543 => x"0c923d0d",
         12544 => x"048b0b84",
         12545 => x"b9c80c92",
         12546 => x"3d0d0475",
         12547 => x"33d01170",
         12548 => x"81ff0656",
         12549 => x"56577389",
         12550 => x"26913882",
         12551 => x"167781ff",
         12552 => x"06d0055c",
         12553 => x"5877792e",
         12554 => x"80f73880",
         12555 => x"7f0883e5",
         12556 => x"b85e5f5b",
         12557 => x"7b087e59",
         12558 => x"5a797081",
         12559 => x"055b3378",
         12560 => x"7081055a",
         12561 => x"33ff9f12",
         12562 => x"59575576",
         12563 => x"99268938",
         12564 => x"e0157081",
         12565 => x"ff065654",
         12566 => x"ff9f1657",
         12567 => x"76992689",
         12568 => x"38e01670",
         12569 => x"81ff0657",
         12570 => x"54743070",
         12571 => x"9f2a5854",
         12572 => x"74762e09",
         12573 => x"81068538",
         12574 => x"76ffbe38",
         12575 => x"77793270",
         12576 => x"30707207",
         12577 => x"9f2a7907",
         12578 => x"5c575479",
         12579 => x"802e9238",
         12580 => x"811b841d",
         12581 => x"5d5b837b",
         12582 => x"25ff9938",
         12583 => x"7f54fe98",
         12584 => x"397a8324",
         12585 => x"f7387a79",
         12586 => x"600c54fe",
         12587 => x"8b39e63d",
         12588 => x"0d6c0284",
         12589 => x"0580fb05",
         12590 => x"33565989",
         12591 => x"5678802e",
         12592 => x"a63874bf",
         12593 => x"0670549d",
         12594 => x"3dcc0553",
         12595 => x"9e3d8405",
         12596 => x"5258ed9f",
         12597 => x"3f84b9c8",
         12598 => x"085784b9",
         12599 => x"c808802e",
         12600 => x"8f388079",
         12601 => x"0c765675",
         12602 => x"84b9c80c",
         12603 => x"9c3d0d04",
         12604 => x"7e406d52",
         12605 => x"903d7052",
         12606 => x"5ae19a3f",
         12607 => x"84b9c808",
         12608 => x"5784b9c8",
         12609 => x"08802e81",
         12610 => x"ba38779c",
         12611 => x"065d7c80",
         12612 => x"2e81ca38",
         12613 => x"76802e83",
         12614 => x"c1387684",
         12615 => x"2e83ea38",
         12616 => x"77880758",
         12617 => x"76ffbb38",
         12618 => x"77832a81",
         12619 => x"065b7a80",
         12620 => x"2e81d138",
         12621 => x"669b1133",
         12622 => x"9a123371",
         12623 => x"882b0761",
         12624 => x"70334258",
         12625 => x"5e5e567d",
         12626 => x"832e84e9",
         12627 => x"38800b8e",
         12628 => x"1734800b",
         12629 => x"8f1734a1",
         12630 => x"0b901734",
         12631 => x"80cc0b91",
         12632 => x"17346656",
         12633 => x"a00b8b17",
         12634 => x"347e6757",
         12635 => x"5e800b9a",
         12636 => x"1734800b",
         12637 => x"9b17347d",
         12638 => x"335d7c83",
         12639 => x"2e84a938",
         12640 => x"665b800b",
         12641 => x"9c1c3480",
         12642 => x"0b9d1c34",
         12643 => x"800b9e1c",
         12644 => x"34800b9f",
         12645 => x"1c347e55",
         12646 => x"810b8316",
         12647 => x"347b802e",
         12648 => x"80e2387e",
         12649 => x"b411087d",
         12650 => x"7c085357",
         12651 => x"5f57817c",
         12652 => x"2789389c",
         12653 => x"17087c26",
         12654 => x"838a3882",
         12655 => x"5780790c",
         12656 => x"fea33902",
         12657 => x"80e70533",
         12658 => x"70982b5d",
         12659 => x"5b7b8025",
         12660 => x"feb83886",
         12661 => x"789c065e",
         12662 => x"577cfeb8",
         12663 => x"3876fe82",
         12664 => x"380280c2",
         12665 => x"05337084",
         12666 => x"2a81065d",
         12667 => x"567b8291",
         12668 => x"3877812a",
         12669 => x"81065e7d",
         12670 => x"802e8938",
         12671 => x"7581065a",
         12672 => x"7981f638",
         12673 => x"77832a81",
         12674 => x"06567580",
         12675 => x"2e863877",
         12676 => x"80c00758",
         12677 => x"7eb41108",
         12678 => x"a01b0c67",
         12679 => x"a41b0c67",
         12680 => x"9b11339a",
         12681 => x"12337188",
         12682 => x"2b077333",
         12683 => x"405e4057",
         12684 => x"5a7b832e",
         12685 => x"81f1387a",
         12686 => x"881a0c9c",
         12687 => x"16831133",
         12688 => x"82123371",
         12689 => x"902b7188",
         12690 => x"2b078114",
         12691 => x"33707207",
         12692 => x"882b7533",
         12693 => x"71077060",
         12694 => x"8c050c60",
         12695 => x"600c5152",
         12696 => x"4159575d",
         12697 => x"5e861a22",
         12698 => x"841a2377",
         12699 => x"901a3480",
         12700 => x"0b911a34",
         12701 => x"800b9c1a",
         12702 => x"0c77852a",
         12703 => x"81065574",
         12704 => x"802e84ac",
         12705 => x"3875802e",
         12706 => x"84f13875",
         12707 => x"941a0c8a",
         12708 => x"1a227089",
         12709 => x"2b7c525b",
         12710 => x"58763070",
         12711 => x"78078025",
         12712 => x"565b7976",
         12713 => x"27849238",
         12714 => x"81707606",
         12715 => x"5f5b7d80",
         12716 => x"2e848638",
         12717 => x"77527851",
         12718 => x"ffacdb3f",
         12719 => x"84b9c808",
         12720 => x"5884b9c8",
         12721 => x"08812683",
         12722 => x"38825784",
         12723 => x"b9c808ff",
         12724 => x"2e80cb38",
         12725 => x"757a3156",
         12726 => x"c0390280",
         12727 => x"c2053391",
         12728 => x"065e7d95",
         12729 => x"3877822a",
         12730 => x"81065574",
         12731 => x"802efcb8",
         12732 => x"38885780",
         12733 => x"790cfbed",
         12734 => x"39875780",
         12735 => x"790cfbe5",
         12736 => x"39845780",
         12737 => x"790cfbdd",
         12738 => x"397951cd",
         12739 => x"ca3f84b9",
         12740 => x"c8087888",
         12741 => x"07595776",
         12742 => x"fbc838fc",
         12743 => x"8b397a76",
         12744 => x"7b315757",
         12745 => x"fef33995",
         12746 => x"16339417",
         12747 => x"3371982b",
         12748 => x"71902b07",
         12749 => x"7d075d5e",
         12750 => x"5cfdfc39",
         12751 => x"7c557c7b",
         12752 => x"2781bd38",
         12753 => x"74527951",
         12754 => x"ffabcb3f",
         12755 => x"84b9c808",
         12756 => x"5d84b9c8",
         12757 => x"08802e81",
         12758 => x"a73884b9",
         12759 => x"c808812e",
         12760 => x"fcd93884",
         12761 => x"b9c808ff",
         12762 => x"2e839938",
         12763 => x"80537452",
         12764 => x"7651ffb2",
         12765 => x"823f84b9",
         12766 => x"c8088390",
         12767 => x"389c1708",
         12768 => x"fe119419",
         12769 => x"0858565b",
         12770 => x"757527ff",
         12771 => x"af388116",
         12772 => x"94180c84",
         12773 => x"17338107",
         12774 => x"55748418",
         12775 => x"347c557a",
         12776 => x"7d26ffa0",
         12777 => x"3880d939",
         12778 => x"800b9417",
         12779 => x"34800b95",
         12780 => x"1734fbcc",
         12781 => x"39951633",
         12782 => x"94173371",
         12783 => x"982b7190",
         12784 => x"2b077e07",
         12785 => x"5e565b80",
         12786 => x"0b8e1734",
         12787 => x"800b8f17",
         12788 => x"34a10b90",
         12789 => x"173480cc",
         12790 => x"0b911734",
         12791 => x"6656a00b",
         12792 => x"8b17347e",
         12793 => x"67575e80",
         12794 => x"0b9a1734",
         12795 => x"800b9b17",
         12796 => x"347d335d",
         12797 => x"7c832e09",
         12798 => x"8106fb84",
         12799 => x"38ffa939",
         12800 => x"807f7f72",
         12801 => x"5e59575d",
         12802 => x"b416087e",
         12803 => x"2eae3883",
         12804 => x"16335a79",
         12805 => x"7d2e0981",
         12806 => x"06b53881",
         12807 => x"547d53b8",
         12808 => x"16528116",
         12809 => x"3351ffa3",
         12810 => x"ba3f84b9",
         12811 => x"c808802e",
         12812 => x"8538ff57",
         12813 => x"815b76b4",
         12814 => x"170c7e56",
         12815 => x"7aff1d90",
         12816 => x"180c577a",
         12817 => x"802efbbc",
         12818 => x"3880790c",
         12819 => x"f9973981",
         12820 => x"54b41608",
         12821 => x"53b81670",
         12822 => x"53811733",
         12823 => x"525affa4",
         12824 => x"813f84b9",
         12825 => x"c8087d2e",
         12826 => x"09810681",
         12827 => x"aa3884b9",
         12828 => x"c8088317",
         12829 => x"34b41608",
         12830 => x"a8170831",
         12831 => x"84b9c808",
         12832 => x"5c5574a0",
         12833 => x"170827ff",
         12834 => x"92388216",
         12835 => x"33557482",
         12836 => x"2e098106",
         12837 => x"ff853881",
         12838 => x"54b41608",
         12839 => x"a0170805",
         12840 => x"53795281",
         12841 => x"163351ff",
         12842 => x"a3b83f7c",
         12843 => x"5bfeec39",
         12844 => x"74941a0c",
         12845 => x"7656f8af",
         12846 => x"3977981a",
         12847 => x"0c76f8a2",
         12848 => x"387583ff",
         12849 => x"065a7980",
         12850 => x"2ef89a38",
         12851 => x"7efe199c",
         12852 => x"1208fe05",
         12853 => x"5f595a77",
         12854 => x"7d27f9df",
         12855 => x"388a1a22",
         12856 => x"787129b0",
         12857 => x"1c080556",
         12858 => x"5c74802e",
         12859 => x"f9cd3875",
         12860 => x"892a159c",
         12861 => x"1a0c7656",
         12862 => x"f7ed3975",
         12863 => x"941a0c76",
         12864 => x"56f7e439",
         12865 => x"81578079",
         12866 => x"0cf7da39",
         12867 => x"84b9c808",
         12868 => x"5780790c",
         12869 => x"f7cf3981",
         12870 => x"7f575bfe",
         12871 => x"9f39f03d",
         12872 => x"0d626567",
         12873 => x"6640405d",
         12874 => x"5a807e0c",
         12875 => x"89577980",
         12876 => x"2e9f3879",
         12877 => x"08567580",
         12878 => x"2e973875",
         12879 => x"33557480",
         12880 => x"2e8f3886",
         12881 => x"1622841b",
         12882 => x"22595978",
         12883 => x"782e84b7",
         12884 => x"38805574",
         12885 => x"41765576",
         12886 => x"828c3891",
         12887 => x"1a335574",
         12888 => x"82843890",
         12889 => x"1a338106",
         12890 => x"57875676",
         12891 => x"802e81ed",
         12892 => x"38941a08",
         12893 => x"8c1b0871",
         12894 => x"3156567b",
         12895 => x"752681ef",
         12896 => x"387b802e",
         12897 => x"81d53860",
         12898 => x"597583ff",
         12899 => x"065b7a81",
         12900 => x"e3388a19",
         12901 => x"22ff0576",
         12902 => x"892a065b",
         12903 => x"7a9b3875",
         12904 => x"83d33888",
         12905 => x"1a085581",
         12906 => x"75278485",
         12907 => x"3874ff2e",
         12908 => x"83f03874",
         12909 => x"981b0c60",
         12910 => x"59981a08",
         12911 => x"fe059c1a",
         12912 => x"08fe0541",
         12913 => x"57766027",
         12914 => x"83e7388a",
         12915 => x"19227078",
         12916 => x"29b01b08",
         12917 => x"05565674",
         12918 => x"802e83d5",
         12919 => x"387a157c",
         12920 => x"892a5957",
         12921 => x"77802e83",
         12922 => x"8138771b",
         12923 => x"55757527",
         12924 => x"8538757b",
         12925 => x"31587754",
         12926 => x"76537c52",
         12927 => x"81193351",
         12928 => x"ff9fe03f",
         12929 => x"84b9c808",
         12930 => x"83983860",
         12931 => x"83113357",
         12932 => x"5975802e",
         12933 => x"a938b419",
         12934 => x"08773156",
         12935 => x"7578279e",
         12936 => x"38848076",
         12937 => x"71291eb8",
         12938 => x"1b585855",
         12939 => x"75708105",
         12940 => x"57337770",
         12941 => x"81055934",
         12942 => x"ff155574",
         12943 => x"ef387789",
         12944 => x"2b587b78",
         12945 => x"317e0819",
         12946 => x"7f0c781e",
         12947 => x"941c081a",
         12948 => x"7059941d",
         12949 => x"0c5e5c7b",
         12950 => x"feaf3880",
         12951 => x"567584b9",
         12952 => x"c80c923d",
         12953 => x"0d047484",
         12954 => x"b9c80c92",
         12955 => x"3d0d0474",
         12956 => x"5cfe8e39",
         12957 => x"9c1a0857",
         12958 => x"7583ff06",
         12959 => x"84807131",
         12960 => x"595b7b78",
         12961 => x"2783387b",
         12962 => x"587656b4",
         12963 => x"1908772e",
         12964 => x"b638800b",
         12965 => x"831a3371",
         12966 => x"5d415f7f",
         12967 => x"7f2e0981",
         12968 => x"0680e438",
         12969 => x"81547653",
         12970 => x"b8195281",
         12971 => x"193351ff",
         12972 => x"9eb13f84",
         12973 => x"b9c80880",
         12974 => x"2e8538ff",
         12975 => x"56815b75",
         12976 => x"b41a0c7a",
         12977 => x"81dc3860",
         12978 => x"941b0883",
         12979 => x"ff061179",
         12980 => x"7f5a58b8",
         12981 => x"05565977",
         12982 => x"802efee6",
         12983 => x"38747081",
         12984 => x"05563377",
         12985 => x"70810559",
         12986 => x"34ff1656",
         12987 => x"75802efe",
         12988 => x"d1387470",
         12989 => x"81055633",
         12990 => x"77708105",
         12991 => x"5934ff16",
         12992 => x"5675da38",
         12993 => x"febc3981",
         12994 => x"54b41908",
         12995 => x"53b81970",
         12996 => x"53811a33",
         12997 => x"5240ff9e",
         12998 => x"c93f815b",
         12999 => x"84b9c808",
         13000 => x"7f2e0981",
         13001 => x"06ff9c38",
         13002 => x"84b9c808",
         13003 => x"831a34b4",
         13004 => x"1908a81a",
         13005 => x"083184b9",
         13006 => x"c8085c55",
         13007 => x"74a01a08",
         13008 => x"27fee138",
         13009 => x"82193355",
         13010 => x"74822e09",
         13011 => x"8106fed4",
         13012 => x"388154b4",
         13013 => x"1908a01a",
         13014 => x"0805537f",
         13015 => x"52811933",
         13016 => x"51ff9dfe",
         13017 => x"3f7e5bfe",
         13018 => x"bb39769c",
         13019 => x"1b0c941a",
         13020 => x"0856fe84",
         13021 => x"39981a08",
         13022 => x"527951ff",
         13023 => x"a3983f84",
         13024 => x"b9c80855",
         13025 => x"fca13981",
         13026 => x"163351ff",
         13027 => x"9c833f84",
         13028 => x"b9c80881",
         13029 => x"065574fb",
         13030 => x"b838747a",
         13031 => x"085657fb",
         13032 => x"b239810b",
         13033 => x"911b3481",
         13034 => x"0b84b9c8",
         13035 => x"0c923d0d",
         13036 => x"04820b91",
         13037 => x"1b34820b",
         13038 => x"84b9c80c",
         13039 => x"923d0d04",
         13040 => x"f03d0d62",
         13041 => x"65676640",
         13042 => x"405c5a80",
         13043 => x"7e0c8957",
         13044 => x"79802e9f",
         13045 => x"38790856",
         13046 => x"75802e97",
         13047 => x"38753355",
         13048 => x"74802e8f",
         13049 => x"38861622",
         13050 => x"841b2259",
         13051 => x"5978782e",
         13052 => x"85fd3880",
         13053 => x"55744176",
         13054 => x"557682c4",
         13055 => x"38911a33",
         13056 => x"557482bc",
         13057 => x"38901a33",
         13058 => x"70812a81",
         13059 => x"06585887",
         13060 => x"5676802e",
         13061 => x"82a13894",
         13062 => x"1a087b11",
         13063 => x"5d577b77",
         13064 => x"27843876",
         13065 => x"095b7a80",
         13066 => x"2e828138",
         13067 => x"7683ff06",
         13068 => x"5f7e82a2",
         13069 => x"38608a11",
         13070 => x"22ff0578",
         13071 => x"892a065a",
         13072 => x"5678aa38",
         13073 => x"76849e38",
         13074 => x"881a0855",
         13075 => x"74802e84",
         13076 => x"b1387481",
         13077 => x"2e86a138",
         13078 => x"74ff2e86",
         13079 => x"8c387498",
         13080 => x"1b0c881a",
         13081 => x"08853874",
         13082 => x"881b0c60",
         13083 => x"56b41608",
         13084 => x"9c1b082e",
         13085 => x"81d33898",
         13086 => x"1a08fe05",
         13087 => x"9c1708fe",
         13088 => x"05585877",
         13089 => x"772785f0",
         13090 => x"388a1622",
         13091 => x"707929b0",
         13092 => x"18080556",
         13093 => x"5774802e",
         13094 => x"85de3878",
         13095 => x"157b892a",
         13096 => x"595c7780",
         13097 => x"2e839838",
         13098 => x"77195f76",
         13099 => x"7f278538",
         13100 => x"76793158",
         13101 => x"77547b53",
         13102 => x"7c528116",
         13103 => x"3351ff9b",
         13104 => x"a13f84b9",
         13105 => x"c80885a1",
         13106 => x"3860b411",
         13107 => x"087d3156",
         13108 => x"57747827",
         13109 => x"a5388480",
         13110 => x"0bb81876",
         13111 => x"72291f57",
         13112 => x"58567470",
         13113 => x"81055633",
         13114 => x"77708105",
         13115 => x"5934ff16",
         13116 => x"5675ef38",
         13117 => x"60597583",
         13118 => x"1a347789",
         13119 => x"2b597a79",
         13120 => x"317e081a",
         13121 => x"7f0c791e",
         13122 => x"941c081b",
         13123 => x"7071941f",
         13124 => x"0c8c1e08",
         13125 => x"5a5a575e",
         13126 => x"5b757527",
         13127 => x"83387456",
         13128 => x"758c1b0c",
         13129 => x"7afe8538",
         13130 => x"901a3358",
         13131 => x"7780c007",
         13132 => x"5b7a901b",
         13133 => x"34805675",
         13134 => x"84b9c80c",
         13135 => x"923d0d04",
         13136 => x"7484b9c8",
         13137 => x"0c923d0d",
         13138 => x"04831633",
         13139 => x"557482c8",
         13140 => x"386056fe",
         13141 => x"a239609c",
         13142 => x"1b085956",
         13143 => x"7683ff06",
         13144 => x"84807131",
         13145 => x"5a5c7a79",
         13146 => x"2783387a",
         13147 => x"597757b4",
         13148 => x"1608782e",
         13149 => x"b638800b",
         13150 => x"83173371",
         13151 => x"5e415f7f",
         13152 => x"7f2e0981",
         13153 => x"0680d538",
         13154 => x"81547753",
         13155 => x"b8165281",
         13156 => x"163351ff",
         13157 => x"98cd3f84",
         13158 => x"b9c80880",
         13159 => x"2e8538ff",
         13160 => x"57815c76",
         13161 => x"b4170c7b",
         13162 => x"83bf3860",
         13163 => x"941b0883",
         13164 => x"ff06117a",
         13165 => x"58b8057e",
         13166 => x"59565878",
         13167 => x"802e9538",
         13168 => x"76708105",
         13169 => x"58337570",
         13170 => x"81055734",
         13171 => x"ff165675",
         13172 => x"ef386058",
         13173 => x"810b8319",
         13174 => x"34fea339",
         13175 => x"8154b416",
         13176 => x"0853b816",
         13177 => x"70538117",
         13178 => x"335240ff",
         13179 => x"98f43f81",
         13180 => x"5c84b9c8",
         13181 => x"087f2e09",
         13182 => x"8106ffab",
         13183 => x"3884b9c8",
         13184 => x"08831734",
         13185 => x"b41608a8",
         13186 => x"17083184",
         13187 => x"b9c8085d",
         13188 => x"5574a017",
         13189 => x"0827fef0",
         13190 => x"38821633",
         13191 => x"5574822e",
         13192 => x"098106fe",
         13193 => x"e3388154",
         13194 => x"b41608a0",
         13195 => x"17080553",
         13196 => x"7f528116",
         13197 => x"3351ff98",
         13198 => x"a93f7e5c",
         13199 => x"feca3994",
         13200 => x"1a08578c",
         13201 => x"1a087726",
         13202 => x"93388316",
         13203 => x"33407f81",
         13204 => x"b938607c",
         13205 => x"b4120c94",
         13206 => x"1b085856",
         13207 => x"7b7c9c1c",
         13208 => x"0c58fdf8",
         13209 => x"39981a08",
         13210 => x"527951ff",
         13211 => x"abe73f84",
         13212 => x"b9c80855",
         13213 => x"84b9c808",
         13214 => x"fbd83890",
         13215 => x"1a3358fd",
         13216 => x"ab397652",
         13217 => x"7951ffab",
         13218 => x"cc3f84b9",
         13219 => x"c8085584",
         13220 => x"b9c808fb",
         13221 => x"bd38e439",
         13222 => x"8154b416",
         13223 => x"0853b816",
         13224 => x"70538117",
         13225 => x"335257ff",
         13226 => x"97b83f84",
         13227 => x"b9c80881",
         13228 => x"b83884b9",
         13229 => x"c8088317",
         13230 => x"34b41608",
         13231 => x"a8170831",
         13232 => x"5877a017",
         13233 => x"0827fd89",
         13234 => x"38821633",
         13235 => x"5c7b822e",
         13236 => x"098106fc",
         13237 => x"fc388154",
         13238 => x"b41608a0",
         13239 => x"17080553",
         13240 => x"76528116",
         13241 => x"3351ff96",
         13242 => x"f93f6056",
         13243 => x"fb893981",
         13244 => x"163351ff",
         13245 => x"959b3f84",
         13246 => x"b9c80881",
         13247 => x"065574f9",
         13248 => x"f238747a",
         13249 => x"085657f9",
         13250 => x"ec398154",
         13251 => x"b4160853",
         13252 => x"b8167053",
         13253 => x"81173352",
         13254 => x"57ff96c6",
         13255 => x"3f84b9c8",
         13256 => x"0880c638",
         13257 => x"84b9c808",
         13258 => x"831734b4",
         13259 => x"1608a817",
         13260 => x"08315574",
         13261 => x"a0170827",
         13262 => x"fe983882",
         13263 => x"16335877",
         13264 => x"822e0981",
         13265 => x"06fe8b38",
         13266 => x"8154b416",
         13267 => x"08a01708",
         13268 => x"05537652",
         13269 => x"81163351",
         13270 => x"ff96873f",
         13271 => x"607cb412",
         13272 => x"0c941b08",
         13273 => x"5856fdf4",
         13274 => x"39810b91",
         13275 => x"1b34810b",
         13276 => x"84b9c80c",
         13277 => x"923d0d04",
         13278 => x"820b911b",
         13279 => x"34820b84",
         13280 => x"b9c80c92",
         13281 => x"3d0d04f5",
         13282 => x"3d0d7d58",
         13283 => x"895a7780",
         13284 => x"2e9f3877",
         13285 => x"08567580",
         13286 => x"2e973875",
         13287 => x"33557480",
         13288 => x"2e8f3886",
         13289 => x"16228419",
         13290 => x"22585978",
         13291 => x"772e83b5",
         13292 => x"38805574",
         13293 => x"5c795679",
         13294 => x"81d83890",
         13295 => x"18337086",
         13296 => x"2a81065c",
         13297 => x"577a802e",
         13298 => x"81c8387b",
         13299 => x"a019085a",
         13300 => x"57b41708",
         13301 => x"792eac38",
         13302 => x"8317335b",
         13303 => x"7a81bc38",
         13304 => x"81547853",
         13305 => x"b8175281",
         13306 => x"173351ff",
         13307 => x"93f53f84",
         13308 => x"b9c80880",
         13309 => x"2e8538ff",
         13310 => x"59815678",
         13311 => x"b4180c75",
         13312 => x"819038a4",
         13313 => x"18088b11",
         13314 => x"33a0075a",
         13315 => x"57788b18",
         13316 => x"34770888",
         13317 => x"19087083",
         13318 => x"ffff065d",
         13319 => x"5a567a9a",
         13320 => x"18347a88",
         13321 => x"2a5a799b",
         13322 => x"18349c17",
         13323 => x"76339619",
         13324 => x"5c565b74",
         13325 => x"832e81c1",
         13326 => x"388c1808",
         13327 => x"55747b34",
         13328 => x"74882a5b",
         13329 => x"7a9d1834",
         13330 => x"74902a56",
         13331 => x"759e1834",
         13332 => x"74982a59",
         13333 => x"789f1834",
         13334 => x"807a3480",
         13335 => x"0b971834",
         13336 => x"a10b9818",
         13337 => x"3480cc0b",
         13338 => x"99183480",
         13339 => x"0b921834",
         13340 => x"800b9318",
         13341 => x"347b5b81",
         13342 => x"0b831c34",
         13343 => x"7b51ff96",
         13344 => x"943f84b9",
         13345 => x"c8089019",
         13346 => x"3381bf06",
         13347 => x"5b567990",
         13348 => x"19347584",
         13349 => x"b9c80c8d",
         13350 => x"3d0d0481",
         13351 => x"54b41708",
         13352 => x"53b81770",
         13353 => x"53811833",
         13354 => x"525bff93",
         13355 => x"b53f8156",
         13356 => x"84b9c808",
         13357 => x"fec93884",
         13358 => x"b9c80883",
         13359 => x"1834b417",
         13360 => x"08a81808",
         13361 => x"3184b9c8",
         13362 => x"08575574",
         13363 => x"a0180827",
         13364 => x"fe8e3882",
         13365 => x"17335574",
         13366 => x"822e0981",
         13367 => x"06fe8138",
         13368 => x"8154b417",
         13369 => x"08a01808",
         13370 => x"05537a52",
         13371 => x"81173351",
         13372 => x"ff92ef3f",
         13373 => x"7956fde8",
         13374 => x"3978902a",
         13375 => x"55749418",
         13376 => x"3474882a",
         13377 => x"56759518",
         13378 => x"348c1808",
         13379 => x"55747b34",
         13380 => x"74882a5b",
         13381 => x"7a9d1834",
         13382 => x"74902a56",
         13383 => x"759e1834",
         13384 => x"74982a59",
         13385 => x"789f1834",
         13386 => x"807a3480",
         13387 => x"0b971834",
         13388 => x"a10b9818",
         13389 => x"3480cc0b",
         13390 => x"99183480",
         13391 => x"0b921834",
         13392 => x"800b9318",
         13393 => x"347b5b81",
         13394 => x"0b831c34",
         13395 => x"7b51ff94",
         13396 => x"c43f84b9",
         13397 => x"c8089019",
         13398 => x"3381bf06",
         13399 => x"5b567990",
         13400 => x"1934feae",
         13401 => x"39811633",
         13402 => x"51ff90a5",
         13403 => x"3f84b9c8",
         13404 => x"08810655",
         13405 => x"74fcba38",
         13406 => x"74780856",
         13407 => x"5afcb439",
         13408 => x"f93d0d79",
         13409 => x"705255fb",
         13410 => x"fe3f84b9",
         13411 => x"c8085484",
         13412 => x"b9c808b1",
         13413 => x"38895674",
         13414 => x"802e9e38",
         13415 => x"74085372",
         13416 => x"802e9638",
         13417 => x"72335271",
         13418 => x"802e8e38",
         13419 => x"86132284",
         13420 => x"16225852",
         13421 => x"71772e96",
         13422 => x"38805271",
         13423 => x"58755475",
         13424 => x"84387575",
         13425 => x"0c7384b9",
         13426 => x"c80c893d",
         13427 => x"0d048113",
         13428 => x"3351ff8f",
         13429 => x"bc3f84b9",
         13430 => x"c8088106",
         13431 => x"5372da38",
         13432 => x"73750853",
         13433 => x"56d539f6",
         13434 => x"3d0dff7d",
         13435 => x"705b575b",
         13436 => x"75802eb2",
         13437 => x"38757081",
         13438 => x"05573370",
         13439 => x"9f265252",
         13440 => x"71ba2eac",
         13441 => x"3870ee38",
         13442 => x"71ba2ea4",
         13443 => x"3884d1a4",
         13444 => x"33518071",
         13445 => x"24903870",
         13446 => x"84d1a434",
         13447 => x"800b84b9",
         13448 => x"c80c8c3d",
         13449 => x"0d048b0b",
         13450 => x"84b9c80c",
         13451 => x"8c3d0d04",
         13452 => x"7833d011",
         13453 => x"7081ff06",
         13454 => x"53535370",
         13455 => x"89269138",
         13456 => x"82197381",
         13457 => x"ff06d005",
         13458 => x"59547376",
         13459 => x"2e80f538",
         13460 => x"800b83e5",
         13461 => x"b85b5879",
         13462 => x"08795657",
         13463 => x"76708105",
         13464 => x"58337570",
         13465 => x"81055733",
         13466 => x"ff9f1253",
         13467 => x"54527099",
         13468 => x"268938e0",
         13469 => x"127081ff",
         13470 => x"065354ff",
         13471 => x"9f135170",
         13472 => x"99268938",
         13473 => x"e0137081",
         13474 => x"ff065454",
         13475 => x"7130709f",
         13476 => x"2a555171",
         13477 => x"732e0981",
         13478 => x"06853873",
         13479 => x"ffbe3874",
         13480 => x"76327030",
         13481 => x"7072079f",
         13482 => x"2a760759",
         13483 => x"52527680",
         13484 => x"2e923881",
         13485 => x"18841b5b",
         13486 => x"58837825",
         13487 => x"ff99387a",
         13488 => x"51fecf39",
         13489 => x"778324f7",
         13490 => x"3877765e",
         13491 => x"51fec339",
         13492 => x"ea3d0d80",
         13493 => x"53983dcc",
         13494 => x"0552993d",
         13495 => x"51d1943f",
         13496 => x"84b9c808",
         13497 => x"5584b9c8",
         13498 => x"08802e8a",
         13499 => x"387484b9",
         13500 => x"c80c983d",
         13501 => x"0d047a5c",
         13502 => x"6852983d",
         13503 => x"d00551c5",
         13504 => x"943f84b9",
         13505 => x"c8085584",
         13506 => x"b9c80880",
         13507 => x"c6380280",
         13508 => x"d7053370",
         13509 => x"982b585a",
         13510 => x"80772480",
         13511 => x"e23802b2",
         13512 => x"05337084",
         13513 => x"2a810657",
         13514 => x"5975802e",
         13515 => x"b2387a63",
         13516 => x"9b11339a",
         13517 => x"12337188",
         13518 => x"2b077333",
         13519 => x"5e5a5b57",
         13520 => x"5879832e",
         13521 => x"a4387698",
         13522 => x"190c7484",
         13523 => x"b9c80c98",
         13524 => x"3d0d0484",
         13525 => x"b9c80884",
         13526 => x"2e098106",
         13527 => x"ff8f3885",
         13528 => x"0b84b9c8",
         13529 => x"0c983d0d",
         13530 => x"04951633",
         13531 => x"94173371",
         13532 => x"982b7190",
         13533 => x"2b077907",
         13534 => x"981b0c5b",
         13535 => x"54cc397a",
         13536 => x"7e98120c",
         13537 => x"587484b9",
         13538 => x"c80c983d",
         13539 => x"0d04ff9e",
         13540 => x"3d0d80e6",
         13541 => x"3d0880e6",
         13542 => x"3d085d40",
         13543 => x"807c3480",
         13544 => x"5380e43d",
         13545 => x"fdb40552",
         13546 => x"80e53d51",
         13547 => x"cfc53f84",
         13548 => x"b9c80859",
         13549 => x"84b9c808",
         13550 => x"83c83860",
         13551 => x"80d93d0c",
         13552 => x"7f619811",
         13553 => x"0880dd3d",
         13554 => x"0c5880db",
         13555 => x"3d085b58",
         13556 => x"79802e82",
         13557 => x"cc3880d8",
         13558 => x"3d983d40",
         13559 => x"5ba0527a",
         13560 => x"51ffa4aa",
         13561 => x"3f84b9c8",
         13562 => x"085984b9",
         13563 => x"c8088392",
         13564 => x"386080df",
         13565 => x"3d085856",
         13566 => x"b4160877",
         13567 => x"2eb13884",
         13568 => x"b9c80883",
         13569 => x"17335f5d",
         13570 => x"7d83c738",
         13571 => x"81547653",
         13572 => x"b8165281",
         13573 => x"163351ff",
         13574 => x"8bc93f84",
         13575 => x"b9c80880",
         13576 => x"2e8538ff",
         13577 => x"57815976",
         13578 => x"b4170c78",
         13579 => x"82d43880",
         13580 => x"df3d089b",
         13581 => x"11339a12",
         13582 => x"3371882b",
         13583 => x"07637033",
         13584 => x"5d405956",
         13585 => x"5678832e",
         13586 => x"82da3876",
         13587 => x"80db3d0c",
         13588 => x"80527a51",
         13589 => x"ffa3b73f",
         13590 => x"84b9c808",
         13591 => x"5984b9c8",
         13592 => x"08829f38",
         13593 => x"80527a51",
         13594 => x"ffa8f53f",
         13595 => x"84b9c808",
         13596 => x"5984b9c8",
         13597 => x"08bb3880",
         13598 => x"df3d089b",
         13599 => x"11339a12",
         13600 => x"3371882b",
         13601 => x"07637033",
         13602 => x"4258595e",
         13603 => x"567d832e",
         13604 => x"81fd3876",
         13605 => x"7a2ea438",
         13606 => x"84b9c808",
         13607 => x"527a51ff",
         13608 => x"a4e23f84",
         13609 => x"b9c80859",
         13610 => x"84b9c808",
         13611 => x"802effb4",
         13612 => x"3878842e",
         13613 => x"83d83878",
         13614 => x"81c83880",
         13615 => x"e43dfdb8",
         13616 => x"05527a51",
         13617 => x"ffbd893f",
         13618 => x"787f8205",
         13619 => x"335b5779",
         13620 => x"802e9038",
         13621 => x"821f5681",
         13622 => x"17811770",
         13623 => x"335f5757",
         13624 => x"7cf53881",
         13625 => x"17567578",
         13626 => x"26819538",
         13627 => x"76802e9c",
         13628 => x"387e1782",
         13629 => x"0556ff18",
         13630 => x"80e63d08",
         13631 => x"11ff19ff",
         13632 => x"19595956",
         13633 => x"58753375",
         13634 => x"3476eb38",
         13635 => x"ff1880e6",
         13636 => x"3d08115f",
         13637 => x"58af7e34",
         13638 => x"80da3d08",
         13639 => x"5a79fdbd",
         13640 => x"3877602e",
         13641 => x"828a3880",
         13642 => x"0b84d1a4",
         13643 => x"33701010",
         13644 => x"83e5b805",
         13645 => x"70087033",
         13646 => x"4359595e",
         13647 => x"5a7e7a2e",
         13648 => x"8d38811a",
         13649 => x"70177033",
         13650 => x"575f5a74",
         13651 => x"f538821a",
         13652 => x"5b7a7826",
         13653 => x"ab388057",
         13654 => x"767a2794",
         13655 => x"3876165f",
         13656 => x"7e337c70",
         13657 => x"81055e34",
         13658 => x"81175779",
         13659 => x"7726ee38",
         13660 => x"ba7c7081",
         13661 => x"055e3476",
         13662 => x"ff2e0981",
         13663 => x"0681df38",
         13664 => x"9159807c",
         13665 => x"347884b9",
         13666 => x"c80c80e4",
         13667 => x"3d0d0495",
         13668 => x"16339417",
         13669 => x"3371982b",
         13670 => x"71902b07",
         13671 => x"79075956",
         13672 => x"5efdf039",
         13673 => x"95163394",
         13674 => x"17337198",
         13675 => x"2b71902b",
         13676 => x"07790780",
         13677 => x"dd3d0c5a",
         13678 => x"5d80527a",
         13679 => x"51ffa0ce",
         13680 => x"3f84b9c8",
         13681 => x"085984b9",
         13682 => x"c808802e",
         13683 => x"fd9638ff",
         13684 => x"b1398154",
         13685 => x"b4160853",
         13686 => x"b8167053",
         13687 => x"81173352",
         13688 => x"5eff88fe",
         13689 => x"3f815984",
         13690 => x"b9c808fc",
         13691 => x"be3884b9",
         13692 => x"c8088317",
         13693 => x"34b41608",
         13694 => x"a8170831",
         13695 => x"84b9c808",
         13696 => x"5a5574a0",
         13697 => x"170827fc",
         13698 => x"83388216",
         13699 => x"33557482",
         13700 => x"2e098106",
         13701 => x"fbf63881",
         13702 => x"54b41608",
         13703 => x"a0170805",
         13704 => x"537d5281",
         13705 => x"163351ff",
         13706 => x"88b83f7c",
         13707 => x"59fbdd39",
         13708 => x"ff1880e6",
         13709 => x"3d08115c",
         13710 => x"58af7b34",
         13711 => x"800b84d1",
         13712 => x"a4337010",
         13713 => x"1083e5b8",
         13714 => x"05700870",
         13715 => x"33435959",
         13716 => x"5e5a7e7a",
         13717 => x"2e098106",
         13718 => x"fde838fd",
         13719 => x"f13980e5",
         13720 => x"3d081881",
         13721 => x"19595a79",
         13722 => x"337c7081",
         13723 => x"055e3477",
         13724 => x"6027fe8e",
         13725 => x"3880e53d",
         13726 => x"08188119",
         13727 => x"595a7933",
         13728 => x"7c708105",
         13729 => x"5e347f78",
         13730 => x"26d438fd",
         13731 => x"f5398259",
         13732 => x"807c3478",
         13733 => x"84b9c80c",
         13734 => x"80e43d0d",
         13735 => x"04f73d0d",
         13736 => x"7b7d5855",
         13737 => x"89567480",
         13738 => x"2e9f3874",
         13739 => x"08547380",
         13740 => x"2e973873",
         13741 => x"33537280",
         13742 => x"2e8f3886",
         13743 => x"14228416",
         13744 => x"22595978",
         13745 => x"782e83a0",
         13746 => x"38805372",
         13747 => x"5a755375",
         13748 => x"81c23891",
         13749 => x"15335372",
         13750 => x"81ba388c",
         13751 => x"15085676",
         13752 => x"762681b9",
         13753 => x"38941508",
         13754 => x"54805876",
         13755 => x"782e81cc",
         13756 => x"38798a11",
         13757 => x"2270892b",
         13758 => x"525a5673",
         13759 => x"782e81f7",
         13760 => x"387552ff",
         13761 => x"1751fdbb",
         13762 => x"9c3f84b9",
         13763 => x"c808ff15",
         13764 => x"77547053",
         13765 => x"5553fdbb",
         13766 => x"8c3f84b9",
         13767 => x"c8087326",
         13768 => x"81d53875",
         13769 => x"30740670",
         13770 => x"94170c77",
         13771 => x"71319817",
         13772 => x"08565859",
         13773 => x"73802e82",
         13774 => x"98387577",
         13775 => x"2781d938",
         13776 => x"76763194",
         13777 => x"16081794",
         13778 => x"170c9016",
         13779 => x"3370812a",
         13780 => x"8106515a",
         13781 => x"5778802e",
         13782 => x"81fe3873",
         13783 => x"527451ff",
         13784 => x"99f33f84",
         13785 => x"b9c80854",
         13786 => x"84b9c808",
         13787 => x"802e81a3",
         13788 => x"3873ff2e",
         13789 => x"98388174",
         13790 => x"2782b438",
         13791 => x"7953739c",
         13792 => x"14082782",
         13793 => x"aa387398",
         13794 => x"160cffae",
         13795 => x"39810b91",
         13796 => x"16348153",
         13797 => x"7284b9c8",
         13798 => x"0c8b3d0d",
         13799 => x"04901533",
         13800 => x"70812a81",
         13801 => x"06555873",
         13802 => x"febb3875",
         13803 => x"94160855",
         13804 => x"57805876",
         13805 => x"782e0981",
         13806 => x"06feb638",
         13807 => x"7794160c",
         13808 => x"94150854",
         13809 => x"75742790",
         13810 => x"38738c16",
         13811 => x"0c901533",
         13812 => x"80c00757",
         13813 => x"76901634",
         13814 => x"7383ff06",
         13815 => x"5978802e",
         13816 => x"8c389c15",
         13817 => x"08782e85",
         13818 => x"38779c16",
         13819 => x"0c800b84",
         13820 => x"b9c80c8b",
         13821 => x"3d0d0480",
         13822 => x"0b94160c",
         13823 => x"88150854",
         13824 => x"73802e80",
         13825 => x"fe387398",
         13826 => x"160c7380",
         13827 => x"2e80c238",
         13828 => x"fea83984",
         13829 => x"b9c80857",
         13830 => x"94150817",
         13831 => x"94160c76",
         13832 => x"83ff0656",
         13833 => x"75802ea9",
         13834 => x"3879fe15",
         13835 => x"9c1208fe",
         13836 => x"055a5556",
         13837 => x"73782780",
         13838 => x"f6388a16",
         13839 => x"22747129",
         13840 => x"b0180805",
         13841 => x"78892a11",
         13842 => x"5a5a5378",
         13843 => x"802e80df",
         13844 => x"388c1508",
         13845 => x"56fee939",
         13846 => x"73527451",
         13847 => x"ff89b73f",
         13848 => x"84b9c808",
         13849 => x"54fe8a39",
         13850 => x"81143351",
         13851 => x"ff82a23f",
         13852 => x"84b9c808",
         13853 => x"81065372",
         13854 => x"fccf3872",
         13855 => x"75085456",
         13856 => x"fcc93973",
         13857 => x"527451ff",
         13858 => x"97cb3f84",
         13859 => x"b9c80854",
         13860 => x"84b9c808",
         13861 => x"812e9838",
         13862 => x"84b9c808",
         13863 => x"ff2efded",
         13864 => x"3884b9c8",
         13865 => x"0888160c",
         13866 => x"7398160c",
         13867 => x"fedc3982",
         13868 => x"0b911634",
         13869 => x"820b84b9",
         13870 => x"c80c8b3d",
         13871 => x"0d04f63d",
         13872 => x"0d7c5689",
         13873 => x"5475802e",
         13874 => x"a2388053",
         13875 => x"8c3dfc05",
         13876 => x"528d3d84",
         13877 => x"0551c59b",
         13878 => x"3f84b9c8",
         13879 => x"085584b9",
         13880 => x"c808802e",
         13881 => x"8f388076",
         13882 => x"0c745473",
         13883 => x"84b9c80c",
         13884 => x"8c3d0d04",
         13885 => x"7a760c7d",
         13886 => x"527551ff",
         13887 => x"b9973f84",
         13888 => x"b9c80855",
         13889 => x"84b9c808",
         13890 => x"80d138ab",
         13891 => x"16337098",
         13892 => x"2b595980",
         13893 => x"7824af38",
         13894 => x"86163370",
         13895 => x"842a8106",
         13896 => x"5b547980",
         13897 => x"2e80c538",
         13898 => x"9c16089b",
         13899 => x"11339a12",
         13900 => x"3371882b",
         13901 => x"077d7033",
         13902 => x"5d5d5a55",
         13903 => x"5778832e",
         13904 => x"b3387788",
         13905 => x"170c7a58",
         13906 => x"86182284",
         13907 => x"17237452",
         13908 => x"7551ff99",
         13909 => x"b93f84b9",
         13910 => x"c8085574",
         13911 => x"842e8d38",
         13912 => x"74802eff",
         13913 => x"84388076",
         13914 => x"0cfefe39",
         13915 => x"85558076",
         13916 => x"0cfef639",
         13917 => x"95173394",
         13918 => x"18337198",
         13919 => x"2b71902b",
         13920 => x"077a0788",
         13921 => x"190c5a5a",
         13922 => x"ffbc39fa",
         13923 => x"3d0d7855",
         13924 => x"89547480",
         13925 => x"2e9e3874",
         13926 => x"08537280",
         13927 => x"2e963872",
         13928 => x"33527180",
         13929 => x"2e8e3886",
         13930 => x"13228416",
         13931 => x"22575271",
         13932 => x"762e9438",
         13933 => x"80527157",
         13934 => x"73843873",
         13935 => x"750c7384",
         13936 => x"b9c80c88",
         13937 => x"3d0d0481",
         13938 => x"133351fe",
         13939 => x"ffc33f84",
         13940 => x"b9c80881",
         13941 => x"065271dc",
         13942 => x"38717508",
         13943 => x"5354d739",
         13944 => x"f83d0d7a",
         13945 => x"7c585589",
         13946 => x"5674802e",
         13947 => x"9f387408",
         13948 => x"5473802e",
         13949 => x"97387333",
         13950 => x"5372802e",
         13951 => x"8f388614",
         13952 => x"22841622",
         13953 => x"59537278",
         13954 => x"2e819738",
         13955 => x"80537259",
         13956 => x"75537580",
         13957 => x"c7387680",
         13958 => x"2e80f338",
         13959 => x"75527451",
         13960 => x"ff9dbd3f",
         13961 => x"84b9c808",
         13962 => x"5384b9c8",
         13963 => x"08842eb5",
         13964 => x"3884b9c8",
         13965 => x"08a63876",
         13966 => x"527451ff",
         13967 => x"b2923f72",
         13968 => x"527451ff",
         13969 => x"99be3f84",
         13970 => x"b9c80884",
         13971 => x"32703070",
         13972 => x"72079f2c",
         13973 => x"84b9c808",
         13974 => x"06555754",
         13975 => x"7284b9c8",
         13976 => x"0c8a3d0d",
         13977 => x"04757753",
         13978 => x"755253ff",
         13979 => x"b1e23f72",
         13980 => x"527451ff",
         13981 => x"998e3f84",
         13982 => x"b9c80884",
         13983 => x"32703070",
         13984 => x"72079f2c",
         13985 => x"84b9c808",
         13986 => x"06555754",
         13987 => x"cf397552",
         13988 => x"7451ff96",
         13989 => x"f93f84b9",
         13990 => x"c80884b9",
         13991 => x"c80c8a3d",
         13992 => x"0d048114",
         13993 => x"3351fefd",
         13994 => x"e83f84b9",
         13995 => x"c8088106",
         13996 => x"5372fed8",
         13997 => x"38727508",
         13998 => x"5456fed2",
         13999 => x"39ed3d0d",
         14000 => x"66578053",
         14001 => x"893d7053",
         14002 => x"973d5256",
         14003 => x"c1a53f84",
         14004 => x"b9c80855",
         14005 => x"84b9c808",
         14006 => x"802e8a38",
         14007 => x"7484b9c8",
         14008 => x"0c953d0d",
         14009 => x"04655275",
         14010 => x"51ffb5a9",
         14011 => x"3f84b9c8",
         14012 => x"085584b9",
         14013 => x"c808e538",
         14014 => x"0280cb05",
         14015 => x"3370982b",
         14016 => x"55588074",
         14017 => x"24973876",
         14018 => x"802ed138",
         14019 => x"76527551",
         14020 => x"ffb0bd3f",
         14021 => x"7484b9c8",
         14022 => x"0c953d0d",
         14023 => x"04860b84",
         14024 => x"b9c80c95",
         14025 => x"3d0d04ed",
         14026 => x"3d0d6668",
         14027 => x"565f8053",
         14028 => x"953dec05",
         14029 => x"52963d51",
         14030 => x"c0b93f84",
         14031 => x"b9c8085a",
         14032 => x"84b9c808",
         14033 => x"9a387f75",
         14034 => x"0c74089c",
         14035 => x"1108fe11",
         14036 => x"94130859",
         14037 => x"57595775",
         14038 => x"75268d38",
         14039 => x"757f0c79",
         14040 => x"84b9c80c",
         14041 => x"953d0d04",
         14042 => x"84b9c808",
         14043 => x"77335a5b",
         14044 => x"78812e82",
         14045 => x"933877a8",
         14046 => x"180884b9",
         14047 => x"c8085a5d",
         14048 => x"597780c1",
         14049 => x"387b811d",
         14050 => x"715c5d56",
         14051 => x"b4170876",
         14052 => x"2e82ef38",
         14053 => x"83173378",
         14054 => x"5f5d7c81",
         14055 => x"8d388154",
         14056 => x"7553b817",
         14057 => x"52811733",
         14058 => x"51fefcb7",
         14059 => x"3f84b9c8",
         14060 => x"08802e85",
         14061 => x"38ff5a81",
         14062 => x"5e79b418",
         14063 => x"0c7f7e5b",
         14064 => x"577d80cc",
         14065 => x"3876335e",
         14066 => x"7d822e82",
         14067 => x"8d387717",
         14068 => x"b8058311",
         14069 => x"33821233",
         14070 => x"71902b71",
         14071 => x"882b0781",
         14072 => x"14337072",
         14073 => x"07882b75",
         14074 => x"337180ff",
         14075 => x"fffe8006",
         14076 => x"07703070",
         14077 => x"80256305",
         14078 => x"60840583",
         14079 => x"ff0662ff",
         14080 => x"05434143",
         14081 => x"53545253",
         14082 => x"58405e56",
         14083 => x"78fef238",
         14084 => x"7a7f0c7a",
         14085 => x"94180c84",
         14086 => x"17338107",
         14087 => x"58778418",
         14088 => x"347984b9",
         14089 => x"c80c953d",
         14090 => x"0d048154",
         14091 => x"b4170853",
         14092 => x"b8177053",
         14093 => x"81183352",
         14094 => x"5dfefca6",
         14095 => x"3f815e84",
         14096 => x"b9c808fe",
         14097 => x"f83884b9",
         14098 => x"c8088318",
         14099 => x"34b41708",
         14100 => x"a8180831",
         14101 => x"84b9c808",
         14102 => x"5f5574a0",
         14103 => x"180827fe",
         14104 => x"bd388217",
         14105 => x"33557482",
         14106 => x"2e098106",
         14107 => x"feb03881",
         14108 => x"54b41708",
         14109 => x"a0180805",
         14110 => x"537c5281",
         14111 => x"173351fe",
         14112 => x"fbe03f77",
         14113 => x"5efe9739",
         14114 => x"82774292",
         14115 => x"3d595675",
         14116 => x"527751ff",
         14117 => x"81803f84",
         14118 => x"b9c808ff",
         14119 => x"2e80e838",
         14120 => x"84b9c808",
         14121 => x"812e80f7",
         14122 => x"3884b9c8",
         14123 => x"08307084",
         14124 => x"b9c80807",
         14125 => x"80257c05",
         14126 => x"8118625a",
         14127 => x"585c5c9c",
         14128 => x"17087626",
         14129 => x"ca387a7f",
         14130 => x"0c7a9418",
         14131 => x"0c841733",
         14132 => x"81075877",
         14133 => x"841834fe",
         14134 => x"c8397717",
         14135 => x"b8058111",
         14136 => x"33713371",
         14137 => x"882b0770",
         14138 => x"30708025",
         14139 => x"1f821d83",
         14140 => x"ff06ff1f",
         14141 => x"5f5d5f59",
         14142 => x"5f5f5578",
         14143 => x"fd8338fe",
         14144 => x"8f39775a",
         14145 => x"fdbf3981",
         14146 => x"60585a7a",
         14147 => x"7f0c7a94",
         14148 => x"180c8417",
         14149 => x"33810758",
         14150 => x"77841834",
         14151 => x"fe833982",
         14152 => x"60585ae7",
         14153 => x"39f73d0d",
         14154 => x"7b578956",
         14155 => x"76802e9f",
         14156 => x"38760855",
         14157 => x"74802e97",
         14158 => x"38743354",
         14159 => x"73802e8f",
         14160 => x"38861522",
         14161 => x"84182259",
         14162 => x"5978782e",
         14163 => x"81da3880",
         14164 => x"54735a75",
         14165 => x"80dc3891",
         14166 => x"17335675",
         14167 => x"80d43890",
         14168 => x"17337081",
         14169 => x"2a810655",
         14170 => x"58875573",
         14171 => x"802e80c4",
         14172 => x"38941708",
         14173 => x"54738c18",
         14174 => x"0827b738",
         14175 => x"7381d538",
         14176 => x"88170877",
         14177 => x"08575481",
         14178 => x"74278838",
         14179 => x"9c160874",
         14180 => x"26b33882",
         14181 => x"56800b88",
         14182 => x"180c9417",
         14183 => x"088c180c",
         14184 => x"7780c007",
         14185 => x"59789018",
         14186 => x"3475802e",
         14187 => x"85387591",
         14188 => x"18347555",
         14189 => x"7484b9c8",
         14190 => x"0c8b3d0d",
         14191 => x"04785478",
         14192 => x"782780ff",
         14193 => x"38735276",
         14194 => x"51fefeca",
         14195 => x"3f84b9c8",
         14196 => x"085984b9",
         14197 => x"c808802e",
         14198 => x"80e93884",
         14199 => x"b9c80881",
         14200 => x"2e82d838",
         14201 => x"84b9c808",
         14202 => x"ff2e82e5",
         14203 => x"38805373",
         14204 => x"527551ff",
         14205 => x"85813f84",
         14206 => x"b9c80882",
         14207 => x"c8389c16",
         14208 => x"08fe1194",
         14209 => x"18085755",
         14210 => x"58747427",
         14211 => x"ffaf3881",
         14212 => x"1594170c",
         14213 => x"84163381",
         14214 => x"07547384",
         14215 => x"17347854",
         14216 => x"777926ff",
         14217 => x"a0389c39",
         14218 => x"81153351",
         14219 => x"fef6e23f",
         14220 => x"84b9c808",
         14221 => x"81065473",
         14222 => x"fe953873",
         14223 => x"77085556",
         14224 => x"fe8f3980",
         14225 => x"0b901833",
         14226 => x"59547356",
         14227 => x"800b8818",
         14228 => x"0cfec739",
         14229 => x"98170852",
         14230 => x"7651fefd",
         14231 => x"b93f84b9",
         14232 => x"c808ff2e",
         14233 => x"81c23884",
         14234 => x"b9c80881",
         14235 => x"2e81be38",
         14236 => x"7581ae38",
         14237 => x"795884b9",
         14238 => x"c8089c19",
         14239 => x"082781a1",
         14240 => x"3884b9c8",
         14241 => x"08981808",
         14242 => x"78085856",
         14243 => x"54810b84",
         14244 => x"b9c80827",
         14245 => x"81a13884",
         14246 => x"b9c8089c",
         14247 => x"17082781",
         14248 => x"96387480",
         14249 => x"2e9738ff",
         14250 => x"53745275",
         14251 => x"51ff83c7",
         14252 => x"3f84b9c8",
         14253 => x"085584b9",
         14254 => x"c80880e3",
         14255 => x"38735276",
         14256 => x"51fefcd2",
         14257 => x"3f84b9c8",
         14258 => x"085984b9",
         14259 => x"c808802e",
         14260 => x"80cb3884",
         14261 => x"b9c80881",
         14262 => x"2e80dc38",
         14263 => x"84b9c808",
         14264 => x"ff2e80fe",
         14265 => x"38805373",
         14266 => x"527551ff",
         14267 => x"83893f84",
         14268 => x"b9c80880",
         14269 => x"e6389c16",
         14270 => x"08fe1194",
         14271 => x"18085755",
         14272 => x"58747427",
         14273 => x"90388115",
         14274 => x"94170c84",
         14275 => x"16338107",
         14276 => x"54738417",
         14277 => x"34785477",
         14278 => x"7926ffa1",
         14279 => x"38805574",
         14280 => x"56901733",
         14281 => x"58fcf339",
         14282 => x"8156febb",
         14283 => x"39820b90",
         14284 => x"18335956",
         14285 => x"fce43982",
         14286 => x"56e73982",
         14287 => x"0b901833",
         14288 => x"5954fe86",
         14289 => x"3984b9c8",
         14290 => x"08901833",
         14291 => x"5954fdfa",
         14292 => x"39810b90",
         14293 => x"18335954",
         14294 => x"fdf03984",
         14295 => x"b9c80856",
         14296 => x"c0398156",
         14297 => x"ffbb39db",
         14298 => x"3d0d8253",
         14299 => x"a73dff9c",
         14300 => x"0552a83d",
         14301 => x"51ffb7fb",
         14302 => x"3f84b9c8",
         14303 => x"085684b9",
         14304 => x"c808802e",
         14305 => x"8a387584",
         14306 => x"b9c80ca7",
         14307 => x"3d0d047d",
         14308 => x"4ba83d08",
         14309 => x"529b3d70",
         14310 => x"5259ffab",
         14311 => x"f83f84b9",
         14312 => x"c8085684",
         14313 => x"b9c808de",
         14314 => x"38028193",
         14315 => x"05337085",
         14316 => x"2a810659",
         14317 => x"57865677",
         14318 => x"cd387698",
         14319 => x"2b5b807b",
         14320 => x"24c43802",
         14321 => x"80ee0533",
         14322 => x"7081065d",
         14323 => x"5787567b",
         14324 => x"ffb4387d",
         14325 => x"a33d089b",
         14326 => x"11339a12",
         14327 => x"3371882b",
         14328 => x"07733341",
         14329 => x"5e5c5758",
         14330 => x"7c832e80",
         14331 => x"d5387684",
         14332 => x"2a810657",
         14333 => x"76802e80",
         14334 => x"ed388756",
         14335 => x"9818087b",
         14336 => x"2eff8338",
         14337 => x"775f7a41",
         14338 => x"84b9c808",
         14339 => x"528f3d70",
         14340 => x"5255ff8b",
         14341 => x"f93f84b9",
         14342 => x"c8085684",
         14343 => x"b9c808fe",
         14344 => x"e53884b9",
         14345 => x"c8085274",
         14346 => x"51ff91b4",
         14347 => x"3f84b9c8",
         14348 => x"085684b9",
         14349 => x"c808a038",
         14350 => x"870b84b9",
         14351 => x"c80ca73d",
         14352 => x"0d049516",
         14353 => x"33941733",
         14354 => x"71982b71",
         14355 => x"902b077d",
         14356 => x"075d5d5d",
         14357 => x"ff983984",
         14358 => x"b9c80884",
         14359 => x"2e883884",
         14360 => x"b9c808fe",
         14361 => x"a1387808",
         14362 => x"6fa83d08",
         14363 => x"575d5774",
         14364 => x"ff2e80d3",
         14365 => x"38745278",
         14366 => x"51ff8b92",
         14367 => x"3f84b9c8",
         14368 => x"085684b9",
         14369 => x"c808802e",
         14370 => x"be387530",
         14371 => x"70770780",
         14372 => x"25565a7a",
         14373 => x"802e9a38",
         14374 => x"74802e95",
         14375 => x"387a7908",
         14376 => x"5855817b",
         14377 => x"2789389c",
         14378 => x"17087b26",
         14379 => x"81fd3882",
         14380 => x"5675fdd2",
         14381 => x"387d51fe",
         14382 => x"f5db3f84",
         14383 => x"b9c80884",
         14384 => x"b9c80ca7",
         14385 => x"3d0d04b8",
         14386 => x"175d9819",
         14387 => x"0856805a",
         14388 => x"b4170876",
         14389 => x"2e82b938",
         14390 => x"8317337a",
         14391 => x"5955747a",
         14392 => x"2e098106",
         14393 => x"80dd3881",
         14394 => x"547553b8",
         14395 => x"17528117",
         14396 => x"3351fef1",
         14397 => x"ee3f84b9",
         14398 => x"c808802e",
         14399 => x"8538ff56",
         14400 => x"815875b4",
         14401 => x"180c7756",
         14402 => x"77ab389c",
         14403 => x"190858e5",
         14404 => x"7834810b",
         14405 => x"83183490",
         14406 => x"19087c27",
         14407 => x"feec3880",
         14408 => x"527851ff",
         14409 => x"8bde3f84",
         14410 => x"b9c80856",
         14411 => x"84b9c808",
         14412 => x"802eff96",
         14413 => x"3875842e",
         14414 => x"098106fe",
         14415 => x"cd388256",
         14416 => x"fec83981",
         14417 => x"54b41708",
         14418 => x"537c5281",
         14419 => x"173351fe",
         14420 => x"f2903f81",
         14421 => x"5884b9c8",
         14422 => x"087a2e09",
         14423 => x"8106ffa6",
         14424 => x"3884b9c8",
         14425 => x"08831834",
         14426 => x"b41708a8",
         14427 => x"18083184",
         14428 => x"b9c80859",
         14429 => x"5574a018",
         14430 => x"0827feeb",
         14431 => x"38821733",
         14432 => x"5574822e",
         14433 => x"098106fe",
         14434 => x"de388154",
         14435 => x"b41708a0",
         14436 => x"18080553",
         14437 => x"7c528117",
         14438 => x"3351fef1",
         14439 => x"c53f7958",
         14440 => x"fec53979",
         14441 => x"55797827",
         14442 => x"80e13874",
         14443 => x"527851fe",
         14444 => x"f6e43f84",
         14445 => x"b9c8085a",
         14446 => x"84b9c808",
         14447 => x"802e80cb",
         14448 => x"3884b9c8",
         14449 => x"08812efd",
         14450 => x"e63884b9",
         14451 => x"c808ff2e",
         14452 => x"80cb3880",
         14453 => x"53745276",
         14454 => x"51fefd9b",
         14455 => x"3f84b9c8",
         14456 => x"08b3389c",
         14457 => x"1708fe11",
         14458 => x"94190858",
         14459 => x"5c58757b",
         14460 => x"27ffb038",
         14461 => x"81169418",
         14462 => x"0c841733",
         14463 => x"81075c7b",
         14464 => x"84183479",
         14465 => x"55777a26",
         14466 => x"ffa13880",
         14467 => x"56fda239",
         14468 => x"7956fdf7",
         14469 => x"3984b9c8",
         14470 => x"0856fd95",
         14471 => x"398156fd",
         14472 => x"9039e33d",
         14473 => x"0d82539f",
         14474 => x"3dffbc05",
         14475 => x"52a03d51",
         14476 => x"ffb2c03f",
         14477 => x"84b9c808",
         14478 => x"5684b9c8",
         14479 => x"08802e8a",
         14480 => x"387584b9",
         14481 => x"c80c9f3d",
         14482 => x"0d047d43",
         14483 => x"6f52933d",
         14484 => x"70525aff",
         14485 => x"a6bf3f84",
         14486 => x"b9c80856",
         14487 => x"84b9c808",
         14488 => x"8b38880b",
         14489 => x"84b9c80c",
         14490 => x"9f3d0d04",
         14491 => x"84b9c808",
         14492 => x"842e0981",
         14493 => x"06cb3802",
         14494 => x"80f30533",
         14495 => x"70852a81",
         14496 => x"06565886",
         14497 => x"5674ffb9",
         14498 => x"387d5f74",
         14499 => x"528f3d70",
         14500 => x"525dff83",
         14501 => x"c03f84b9",
         14502 => x"c8087557",
         14503 => x"5c84b9c8",
         14504 => x"08833887",
         14505 => x"5684b9c8",
         14506 => x"08812e80",
         14507 => x"f93884b9",
         14508 => x"c808ff2e",
         14509 => x"81cb3875",
         14510 => x"81c9387d",
         14511 => x"84b9c808",
         14512 => x"8312335d",
         14513 => x"5a577a80",
         14514 => x"e238fe19",
         14515 => x"9c1808fe",
         14516 => x"055a5680",
         14517 => x"5b757927",
         14518 => x"8d388a17",
         14519 => x"22767129",
         14520 => x"b0190805",
         14521 => x"5c587ab4",
         14522 => x"180cb817",
         14523 => x"59848079",
         14524 => x"57558076",
         14525 => x"70810558",
         14526 => x"34ff1555",
         14527 => x"74f43874",
         14528 => x"588a1722",
         14529 => x"55777527",
         14530 => x"81f93881",
         14531 => x"54771b53",
         14532 => x"78528117",
         14533 => x"3351feee",
         14534 => x"c93f84b9",
         14535 => x"c80881df",
         14536 => x"38811858",
         14537 => x"dc398256",
         14538 => x"ff843981",
         14539 => x"54b41708",
         14540 => x"53b81770",
         14541 => x"53811833",
         14542 => x"5258feee",
         14543 => x"a53f8156",
         14544 => x"84b9c808",
         14545 => x"be3884b9",
         14546 => x"c8088318",
         14547 => x"34b41708",
         14548 => x"a8180831",
         14549 => x"5574a018",
         14550 => x"0827feee",
         14551 => x"38821733",
         14552 => x"5b7a822e",
         14553 => x"098106fe",
         14554 => x"e1387554",
         14555 => x"b41708a0",
         14556 => x"18080553",
         14557 => x"77528117",
         14558 => x"3351feed",
         14559 => x"e53ffeca",
         14560 => x"3981567b",
         14561 => x"7d085855",
         14562 => x"817c27fd",
         14563 => x"b4387b9c",
         14564 => x"180827fd",
         14565 => x"ac387452",
         14566 => x"7c51fef2",
         14567 => x"f93f84b9",
         14568 => x"c8085a84",
         14569 => x"b9c80880",
         14570 => x"2efd9638",
         14571 => x"84b9c808",
         14572 => x"812efd8d",
         14573 => x"3884b9c8",
         14574 => x"08ff2efd",
         14575 => x"84388053",
         14576 => x"74527651",
         14577 => x"fef9b03f",
         14578 => x"84b9c808",
         14579 => x"fcf3389c",
         14580 => x"1708fe11",
         14581 => x"9419085a",
         14582 => x"5c59777b",
         14583 => x"27903881",
         14584 => x"1894180c",
         14585 => x"84173381",
         14586 => x"075c7b84",
         14587 => x"18347955",
         14588 => x"787a26ff",
         14589 => x"a1387584",
         14590 => x"b9c80c9f",
         14591 => x"3d0d048a",
         14592 => x"17225574",
         14593 => x"83ffff06",
         14594 => x"57815676",
         14595 => x"782e0981",
         14596 => x"06fef038",
         14597 => x"8b0bb81f",
         14598 => x"5656a075",
         14599 => x"70810557",
         14600 => x"34ff1656",
         14601 => x"75f4387d",
         14602 => x"57ae0bb8",
         14603 => x"18347d58",
         14604 => x"900b80c3",
         14605 => x"19347d59",
         14606 => x"7580ce1a",
         14607 => x"347580cf",
         14608 => x"1a34a10b",
         14609 => x"80d01a34",
         14610 => x"80cc0b80",
         14611 => x"d11a347d",
         14612 => x"7c83ffff",
         14613 => x"06595677",
         14614 => x"80d21734",
         14615 => x"77882a5b",
         14616 => x"7a80d317",
         14617 => x"34753355",
         14618 => x"74832e81",
         14619 => x"cc387d59",
         14620 => x"a00b80d8",
         14621 => x"1ab81b57",
         14622 => x"58567470",
         14623 => x"81055633",
         14624 => x"77708105",
         14625 => x"5934ff16",
         14626 => x"5675ef38",
         14627 => x"7d56ae0b",
         14628 => x"80d91734",
         14629 => x"647e7183",
         14630 => x"ffff065b",
         14631 => x"57577880",
         14632 => x"f2173478",
         14633 => x"882a5b7a",
         14634 => x"80f31734",
         14635 => x"75335574",
         14636 => x"832e80f0",
         14637 => x"387d5b81",
         14638 => x"0b831c34",
         14639 => x"7951ff92",
         14640 => x"963f84b9",
         14641 => x"c8085684",
         14642 => x"b9c808fd",
         14643 => x"b6386956",
         14644 => x"84b9c808",
         14645 => x"96173484",
         14646 => x"b9c80897",
         14647 => x"1734a10b",
         14648 => x"98173480",
         14649 => x"cc0b9917",
         14650 => x"347d6a58",
         14651 => x"5d779a18",
         14652 => x"3477882a",
         14653 => x"59789b18",
         14654 => x"347c335a",
         14655 => x"79832e80",
         14656 => x"d9386955",
         14657 => x"900b8b16",
         14658 => x"347d5781",
         14659 => x"0b831834",
         14660 => x"7d51feed",
         14661 => x"803f84b9",
         14662 => x"c8085675",
         14663 => x"84b9c80c",
         14664 => x"9f3d0d04",
         14665 => x"76902a55",
         14666 => x"7480ec17",
         14667 => x"3474882a",
         14668 => x"577680ed",
         14669 => x"1734fefd",
         14670 => x"397b902a",
         14671 => x"5b7a80cc",
         14672 => x"17347a88",
         14673 => x"2a557480",
         14674 => x"cd17347d",
         14675 => x"59a00b80",
         14676 => x"d81ab81b",
         14677 => x"575856fe",
         14678 => x"a1397b90",
         14679 => x"2a587794",
         14680 => x"18347788",
         14681 => x"2a5c7b95",
         14682 => x"18346955",
         14683 => x"900b8b16",
         14684 => x"347d5781",
         14685 => x"0b831834",
         14686 => x"7d51feec",
         14687 => x"983f84b9",
         14688 => x"c80856ff",
         14689 => x"9639d13d",
         14690 => x"0db33db4",
         14691 => x"3d087059",
         14692 => x"5b5f7980",
         14693 => x"2e9b3879",
         14694 => x"7081055b",
         14695 => x"33709f26",
         14696 => x"565675ba",
         14697 => x"2e81b838",
         14698 => x"74ed3875",
         14699 => x"ba2e81af",
         14700 => x"388253b1",
         14701 => x"3dfefc05",
         14702 => x"52b23d51",
         14703 => x"ffabb43f",
         14704 => x"84b9c808",
         14705 => x"5684b9c8",
         14706 => x"08802e8a",
         14707 => x"387584b9",
         14708 => x"c80cb13d",
         14709 => x"0d047fa6",
         14710 => x"3d0cb23d",
         14711 => x"0852a53d",
         14712 => x"705259ff",
         14713 => x"9faf3f84",
         14714 => x"b9c80856",
         14715 => x"84b9c808",
         14716 => x"dc380281",
         14717 => x"bb053381",
         14718 => x"a0065d86",
         14719 => x"567cce38",
         14720 => x"a00b923d",
         14721 => x"ae3d0858",
         14722 => x"58557570",
         14723 => x"81055733",
         14724 => x"77708105",
         14725 => x"5934ff15",
         14726 => x"5574ef38",
         14727 => x"993d58b0",
         14728 => x"787a5858",
         14729 => x"55757081",
         14730 => x"05573377",
         14731 => x"70810559",
         14732 => x"34ff1555",
         14733 => x"74ef38b3",
         14734 => x"3d085277",
         14735 => x"51ff9ed5",
         14736 => x"3f84b9c8",
         14737 => x"085684b9",
         14738 => x"c80885d8",
         14739 => x"386aa83d",
         14740 => x"082e81cb",
         14741 => x"38880b84",
         14742 => x"b9c80cb1",
         14743 => x"3d0d0476",
         14744 => x"33d01170",
         14745 => x"81ff0657",
         14746 => x"57587489",
         14747 => x"26913882",
         14748 => x"177881ff",
         14749 => x"06d0055d",
         14750 => x"59787a2e",
         14751 => x"80fa3880",
         14752 => x"7f0883e5",
         14753 => x"b8700872",
         14754 => x"5d5e5f5f",
         14755 => x"5c7a7081",
         14756 => x"055c3379",
         14757 => x"7081055b",
         14758 => x"33ff9f12",
         14759 => x"5a585677",
         14760 => x"99268938",
         14761 => x"e0167081",
         14762 => x"ff065755",
         14763 => x"ff9f1758",
         14764 => x"77992689",
         14765 => x"38e01770",
         14766 => x"81ff0658",
         14767 => x"55753070",
         14768 => x"9f2a5955",
         14769 => x"75772e09",
         14770 => x"81068538",
         14771 => x"77ffbe38",
         14772 => x"787a3270",
         14773 => x"30707207",
         14774 => x"9f2a7a07",
         14775 => x"5d58557a",
         14776 => x"802e9538",
         14777 => x"811c841e",
         14778 => x"5e5c7b83",
         14779 => x"24fdc238",
         14780 => x"7c087e5a",
         14781 => x"5bff9639",
         14782 => x"7b8324fd",
         14783 => x"b438797f",
         14784 => x"0c8253b1",
         14785 => x"3dfefc05",
         14786 => x"52b23d51",
         14787 => x"ffa8e43f",
         14788 => x"84b9c808",
         14789 => x"5684b9c8",
         14790 => x"08fdb238",
         14791 => x"fdb8396c",
         14792 => x"aa3d082e",
         14793 => x"098106fe",
         14794 => x"ac387751",
         14795 => x"ff8da83f",
         14796 => x"84b9c808",
         14797 => x"5684b9c8",
         14798 => x"08fd9238",
         14799 => x"6f58930b",
         14800 => x"8d190288",
         14801 => x"0580cd05",
         14802 => x"58565a75",
         14803 => x"70810557",
         14804 => x"33757081",
         14805 => x"055734ff",
         14806 => x"1a5a79ef",
         14807 => x"380280cb",
         14808 => x"05338b19",
         14809 => x"348b1833",
         14810 => x"70842a81",
         14811 => x"0640567e",
         14812 => x"893875a0",
         14813 => x"0757768b",
         14814 => x"19347f5d",
         14815 => x"810b831e",
         14816 => x"348b1833",
         14817 => x"70842a81",
         14818 => x"06575c75",
         14819 => x"802e81c5",
         14820 => x"38a73d08",
         14821 => x"6b2e81bd",
         14822 => x"387f9b19",
         14823 => x"339a1a33",
         14824 => x"71882b07",
         14825 => x"72334158",
         14826 => x"5c577d83",
         14827 => x"2e82e038",
         14828 => x"fe169c18",
         14829 => x"08fe055e",
         14830 => x"56757d27",
         14831 => x"82c7388a",
         14832 => x"17227671",
         14833 => x"29b01908",
         14834 => x"05575e75",
         14835 => x"802e82b5",
         14836 => x"38757a5d",
         14837 => x"58b41708",
         14838 => x"762eaa38",
         14839 => x"8317335f",
         14840 => x"7e83bc38",
         14841 => x"81547553",
         14842 => x"b8175281",
         14843 => x"173351fe",
         14844 => x"e3f13f84",
         14845 => x"b9c80880",
         14846 => x"2e8538ff",
         14847 => x"58815c77",
         14848 => x"b4180c7f",
         14849 => x"577b80d8",
         14850 => x"1856567b",
         14851 => x"fbbf3881",
         14852 => x"15335a79",
         14853 => x"ae2e0981",
         14854 => x"06bb386a",
         14855 => x"7083ffff",
         14856 => x"065d567b",
         14857 => x"80f21834",
         14858 => x"7b882a58",
         14859 => x"7780f318",
         14860 => x"3476335b",
         14861 => x"7a832e09",
         14862 => x"81069338",
         14863 => x"75902a5e",
         14864 => x"7d80ec18",
         14865 => x"347d882a",
         14866 => x"567580ed",
         14867 => x"18347f57",
         14868 => x"810b8318",
         14869 => x"347808aa",
         14870 => x"3d08b23d",
         14871 => x"08575c56",
         14872 => x"74ff2e95",
         14873 => x"38745278",
         14874 => x"51fefba2",
         14875 => x"3f84b9c8",
         14876 => x"085584b9",
         14877 => x"c80880f5",
         14878 => x"38b8165c",
         14879 => x"98190857",
         14880 => x"805ab416",
         14881 => x"08772eb4",
         14882 => x"38831633",
         14883 => x"7a595f7e",
         14884 => x"7a2e0981",
         14885 => x"0681a838",
         14886 => x"81547653",
         14887 => x"b8165281",
         14888 => x"163351fe",
         14889 => x"e2bd3f84",
         14890 => x"b9c80880",
         14891 => x"2e8538ff",
         14892 => x"57815876",
         14893 => x"b4170c77",
         14894 => x"5577aa38",
         14895 => x"9c19085a",
         14896 => x"e57a3481",
         14897 => x"0b831734",
         14898 => x"9019087b",
         14899 => x"27a53880",
         14900 => x"527851fe",
         14901 => x"fcae3f84",
         14902 => x"b9c80855",
         14903 => x"84b9c808",
         14904 => x"802eff98",
         14905 => x"38825674",
         14906 => x"842ef9e1",
         14907 => x"38745674",
         14908 => x"f9db387f",
         14909 => x"51fee59d",
         14910 => x"3f84b9c8",
         14911 => x"0884b9c8",
         14912 => x"0cb13d0d",
         14913 => x"04820b84",
         14914 => x"b9c80cb1",
         14915 => x"3d0d0495",
         14916 => x"18339419",
         14917 => x"3371982b",
         14918 => x"71902b07",
         14919 => x"78075856",
         14920 => x"5cfd8d39",
         14921 => x"84b9c808",
         14922 => x"842efbfe",
         14923 => x"3884b9c8",
         14924 => x"08802efe",
         14925 => x"a0387584",
         14926 => x"b9c80cb1",
         14927 => x"3d0d0481",
         14928 => x"54b41608",
         14929 => x"537b5281",
         14930 => x"163351fe",
         14931 => x"e2943f81",
         14932 => x"5884b9c8",
         14933 => x"087a2e09",
         14934 => x"8106fedb",
         14935 => x"3884b9c8",
         14936 => x"08831734",
         14937 => x"b41608a8",
         14938 => x"17083184",
         14939 => x"b9c80859",
         14940 => x"5574a017",
         14941 => x"0827fea0",
         14942 => x"38821633",
         14943 => x"5d7c822e",
         14944 => x"098106fe",
         14945 => x"93388154",
         14946 => x"b41608a0",
         14947 => x"17080553",
         14948 => x"7b528116",
         14949 => x"3351fee1",
         14950 => x"c93f7958",
         14951 => x"fdfa3981",
         14952 => x"54b41708",
         14953 => x"53b81770",
         14954 => x"53811833",
         14955 => x"525bfee1",
         14956 => x"b13f815c",
         14957 => x"84b9c808",
         14958 => x"fcc93884",
         14959 => x"b9c80883",
         14960 => x"1834b417",
         14961 => x"08a81808",
         14962 => x"3184b9c8",
         14963 => x"085d5574",
         14964 => x"a0180827",
         14965 => x"fc8e3882",
         14966 => x"17335d7c",
         14967 => x"822e0981",
         14968 => x"06fc8138",
         14969 => x"8154b417",
         14970 => x"08a01808",
         14971 => x"05537a52",
         14972 => x"81173351",
         14973 => x"fee0eb3f",
         14974 => x"795cfbe8",
         14975 => x"39ec3d0d",
         14976 => x"0280df05",
         14977 => x"33028405",
         14978 => x"80e30533",
         14979 => x"56578253",
         14980 => x"963dcc05",
         14981 => x"52973d51",
         14982 => x"ffa2d83f",
         14983 => x"84b9c808",
         14984 => x"5684b9c8",
         14985 => x"08802e8a",
         14986 => x"387584b9",
         14987 => x"c80c963d",
         14988 => x"0d04785a",
         14989 => x"6652963d",
         14990 => x"d00551ff",
         14991 => x"96d73f84",
         14992 => x"b9c80856",
         14993 => x"84b9c808",
         14994 => x"e0380280",
         14995 => x"cf053381",
         14996 => x"a0065486",
         14997 => x"5673d238",
         14998 => x"74a70661",
         14999 => x"71098b12",
         15000 => x"3371067a",
         15001 => x"74060751",
         15002 => x"56575573",
         15003 => x"8b173478",
         15004 => x"55810b83",
         15005 => x"16347851",
         15006 => x"fee29a3f",
         15007 => x"84b9c808",
         15008 => x"84b9c80c",
         15009 => x"963d0d04",
         15010 => x"ec3d0d67",
         15011 => x"57825396",
         15012 => x"3dcc0552",
         15013 => x"973d51ff",
         15014 => x"a1d93f84",
         15015 => x"b9c80855",
         15016 => x"84b9c808",
         15017 => x"802e8a38",
         15018 => x"7484b9c8",
         15019 => x"0c963d0d",
         15020 => x"04785a66",
         15021 => x"52963dd0",
         15022 => x"0551ff95",
         15023 => x"d83f84b9",
         15024 => x"c8085584",
         15025 => x"b9c808e0",
         15026 => x"380280cf",
         15027 => x"053381a0",
         15028 => x"06568655",
         15029 => x"75d23860",
         15030 => x"84182286",
         15031 => x"19227190",
         15032 => x"2b075959",
         15033 => x"56769617",
         15034 => x"3476882a",
         15035 => x"55749717",
         15036 => x"3476902a",
         15037 => x"58779817",
         15038 => x"3476982a",
         15039 => x"54739917",
         15040 => x"34785781",
         15041 => x"0b831834",
         15042 => x"7851fee1",
         15043 => x"883f84b9",
         15044 => x"c80884b9",
         15045 => x"c80c963d",
         15046 => x"0d04e83d",
         15047 => x"0d6b6d5d",
         15048 => x"5b80539a",
         15049 => x"3dcc0552",
         15050 => x"9b3d51ff",
         15051 => x"a0c53f84",
         15052 => x"b9c80884",
         15053 => x"b9c80830",
         15054 => x"7084b9c8",
         15055 => x"08078025",
         15056 => x"5156577a",
         15057 => x"802e8b38",
         15058 => x"81707606",
         15059 => x"5a567881",
         15060 => x"a4387630",
         15061 => x"70780780",
         15062 => x"25565b7b",
         15063 => x"802e818c",
         15064 => x"38817076",
         15065 => x"065a5878",
         15066 => x"802e8180",
         15067 => x"387ca411",
         15068 => x"08585680",
         15069 => x"5ab41608",
         15070 => x"772e82f6",
         15071 => x"38831633",
         15072 => x"7a5a5574",
         15073 => x"7a2e0981",
         15074 => x"06819838",
         15075 => x"81547653",
         15076 => x"b8165281",
         15077 => x"163351fe",
         15078 => x"dcc93f84",
         15079 => x"b9c80880",
         15080 => x"2e8538ff",
         15081 => x"57815976",
         15082 => x"b4170c78",
         15083 => x"5778bd38",
         15084 => x"7c703356",
         15085 => x"5880c356",
         15086 => x"74832e8b",
         15087 => x"3880e456",
         15088 => x"74842e83",
         15089 => x"38a75675",
         15090 => x"18b80583",
         15091 => x"11338212",
         15092 => x"3371902b",
         15093 => x"71882b07",
         15094 => x"81143370",
         15095 => x"7207882b",
         15096 => x"75337107",
         15097 => x"620c5f5d",
         15098 => x"5e575956",
         15099 => x"7684b9c8",
         15100 => x"0c9a3d0d",
         15101 => x"047c5e80",
         15102 => x"4080528e",
         15103 => x"3d705255",
         15104 => x"fef48b3f",
         15105 => x"84b9c808",
         15106 => x"5784b9c8",
         15107 => x"08802e81",
         15108 => x"8d387684",
         15109 => x"2e098106",
         15110 => x"feb83880",
         15111 => x"7b348057",
         15112 => x"feb03977",
         15113 => x"54b41608",
         15114 => x"53b81670",
         15115 => x"53811733",
         15116 => x"525bfedc",
         15117 => x"ad3f7759",
         15118 => x"84b9c808",
         15119 => x"7a2e0981",
         15120 => x"06fee838",
         15121 => x"84b9c808",
         15122 => x"831734b4",
         15123 => x"1608a817",
         15124 => x"083184b9",
         15125 => x"c8085a55",
         15126 => x"74a01708",
         15127 => x"27fead38",
         15128 => x"82163355",
         15129 => x"74822e09",
         15130 => x"8106fea0",
         15131 => x"387754b4",
         15132 => x"1608a017",
         15133 => x"0805537a",
         15134 => x"52811633",
         15135 => x"51fedbe2",
         15136 => x"3f795981",
         15137 => x"547653b8",
         15138 => x"16528116",
         15139 => x"3351feda",
         15140 => x"d23f84b9",
         15141 => x"c808802e",
         15142 => x"fe8d38fe",
         15143 => x"86397552",
         15144 => x"7451fef8",
         15145 => x"bb3f84b9",
         15146 => x"c8085784",
         15147 => x"b9c808fe",
         15148 => x"e13884b9",
         15149 => x"c80884b9",
         15150 => x"c808665c",
         15151 => x"59597918",
         15152 => x"81197c1b",
         15153 => x"57595675",
         15154 => x"33753481",
         15155 => x"19598a78",
         15156 => x"27ec388b",
         15157 => x"701c5758",
         15158 => x"80763477",
         15159 => x"802efcf2",
         15160 => x"38ff187b",
         15161 => x"1170335c",
         15162 => x"575879a0",
         15163 => x"2eea38fc",
         15164 => x"e1397957",
         15165 => x"fdba39e1",
         15166 => x"3d0d8253",
         15167 => x"a13dffb4",
         15168 => x"0552a23d",
         15169 => x"51ff9ceb",
         15170 => x"3f84b9c8",
         15171 => x"085684b9",
         15172 => x"c80882a6",
         15173 => x"388f3d5d",
         15174 => x"8b7d5755",
         15175 => x"a0767081",
         15176 => x"055834ff",
         15177 => x"155574f4",
         15178 => x"3874a33d",
         15179 => x"08703370",
         15180 => x"81ff065b",
         15181 => x"58585a9f",
         15182 => x"782781b7",
         15183 => x"38a23d90",
         15184 => x"3d5c5c75",
         15185 => x"81ff0681",
         15186 => x"18575574",
         15187 => x"81f53875",
         15188 => x"7c0c7483",
         15189 => x"ffff2681",
         15190 => x"ff387451",
         15191 => x"a1953f83",
         15192 => x"b55284b9",
         15193 => x"c808519f",
         15194 => x"dc3f84b9",
         15195 => x"c80883ff",
         15196 => x"ff065776",
         15197 => x"802e81e0",
         15198 => x"3883e6d8",
         15199 => x"0b83e6d8",
         15200 => x"337081ff",
         15201 => x"065b5658",
         15202 => x"78802e81",
         15203 => x"d6387456",
         15204 => x"78772e99",
         15205 => x"38811870",
         15206 => x"337081ff",
         15207 => x"06575758",
         15208 => x"74802e89",
         15209 => x"3874772e",
         15210 => x"098106e9",
         15211 => x"387581ff",
         15212 => x"06597881",
         15213 => x"a33881ff",
         15214 => x"772781f8",
         15215 => x"38798926",
         15216 => x"81963881",
         15217 => x"ff77278f",
         15218 => x"3876882a",
         15219 => x"55747b70",
         15220 => x"81055d34",
         15221 => x"811a5a76",
         15222 => x"7b708105",
         15223 => x"5d34811a",
         15224 => x"a33d0870",
         15225 => x"337081ff",
         15226 => x"065b5858",
         15227 => x"5a779f26",
         15228 => x"fed1388f",
         15229 => x"3d335786",
         15230 => x"567681e5",
         15231 => x"2ebc3879",
         15232 => x"802e9938",
         15233 => x"02b70556",
         15234 => x"79167033",
         15235 => x"5c5c7aa0",
         15236 => x"2e098106",
         15237 => x"8738ff1a",
         15238 => x"5a79ed38",
         15239 => x"7d458047",
         15240 => x"8052953d",
         15241 => x"705256fe",
         15242 => x"efe43f84",
         15243 => x"b9c80855",
         15244 => x"84b9c808",
         15245 => x"802eb438",
         15246 => x"74567584",
         15247 => x"b9c80ca1",
         15248 => x"3d0d0483",
         15249 => x"b5527451",
         15250 => x"9ee73f84",
         15251 => x"b9c80883",
         15252 => x"ffff0655",
         15253 => x"74fdf838",
         15254 => x"86567584",
         15255 => x"b9c80ca1",
         15256 => x"3d0d0483",
         15257 => x"e6d83356",
         15258 => x"fec33981",
         15259 => x"527551fe",
         15260 => x"f4ee3f84",
         15261 => x"b9c80855",
         15262 => x"84b9c808",
         15263 => x"80c13879",
         15264 => x"802e82c4",
         15265 => x"388b6c7e",
         15266 => x"59575576",
         15267 => x"70810558",
         15268 => x"33767081",
         15269 => x"055834ff",
         15270 => x"155574ef",
         15271 => x"387d5d81",
         15272 => x"0b831e34",
         15273 => x"7d51fed9",
         15274 => x"ec3f84b9",
         15275 => x"c8085574",
         15276 => x"56ff8739",
         15277 => x"8a7a27fe",
         15278 => x"8a388656",
         15279 => x"ff9c3984",
         15280 => x"b9c80884",
         15281 => x"2e098106",
         15282 => x"feee3880",
         15283 => x"5579752e",
         15284 => x"fee63875",
         15285 => x"08755376",
         15286 => x"5258feee",
         15287 => x"b13f84b9",
         15288 => x"c8085784",
         15289 => x"b9c80875",
         15290 => x"2e098106",
         15291 => x"81843884",
         15292 => x"b9c808b8",
         15293 => x"195c5a98",
         15294 => x"16085780",
         15295 => x"59b41808",
         15296 => x"772eb238",
         15297 => x"83183355",
         15298 => x"74792e09",
         15299 => x"810681d7",
         15300 => x"38815476",
         15301 => x"53b81852",
         15302 => x"81183351",
         15303 => x"fed5c43f",
         15304 => x"84b9c808",
         15305 => x"802e8538",
         15306 => x"ff578159",
         15307 => x"76b4190c",
         15308 => x"785778be",
         15309 => x"38789c17",
         15310 => x"08703357",
         15311 => x"5a577481",
         15312 => x"e52e819e",
         15313 => x"38743070",
         15314 => x"80257807",
         15315 => x"565c7480",
         15316 => x"2e81d738",
         15317 => x"811a5a79",
         15318 => x"812ea538",
         15319 => x"81527551",
         15320 => x"feefa13f",
         15321 => x"84b9c808",
         15322 => x"5784b9c8",
         15323 => x"08802eff",
         15324 => x"86388755",
         15325 => x"76842efd",
         15326 => x"bf387655",
         15327 => x"76fdb938",
         15328 => x"a06c5755",
         15329 => x"80767081",
         15330 => x"055834ff",
         15331 => x"155574f4",
         15332 => x"386b5688",
         15333 => x"0b8b1734",
         15334 => x"8b6c7e59",
         15335 => x"57557670",
         15336 => x"81055833",
         15337 => x"76708105",
         15338 => x"5834ff15",
         15339 => x"5574802e",
         15340 => x"fdeb3876",
         15341 => x"70810558",
         15342 => x"33767081",
         15343 => x"055834ff",
         15344 => x"155574da",
         15345 => x"38fdd639",
         15346 => x"6b5ae57a",
         15347 => x"347d5d81",
         15348 => x"0b831e34",
         15349 => x"7d51fed7",
         15350 => x"bc3f84b9",
         15351 => x"c80855fd",
         15352 => x"ce398157",
         15353 => x"fedf3981",
         15354 => x"54b41808",
         15355 => x"537a5281",
         15356 => x"183351fe",
         15357 => x"d4ec3f84",
         15358 => x"b9c80879",
         15359 => x"2e098106",
         15360 => x"80c33884",
         15361 => x"b9c80883",
         15362 => x"1934b418",
         15363 => x"08a81908",
         15364 => x"315c7ba0",
         15365 => x"1908278a",
         15366 => x"38821833",
         15367 => x"5574822e",
         15368 => x"b13884b9",
         15369 => x"c80859fd",
         15370 => x"e839745a",
         15371 => x"81527551",
         15372 => x"feedd13f",
         15373 => x"84b9c808",
         15374 => x"5784b9c8",
         15375 => x"08802efd",
         15376 => x"b638feae",
         15377 => x"39817058",
         15378 => x"5978802e",
         15379 => x"fde738fe",
         15380 => x"a1398154",
         15381 => x"b41808a0",
         15382 => x"19080553",
         15383 => x"7a528118",
         15384 => x"3351fed3",
         15385 => x"fd3ffda9",
         15386 => x"39f23d0d",
         15387 => x"60620288",
         15388 => x"0580cb05",
         15389 => x"335e5b57",
         15390 => x"89567680",
         15391 => x"2e9f3876",
         15392 => x"08557480",
         15393 => x"2e973874",
         15394 => x"33547380",
         15395 => x"2e8f3886",
         15396 => x"15228418",
         15397 => x"22595978",
         15398 => x"782e81c2",
         15399 => x"38805473",
         15400 => x"5f7581a5",
         15401 => x"38911733",
         15402 => x"5675819d",
         15403 => x"3879802e",
         15404 => x"81a2388c",
         15405 => x"1708819c",
         15406 => x"38901733",
         15407 => x"70812a81",
         15408 => x"06565d74",
         15409 => x"802e818c",
         15410 => x"387e8a11",
         15411 => x"2270892b",
         15412 => x"70557c54",
         15413 => x"575c59fd",
         15414 => x"87cb3fff",
         15415 => x"157a0670",
         15416 => x"30707207",
         15417 => x"9f2a84b9",
         15418 => x"c8080590",
         15419 => x"1c087942",
         15420 => x"535f5558",
         15421 => x"81782788",
         15422 => x"389c1908",
         15423 => x"78268338",
         15424 => x"82587778",
         15425 => x"565b8059",
         15426 => x"74527651",
         15427 => x"fed8873f",
         15428 => x"81157f55",
         15429 => x"559c1408",
         15430 => x"75268338",
         15431 => x"825584b9",
         15432 => x"c808812e",
         15433 => x"81dc3884",
         15434 => x"b9c808ff",
         15435 => x"2e81d838",
         15436 => x"84b9c808",
         15437 => x"81c53881",
         15438 => x"1959787d",
         15439 => x"2ebb3874",
         15440 => x"782e0981",
         15441 => x"06c23887",
         15442 => x"56755473",
         15443 => x"84b9c80c",
         15444 => x"903d0d04",
         15445 => x"870b84b9",
         15446 => x"c80c903d",
         15447 => x"0d048115",
         15448 => x"3351fed0",
         15449 => x"ac3f84b9",
         15450 => x"c8088106",
         15451 => x"5473fead",
         15452 => x"38737708",
         15453 => x"5556fea7",
         15454 => x"397b802e",
         15455 => x"818e387a",
         15456 => x"7d56587c",
         15457 => x"802eab38",
         15458 => x"81185474",
         15459 => x"812e80e6",
         15460 => x"38735377",
         15461 => x"527e51fe",
         15462 => x"dddd3f84",
         15463 => x"b9c80856",
         15464 => x"84b9c808",
         15465 => x"ffa33877",
         15466 => x"8119ff17",
         15467 => x"57595e74",
         15468 => x"d7387e7e",
         15469 => x"90120c55",
         15470 => x"7b802eff",
         15471 => x"8c387a88",
         15472 => x"180c798c",
         15473 => x"180c9017",
         15474 => x"3380c007",
         15475 => x"5c7b9018",
         15476 => x"349c1508",
         15477 => x"fe059416",
         15478 => x"08585a76",
         15479 => x"7a26fee9",
         15480 => x"38767d31",
         15481 => x"94160c84",
         15482 => x"15338107",
         15483 => x"5d7c8416",
         15484 => x"347554fe",
         15485 => x"d639ff54",
         15486 => x"ff973974",
         15487 => x"5b8059fe",
         15488 => x"be398254",
         15489 => x"fec53981",
         15490 => x"54fec039",
         15491 => x"ff1b5eff",
         15492 => x"a13984b9",
         15493 => x"d408e33d",
         15494 => x"0da33d08",
         15495 => x"a53d0802",
         15496 => x"88058187",
         15497 => x"05334442",
         15498 => x"5fff0ba2",
         15499 => x"3d08705f",
         15500 => x"5b407980",
         15501 => x"2e858a38",
         15502 => x"79708105",
         15503 => x"5b33709f",
         15504 => x"26565675",
         15505 => x"ba2e859b",
         15506 => x"3874ed38",
         15507 => x"75ba2e85",
         15508 => x"923884d1",
         15509 => x"a4335680",
         15510 => x"762484e5",
         15511 => x"38751010",
         15512 => x"84d19005",
         15513 => x"7008565a",
         15514 => x"74802e84",
         15515 => x"38807534",
         15516 => x"751684b9",
         15517 => x"bc113384",
         15518 => x"b9bd1233",
         15519 => x"405b5d81",
         15520 => x"527951fe",
         15521 => x"cea93f84",
         15522 => x"b9c80881",
         15523 => x"ff067081",
         15524 => x"065d5683",
         15525 => x"577b84ab",
         15526 => x"3875822a",
         15527 => x"8106408a",
         15528 => x"577f849f",
         15529 => x"389f3dfc",
         15530 => x"05538352",
         15531 => x"7951fed0",
         15532 => x"b03f84b9",
         15533 => x"c8088498",
         15534 => x"386d5574",
         15535 => x"802e8490",
         15536 => x"38748280",
         15537 => x"80268488",
         15538 => x"38ff1575",
         15539 => x"06557483",
         15540 => x"ff387e80",
         15541 => x"2e883884",
         15542 => x"807f2683",
         15543 => x"f8387e81",
         15544 => x"800a2683",
         15545 => x"f038ff1f",
         15546 => x"7f065574",
         15547 => x"83e7387e",
         15548 => x"892aa63d",
         15549 => x"08892a70",
         15550 => x"892b7759",
         15551 => x"4c475b60",
         15552 => x"802e85ab",
         15553 => x"38653070",
         15554 => x"80257707",
         15555 => x"565f9157",
         15556 => x"7483b038",
         15557 => x"7d802e84",
         15558 => x"df388154",
         15559 => x"74536052",
         15560 => x"7951fecd",
         15561 => x"be3f8157",
         15562 => x"84b9c808",
         15563 => x"83953860",
         15564 => x"83ff0533",
         15565 => x"6183fe05",
         15566 => x"3371882b",
         15567 => x"0759568e",
         15568 => x"577782d4",
         15569 => x"d52e0981",
         15570 => x"0682f838",
         15571 => x"7d902961",
         15572 => x"0583b211",
         15573 => x"33445862",
         15574 => x"802e82e7",
         15575 => x"3883b618",
         15576 => x"83113382",
         15577 => x"12337190",
         15578 => x"2b71882b",
         15579 => x"07811433",
         15580 => x"70720788",
         15581 => x"2b753371",
         15582 => x"0783ba1f",
         15583 => x"83113382",
         15584 => x"12337190",
         15585 => x"2b71882b",
         15586 => x"07811433",
         15587 => x"70720788",
         15588 => x"2b753371",
         15589 => x"075ca23d",
         15590 => x"0c42a33d",
         15591 => x"0ca33d0c",
         15592 => x"444e5445",
         15593 => x"594f415a",
         15594 => x"4b784d8e",
         15595 => x"5780ff79",
         15596 => x"27829038",
         15597 => x"93577a81",
         15598 => x"80268287",
         15599 => x"3861812a",
         15600 => x"70810645",
         15601 => x"4963802e",
         15602 => x"83f93861",
         15603 => x"87064564",
         15604 => x"822e8938",
         15605 => x"61810647",
         15606 => x"6683f438",
         15607 => x"836e7030",
         15608 => x"4a46437a",
         15609 => x"5862832e",
         15610 => x"8ac2387a",
         15611 => x"ae38788c",
         15612 => x"2a57810b",
         15613 => x"83e6ec22",
         15614 => x"56587480",
         15615 => x"2e9d3874",
         15616 => x"77269838",
         15617 => x"83e6ec56",
         15618 => x"77108217",
         15619 => x"70225757",
         15620 => x"5874802e",
         15621 => x"86387675",
         15622 => x"27ee3877",
         15623 => x"527851fd",
         15624 => x"81833f84",
         15625 => x"b9c80810",
         15626 => x"84055584",
         15627 => x"b9c8089f",
         15628 => x"f5269638",
         15629 => x"810b84b9",
         15630 => x"c8081084",
         15631 => x"b9c80805",
         15632 => x"7111722a",
         15633 => x"8305574c",
         15634 => x"4383ff15",
         15635 => x"892a5d81",
         15636 => x"5ca0477b",
         15637 => x"1f7d1168",
         15638 => x"056611ff",
         15639 => x"05706b06",
         15640 => x"7231584e",
         15641 => x"57446283",
         15642 => x"2e89b838",
         15643 => x"741d5d77",
         15644 => x"90291670",
         15645 => x"60315657",
         15646 => x"74792682",
         15647 => x"f238787c",
         15648 => x"317d3178",
         15649 => x"53706831",
         15650 => x"5256fd80",
         15651 => x"983f84b9",
         15652 => x"c8084062",
         15653 => x"832e89f6",
         15654 => x"3862822e",
         15655 => x"09810682",
         15656 => x"dd3883ff",
         15657 => x"f50b84b9",
         15658 => x"c8082782",
         15659 => x"ac387a89",
         15660 => x"f9387718",
         15661 => x"557480c0",
         15662 => x"2689ef38",
         15663 => x"745bfea3",
         15664 => x"398b5776",
         15665 => x"84b9c80c",
         15666 => x"9f3d0d84",
         15667 => x"b9d40c04",
         15668 => x"814efbfe",
         15669 => x"39930b84",
         15670 => x"b9c80c9f",
         15671 => x"3d0d84b9",
         15672 => x"d40c047c",
         15673 => x"33d01170",
         15674 => x"81ff0657",
         15675 => x"57577489",
         15676 => x"26913882",
         15677 => x"1d7781ff",
         15678 => x"06d0055d",
         15679 => x"58777a2e",
         15680 => x"81b23880",
         15681 => x"0b83e5b8",
         15682 => x"5f5c7d08",
         15683 => x"7d575b7a",
         15684 => x"7081055c",
         15685 => x"33767081",
         15686 => x"055833ff",
         15687 => x"9f124559",
         15688 => x"57629926",
         15689 => x"8938e017",
         15690 => x"7081ff06",
         15691 => x"5844ff9f",
         15692 => x"18456499",
         15693 => x"268938e0",
         15694 => x"187081ff",
         15695 => x"06594676",
         15696 => x"30709f2a",
         15697 => x"5a477678",
         15698 => x"2e098106",
         15699 => x"853878ff",
         15700 => x"be38757a",
         15701 => x"32703070",
         15702 => x"72079f2a",
         15703 => x"7b075d4a",
         15704 => x"4a7a802e",
         15705 => x"80ce3881",
         15706 => x"1c841f5f",
         15707 => x"5c837c25",
         15708 => x"ff98387f",
         15709 => x"56f9e039",
         15710 => x"9f3df805",
         15711 => x"53815279",
         15712 => x"51fecadd",
         15713 => x"3f815784",
         15714 => x"b9c808fe",
         15715 => x"b6386183",
         15716 => x"2a770684",
         15717 => x"b9c80840",
         15718 => x"56758338",
         15719 => x"bf5f6c55",
         15720 => x"8e577e75",
         15721 => x"26fe9c38",
         15722 => x"747f3159",
         15723 => x"fbfb3981",
         15724 => x"56fad239",
         15725 => x"7b8324ff",
         15726 => x"ba387b7a",
         15727 => x"a33d0c56",
         15728 => x"f9953961",
         15729 => x"81064893",
         15730 => x"5767802e",
         15731 => x"fdf53882",
         15732 => x"6e70304a",
         15733 => x"4643fc8b",
         15734 => x"3984b9c8",
         15735 => x"089ff526",
         15736 => x"9d387a8b",
         15737 => x"3877185b",
         15738 => x"81807b27",
         15739 => x"fbf5388e",
         15740 => x"577684b9",
         15741 => x"c80c9f3d",
         15742 => x"0d84b9d4",
         15743 => x"0c048055",
         15744 => x"62812e86",
         15745 => x"99389ff5",
         15746 => x"60278b38",
         15747 => x"7481065b",
         15748 => x"8e577afd",
         15749 => x"ae388480",
         15750 => x"61575580",
         15751 => x"76708105",
         15752 => x"5834ff15",
         15753 => x"5574f438",
         15754 => x"8b6183e5",
         15755 => x"84595755",
         15756 => x"76708105",
         15757 => x"58337670",
         15758 => x"81055834",
         15759 => x"ff155574",
         15760 => x"ef38608b",
         15761 => x"05457465",
         15762 => x"3482618c",
         15763 => x"05347761",
         15764 => x"8d05347b",
         15765 => x"83ffff06",
         15766 => x"4b6a618e",
         15767 => x"05346a88",
         15768 => x"2a5c7b61",
         15769 => x"8f053481",
         15770 => x"61900534",
         15771 => x"62833270",
         15772 => x"305a4880",
         15773 => x"61910534",
         15774 => x"789e2a82",
         15775 => x"06496861",
         15776 => x"9205346c",
         15777 => x"567583ff",
         15778 => x"ff2686ad",
         15779 => x"387583ff",
         15780 => x"ff065574",
         15781 => x"61930534",
         15782 => x"74882a4c",
         15783 => x"6b619405",
         15784 => x"34f86195",
         15785 => x"0534bf61",
         15786 => x"98053480",
         15787 => x"61990534",
         15788 => x"ff619a05",
         15789 => x"3480619b",
         15790 => x"05347e61",
         15791 => x"9c05347e",
         15792 => x"882a4867",
         15793 => x"619d0534",
         15794 => x"7e902a4c",
         15795 => x"6b619e05",
         15796 => x"347e982a",
         15797 => x"84b9d40c",
         15798 => x"84b9d408",
         15799 => x"619f0534",
         15800 => x"62832e85",
         15801 => x"f7388061",
         15802 => x"a7053480",
         15803 => x"61a80534",
         15804 => x"a161a905",
         15805 => x"3480cc61",
         15806 => x"aa05347c",
         15807 => x"83ffff06",
         15808 => x"55746196",
         15809 => x"05347488",
         15810 => x"2a4b6a61",
         15811 => x"970534ff",
         15812 => x"8061a405",
         15813 => x"34a961a6",
         15814 => x"05349361",
         15815 => x"ab0583e5",
         15816 => x"90595755",
         15817 => x"76708105",
         15818 => x"58337670",
         15819 => x"81055834",
         15820 => x"ff155574",
         15821 => x"ef386083",
         15822 => x"fe054980",
         15823 => x"d5693460",
         15824 => x"83ff054b",
         15825 => x"ffaa6b34",
         15826 => x"81547e53",
         15827 => x"60527951",
         15828 => x"fec68f3f",
         15829 => x"815784b9",
         15830 => x"c808fae7",
         15831 => x"3860175c",
         15832 => x"62832e87",
         15833 => x"9c386961",
         15834 => x"57558076",
         15835 => x"70810558",
         15836 => x"34ff1555",
         15837 => x"74f43863",
         15838 => x"75415b62",
         15839 => x"832e86c0",
         15840 => x"3887ffff",
         15841 => x"f8576281",
         15842 => x"2e8338f8",
         15843 => x"57766134",
         15844 => x"76882a7c",
         15845 => x"45557464",
         15846 => x"70810546",
         15847 => x"3476902a",
         15848 => x"59786470",
         15849 => x"81054634",
         15850 => x"76982a56",
         15851 => x"7564347c",
         15852 => x"57655976",
         15853 => x"66268338",
         15854 => x"76597854",
         15855 => x"7a536052",
         15856 => x"7951fec5",
         15857 => x"9d3f84b9",
         15858 => x"c80885e6",
         15859 => x"38848061",
         15860 => x"57558076",
         15861 => x"70810558",
         15862 => x"34ff1555",
         15863 => x"74f43878",
         15864 => x"1b777a31",
         15865 => x"585b76c9",
         15866 => x"387f8105",
         15867 => x"407f802e",
         15868 => x"ff893877",
         15869 => x"5662832e",
         15870 => x"83386656",
         15871 => x"65557566",
         15872 => x"26833875",
         15873 => x"5574547a",
         15874 => x"53605279",
         15875 => x"51fec4d2",
         15876 => x"3f84b9c8",
         15877 => x"08859b38",
         15878 => x"741b7676",
         15879 => x"31575b75",
         15880 => x"db388c58",
         15881 => x"62832e93",
         15882 => x"3886586c",
         15883 => x"83ffff26",
         15884 => x"8a388458",
         15885 => x"62822e83",
         15886 => x"3881587d",
         15887 => x"84c13861",
         15888 => x"832a8106",
         15889 => x"5e7d81b3",
         15890 => x"38848061",
         15891 => x"56598075",
         15892 => x"70810557",
         15893 => x"34ff1959",
         15894 => x"78f43880",
         15895 => x"d56934ff",
         15896 => x"aa6b3460",
         15897 => x"83be0547",
         15898 => x"78673481",
         15899 => x"67810534",
         15900 => x"81678205",
         15901 => x"34786783",
         15902 => x"05347767",
         15903 => x"8405346c",
         15904 => x"4380fdc1",
         15905 => x"52621f51",
         15906 => x"fcf89a3f",
         15907 => x"fe678505",
         15908 => x"3484b9c8",
         15909 => x"08822abf",
         15910 => x"07577667",
         15911 => x"86053484",
         15912 => x"b9c80867",
         15913 => x"8705347e",
         15914 => x"6183c605",
         15915 => x"34676183",
         15916 => x"c705346b",
         15917 => x"6183c805",
         15918 => x"3484b9d4",
         15919 => x"086183c9",
         15920 => x"05346261",
         15921 => x"83ca0534",
         15922 => x"62882a45",
         15923 => x"646183cb",
         15924 => x"05346290",
         15925 => x"2a587761",
         15926 => x"83cc0534",
         15927 => x"62982a5f",
         15928 => x"7e6183cd",
         15929 => x"05348154",
         15930 => x"78536052",
         15931 => x"7951fec2",
         15932 => x"f13f8157",
         15933 => x"84b9c808",
         15934 => x"f7c93880",
         15935 => x"53805279",
         15936 => x"51fec3dd",
         15937 => x"3f815784",
         15938 => x"b9c808f7",
         15939 => x"b63884b9",
         15940 => x"c80884b9",
         15941 => x"c80c9f3d",
         15942 => x"0d84b9d4",
         15943 => x"0c046255",
         15944 => x"f9e43974",
         15945 => x"1c641645",
         15946 => x"5cf6c439",
         15947 => x"7aae3878",
         15948 => x"912a5781",
         15949 => x"0b83e6fc",
         15950 => x"22565874",
         15951 => x"802e9d38",
         15952 => x"74772698",
         15953 => x"3883e6fc",
         15954 => x"56771082",
         15955 => x"17702257",
         15956 => x"57587480",
         15957 => x"2e863876",
         15958 => x"7527ee38",
         15959 => x"77527851",
         15960 => x"fcf6c23f",
         15961 => x"84b9c808",
         15962 => x"10108487",
         15963 => x"0570892a",
         15964 => x"5e5ca05c",
         15965 => x"800b84b9",
         15966 => x"c808fc80",
         15967 => x"8a055847",
         15968 => x"fdfff00a",
         15969 => x"7727f5cb",
         15970 => x"388e57f8",
         15971 => x"e43984b9",
         15972 => x"c80883ff",
         15973 => x"f526f8e6",
         15974 => x"387af8d3",
         15975 => x"3877812a",
         15976 => x"5b7af4bf",
         15977 => x"388e57f8",
         15978 => x"c8396881",
         15979 => x"06446380",
         15980 => x"2ef8af38",
         15981 => x"8343f4ab",
         15982 => x"397561a0",
         15983 => x"05347588",
         15984 => x"2a496861",
         15985 => x"a1053475",
         15986 => x"902a5b7a",
         15987 => x"61a20534",
         15988 => x"75982a57",
         15989 => x"7661a305",
         15990 => x"34f9c639",
         15991 => x"806180c3",
         15992 => x"05348061",
         15993 => x"80c40534",
         15994 => x"a16180c5",
         15995 => x"053480cc",
         15996 => x"6180c605",
         15997 => x"347c61a4",
         15998 => x"05347c88",
         15999 => x"2a5c7b61",
         16000 => x"a505347c",
         16001 => x"902a5978",
         16002 => x"61a60534",
         16003 => x"7c982a56",
         16004 => x"7561a705",
         16005 => x"348261ac",
         16006 => x"05348061",
         16007 => x"ad053480",
         16008 => x"61ae0534",
         16009 => x"8061af05",
         16010 => x"348161b0",
         16011 => x"05348061",
         16012 => x"b1053486",
         16013 => x"61b20534",
         16014 => x"8061b305",
         16015 => x"34ff8061",
         16016 => x"80c00534",
         16017 => x"a96180c2",
         16018 => x"05349361",
         16019 => x"80c70583",
         16020 => x"e5a45957",
         16021 => x"55767081",
         16022 => x"05583376",
         16023 => x"70810558",
         16024 => x"34ff1555",
         16025 => x"74802ef9",
         16026 => x"cd387670",
         16027 => x"81055833",
         16028 => x"76708105",
         16029 => x"5834ff15",
         16030 => x"5574da38",
         16031 => x"f9b83981",
         16032 => x"54805360",
         16033 => x"527951fe",
         16034 => x"bed93f81",
         16035 => x"5784b9c8",
         16036 => x"08f4b038",
         16037 => x"7d902961",
         16038 => x"05427762",
         16039 => x"83b20534",
         16040 => x"765484b9",
         16041 => x"c8085360",
         16042 => x"527951fe",
         16043 => x"bfb43ffc",
         16044 => x"c339810b",
         16045 => x"84b9c80c",
         16046 => x"9f3d0d84",
         16047 => x"b9d40c04",
         16048 => x"f861347b",
         16049 => x"4aff6a70",
         16050 => x"81054c34",
         16051 => x"ff6a7081",
         16052 => x"054c34ff",
         16053 => x"6a34ff61",
         16054 => x"840534ff",
         16055 => x"61850534",
         16056 => x"ff618605",
         16057 => x"34ff6187",
         16058 => x"0534ff61",
         16059 => x"880534ff",
         16060 => x"61890534",
         16061 => x"ff618a05",
         16062 => x"348f6534",
         16063 => x"7c57f9b1",
         16064 => x"39765486",
         16065 => x"1f536052",
         16066 => x"7951febe",
         16067 => x"d53f8480",
         16068 => x"61565780",
         16069 => x"75708105",
         16070 => x"5734ff17",
         16071 => x"5776f438",
         16072 => x"605c80d2",
         16073 => x"7c708105",
         16074 => x"5e347b55",
         16075 => x"80d27570",
         16076 => x"81055734",
         16077 => x"80e17570",
         16078 => x"81055734",
         16079 => x"80c17534",
         16080 => x"80f26183",
         16081 => x"e4053480",
         16082 => x"f26183e5",
         16083 => x"053480c1",
         16084 => x"6183e605",
         16085 => x"3480e161",
         16086 => x"83e70534",
         16087 => x"7fff055b",
         16088 => x"7a6183e8",
         16089 => x"05347a88",
         16090 => x"2a597861",
         16091 => x"83e90534",
         16092 => x"7a902a56",
         16093 => x"756183ea",
         16094 => x"05347a98",
         16095 => x"2a407f61",
         16096 => x"83eb0534",
         16097 => x"826183ec",
         16098 => x"05347661",
         16099 => x"83ed0534",
         16100 => x"766183ee",
         16101 => x"05347661",
         16102 => x"83ef0534",
         16103 => x"80d56934",
         16104 => x"ffaa6b34",
         16105 => x"8154871f",
         16106 => x"53605279",
         16107 => x"51febdb2",
         16108 => x"3f815481",
         16109 => x"1f536052",
         16110 => x"7951febd",
         16111 => x"a53f6961",
         16112 => x"5755f7a6",
         16113 => x"39f43d0d",
         16114 => x"7e615b5b",
         16115 => x"807b61ff",
         16116 => x"055a5757",
         16117 => x"767825b8",
         16118 => x"388d3d59",
         16119 => x"8e3df805",
         16120 => x"54815378",
         16121 => x"527951ff",
         16122 => x"9ab43f7b",
         16123 => x"812e0981",
         16124 => x"069e388d",
         16125 => x"3d335574",
         16126 => x"8d2e9038",
         16127 => x"74767081",
         16128 => x"05583481",
         16129 => x"1757748a",
         16130 => x"2e863877",
         16131 => x"7724cd38",
         16132 => x"8076347a",
         16133 => x"55768338",
         16134 => x"76557484",
         16135 => x"b9c80c8e",
         16136 => x"3d0d04f7",
         16137 => x"3d0d7b02",
         16138 => x"8405b305",
         16139 => x"33595777",
         16140 => x"8a2e80d5",
         16141 => x"38841708",
         16142 => x"56807624",
         16143 => x"9e388817",
         16144 => x"0877178c",
         16145 => x"05565977",
         16146 => x"75348116",
         16147 => x"5574bb24",
         16148 => x"8e387484",
         16149 => x"180c8119",
         16150 => x"88180c8b",
         16151 => x"3d0d048b",
         16152 => x"3dfc0554",
         16153 => x"74538c17",
         16154 => x"52760851",
         16155 => x"ff9ed13f",
         16156 => x"747a3270",
         16157 => x"30707207",
         16158 => x"9f2a7030",
         16159 => x"841b0c81",
         16160 => x"1c881b0c",
         16161 => x"5a5656d3",
         16162 => x"398d5276",
         16163 => x"51ff943f",
         16164 => x"ffa339e3",
         16165 => x"3d0d0280",
         16166 => x"ff05338d",
         16167 => x"3d585880",
         16168 => x"cc775755",
         16169 => x"80767081",
         16170 => x"055834ff",
         16171 => x"155574f4",
         16172 => x"38a13d08",
         16173 => x"770c778a",
         16174 => x"2e80f738",
         16175 => x"7c568076",
         16176 => x"2480c038",
         16177 => x"7d77178c",
         16178 => x"05565977",
         16179 => x"75348116",
         16180 => x"5574bb24",
         16181 => x"b8387484",
         16182 => x"180c8119",
         16183 => x"88180c7c",
         16184 => x"55807524",
         16185 => x"9e389f3d",
         16186 => x"ffac1155",
         16187 => x"7554c005",
         16188 => x"52760851",
         16189 => x"ff9dc93f",
         16190 => x"84b9c808",
         16191 => x"86387c7a",
         16192 => x"2eba38ff",
         16193 => x"0b84b9c8",
         16194 => x"0c9f3d0d",
         16195 => x"049f3dff",
         16196 => x"b0115575",
         16197 => x"54c00552",
         16198 => x"760851ff",
         16199 => x"9da23f74",
         16200 => x"7b327030",
         16201 => x"7072079f",
         16202 => x"2a703052",
         16203 => x"5a5656ff",
         16204 => x"a5398d52",
         16205 => x"7651fdeb",
         16206 => x"3fff8139",
         16207 => x"7d84b9c8",
         16208 => x"0c9f3d0d",
         16209 => x"04fd3d0d",
         16210 => x"75028405",
         16211 => x"9a052252",
         16212 => x"53805272",
         16213 => x"80ff2690",
         16214 => x"387283ff",
         16215 => x"ff065271",
         16216 => x"84b9c80c",
         16217 => x"853d0d04",
         16218 => x"83ffff73",
         16219 => x"27547083",
         16220 => x"b52e0981",
         16221 => x"06e93873",
         16222 => x"802ee438",
         16223 => x"83e78c22",
         16224 => x"5172712e",
         16225 => x"9c388112",
         16226 => x"7083ffff",
         16227 => x"06535471",
         16228 => x"80ff268d",
         16229 => x"38711083",
         16230 => x"e78c0570",
         16231 => x"225151e1",
         16232 => x"39818012",
         16233 => x"7081ff06",
         16234 => x"84b9c80c",
         16235 => x"53853d0d",
         16236 => x"04fe3d0d",
         16237 => x"02920522",
         16238 => x"02840596",
         16239 => x"05225351",
         16240 => x"80537080",
         16241 => x"ff268c38",
         16242 => x"70537284",
         16243 => x"b9c80c84",
         16244 => x"3d0d0471",
         16245 => x"83b52e09",
         16246 => x"8106ef38",
         16247 => x"7081ff26",
         16248 => x"e9387010",
         16249 => x"83e58c05",
         16250 => x"702284b9",
         16251 => x"c80c5184",
         16252 => x"3d0d04fb",
         16253 => x"3d0d7751",
         16254 => x"7083ffff",
         16255 => x"2680e138",
         16256 => x"7083ffff",
         16257 => x"0683e98c",
         16258 => x"5656759f",
         16259 => x"ff2680d9",
         16260 => x"38747082",
         16261 => x"05562275",
         16262 => x"71307080",
         16263 => x"25737a26",
         16264 => x"07545653",
         16265 => x"5370b738",
         16266 => x"71708205",
         16267 => x"53227271",
         16268 => x"882a5456",
         16269 => x"81ff0670",
         16270 => x"14525470",
         16271 => x"7624b138",
         16272 => x"71cf3873",
         16273 => x"10157070",
         16274 => x"82055222",
         16275 => x"54733070",
         16276 => x"80257579",
         16277 => x"26075355",
         16278 => x"5270802e",
         16279 => x"cb387551",
         16280 => x"7084b9c8",
         16281 => x"0c873d0d",
         16282 => x"0483ed80",
         16283 => x"55ffa239",
         16284 => x"718826ea",
         16285 => x"38711010",
         16286 => x"83c9e005",
         16287 => x"54730804",
         16288 => x"c7a01670",
         16289 => x"83ffff06",
         16290 => x"57517551",
         16291 => x"d339ffb0",
         16292 => x"167083ff",
         16293 => x"ff065751",
         16294 => x"f1398816",
         16295 => x"7083ffff",
         16296 => x"065751e6",
         16297 => x"39e61670",
         16298 => x"83ffff06",
         16299 => x"5751db39",
         16300 => x"d0167083",
         16301 => x"ffff0657",
         16302 => x"51d039e0",
         16303 => x"167083ff",
         16304 => x"ff065751",
         16305 => x"c539f016",
         16306 => x"7083ffff",
         16307 => x"065751ff",
         16308 => x"b9397573",
         16309 => x"31810676",
         16310 => x"71317083",
         16311 => x"ffff0658",
         16312 => x"5255ffa6",
         16313 => x"39757331",
         16314 => x"10750570",
         16315 => x"225252fe",
         16316 => x"ef390000",
         16317 => x"00ffffff",
         16318 => x"ff00ffff",
         16319 => x"ffff00ff",
         16320 => x"ffffff00",
         16321 => x"0000198b",
         16322 => x"00001980",
         16323 => x"00001975",
         16324 => x"0000196a",
         16325 => x"0000195f",
         16326 => x"00001954",
         16327 => x"00001949",
         16328 => x"0000193e",
         16329 => x"00001933",
         16330 => x"00001928",
         16331 => x"0000191d",
         16332 => x"00001912",
         16333 => x"00001907",
         16334 => x"000018fc",
         16335 => x"000018f1",
         16336 => x"000018e6",
         16337 => x"000018db",
         16338 => x"000018d0",
         16339 => x"000018c5",
         16340 => x"000018ba",
         16341 => x"00001ebf",
         16342 => x"00001f59",
         16343 => x"00001f59",
         16344 => x"00001f59",
         16345 => x"00001f59",
         16346 => x"00001f59",
         16347 => x"00001f59",
         16348 => x"00001f59",
         16349 => x"00001f59",
         16350 => x"00001f59",
         16351 => x"00001f59",
         16352 => x"00001f59",
         16353 => x"00001f59",
         16354 => x"00001f59",
         16355 => x"00001f59",
         16356 => x"00001f59",
         16357 => x"00001f59",
         16358 => x"00001f59",
         16359 => x"00001f59",
         16360 => x"00001f59",
         16361 => x"00001f59",
         16362 => x"00001f59",
         16363 => x"00001f59",
         16364 => x"00001f59",
         16365 => x"00001f59",
         16366 => x"00001f59",
         16367 => x"00001f59",
         16368 => x"00001f59",
         16369 => x"00001f59",
         16370 => x"00001f59",
         16371 => x"00001f59",
         16372 => x"00001f59",
         16373 => x"00001f59",
         16374 => x"00001f59",
         16375 => x"00001f59",
         16376 => x"00001f59",
         16377 => x"00001f59",
         16378 => x"00001f59",
         16379 => x"00001f59",
         16380 => x"00001f59",
         16381 => x"00001f59",
         16382 => x"00001f59",
         16383 => x"00001f59",
         16384 => x"00002471",
         16385 => x"00001f59",
         16386 => x"00001f59",
         16387 => x"00001f59",
         16388 => x"00001f59",
         16389 => x"00001f59",
         16390 => x"00001f59",
         16391 => x"00001f59",
         16392 => x"00001f59",
         16393 => x"00001f59",
         16394 => x"00001f59",
         16395 => x"00001f59",
         16396 => x"00001f59",
         16397 => x"00001f59",
         16398 => x"00001f59",
         16399 => x"00001f59",
         16400 => x"00001f59",
         16401 => x"00002407",
         16402 => x"00002306",
         16403 => x"00001f59",
         16404 => x"0000228a",
         16405 => x"000024a8",
         16406 => x"00002367",
         16407 => x"0000222c",
         16408 => x"000021ce",
         16409 => x"00001f59",
         16410 => x"00001f59",
         16411 => x"00001f59",
         16412 => x"00001f59",
         16413 => x"00001f59",
         16414 => x"00001f59",
         16415 => x"00001f59",
         16416 => x"00001f59",
         16417 => x"00001f59",
         16418 => x"00001f59",
         16419 => x"00001f59",
         16420 => x"00001f59",
         16421 => x"00001f59",
         16422 => x"00001f59",
         16423 => x"00001f59",
         16424 => x"00001f59",
         16425 => x"00001f59",
         16426 => x"00001f59",
         16427 => x"00001f59",
         16428 => x"00001f59",
         16429 => x"00001f59",
         16430 => x"00001f59",
         16431 => x"00001f59",
         16432 => x"00001f59",
         16433 => x"00001f59",
         16434 => x"00001f59",
         16435 => x"00001f59",
         16436 => x"00001f59",
         16437 => x"00001f59",
         16438 => x"00001f59",
         16439 => x"00001f59",
         16440 => x"00001f59",
         16441 => x"00001f59",
         16442 => x"00001f59",
         16443 => x"00001f59",
         16444 => x"00001f59",
         16445 => x"00001f59",
         16446 => x"00001f59",
         16447 => x"00001f59",
         16448 => x"00001f59",
         16449 => x"00001f59",
         16450 => x"00001f59",
         16451 => x"00001f59",
         16452 => x"00001f59",
         16453 => x"00001f59",
         16454 => x"00001f59",
         16455 => x"00001f59",
         16456 => x"00001f59",
         16457 => x"00001f59",
         16458 => x"00001f59",
         16459 => x"00001f59",
         16460 => x"00001f59",
         16461 => x"000021ab",
         16462 => x"00002170",
         16463 => x"00001f59",
         16464 => x"00001f59",
         16465 => x"00001f59",
         16466 => x"00001f59",
         16467 => x"00001f59",
         16468 => x"00001f59",
         16469 => x"00001f59",
         16470 => x"00001f59",
         16471 => x"00002163",
         16472 => x"00002158",
         16473 => x"00001f59",
         16474 => x"00002141",
         16475 => x"00001f59",
         16476 => x"00002151",
         16477 => x"00002147",
         16478 => x"0000213a",
         16479 => x"00003222",
         16480 => x"0000323a",
         16481 => x"00003246",
         16482 => x"00003252",
         16483 => x"0000325e",
         16484 => x"0000322e",
         16485 => x"00003b97",
         16486 => x"00003a85",
         16487 => x"00003901",
         16488 => x"0000364f",
         16489 => x"00003a21",
         16490 => x"000034de",
         16491 => x"0000379b",
         16492 => x"00003674",
         16493 => x"000039cb",
         16494 => x"000036a3",
         16495 => x"00003712",
         16496 => x"0000392a",
         16497 => x"000034de",
         16498 => x"00003901",
         16499 => x"0000380b",
         16500 => x"0000379b",
         16501 => x"000034de",
         16502 => x"000034de",
         16503 => x"00003712",
         16504 => x"000036a3",
         16505 => x"00003674",
         16506 => x"0000364f",
         16507 => x"0000467c",
         16508 => x"00004695",
         16509 => x"000046ba",
         16510 => x"000046db",
         16511 => x"0000463c",
         16512 => x"00004700",
         16513 => x"00004655",
         16514 => x"000047a5",
         16515 => x"00004762",
         16516 => x"00004762",
         16517 => x"00004762",
         16518 => x"00004762",
         16519 => x"00004762",
         16520 => x"00004762",
         16521 => x"0000473b",
         16522 => x"00004762",
         16523 => x"00004762",
         16524 => x"00004762",
         16525 => x"00004762",
         16526 => x"00004762",
         16527 => x"00004762",
         16528 => x"00004762",
         16529 => x"00004762",
         16530 => x"00004762",
         16531 => x"00004762",
         16532 => x"00004762",
         16533 => x"00004762",
         16534 => x"00004762",
         16535 => x"00004762",
         16536 => x"00004762",
         16537 => x"00004762",
         16538 => x"00004762",
         16539 => x"00004762",
         16540 => x"00004762",
         16541 => x"00004762",
         16542 => x"00004762",
         16543 => x"00004762",
         16544 => x"0000487a",
         16545 => x"00004868",
         16546 => x"00004855",
         16547 => x"00004842",
         16548 => x"0000476c",
         16549 => x"00004830",
         16550 => x"0000481d",
         16551 => x"00004785",
         16552 => x"00004762",
         16553 => x"00004785",
         16554 => x"0000480d",
         16555 => x"0000488a",
         16556 => x"000047b6",
         16557 => x"00004794",
         16558 => x"000047fb",
         16559 => x"000047e9",
         16560 => x"000047d7",
         16561 => x"000047c8",
         16562 => x"00004762",
         16563 => x"0000476c",
         16564 => x"00005408",
         16565 => x"00005577",
         16566 => x"00005549",
         16567 => x"000054a0",
         16568 => x"0000547d",
         16569 => x"0000545c",
         16570 => x"00005432",
         16571 => x"00005602",
         16572 => x"00005289",
         16573 => x"000055dc",
         16574 => x"000057cb",
         16575 => x"00005289",
         16576 => x"00005289",
         16577 => x"00005289",
         16578 => x"00005289",
         16579 => x"00005289",
         16580 => x"00005289",
         16581 => x"000055a5",
         16582 => x"000057b3",
         16583 => x"0000566a",
         16584 => x"00005289",
         16585 => x"00005289",
         16586 => x"00005289",
         16587 => x"00005289",
         16588 => x"00005289",
         16589 => x"00005289",
         16590 => x"00005289",
         16591 => x"00005289",
         16592 => x"00005289",
         16593 => x"00005289",
         16594 => x"00005289",
         16595 => x"00005289",
         16596 => x"00005289",
         16597 => x"00005289",
         16598 => x"00005289",
         16599 => x"00005289",
         16600 => x"00005289",
         16601 => x"00005289",
         16602 => x"00005289",
         16603 => x"00005527",
         16604 => x"00005289",
         16605 => x"00005289",
         16606 => x"00005289",
         16607 => x"000054ca",
         16608 => x"000053d9",
         16609 => x"0000537b",
         16610 => x"00005289",
         16611 => x"00005289",
         16612 => x"00005289",
         16613 => x"00005289",
         16614 => x"00005360",
         16615 => x"00005289",
         16616 => x"00005343",
         16617 => x"000059ac",
         16618 => x"00005921",
         16619 => x"00005921",
         16620 => x"00005921",
         16621 => x"00005921",
         16622 => x"00005921",
         16623 => x"00005921",
         16624 => x"000058fc",
         16625 => x"00005921",
         16626 => x"00005921",
         16627 => x"00005921",
         16628 => x"00005921",
         16629 => x"00005921",
         16630 => x"00005921",
         16631 => x"00005921",
         16632 => x"00005921",
         16633 => x"00005921",
         16634 => x"00005921",
         16635 => x"00005921",
         16636 => x"00005921",
         16637 => x"00005921",
         16638 => x"00005921",
         16639 => x"00005921",
         16640 => x"00005921",
         16641 => x"00005921",
         16642 => x"00005921",
         16643 => x"00005921",
         16644 => x"00005921",
         16645 => x"00005921",
         16646 => x"00005921",
         16647 => x"000059be",
         16648 => x"00005a06",
         16649 => x"000059f3",
         16650 => x"000059e0",
         16651 => x"000059ce",
         16652 => x"00005a91",
         16653 => x"00005a7e",
         16654 => x"00005a6e",
         16655 => x"00005921",
         16656 => x"00005a5e",
         16657 => x"00005a4e",
         16658 => x"00005a3c",
         16659 => x"00005a2a",
         16660 => x"00005a18",
         16661 => x"00005989",
         16662 => x"00005978",
         16663 => x"00005967",
         16664 => x"00005950",
         16665 => x"00005921",
         16666 => x"0000599a",
         16667 => x"0000637b",
         16668 => x"000061d7",
         16669 => x"000061d7",
         16670 => x"000061d7",
         16671 => x"000061d7",
         16672 => x"000061d7",
         16673 => x"000061d7",
         16674 => x"000061d7",
         16675 => x"000061d7",
         16676 => x"000061d7",
         16677 => x"000061d7",
         16678 => x"000061d7",
         16679 => x"000061d7",
         16680 => x"000061d7",
         16681 => x"00005ef9",
         16682 => x"000061d7",
         16683 => x"000061d7",
         16684 => x"000061d7",
         16685 => x"000061d7",
         16686 => x"000061d7",
         16687 => x"000061d7",
         16688 => x"000063c5",
         16689 => x"000061d7",
         16690 => x"000061d7",
         16691 => x"00006350",
         16692 => x"000061d7",
         16693 => x"00006367",
         16694 => x"00005ed8",
         16695 => x"00006339",
         16696 => x"0000dee5",
         16697 => x"0000ded2",
         16698 => x"0000dec6",
         16699 => x"0000debb",
         16700 => x"0000deb0",
         16701 => x"0000dea5",
         16702 => x"0000de9a",
         16703 => x"0000de8e",
         16704 => x"0000de80",
         16705 => x"00000e01",
         16706 => x"00000bfd",
         16707 => x"00000bfd",
         16708 => x"00000f49",
         16709 => x"00000bfd",
         16710 => x"00000bfd",
         16711 => x"00000bfd",
         16712 => x"00000bfd",
         16713 => x"00000bfd",
         16714 => x"00000bfd",
         16715 => x"00000bfd",
         16716 => x"00000dfd",
         16717 => x"00000bfd",
         16718 => x"00000f7f",
         16719 => x"00000f0d",
         16720 => x"00000bfd",
         16721 => x"00000bfd",
         16722 => x"00000bfd",
         16723 => x"00000bfd",
         16724 => x"00000bfd",
         16725 => x"00000bfd",
         16726 => x"00000bfd",
         16727 => x"00000bfd",
         16728 => x"00000bfd",
         16729 => x"00000bfd",
         16730 => x"00000bfd",
         16731 => x"00000bfd",
         16732 => x"00000bfd",
         16733 => x"00000bfd",
         16734 => x"00000bfd",
         16735 => x"00000bfd",
         16736 => x"00000bfd",
         16737 => x"00000bfd",
         16738 => x"00000bfd",
         16739 => x"00000bfd",
         16740 => x"00000bfd",
         16741 => x"00000bfd",
         16742 => x"00000bfd",
         16743 => x"00000bfd",
         16744 => x"00000bfd",
         16745 => x"00000bfd",
         16746 => x"00000bfd",
         16747 => x"00000bfd",
         16748 => x"00000bfd",
         16749 => x"00000bfd",
         16750 => x"00000bfd",
         16751 => x"00000bfd",
         16752 => x"00000bfd",
         16753 => x"00000bfd",
         16754 => x"00000bfd",
         16755 => x"00000bfd",
         16756 => x"00000f1d",
         16757 => x"00000bfd",
         16758 => x"00000bfd",
         16759 => x"00000bfd",
         16760 => x"00000bfd",
         16761 => x"00000e17",
         16762 => x"00000bfd",
         16763 => x"00000bfd",
         16764 => x"00000bfd",
         16765 => x"00000bfd",
         16766 => x"00000bfd",
         16767 => x"00000bfd",
         16768 => x"00000bfd",
         16769 => x"00000bfd",
         16770 => x"00000bfd",
         16771 => x"00000bfd",
         16772 => x"00000e2b",
         16773 => x"00000ee1",
         16774 => x"00000eb8",
         16775 => x"00000eb8",
         16776 => x"00000eb8",
         16777 => x"00000bfd",
         16778 => x"00000ee1",
         16779 => x"00000bfd",
         16780 => x"00000bfd",
         16781 => x"00000eff",
         16782 => x"00000bfd",
         16783 => x"00000bfd",
         16784 => x"00000c16",
         16785 => x"00000e0f",
         16786 => x"00000bfd",
         16787 => x"00000bfd",
         16788 => x"00000f58",
         16789 => x"00000bfd",
         16790 => x"00000c18",
         16791 => x"00000bfd",
         16792 => x"00000bfd",
         16793 => x"00000e17",
         16794 => x"64696e69",
         16795 => x"74000000",
         16796 => x"64696f63",
         16797 => x"746c0000",
         16798 => x"66696e69",
         16799 => x"74000000",
         16800 => x"666c6f61",
         16801 => x"64000000",
         16802 => x"66657865",
         16803 => x"63000000",
         16804 => x"6d636c65",
         16805 => x"61720000",
         16806 => x"6d636f70",
         16807 => x"79000000",
         16808 => x"6d646966",
         16809 => x"66000000",
         16810 => x"6d64756d",
         16811 => x"70000000",
         16812 => x"6d656200",
         16813 => x"6d656800",
         16814 => x"6d657700",
         16815 => x"68696400",
         16816 => x"68696500",
         16817 => x"68666400",
         16818 => x"68666500",
         16819 => x"63616c6c",
         16820 => x"00000000",
         16821 => x"6a6d7000",
         16822 => x"72657374",
         16823 => x"61727400",
         16824 => x"72657365",
         16825 => x"74000000",
         16826 => x"696e666f",
         16827 => x"00000000",
         16828 => x"74657374",
         16829 => x"00000000",
         16830 => x"636c7300",
         16831 => x"7a383000",
         16832 => x"74626173",
         16833 => x"69630000",
         16834 => x"6d626173",
         16835 => x"69630000",
         16836 => x"6b696c6f",
         16837 => x"00000000",
         16838 => x"65640000",
         16839 => x"556e6b6e",
         16840 => x"6f776e20",
         16841 => x"6572726f",
         16842 => x"722e0000",
         16843 => x"50617261",
         16844 => x"6d657465",
         16845 => x"72732069",
         16846 => x"6e636f72",
         16847 => x"72656374",
         16848 => x"2e000000",
         16849 => x"546f6f20",
         16850 => x"6d616e79",
         16851 => x"206f7065",
         16852 => x"6e206669",
         16853 => x"6c65732e",
         16854 => x"00000000",
         16855 => x"496e7375",
         16856 => x"66666963",
         16857 => x"69656e74",
         16858 => x"206d656d",
         16859 => x"6f72792e",
         16860 => x"00000000",
         16861 => x"46696c65",
         16862 => x"20697320",
         16863 => x"6c6f636b",
         16864 => x"65642e00",
         16865 => x"54696d65",
         16866 => x"6f75742c",
         16867 => x"206f7065",
         16868 => x"72617469",
         16869 => x"6f6e2063",
         16870 => x"616e6365",
         16871 => x"6c6c6564",
         16872 => x"2e000000",
         16873 => x"466f726d",
         16874 => x"61742061",
         16875 => x"626f7274",
         16876 => x"65642e00",
         16877 => x"4e6f2063",
         16878 => x"6f6d7061",
         16879 => x"7469626c",
         16880 => x"65206669",
         16881 => x"6c657379",
         16882 => x"7374656d",
         16883 => x"20666f75",
         16884 => x"6e64206f",
         16885 => x"6e206469",
         16886 => x"736b2e00",
         16887 => x"4469736b",
         16888 => x"206e6f74",
         16889 => x"20656e61",
         16890 => x"626c6564",
         16891 => x"2e000000",
         16892 => x"44726976",
         16893 => x"65206e75",
         16894 => x"6d626572",
         16895 => x"20697320",
         16896 => x"696e7661",
         16897 => x"6c69642e",
         16898 => x"00000000",
         16899 => x"53442069",
         16900 => x"73207772",
         16901 => x"69746520",
         16902 => x"70726f74",
         16903 => x"65637465",
         16904 => x"642e0000",
         16905 => x"46696c65",
         16906 => x"2068616e",
         16907 => x"646c6520",
         16908 => x"696e7661",
         16909 => x"6c69642e",
         16910 => x"00000000",
         16911 => x"46696c65",
         16912 => x"20616c72",
         16913 => x"65616479",
         16914 => x"20657869",
         16915 => x"7374732e",
         16916 => x"00000000",
         16917 => x"41636365",
         16918 => x"73732064",
         16919 => x"656e6965",
         16920 => x"642e0000",
         16921 => x"496e7661",
         16922 => x"6c696420",
         16923 => x"66696c65",
         16924 => x"6e616d65",
         16925 => x"2e000000",
         16926 => x"4e6f2070",
         16927 => x"61746820",
         16928 => x"666f756e",
         16929 => x"642e0000",
         16930 => x"4e6f2066",
         16931 => x"696c6520",
         16932 => x"666f756e",
         16933 => x"642e0000",
         16934 => x"4469736b",
         16935 => x"206e6f74",
         16936 => x"20726561",
         16937 => x"64792e00",
         16938 => x"496e7465",
         16939 => x"726e616c",
         16940 => x"20657272",
         16941 => x"6f722e00",
         16942 => x"4469736b",
         16943 => x"20457272",
         16944 => x"6f720000",
         16945 => x"53756363",
         16946 => x"6573732e",
         16947 => x"00000000",
         16948 => x"0a256c75",
         16949 => x"20627974",
         16950 => x"65732025",
         16951 => x"73206174",
         16952 => x"20256c75",
         16953 => x"20627974",
         16954 => x"65732f73",
         16955 => x"65632e0a",
         16956 => x"00000000",
         16957 => x"72656164",
         16958 => x"00000000",
         16959 => x"2530386c",
         16960 => x"58000000",
         16961 => x"3a202000",
         16962 => x"25303258",
         16963 => x"00000000",
         16964 => x"207c0000",
         16965 => x"7c000000",
         16966 => x"20200000",
         16967 => x"25303458",
         16968 => x"00000000",
         16969 => x"20202020",
         16970 => x"20202020",
         16971 => x"00000000",
         16972 => x"7a4f5300",
         16973 => x"2a2a2025",
         16974 => x"73202800",
         16975 => x"31372f30",
         16976 => x"342f3230",
         16977 => x"32310000",
         16978 => x"76312e32",
         16979 => x"00000000",
         16980 => x"205a5055",
         16981 => x"2c207265",
         16982 => x"76202530",
         16983 => x"32782920",
         16984 => x"25732025",
         16985 => x"73202a2a",
         16986 => x"0a0a0000",
         16987 => x"4f533a00",
         16988 => x"20202020",
         16989 => x"42617365",
         16990 => x"20416464",
         16991 => x"72657373",
         16992 => x"20202020",
         16993 => x"20202020",
         16994 => x"20202020",
         16995 => x"203d2025",
         16996 => x"30386c78",
         16997 => x"0a000000",
         16998 => x"20202020",
         16999 => x"41707020",
         17000 => x"41646472",
         17001 => x"65737320",
         17002 => x"20202020",
         17003 => x"20202020",
         17004 => x"20202020",
         17005 => x"203d2025",
         17006 => x"30386c78",
         17007 => x"0a000000",
         17008 => x"5a505520",
         17009 => x"496e7465",
         17010 => x"72727570",
         17011 => x"74204861",
         17012 => x"6e646c65",
         17013 => x"72000000",
         17014 => x"55415254",
         17015 => x"31205458",
         17016 => x"20696e74",
         17017 => x"65727275",
         17018 => x"70740000",
         17019 => x"55415254",
         17020 => x"31205258",
         17021 => x"20696e74",
         17022 => x"65727275",
         17023 => x"70740000",
         17024 => x"55415254",
         17025 => x"30205458",
         17026 => x"20696e74",
         17027 => x"65727275",
         17028 => x"70740000",
         17029 => x"55415254",
         17030 => x"30205258",
         17031 => x"20696e74",
         17032 => x"65727275",
         17033 => x"70740000",
         17034 => x"494f4354",
         17035 => x"4c205752",
         17036 => x"20696e74",
         17037 => x"65727275",
         17038 => x"70740000",
         17039 => x"494f4354",
         17040 => x"4c205244",
         17041 => x"20696e74",
         17042 => x"65727275",
         17043 => x"70740000",
         17044 => x"50533220",
         17045 => x"696e7465",
         17046 => x"72727570",
         17047 => x"74000000",
         17048 => x"54696d65",
         17049 => x"7220696e",
         17050 => x"74657272",
         17051 => x"75707400",
         17052 => x"53657474",
         17053 => x"696e6720",
         17054 => x"75702074",
         17055 => x"696d6572",
         17056 => x"2e2e2e00",
         17057 => x"456e6162",
         17058 => x"6c696e67",
         17059 => x"2074696d",
         17060 => x"65722e2e",
         17061 => x"2e000000",
         17062 => x"6175746f",
         17063 => x"65786563",
         17064 => x"2e626174",
         17065 => x"00000000",
         17066 => x"7a4f535f",
         17067 => x"7a70752e",
         17068 => x"68737400",
         17069 => x"4661696c",
         17070 => x"65642074",
         17071 => x"6f20696e",
         17072 => x"69746961",
         17073 => x"6c697365",
         17074 => x"20736420",
         17075 => x"63617264",
         17076 => x"20302c20",
         17077 => x"706c6561",
         17078 => x"73652069",
         17079 => x"6e697420",
         17080 => x"6d616e75",
         17081 => x"616c6c79",
         17082 => x"2e000000",
         17083 => x"2a200000",
         17084 => x"25643a5c",
         17085 => x"25730000",
         17086 => x"303a0000",
         17087 => x"42616420",
         17088 => x"636f6d6d",
         17089 => x"616e642e",
         17090 => x"00000000",
         17091 => x"5a505500",
         17092 => x"62696e00",
         17093 => x"25643a5c",
         17094 => x"25735c25",
         17095 => x"732e2573",
         17096 => x"00000000",
         17097 => x"436f6c64",
         17098 => x"20726562",
         17099 => x"6f6f7469",
         17100 => x"6e672e2e",
         17101 => x"2e000000",
         17102 => x"52657374",
         17103 => x"61727469",
         17104 => x"6e672061",
         17105 => x"70706c69",
         17106 => x"63617469",
         17107 => x"6f6e2e2e",
         17108 => x"2e000000",
         17109 => x"43616c6c",
         17110 => x"696e6720",
         17111 => x"636f6465",
         17112 => x"20402025",
         17113 => x"30386c78",
         17114 => x"202e2e2e",
         17115 => x"0a000000",
         17116 => x"43616c6c",
         17117 => x"20726574",
         17118 => x"75726e65",
         17119 => x"6420636f",
         17120 => x"64652028",
         17121 => x"2564292e",
         17122 => x"0a000000",
         17123 => x"45786563",
         17124 => x"7574696e",
         17125 => x"6720636f",
         17126 => x"64652040",
         17127 => x"20253038",
         17128 => x"6c78202e",
         17129 => x"2e2e0a00",
         17130 => x"2530386c",
         17131 => x"58202530",
         17132 => x"386c582d",
         17133 => x"00000000",
         17134 => x"2530386c",
         17135 => x"58202530",
         17136 => x"34582d00",
         17137 => x"436f6d70",
         17138 => x"6172696e",
         17139 => x"672e2e2e",
         17140 => x"00000000",
         17141 => x"2530386c",
         17142 => x"78282530",
         17143 => x"3878292d",
         17144 => x"3e253038",
         17145 => x"6c782825",
         17146 => x"30387829",
         17147 => x"0a000000",
         17148 => x"436f7079",
         17149 => x"696e672e",
         17150 => x"2e2e0000",
         17151 => x"2530386c",
         17152 => x"58202530",
         17153 => x"32582d00",
         17154 => x"436c6561",
         17155 => x"72696e67",
         17156 => x"2e2e2e2e",
         17157 => x"00000000",
         17158 => x"44756d70",
         17159 => x"204d656d",
         17160 => x"6f727900",
         17161 => x"0a436f6d",
         17162 => x"706c6574",
         17163 => x"652e0000",
         17164 => x"25643a5c",
         17165 => x"25735c25",
         17166 => x"73000000",
         17167 => x"4d656d6f",
         17168 => x"72792065",
         17169 => x"78686175",
         17170 => x"73746564",
         17171 => x"2c206361",
         17172 => x"6e6e6f74",
         17173 => x"2070726f",
         17174 => x"63657373",
         17175 => x"20636f6d",
         17176 => x"6d616e64",
         17177 => x"2e000000",
         17178 => x"3f3f3f00",
         17179 => x"25642f25",
         17180 => x"642f2564",
         17181 => x"2025643a",
         17182 => x"25643a25",
         17183 => x"642e2564",
         17184 => x"25640a00",
         17185 => x"536f4320",
         17186 => x"436f6e66",
         17187 => x"69677572",
         17188 => x"6174696f",
         17189 => x"6e000000",
         17190 => x"3a0a4465",
         17191 => x"76696365",
         17192 => x"7320696d",
         17193 => x"706c656d",
         17194 => x"656e7465",
         17195 => x"643a0000",
         17196 => x"41646472",
         17197 => x"65737365",
         17198 => x"733a0000",
         17199 => x"20202020",
         17200 => x"43505520",
         17201 => x"52657365",
         17202 => x"74205665",
         17203 => x"63746f72",
         17204 => x"20416464",
         17205 => x"72657373",
         17206 => x"203d2025",
         17207 => x"3038580a",
         17208 => x"00000000",
         17209 => x"20202020",
         17210 => x"43505520",
         17211 => x"4d656d6f",
         17212 => x"72792053",
         17213 => x"74617274",
         17214 => x"20416464",
         17215 => x"72657373",
         17216 => x"203d2025",
         17217 => x"3038580a",
         17218 => x"00000000",
         17219 => x"20202020",
         17220 => x"53746163",
         17221 => x"6b205374",
         17222 => x"61727420",
         17223 => x"41646472",
         17224 => x"65737320",
         17225 => x"20202020",
         17226 => x"203d2025",
         17227 => x"3038580a",
         17228 => x"00000000",
         17229 => x"4d697363",
         17230 => x"3a000000",
         17231 => x"20202020",
         17232 => x"5a505520",
         17233 => x"49642020",
         17234 => x"20202020",
         17235 => x"20202020",
         17236 => x"20202020",
         17237 => x"20202020",
         17238 => x"203d2025",
         17239 => x"3034580a",
         17240 => x"00000000",
         17241 => x"20202020",
         17242 => x"53797374",
         17243 => x"656d2043",
         17244 => x"6c6f636b",
         17245 => x"20467265",
         17246 => x"71202020",
         17247 => x"20202020",
         17248 => x"203d2025",
         17249 => x"642e2530",
         17250 => x"34644d48",
         17251 => x"7a0a0000",
         17252 => x"20202020",
         17253 => x"57697368",
         17254 => x"626f6e65",
         17255 => x"20534452",
         17256 => x"414d2043",
         17257 => x"6c6f636b",
         17258 => x"20467265",
         17259 => x"713d2025",
         17260 => x"642e2530",
         17261 => x"34644d48",
         17262 => x"7a0a0000",
         17263 => x"20202020",
         17264 => x"53445241",
         17265 => x"4d20436c",
         17266 => x"6f636b20",
         17267 => x"46726571",
         17268 => x"20202020",
         17269 => x"20202020",
         17270 => x"203d2025",
         17271 => x"642e2530",
         17272 => x"34644d48",
         17273 => x"7a0a0000",
         17274 => x"20202020",
         17275 => x"53504900",
         17276 => x"20202020",
         17277 => x"50533200",
         17278 => x"20202020",
         17279 => x"494f4354",
         17280 => x"4c000000",
         17281 => x"20202020",
         17282 => x"57422049",
         17283 => x"32430000",
         17284 => x"20202020",
         17285 => x"57495348",
         17286 => x"424f4e45",
         17287 => x"20425553",
         17288 => x"00000000",
         17289 => x"20202020",
         17290 => x"494e5452",
         17291 => x"20435452",
         17292 => x"4c202843",
         17293 => x"68616e6e",
         17294 => x"656c733d",
         17295 => x"25303264",
         17296 => x"292e0a00",
         17297 => x"20202020",
         17298 => x"54494d45",
         17299 => x"52312020",
         17300 => x"20202854",
         17301 => x"696d6572",
         17302 => x"7320203d",
         17303 => x"25303264",
         17304 => x"292e0a00",
         17305 => x"20202020",
         17306 => x"53442043",
         17307 => x"41524420",
         17308 => x"20202844",
         17309 => x"65766963",
         17310 => x"6573203d",
         17311 => x"25303264",
         17312 => x"292e0a00",
         17313 => x"20202020",
         17314 => x"52414d20",
         17315 => x"20202020",
         17316 => x"20202825",
         17317 => x"3038583a",
         17318 => x"25303858",
         17319 => x"292e0a00",
         17320 => x"20202020",
         17321 => x"4252414d",
         17322 => x"20202020",
         17323 => x"20202825",
         17324 => x"3038583a",
         17325 => x"25303858",
         17326 => x"292e0a00",
         17327 => x"20202020",
         17328 => x"494e534e",
         17329 => x"20425241",
         17330 => x"4d202825",
         17331 => x"3038583a",
         17332 => x"25303858",
         17333 => x"292e0a00",
         17334 => x"20202020",
         17335 => x"53445241",
         17336 => x"4d202020",
         17337 => x"20202825",
         17338 => x"3038583a",
         17339 => x"25303858",
         17340 => x"292e0a00",
         17341 => x"20202020",
         17342 => x"57422053",
         17343 => x"4452414d",
         17344 => x"20202825",
         17345 => x"3038583a",
         17346 => x"25303858",
         17347 => x"292e0a00",
         17348 => x"20286672",
         17349 => x"6f6d2053",
         17350 => x"6f432063",
         17351 => x"6f6e6669",
         17352 => x"67290000",
         17353 => x"556e6b6e",
         17354 => x"6f776e00",
         17355 => x"45564f6d",
         17356 => x"00000000",
         17357 => x"536d616c",
         17358 => x"6c000000",
         17359 => x"4d656469",
         17360 => x"756d0000",
         17361 => x"466c6578",
         17362 => x"00000000",
         17363 => x"45564f00",
         17364 => x"0000f0ac",
         17365 => x"01000000",
         17366 => x"00000002",
         17367 => x"0000f0a8",
         17368 => x"01000000",
         17369 => x"00000003",
         17370 => x"0000f0a4",
         17371 => x"01000000",
         17372 => x"00000004",
         17373 => x"0000f0a0",
         17374 => x"01000000",
         17375 => x"00000005",
         17376 => x"0000f09c",
         17377 => x"01000000",
         17378 => x"00000006",
         17379 => x"0000f098",
         17380 => x"01000000",
         17381 => x"00000007",
         17382 => x"0000f094",
         17383 => x"01000000",
         17384 => x"00000001",
         17385 => x"0000f090",
         17386 => x"01000000",
         17387 => x"00000008",
         17388 => x"0000f08c",
         17389 => x"01000000",
         17390 => x"0000000b",
         17391 => x"0000f088",
         17392 => x"01000000",
         17393 => x"00000009",
         17394 => x"0000f084",
         17395 => x"01000000",
         17396 => x"0000000a",
         17397 => x"0000f080",
         17398 => x"04000000",
         17399 => x"0000000d",
         17400 => x"0000f07c",
         17401 => x"04000000",
         17402 => x"0000000c",
         17403 => x"0000f078",
         17404 => x"04000000",
         17405 => x"0000000e",
         17406 => x"0000f074",
         17407 => x"03000000",
         17408 => x"0000000f",
         17409 => x"0000f070",
         17410 => x"04000000",
         17411 => x"0000000f",
         17412 => x"0000f06c",
         17413 => x"04000000",
         17414 => x"00000010",
         17415 => x"0000f068",
         17416 => x"04000000",
         17417 => x"00000011",
         17418 => x"0000f064",
         17419 => x"03000000",
         17420 => x"00000012",
         17421 => x"0000f060",
         17422 => x"03000000",
         17423 => x"00000013",
         17424 => x"0000f05c",
         17425 => x"03000000",
         17426 => x"00000014",
         17427 => x"0000f058",
         17428 => x"03000000",
         17429 => x"00000015",
         17430 => x"1b5b4400",
         17431 => x"1b5b4300",
         17432 => x"1b5b4200",
         17433 => x"1b5b4100",
         17434 => x"1b5b367e",
         17435 => x"1b5b357e",
         17436 => x"1b5b347e",
         17437 => x"1b304600",
         17438 => x"1b5b337e",
         17439 => x"1b5b327e",
         17440 => x"1b5b317e",
         17441 => x"10000000",
         17442 => x"0e000000",
         17443 => x"0d000000",
         17444 => x"0b000000",
         17445 => x"08000000",
         17446 => x"06000000",
         17447 => x"05000000",
         17448 => x"04000000",
         17449 => x"03000000",
         17450 => x"02000000",
         17451 => x"01000000",
         17452 => x"43616e6e",
         17453 => x"6f74206f",
         17454 => x"70656e2f",
         17455 => x"63726561",
         17456 => x"74652068",
         17457 => x"6973746f",
         17458 => x"72792066",
         17459 => x"696c652c",
         17460 => x"20646973",
         17461 => x"61626c69",
         17462 => x"6e672e00",
         17463 => x"68697374",
         17464 => x"6f727900",
         17465 => x"68697374",
         17466 => x"00000000",
         17467 => x"21000000",
         17468 => x"2530366c",
         17469 => x"75202025",
         17470 => x"730a0000",
         17471 => x"4661696c",
         17472 => x"65642074",
         17473 => x"6f207265",
         17474 => x"73657420",
         17475 => x"74686520",
         17476 => x"68697374",
         17477 => x"6f727920",
         17478 => x"66696c65",
         17479 => x"20746f20",
         17480 => x"454f462e",
         17481 => x"00000000",
         17482 => x"3e25730a",
         17483 => x"00000000",
         17484 => x"1b5b317e",
         17485 => x"00000000",
         17486 => x"1b5b4100",
         17487 => x"1b5b4200",
         17488 => x"1b5b4300",
         17489 => x"1b5b4400",
         17490 => x"1b5b3130",
         17491 => x"7e000000",
         17492 => x"1b5b3131",
         17493 => x"7e000000",
         17494 => x"1b5b3132",
         17495 => x"7e000000",
         17496 => x"1b5b3133",
         17497 => x"7e000000",
         17498 => x"1b5b3134",
         17499 => x"7e000000",
         17500 => x"1b5b3135",
         17501 => x"7e000000",
         17502 => x"1b5b3137",
         17503 => x"7e000000",
         17504 => x"1b5b3138",
         17505 => x"7e000000",
         17506 => x"1b5b3139",
         17507 => x"7e000000",
         17508 => x"1b5b3230",
         17509 => x"7e000000",
         17510 => x"1b5b327e",
         17511 => x"00000000",
         17512 => x"1b5b337e",
         17513 => x"00000000",
         17514 => x"1b5b4600",
         17515 => x"1b5b357e",
         17516 => x"00000000",
         17517 => x"1b5b367e",
         17518 => x"00000000",
         17519 => x"583a2564",
         17520 => x"2c25642c",
         17521 => x"25642c25",
         17522 => x"642c2564",
         17523 => x"2c25643a",
         17524 => x"25303278",
         17525 => x"00000000",
         17526 => x"443a2564",
         17527 => x"2d25642d",
         17528 => x"25643a25",
         17529 => x"633a2564",
         17530 => x"2c25642c",
         17531 => x"25643a00",
         17532 => x"25642c00",
         17533 => x"4b3a2564",
         17534 => x"3a000000",
         17535 => x"25303278",
         17536 => x"2c000000",
         17537 => x"25635b25",
         17538 => x"643b2564",
         17539 => x"52000000",
         17540 => x"5265706f",
         17541 => x"72742043",
         17542 => x"7572736f",
         17543 => x"723a0000",
         17544 => x"55703a25",
         17545 => x"30327820",
         17546 => x"25303278",
         17547 => x"00000000",
         17548 => x"44773a25",
         17549 => x"30327820",
         17550 => x"25303278",
         17551 => x"00000000",
         17552 => x"48643a25",
         17553 => x"30327820",
         17554 => x"00000000",
         17555 => x"4e6f2074",
         17556 => x"65737420",
         17557 => x"64656669",
         17558 => x"6e65642e",
         17559 => x"00000000",
         17560 => x"53440000",
         17561 => x"222a3a3c",
         17562 => x"3e3f7c7f",
         17563 => x"00000000",
         17564 => x"2b2c3b3d",
         17565 => x"5b5d0000",
         17566 => x"46415400",
         17567 => x"46415433",
         17568 => x"32000000",
         17569 => x"ebfe904d",
         17570 => x"53444f53",
         17571 => x"352e3000",
         17572 => x"4e4f204e",
         17573 => x"414d4520",
         17574 => x"20202046",
         17575 => x"41542020",
         17576 => x"20202000",
         17577 => x"4e4f204e",
         17578 => x"414d4520",
         17579 => x"20202046",
         17580 => x"41543332",
         17581 => x"20202000",
         17582 => x"0000f260",
         17583 => x"00000000",
         17584 => x"00000000",
         17585 => x"00000000",
         17586 => x"01030507",
         17587 => x"090e1012",
         17588 => x"1416181c",
         17589 => x"1e000000",
         17590 => x"809a4541",
         17591 => x"8e418f80",
         17592 => x"45454549",
         17593 => x"49498e8f",
         17594 => x"9092924f",
         17595 => x"994f5555",
         17596 => x"59999a9b",
         17597 => x"9c9d9e9f",
         17598 => x"41494f55",
         17599 => x"a5a5a6a7",
         17600 => x"a8a9aaab",
         17601 => x"acadaeaf",
         17602 => x"b0b1b2b3",
         17603 => x"b4b5b6b7",
         17604 => x"b8b9babb",
         17605 => x"bcbdbebf",
         17606 => x"c0c1c2c3",
         17607 => x"c4c5c6c7",
         17608 => x"c8c9cacb",
         17609 => x"cccdcecf",
         17610 => x"d0d1d2d3",
         17611 => x"d4d5d6d7",
         17612 => x"d8d9dadb",
         17613 => x"dcdddedf",
         17614 => x"e0e1e2e3",
         17615 => x"e4e5e6e7",
         17616 => x"e8e9eaeb",
         17617 => x"ecedeeef",
         17618 => x"f0f1f2f3",
         17619 => x"f4f5f6f7",
         17620 => x"f8f9fafb",
         17621 => x"fcfdfeff",
         17622 => x"2b2e2c3b",
         17623 => x"3d5b5d2f",
         17624 => x"5c222a3a",
         17625 => x"3c3e3f7c",
         17626 => x"7f000000",
         17627 => x"00010004",
         17628 => x"00100040",
         17629 => x"01000200",
         17630 => x"00000000",
         17631 => x"00010002",
         17632 => x"00040008",
         17633 => x"00100020",
         17634 => x"00000000",
         17635 => x"00c700fc",
         17636 => x"00e900e2",
         17637 => x"00e400e0",
         17638 => x"00e500e7",
         17639 => x"00ea00eb",
         17640 => x"00e800ef",
         17641 => x"00ee00ec",
         17642 => x"00c400c5",
         17643 => x"00c900e6",
         17644 => x"00c600f4",
         17645 => x"00f600f2",
         17646 => x"00fb00f9",
         17647 => x"00ff00d6",
         17648 => x"00dc00a2",
         17649 => x"00a300a5",
         17650 => x"20a70192",
         17651 => x"00e100ed",
         17652 => x"00f300fa",
         17653 => x"00f100d1",
         17654 => x"00aa00ba",
         17655 => x"00bf2310",
         17656 => x"00ac00bd",
         17657 => x"00bc00a1",
         17658 => x"00ab00bb",
         17659 => x"25912592",
         17660 => x"25932502",
         17661 => x"25242561",
         17662 => x"25622556",
         17663 => x"25552563",
         17664 => x"25512557",
         17665 => x"255d255c",
         17666 => x"255b2510",
         17667 => x"25142534",
         17668 => x"252c251c",
         17669 => x"2500253c",
         17670 => x"255e255f",
         17671 => x"255a2554",
         17672 => x"25692566",
         17673 => x"25602550",
         17674 => x"256c2567",
         17675 => x"25682564",
         17676 => x"25652559",
         17677 => x"25582552",
         17678 => x"2553256b",
         17679 => x"256a2518",
         17680 => x"250c2588",
         17681 => x"2584258c",
         17682 => x"25902580",
         17683 => x"03b100df",
         17684 => x"039303c0",
         17685 => x"03a303c3",
         17686 => x"00b503c4",
         17687 => x"03a60398",
         17688 => x"03a903b4",
         17689 => x"221e03c6",
         17690 => x"03b52229",
         17691 => x"226100b1",
         17692 => x"22652264",
         17693 => x"23202321",
         17694 => x"00f72248",
         17695 => x"00b02219",
         17696 => x"00b7221a",
         17697 => x"207f00b2",
         17698 => x"25a000a0",
         17699 => x"0061031a",
         17700 => x"00e00317",
         17701 => x"00f80307",
         17702 => x"00ff0001",
         17703 => x"01780100",
         17704 => x"01300132",
         17705 => x"01060139",
         17706 => x"0110014a",
         17707 => x"012e0179",
         17708 => x"01060180",
         17709 => x"004d0243",
         17710 => x"01810182",
         17711 => x"01820184",
         17712 => x"01840186",
         17713 => x"01870187",
         17714 => x"0189018a",
         17715 => x"018b018b",
         17716 => x"018d018e",
         17717 => x"018f0190",
         17718 => x"01910191",
         17719 => x"01930194",
         17720 => x"01f60196",
         17721 => x"01970198",
         17722 => x"0198023d",
         17723 => x"019b019c",
         17724 => x"019d0220",
         17725 => x"019f01a0",
         17726 => x"01a001a2",
         17727 => x"01a201a4",
         17728 => x"01a401a6",
         17729 => x"01a701a7",
         17730 => x"01a901aa",
         17731 => x"01ab01ac",
         17732 => x"01ac01ae",
         17733 => x"01af01af",
         17734 => x"01b101b2",
         17735 => x"01b301b3",
         17736 => x"01b501b5",
         17737 => x"01b701b8",
         17738 => x"01b801ba",
         17739 => x"01bb01bc",
         17740 => x"01bc01be",
         17741 => x"01f701c0",
         17742 => x"01c101c2",
         17743 => x"01c301c4",
         17744 => x"01c501c4",
         17745 => x"01c701c8",
         17746 => x"01c701ca",
         17747 => x"01cb01ca",
         17748 => x"01cd0110",
         17749 => x"01dd0001",
         17750 => x"018e01de",
         17751 => x"011201f3",
         17752 => x"000301f1",
         17753 => x"01f401f4",
         17754 => x"01f80128",
         17755 => x"02220112",
         17756 => x"023a0009",
         17757 => x"2c65023b",
         17758 => x"023b023d",
         17759 => x"2c66023f",
         17760 => x"02400241",
         17761 => x"02410246",
         17762 => x"010a0253",
         17763 => x"00400181",
         17764 => x"01860255",
         17765 => x"0189018a",
         17766 => x"0258018f",
         17767 => x"025a0190",
         17768 => x"025c025d",
         17769 => x"025e025f",
         17770 => x"01930261",
         17771 => x"02620194",
         17772 => x"02640265",
         17773 => x"02660267",
         17774 => x"01970196",
         17775 => x"026a2c62",
         17776 => x"026c026d",
         17777 => x"026e019c",
         17778 => x"02700271",
         17779 => x"019d0273",
         17780 => x"0274019f",
         17781 => x"02760277",
         17782 => x"02780279",
         17783 => x"027a027b",
         17784 => x"027c2c64",
         17785 => x"027e027f",
         17786 => x"01a60281",
         17787 => x"028201a9",
         17788 => x"02840285",
         17789 => x"02860287",
         17790 => x"01ae0244",
         17791 => x"01b101b2",
         17792 => x"0245028d",
         17793 => x"028e028f",
         17794 => x"02900291",
         17795 => x"01b7037b",
         17796 => x"000303fd",
         17797 => x"03fe03ff",
         17798 => x"03ac0004",
         17799 => x"03860388",
         17800 => x"0389038a",
         17801 => x"03b10311",
         17802 => x"03c20002",
         17803 => x"03a303a3",
         17804 => x"03c40308",
         17805 => x"03cc0003",
         17806 => x"038c038e",
         17807 => x"038f03d8",
         17808 => x"011803f2",
         17809 => x"000a03f9",
         17810 => x"03f303f4",
         17811 => x"03f503f6",
         17812 => x"03f703f7",
         17813 => x"03f903fa",
         17814 => x"03fa0430",
         17815 => x"03200450",
         17816 => x"07100460",
         17817 => x"0122048a",
         17818 => x"013604c1",
         17819 => x"010e04cf",
         17820 => x"000104c0",
         17821 => x"04d00144",
         17822 => x"05610426",
         17823 => x"00000000",
         17824 => x"1d7d0001",
         17825 => x"2c631e00",
         17826 => x"01961ea0",
         17827 => x"015a1f00",
         17828 => x"06081f10",
         17829 => x"06061f20",
         17830 => x"06081f30",
         17831 => x"06081f40",
         17832 => x"06061f51",
         17833 => x"00071f59",
         17834 => x"1f521f5b",
         17835 => x"1f541f5d",
         17836 => x"1f561f5f",
         17837 => x"1f600608",
         17838 => x"1f70000e",
         17839 => x"1fba1fbb",
         17840 => x"1fc81fc9",
         17841 => x"1fca1fcb",
         17842 => x"1fda1fdb",
         17843 => x"1ff81ff9",
         17844 => x"1fea1feb",
         17845 => x"1ffa1ffb",
         17846 => x"1f800608",
         17847 => x"1f900608",
         17848 => x"1fa00608",
         17849 => x"1fb00004",
         17850 => x"1fb81fb9",
         17851 => x"1fb21fbc",
         17852 => x"1fcc0001",
         17853 => x"1fc31fd0",
         17854 => x"06021fe0",
         17855 => x"06021fe5",
         17856 => x"00011fec",
         17857 => x"1ff30001",
         17858 => x"1ffc214e",
         17859 => x"00012132",
         17860 => x"21700210",
         17861 => x"21840001",
         17862 => x"218324d0",
         17863 => x"051a2c30",
         17864 => x"042f2c60",
         17865 => x"01022c67",
         17866 => x"01062c75",
         17867 => x"01022c80",
         17868 => x"01642d00",
         17869 => x"0826ff41",
         17870 => x"031a0000",
         17871 => x"00000000",
         17872 => x"0000e668",
         17873 => x"01020100",
         17874 => x"00000000",
         17875 => x"00000000",
         17876 => x"0000e670",
         17877 => x"01040100",
         17878 => x"00000000",
         17879 => x"00000000",
         17880 => x"0000e678",
         17881 => x"01140300",
         17882 => x"00000000",
         17883 => x"00000000",
         17884 => x"0000e680",
         17885 => x"012b0300",
         17886 => x"00000000",
         17887 => x"00000000",
         17888 => x"0000e688",
         17889 => x"01300300",
         17890 => x"00000000",
         17891 => x"00000000",
         17892 => x"0000e690",
         17893 => x"013c0400",
         17894 => x"00000000",
         17895 => x"00000000",
         17896 => x"0000e698",
         17897 => x"013d0400",
         17898 => x"00000000",
         17899 => x"00000000",
         17900 => x"0000e6a0",
         17901 => x"013f0400",
         17902 => x"00000000",
         17903 => x"00000000",
         17904 => x"0000e6a8",
         17905 => x"01400400",
         17906 => x"00000000",
         17907 => x"00000000",
         17908 => x"0000e6b0",
         17909 => x"01410400",
         17910 => x"00000000",
         17911 => x"00000000",
         17912 => x"0000e6b4",
         17913 => x"01420400",
         17914 => x"00000000",
         17915 => x"00000000",
         17916 => x"0000e6b8",
         17917 => x"01430400",
         17918 => x"00000000",
         17919 => x"00000000",
         17920 => x"0000e6bc",
         17921 => x"01500500",
         17922 => x"00000000",
         17923 => x"00000000",
         17924 => x"0000e6c0",
         17925 => x"01510500",
         17926 => x"00000000",
         17927 => x"00000000",
         17928 => x"0000e6c4",
         17929 => x"01540500",
         17930 => x"00000000",
         17931 => x"00000000",
         17932 => x"0000e6c8",
         17933 => x"01550500",
         17934 => x"00000000",
         17935 => x"00000000",
         17936 => x"0000e6cc",
         17937 => x"01790700",
         17938 => x"00000000",
         17939 => x"00000000",
         17940 => x"0000e6d4",
         17941 => x"01780700",
         17942 => x"00000000",
         17943 => x"00000000",
         17944 => x"0000e6d8",
         17945 => x"01820800",
         17946 => x"00000000",
         17947 => x"00000000",
         17948 => x"0000e6e0",
         17949 => x"01830800",
         17950 => x"00000000",
         17951 => x"00000000",
         17952 => x"0000e6e8",
         17953 => x"01850800",
         17954 => x"00000000",
         17955 => x"00000000",
         17956 => x"0000e6f0",
         17957 => x"01870800",
         17958 => x"00000000",
         17959 => x"00000000",
         17960 => x"0000e6f8",
         17961 => x"01880800",
         17962 => x"00000000",
         17963 => x"00000000",
         17964 => x"0000e6fc",
         17965 => x"01890800",
         17966 => x"00000000",
         17967 => x"00000000",
         17968 => x"0000e700",
         17969 => x"018c0900",
         17970 => x"00000000",
         17971 => x"00000000",
         17972 => x"0000e708",
         17973 => x"018d0900",
         17974 => x"00000000",
         17975 => x"00000000",
         17976 => x"0000e710",
         17977 => x"018e0900",
         17978 => x"00000000",
         17979 => x"00000000",
         17980 => x"0000e718",
         17981 => x"018f0900",
         17982 => x"00000000",
         17983 => x"00000000",
         17984 => x"00000000",
         17985 => x"00000000",
         17986 => x"00007fff",
         17987 => x"00000000",
         17988 => x"00007fff",
         17989 => x"00010000",
         17990 => x"00007fff",
         17991 => x"00010000",
         17992 => x"00810000",
         17993 => x"01000000",
         17994 => x"017fffff",
         17995 => x"00000000",
         17996 => x"00000000",
         17997 => x"00007800",
         17998 => x"00000000",
         17999 => x"05f5e100",
         18000 => x"05f5e100",
         18001 => x"05f5e100",
         18002 => x"00000000",
         18003 => x"01010101",
         18004 => x"01010101",
         18005 => x"01011001",
         18006 => x"01000000",
         18007 => x"00000000",
         18008 => x"00000000",
         18009 => x"00000000",
         18010 => x"00000000",
         18011 => x"00000000",
         18012 => x"00000000",
         18013 => x"00000000",
         18014 => x"00000000",
         18015 => x"00000000",
         18016 => x"00000000",
         18017 => x"00000000",
         18018 => x"00000000",
         18019 => x"00000000",
         18020 => x"00000000",
         18021 => x"00000000",
         18022 => x"00000000",
         18023 => x"00000000",
         18024 => x"00000000",
         18025 => x"00000000",
         18026 => x"00000000",
         18027 => x"00000000",
         18028 => x"00000000",
         18029 => x"00000000",
         18030 => x"00000000",
         18031 => x"0000f0dc",
         18032 => x"01000000",
         18033 => x"0000f0e4",
         18034 => x"01000000",
         18035 => x"0000f0ec",
         18036 => x"02000000",
         18037 => x"0001fd80",
         18038 => x"1bfc5ffd",
         18039 => x"f03b3a0d",
         18040 => x"797a405b",
         18041 => x"5df0f0f0",
         18042 => x"71727374",
         18043 => x"75767778",
         18044 => x"696a6b6c",
         18045 => x"6d6e6f70",
         18046 => x"61626364",
         18047 => x"65666768",
         18048 => x"31323334",
         18049 => x"35363738",
         18050 => x"5cf32d20",
         18051 => x"30392c2e",
         18052 => x"f67ff3f4",
         18053 => x"f1f23f2f",
         18054 => x"08f0f0f0",
         18055 => x"f0f0f0f0",
         18056 => x"80818283",
         18057 => x"84f0f0f0",
         18058 => x"1bfc58fd",
         18059 => x"f03a3b0d",
         18060 => x"595a405b",
         18061 => x"5df0f0f0",
         18062 => x"51525354",
         18063 => x"55565758",
         18064 => x"494a4b4c",
         18065 => x"4d4e4f50",
         18066 => x"41424344",
         18067 => x"45464748",
         18068 => x"31323334",
         18069 => x"35363738",
         18070 => x"5cf32d20",
         18071 => x"30392c2e",
         18072 => x"f67ff3f4",
         18073 => x"f1f23f2f",
         18074 => x"08f0f0f0",
         18075 => x"f0f0f0f0",
         18076 => x"80818283",
         18077 => x"84f0f0f0",
         18078 => x"1bfc58fd",
         18079 => x"f02b2a0d",
         18080 => x"595a607b",
         18081 => x"7df0f0f0",
         18082 => x"51525354",
         18083 => x"55565758",
         18084 => x"494a4b4c",
         18085 => x"4d4e4f50",
         18086 => x"41424344",
         18087 => x"45464748",
         18088 => x"21222324",
         18089 => x"25262728",
         18090 => x"7c7e3d20",
         18091 => x"20293c3e",
         18092 => x"f7e2e0e1",
         18093 => x"f9f83f2f",
         18094 => x"fbf0f0f0",
         18095 => x"f0f0f0f0",
         18096 => x"85868788",
         18097 => x"89f0f0f0",
         18098 => x"1bfe1efa",
         18099 => x"f0f0f0f0",
         18100 => x"191a001b",
         18101 => x"1df0f0f0",
         18102 => x"11121314",
         18103 => x"15161718",
         18104 => x"090a0b0c",
         18105 => x"0d0e0f10",
         18106 => x"01020304",
         18107 => x"05060708",
         18108 => x"f0f0f0f0",
         18109 => x"f0f0f0f0",
         18110 => x"f01ef0f0",
         18111 => x"f01ff0f0",
         18112 => x"f0f0f0f0",
         18113 => x"f0f0f01c",
         18114 => x"f0f0f0f0",
         18115 => x"f0f0f0f0",
         18116 => x"80818283",
         18117 => x"84f0f0f0",
         18118 => x"bff0cfc9",
         18119 => x"f0b54dcd",
         18120 => x"3577d7b3",
         18121 => x"b7f0f0f0",
         18122 => x"7c704131",
         18123 => x"39a678dd",
         18124 => x"3d5d6c56",
         18125 => x"1d33d5b1",
         18126 => x"466ed948",
         18127 => x"74434c73",
         18128 => x"3f367e3b",
         18129 => x"7a1e5fa2",
         18130 => x"d39fd100",
         18131 => x"9da3d0b9",
         18132 => x"c6c5c2c1",
         18133 => x"c3c4bbbe",
         18134 => x"f0f0f0f0",
         18135 => x"f0f0f0f0",
         18136 => x"80818283",
         18137 => x"84f0f0f0",
         18138 => x"00000000",
         18139 => x"00000000",
         18140 => x"00000000",
         18141 => x"00000000",
         18142 => x"00000000",
         18143 => x"00000000",
         18144 => x"00000000",
         18145 => x"00000000",
         18146 => x"00000000",
         18147 => x"00000000",
         18148 => x"00000000",
         18149 => x"00000000",
         18150 => x"00000000",
         18151 => x"00000000",
         18152 => x"00000000",
         18153 => x"00000000",
         18154 => x"00000000",
         18155 => x"00000000",
         18156 => x"00000000",
         18157 => x"00000000",
         18158 => x"00000000",
         18159 => x"00000000",
         18160 => x"00000000",
         18161 => x"00000000",
         18162 => x"00000000",
         18163 => x"00010000",
         18164 => x"00000000",
         18165 => x"f8000000",
         18166 => x"0000f130",
         18167 => x"f3000000",
         18168 => x"0000f138",
         18169 => x"f4000000",
         18170 => x"0000f13c",
         18171 => x"f1000000",
         18172 => x"0000f140",
         18173 => x"f2000000",
         18174 => x"0000f144",
         18175 => x"80000000",
         18176 => x"0000f148",
         18177 => x"81000000",
         18178 => x"0000f150",
         18179 => x"82000000",
         18180 => x"0000f158",
         18181 => x"83000000",
         18182 => x"0000f160",
         18183 => x"84000000",
         18184 => x"0000f168",
         18185 => x"85000000",
         18186 => x"0000f170",
         18187 => x"86000000",
         18188 => x"0000f178",
         18189 => x"87000000",
         18190 => x"0000f180",
         18191 => x"88000000",
         18192 => x"0000f188",
         18193 => x"89000000",
         18194 => x"0000f190",
         18195 => x"f6000000",
         18196 => x"0000f198",
         18197 => x"7f000000",
         18198 => x"0000f1a0",
         18199 => x"f9000000",
         18200 => x"0000f1a8",
         18201 => x"e0000000",
         18202 => x"0000f1ac",
         18203 => x"e1000000",
         18204 => x"0000f1b4",
         18205 => x"71000000",
         18206 => x"00000000",
         18207 => x"00000000",
         18208 => x"00000000",
         18209 => x"00000000",
         18210 => x"00000000",
         18211 => x"00000000",
         18212 => x"00000000",
         18213 => x"00000000",
         18214 => x"00000000",
         18215 => x"00000000",
         18216 => x"00000000",
         18217 => x"00000000",
         18218 => x"00000000",
         18219 => x"00000000",
         18220 => x"00000000",
         18221 => x"00000000",
         18222 => x"00000000",
         18223 => x"00000000",
         18224 => x"00000000",
         18225 => x"00000000",
         18226 => x"00000000",
         18227 => x"00000000",
         18228 => x"00000000",
         18229 => x"00000000",
         18230 => x"00000000",
         18231 => x"00000000",
         18232 => x"00000000",
         18233 => x"00000000",
         18234 => x"00000000",
         18235 => x"00000000",
         18236 => x"00000000",
         18237 => x"00000000",
         18238 => x"00000000",
         18239 => x"00000000",
         18240 => x"00000000",
         18241 => x"00000000",
         18242 => x"00000000",
         18243 => x"00000000",
         18244 => x"00000000",
         18245 => x"00000000",
         18246 => x"00000000",
         18247 => x"00000000",
         18248 => x"00000000",
         18249 => x"00000000",
         18250 => x"00000000",
         18251 => x"00000000",
         18252 => x"00000000",
         18253 => x"00000000",
         18254 => x"00000000",
         18255 => x"00000000",
         18256 => x"00000000",
         18257 => x"00000000",
         18258 => x"00000000",
         18259 => x"00000000",
         18260 => x"00000000",
         18261 => x"00000000",
         18262 => x"00000000",
         18263 => x"00000000",
         18264 => x"00000000",
         18265 => x"00000000",
         18266 => x"00000000",
         18267 => x"00000000",
         18268 => x"00000000",
         18269 => x"00000000",
         18270 => x"00000000",
         18271 => x"00000000",
         18272 => x"00000000",
         18273 => x"00000000",
         18274 => x"00000000",
         18275 => x"00000000",
         18276 => x"00000000",
         18277 => x"00000000",
         18278 => x"00000000",
         18279 => x"00000000",
         18280 => x"00000000",
         18281 => x"00000000",
         18282 => x"00000000",
         18283 => x"00000000",
         18284 => x"00000000",
         18285 => x"00000000",
         18286 => x"00000000",
         18287 => x"00000000",
         18288 => x"00000000",
         18289 => x"00000000",
         18290 => x"00000000",
         18291 => x"00000000",
         18292 => x"00000000",
         18293 => x"00000000",
         18294 => x"00000000",
         18295 => x"00000000",
         18296 => x"00000000",
         18297 => x"00000000",
         18298 => x"00000000",
         18299 => x"00000000",
         18300 => x"00000000",
         18301 => x"00000000",
         18302 => x"00000000",
         18303 => x"00000000",
         18304 => x"00000000",
         18305 => x"00000000",
         18306 => x"00000000",
         18307 => x"00000000",
         18308 => x"00000000",
         18309 => x"00000000",
         18310 => x"00000000",
         18311 => x"00000000",
         18312 => x"00000000",
         18313 => x"00000000",
         18314 => x"00000000",
         18315 => x"00000000",
         18316 => x"00000000",
         18317 => x"00000000",
         18318 => x"00000000",
         18319 => x"00000000",
         18320 => x"00000000",
         18321 => x"00000000",
         18322 => x"00000000",
         18323 => x"00000000",
         18324 => x"00000000",
         18325 => x"00000000",
         18326 => x"00000000",
         18327 => x"00000000",
         18328 => x"00000000",
         18329 => x"00000000",
         18330 => x"00000000",
         18331 => x"00000000",
         18332 => x"00000000",
         18333 => x"00000000",
         18334 => x"00000000",
         18335 => x"00000000",
         18336 => x"00000000",
         18337 => x"00000000",
         18338 => x"00000000",
         18339 => x"00000000",
         18340 => x"00000000",
         18341 => x"00000000",
         18342 => x"00000000",
         18343 => x"00000000",
         18344 => x"00000000",
         18345 => x"00000000",
         18346 => x"00000000",
         18347 => x"00000000",
         18348 => x"00000000",
         18349 => x"00000000",
         18350 => x"00000000",
         18351 => x"00000000",
         18352 => x"00000000",
         18353 => x"00000000",
         18354 => x"00000000",
         18355 => x"00000000",
         18356 => x"00000000",
         18357 => x"00000000",
         18358 => x"00000000",
         18359 => x"00000000",
         18360 => x"00000000",
         18361 => x"00000000",
         18362 => x"00000000",
         18363 => x"00000000",
         18364 => x"00000000",
         18365 => x"00000000",
         18366 => x"00000000",
         18367 => x"00000000",
         18368 => x"00000000",
         18369 => x"00000000",
         18370 => x"00000000",
         18371 => x"00000000",
         18372 => x"00000000",
         18373 => x"00000000",
         18374 => x"00000000",
         18375 => x"00000000",
         18376 => x"00000000",
         18377 => x"00000000",
         18378 => x"00000000",
         18379 => x"00000000",
         18380 => x"00000000",
         18381 => x"00000000",
         18382 => x"00000000",
         18383 => x"00000000",
         18384 => x"00000000",
         18385 => x"00000000",
         18386 => x"00000000",
         18387 => x"00000000",
         18388 => x"00000000",
         18389 => x"00000000",
         18390 => x"00000000",
         18391 => x"00000000",
         18392 => x"00000000",
         18393 => x"00000000",
         18394 => x"00000000",
         18395 => x"00000000",
         18396 => x"00000000",
         18397 => x"00000000",
         18398 => x"00000000",
         18399 => x"00000000",
         18400 => x"00000000",
         18401 => x"00000000",
         18402 => x"00000000",
         18403 => x"00000000",
         18404 => x"00000000",
         18405 => x"00000000",
         18406 => x"00000000",
         18407 => x"00000000",
         18408 => x"00000000",
         18409 => x"00000000",
         18410 => x"00000000",
         18411 => x"00000000",
         18412 => x"00000000",
         18413 => x"00000000",
         18414 => x"00000000",
         18415 => x"00000000",
         18416 => x"00000000",
         18417 => x"00000000",
         18418 => x"00000000",
         18419 => x"00000000",
         18420 => x"00000000",
         18421 => x"00000000",
         18422 => x"00000000",
         18423 => x"00000000",
         18424 => x"00000000",
         18425 => x"00000000",
         18426 => x"00000000",
         18427 => x"00000000",
         18428 => x"00000000",
         18429 => x"00000000",
         18430 => x"00000000",
         18431 => x"00000000",
         18432 => x"00000000",
         18433 => x"00000000",
         18434 => x"00000000",
         18435 => x"00000000",
         18436 => x"00000000",
         18437 => x"00000000",
         18438 => x"00000000",
         18439 => x"00000000",
         18440 => x"00000000",
         18441 => x"00000000",
         18442 => x"00000000",
         18443 => x"00000000",
         18444 => x"00000000",
         18445 => x"00000000",
         18446 => x"00000000",
         18447 => x"00000000",
         18448 => x"00000000",
         18449 => x"00000000",
         18450 => x"00000000",
         18451 => x"00000000",
         18452 => x"00000000",
         18453 => x"00000000",
         18454 => x"00000000",
         18455 => x"00000000",
         18456 => x"00000000",
         18457 => x"00000000",
         18458 => x"00000000",
         18459 => x"00000000",
         18460 => x"00000000",
         18461 => x"00000000",
         18462 => x"00000000",
         18463 => x"00000000",
         18464 => x"00000000",
         18465 => x"00000000",
         18466 => x"00000000",
         18467 => x"00000000",
         18468 => x"00000000",
         18469 => x"00000000",
         18470 => x"00000000",
         18471 => x"00000000",
         18472 => x"00000000",
         18473 => x"00000000",
         18474 => x"00000000",
         18475 => x"00000000",
         18476 => x"00000000",
         18477 => x"00000000",
         18478 => x"00000000",
         18479 => x"00000000",
         18480 => x"00000000",
         18481 => x"00000000",
         18482 => x"00000000",
         18483 => x"00000000",
         18484 => x"00000000",
         18485 => x"00000000",
         18486 => x"00000000",
         18487 => x"00000000",
         18488 => x"00000000",
         18489 => x"00000000",
         18490 => x"00000000",
         18491 => x"00000000",
         18492 => x"00000000",
         18493 => x"00000000",
         18494 => x"00000000",
         18495 => x"00000000",
         18496 => x"00000000",
         18497 => x"00000000",
         18498 => x"00000000",
         18499 => x"00000000",
         18500 => x"00000000",
         18501 => x"00000000",
         18502 => x"00000000",
         18503 => x"00000000",
         18504 => x"00000000",
         18505 => x"00000000",
         18506 => x"00000000",
         18507 => x"00000000",
         18508 => x"00000000",
         18509 => x"00000000",
         18510 => x"00000000",
         18511 => x"00000000",
         18512 => x"00000000",
         18513 => x"00000000",
         18514 => x"00000000",
         18515 => x"00000000",
         18516 => x"00000000",
         18517 => x"00000000",
         18518 => x"00000000",
         18519 => x"00000000",
         18520 => x"00000000",
         18521 => x"00000000",
         18522 => x"00000000",
         18523 => x"00000000",
         18524 => x"00000000",
         18525 => x"00000000",
         18526 => x"00000000",
         18527 => x"00000000",
         18528 => x"00000000",
         18529 => x"00000000",
         18530 => x"00000000",
         18531 => x"00000000",
         18532 => x"00000000",
         18533 => x"00000000",
         18534 => x"00000000",
         18535 => x"00000000",
         18536 => x"00000000",
         18537 => x"00000000",
         18538 => x"00000000",
         18539 => x"00000000",
         18540 => x"00000000",
         18541 => x"00000000",
         18542 => x"00000000",
         18543 => x"00000000",
         18544 => x"00000000",
         18545 => x"00000000",
         18546 => x"00000000",
         18547 => x"00000000",
         18548 => x"00000000",
         18549 => x"00000000",
         18550 => x"00000000",
         18551 => x"00000000",
         18552 => x"00000000",
         18553 => x"00000000",
         18554 => x"00000000",
         18555 => x"00000000",
         18556 => x"00000000",
         18557 => x"00000000",
         18558 => x"00000000",
         18559 => x"00000000",
         18560 => x"00000000",
         18561 => x"00000000",
         18562 => x"00000000",
         18563 => x"00000000",
         18564 => x"00000000",
         18565 => x"00000000",
         18566 => x"00000000",
         18567 => x"00000000",
         18568 => x"00000000",
         18569 => x"00000000",
         18570 => x"00000000",
         18571 => x"00000000",
         18572 => x"00000000",
         18573 => x"00000000",
         18574 => x"00000000",
         18575 => x"00000000",
         18576 => x"00000000",
         18577 => x"00000000",
         18578 => x"00000000",
         18579 => x"00000000",
         18580 => x"00000000",
         18581 => x"00000000",
         18582 => x"00000000",
         18583 => x"00000000",
         18584 => x"00000000",
         18585 => x"00000000",
         18586 => x"00000000",
         18587 => x"00000000",
         18588 => x"00000000",
         18589 => x"00000000",
         18590 => x"00000000",
         18591 => x"00000000",
         18592 => x"00000000",
         18593 => x"00000000",
         18594 => x"00000000",
         18595 => x"00000000",
         18596 => x"00000000",
         18597 => x"00000000",
         18598 => x"00000000",
         18599 => x"00000000",
         18600 => x"00000000",
         18601 => x"00000000",
         18602 => x"00000000",
         18603 => x"00000000",
         18604 => x"00000000",
         18605 => x"00000000",
         18606 => x"00000000",
         18607 => x"00000000",
         18608 => x"00000000",
         18609 => x"00000000",
         18610 => x"00000000",
         18611 => x"00000000",
         18612 => x"00000000",
         18613 => x"00000000",
         18614 => x"00000000",
         18615 => x"00000000",
         18616 => x"00000000",
         18617 => x"00000000",
         18618 => x"00000000",
         18619 => x"00000000",
         18620 => x"00000000",
         18621 => x"00000000",
         18622 => x"00000000",
         18623 => x"00000000",
         18624 => x"00000000",
         18625 => x"00000000",
         18626 => x"00000000",
         18627 => x"00000000",
         18628 => x"00000000",
         18629 => x"00000000",
         18630 => x"00000000",
         18631 => x"00000000",
         18632 => x"00000000",
         18633 => x"00000000",
         18634 => x"00000000",
         18635 => x"00000000",
         18636 => x"00000000",
         18637 => x"00000000",
         18638 => x"00000000",
         18639 => x"00000000",
         18640 => x"00000000",
         18641 => x"00000000",
         18642 => x"00000000",
         18643 => x"00000000",
         18644 => x"00000000",
         18645 => x"00000000",
         18646 => x"00000000",
         18647 => x"00000000",
         18648 => x"00000000",
         18649 => x"00000000",
         18650 => x"00000000",
         18651 => x"00000000",
         18652 => x"00000000",
         18653 => x"00000000",
         18654 => x"00000000",
         18655 => x"00000000",
         18656 => x"00000000",
         18657 => x"00000000",
         18658 => x"00000000",
         18659 => x"00000000",
         18660 => x"00000000",
         18661 => x"00000000",
         18662 => x"00000000",
         18663 => x"00000000",
         18664 => x"00000000",
         18665 => x"00000000",
         18666 => x"00000000",
         18667 => x"00000000",
         18668 => x"00000000",
         18669 => x"00000000",
         18670 => x"00000000",
         18671 => x"00000000",
         18672 => x"00000000",
         18673 => x"00000000",
         18674 => x"00000000",
         18675 => x"00000000",
         18676 => x"00000000",
         18677 => x"00000000",
         18678 => x"00000000",
         18679 => x"00000000",
         18680 => x"00000000",
         18681 => x"00000000",
         18682 => x"00000000",
         18683 => x"00000000",
         18684 => x"00000000",
         18685 => x"00000000",
         18686 => x"00000000",
         18687 => x"00000000",
         18688 => x"00000000",
         18689 => x"00000000",
         18690 => x"00000000",
         18691 => x"00000000",
         18692 => x"00000000",
         18693 => x"00000000",
         18694 => x"00000000",
         18695 => x"00000000",
         18696 => x"00000000",
         18697 => x"00000000",
         18698 => x"00000000",
         18699 => x"00000000",
         18700 => x"00000000",
         18701 => x"00000000",
         18702 => x"00000000",
         18703 => x"00000000",
         18704 => x"00000000",
         18705 => x"00000000",
         18706 => x"00000000",
         18707 => x"00000000",
         18708 => x"00000000",
         18709 => x"00000000",
         18710 => x"00000000",
         18711 => x"00000000",
         18712 => x"00000000",
         18713 => x"00000000",
         18714 => x"00000000",
         18715 => x"00000000",
         18716 => x"00000000",
         18717 => x"00000000",
         18718 => x"00000000",
         18719 => x"00000000",
         18720 => x"00000000",
         18721 => x"00000000",
         18722 => x"00000000",
         18723 => x"00000000",
         18724 => x"00000000",
         18725 => x"00000000",
         18726 => x"00000000",
         18727 => x"00000000",
         18728 => x"00000000",
         18729 => x"00000000",
         18730 => x"00000000",
         18731 => x"00000000",
         18732 => x"00000000",
         18733 => x"00000000",
         18734 => x"00000000",
         18735 => x"00000000",
         18736 => x"00000000",
         18737 => x"00000000",
         18738 => x"00000000",
         18739 => x"00000000",
         18740 => x"00000000",
         18741 => x"00000000",
         18742 => x"00000000",
         18743 => x"00000000",
         18744 => x"00000000",
         18745 => x"00000000",
         18746 => x"00000000",
         18747 => x"00000000",
         18748 => x"00000000",
         18749 => x"00000000",
         18750 => x"00000000",
         18751 => x"00000000",
         18752 => x"00000000",
         18753 => x"00000000",
         18754 => x"00000000",
         18755 => x"00000000",
         18756 => x"00000000",
         18757 => x"00000000",
         18758 => x"00000000",
         18759 => x"00000000",
         18760 => x"00000000",
         18761 => x"00000000",
         18762 => x"00000000",
         18763 => x"00000000",
         18764 => x"00000000",
         18765 => x"00000000",
         18766 => x"00000000",
         18767 => x"00000000",
         18768 => x"00000000",
         18769 => x"00000000",
         18770 => x"00000000",
         18771 => x"00000000",
         18772 => x"00000000",
         18773 => x"00000000",
         18774 => x"00000000",
         18775 => x"00000000",
         18776 => x"00000000",
         18777 => x"00000000",
         18778 => x"00000000",
         18779 => x"00000000",
         18780 => x"00000000",
         18781 => x"00000000",
         18782 => x"00000000",
         18783 => x"00000000",
         18784 => x"00000000",
         18785 => x"00000000",
         18786 => x"00000000",
         18787 => x"00000000",
         18788 => x"00000000",
         18789 => x"00000000",
         18790 => x"00000000",
         18791 => x"00000000",
         18792 => x"00000000",
         18793 => x"00000000",
         18794 => x"00000000",
         18795 => x"00000000",
         18796 => x"00000000",
         18797 => x"00000000",
         18798 => x"00000000",
         18799 => x"00000000",
         18800 => x"00000000",
         18801 => x"00000000",
         18802 => x"00000000",
         18803 => x"00000000",
         18804 => x"00000000",
         18805 => x"00000000",
         18806 => x"00000000",
         18807 => x"00000000",
         18808 => x"00000000",
         18809 => x"00000000",
         18810 => x"00000000",
         18811 => x"00000000",
         18812 => x"00000000",
         18813 => x"00000000",
         18814 => x"00000000",
         18815 => x"00000000",
         18816 => x"00000000",
         18817 => x"00000000",
         18818 => x"00000000",
         18819 => x"00000000",
         18820 => x"00000000",
         18821 => x"00000000",
         18822 => x"00000000",
         18823 => x"00000000",
         18824 => x"00000000",
         18825 => x"00000000",
         18826 => x"00000000",
         18827 => x"00000000",
         18828 => x"00000000",
         18829 => x"00000000",
         18830 => x"00000000",
         18831 => x"00000000",
         18832 => x"00000000",
         18833 => x"00000000",
         18834 => x"00000000",
         18835 => x"00000000",
         18836 => x"00000000",
         18837 => x"00000000",
         18838 => x"00000000",
         18839 => x"00000000",
         18840 => x"00000000",
         18841 => x"00000000",
         18842 => x"00000000",
         18843 => x"00000000",
         18844 => x"00000000",
         18845 => x"00000000",
         18846 => x"00000000",
         18847 => x"00000000",
         18848 => x"00000000",
         18849 => x"00000000",
         18850 => x"00000000",
         18851 => x"00000000",
         18852 => x"00000000",
         18853 => x"00000000",
         18854 => x"00000000",
         18855 => x"00000000",
         18856 => x"00000000",
         18857 => x"00000000",
         18858 => x"00000000",
         18859 => x"00000000",
         18860 => x"00000000",
         18861 => x"00000000",
         18862 => x"00000000",
         18863 => x"00000000",
         18864 => x"00000000",
         18865 => x"00000000",
         18866 => x"00000000",
         18867 => x"00000000",
         18868 => x"00000000",
         18869 => x"00000000",
         18870 => x"00000000",
         18871 => x"00000000",
         18872 => x"00000000",
         18873 => x"00000000",
         18874 => x"00000000",
         18875 => x"00000000",
         18876 => x"00000000",
         18877 => x"00000000",
         18878 => x"00000000",
         18879 => x"00000000",
         18880 => x"00000000",
         18881 => x"00000000",
         18882 => x"00000000",
         18883 => x"00000000",
         18884 => x"00000000",
         18885 => x"00000000",
         18886 => x"00000000",
         18887 => x"00000000",
         18888 => x"00000000",
         18889 => x"00000000",
         18890 => x"00000000",
         18891 => x"00000000",
         18892 => x"00000000",
         18893 => x"00000000",
         18894 => x"00000000",
         18895 => x"00000000",
         18896 => x"00000000",
         18897 => x"00000000",
         18898 => x"00000000",
         18899 => x"00000000",
         18900 => x"00000000",
         18901 => x"00000000",
         18902 => x"00000000",
         18903 => x"00000000",
         18904 => x"00000000",
         18905 => x"00000000",
         18906 => x"00000000",
         18907 => x"00000000",
         18908 => x"00000000",
         18909 => x"00000000",
         18910 => x"00000000",
         18911 => x"00000000",
         18912 => x"00000000",
         18913 => x"00000000",
         18914 => x"00000000",
         18915 => x"00000000",
         18916 => x"00000000",
         18917 => x"00000000",
         18918 => x"00000000",
         18919 => x"00000000",
         18920 => x"00000000",
         18921 => x"00000000",
         18922 => x"00000000",
         18923 => x"00000000",
         18924 => x"00000000",
         18925 => x"00000000",
         18926 => x"00000000",
         18927 => x"00000000",
         18928 => x"00000000",
         18929 => x"00000000",
         18930 => x"00000000",
         18931 => x"00000000",
         18932 => x"00000000",
         18933 => x"00000000",
         18934 => x"00000000",
         18935 => x"00000000",
         18936 => x"00000000",
         18937 => x"00000000",
         18938 => x"00000000",
         18939 => x"00000000",
         18940 => x"00000000",
         18941 => x"00000000",
         18942 => x"00000000",
         18943 => x"00000000",
         18944 => x"00000000",
         18945 => x"00000000",
         18946 => x"00000000",
         18947 => x"00000000",
         18948 => x"00000000",
         18949 => x"00000000",
         18950 => x"00000000",
         18951 => x"00000000",
         18952 => x"00000000",
         18953 => x"00000000",
         18954 => x"00000000",
         18955 => x"00000000",
         18956 => x"00000000",
         18957 => x"00000000",
         18958 => x"00000000",
         18959 => x"00000000",
         18960 => x"00000000",
         18961 => x"00000000",
         18962 => x"00000000",
         18963 => x"00000000",
         18964 => x"00000000",
         18965 => x"00000000",
         18966 => x"00000000",
         18967 => x"00000000",
         18968 => x"00000000",
         18969 => x"00000000",
         18970 => x"00000000",
         18971 => x"00000000",
         18972 => x"00000000",
         18973 => x"00000000",
         18974 => x"00000000",
         18975 => x"00000000",
         18976 => x"00000000",
         18977 => x"00000000",
         18978 => x"00000000",
         18979 => x"00000000",
         18980 => x"00000000",
         18981 => x"00000000",
         18982 => x"00000000",
         18983 => x"00000000",
         18984 => x"00000000",
         18985 => x"00000000",
         18986 => x"00000000",
         18987 => x"00000000",
         18988 => x"00000000",
         18989 => x"00000000",
         18990 => x"00000000",
         18991 => x"00000000",
         18992 => x"00000000",
         18993 => x"00000000",
         18994 => x"00000000",
         18995 => x"00000000",
         18996 => x"00000000",
         18997 => x"00000000",
         18998 => x"00000000",
         18999 => x"00000000",
         19000 => x"00000000",
         19001 => x"00000000",
         19002 => x"00000000",
         19003 => x"00000000",
         19004 => x"00000000",
         19005 => x"00000000",
         19006 => x"00000000",
         19007 => x"00000000",
         19008 => x"00000000",
         19009 => x"00000000",
         19010 => x"00000000",
         19011 => x"00000000",
         19012 => x"00000000",
         19013 => x"00000000",
         19014 => x"00000000",
         19015 => x"00000000",
         19016 => x"00000000",
         19017 => x"00000000",
         19018 => x"00000000",
         19019 => x"00000000",
         19020 => x"00000000",
         19021 => x"00000000",
         19022 => x"00000000",
         19023 => x"00000000",
         19024 => x"00000000",
         19025 => x"00000000",
         19026 => x"00000000",
         19027 => x"00000000",
         19028 => x"00000000",
         19029 => x"00000000",
         19030 => x"00000000",
         19031 => x"00000000",
         19032 => x"00000000",
         19033 => x"00000000",
         19034 => x"00000000",
         19035 => x"00000000",
         19036 => x"00000000",
         19037 => x"00000000",
         19038 => x"00000000",
         19039 => x"00000000",
         19040 => x"00000000",
         19041 => x"00000000",
         19042 => x"00000000",
         19043 => x"00000000",
         19044 => x"00000000",
         19045 => x"00000000",
         19046 => x"00000000",
         19047 => x"00000000",
         19048 => x"00000000",
         19049 => x"00000000",
         19050 => x"00000000",
         19051 => x"00000000",
         19052 => x"00000000",
         19053 => x"00000000",
         19054 => x"00000000",
         19055 => x"00000000",
         19056 => x"00000000",
         19057 => x"00000000",
         19058 => x"00000000",
         19059 => x"00000000",
         19060 => x"00000000",
         19061 => x"00000000",
         19062 => x"00000000",
         19063 => x"00000000",
         19064 => x"00000000",
         19065 => x"00000000",
         19066 => x"00000000",
         19067 => x"00000000",
         19068 => x"00000000",
         19069 => x"00000000",
         19070 => x"00000000",
         19071 => x"00000000",
         19072 => x"00000000",
         19073 => x"00000000",
         19074 => x"00000000",
         19075 => x"00000000",
         19076 => x"00000000",
         19077 => x"00000000",
         19078 => x"00000000",
         19079 => x"00000000",
         19080 => x"00000000",
         19081 => x"00000000",
         19082 => x"00000000",
         19083 => x"00000000",
         19084 => x"00000000",
         19085 => x"00000000",
         19086 => x"00000000",
         19087 => x"00000000",
         19088 => x"00000000",
         19089 => x"00000000",
         19090 => x"00000000",
         19091 => x"00000000",
         19092 => x"00000000",
         19093 => x"00000000",
         19094 => x"00000000",
         19095 => x"00000000",
         19096 => x"00000000",
         19097 => x"00000000",
         19098 => x"00000000",
         19099 => x"00000000",
         19100 => x"00000000",
         19101 => x"00000000",
         19102 => x"00000000",
         19103 => x"00000000",
         19104 => x"00000000",
         19105 => x"00000000",
         19106 => x"00000000",
         19107 => x"00000000",
         19108 => x"00000000",
         19109 => x"00000000",
         19110 => x"00000000",
         19111 => x"00000000",
         19112 => x"00000000",
         19113 => x"00000000",
         19114 => x"00000000",
         19115 => x"00000000",
         19116 => x"00000000",
         19117 => x"00000000",
         19118 => x"00000000",
         19119 => x"00000000",
         19120 => x"00000000",
         19121 => x"00000000",
         19122 => x"00000000",
         19123 => x"00000000",
         19124 => x"00000000",
         19125 => x"00000000",
         19126 => x"00000000",
         19127 => x"00000000",
         19128 => x"00000000",
         19129 => x"00000000",
         19130 => x"00000000",
         19131 => x"00000000",
         19132 => x"00000000",
         19133 => x"00000000",
         19134 => x"00000000",
         19135 => x"00000000",
         19136 => x"00000000",
         19137 => x"00000000",
         19138 => x"00000000",
         19139 => x"00000000",
         19140 => x"00000000",
         19141 => x"00000000",
         19142 => x"00000000",
         19143 => x"00000000",
         19144 => x"00000000",
         19145 => x"00000000",
         19146 => x"00000000",
         19147 => x"00000000",
         19148 => x"00000000",
         19149 => x"00000000",
         19150 => x"00000000",
         19151 => x"00000000",
         19152 => x"00000000",
         19153 => x"00000000",
         19154 => x"00000000",
         19155 => x"00000000",
         19156 => x"00000000",
         19157 => x"00000000",
         19158 => x"00000000",
         19159 => x"00000000",
         19160 => x"00000000",
         19161 => x"00000000",
         19162 => x"00000000",
         19163 => x"00000000",
         19164 => x"00000000",
         19165 => x"00000000",
         19166 => x"00000000",
         19167 => x"00000000",
         19168 => x"00000000",
         19169 => x"00000000",
         19170 => x"00000000",
         19171 => x"00000000",
         19172 => x"00000000",
         19173 => x"00000000",
         19174 => x"00000000",
         19175 => x"00000000",
         19176 => x"00000000",
         19177 => x"00000000",
         19178 => x"00000000",
         19179 => x"00000000",
         19180 => x"00000000",
         19181 => x"00000000",
         19182 => x"00000000",
         19183 => x"00000000",
         19184 => x"00000000",
         19185 => x"00000000",
         19186 => x"00000000",
         19187 => x"00000000",
         19188 => x"00000000",
         19189 => x"00000000",
         19190 => x"00000000",
         19191 => x"00000000",
         19192 => x"00000000",
         19193 => x"00000000",
         19194 => x"00000000",
         19195 => x"00000000",
         19196 => x"00000000",
         19197 => x"00000000",
         19198 => x"00000000",
         19199 => x"00000000",
         19200 => x"00000000",
         19201 => x"00000000",
         19202 => x"00000000",
         19203 => x"00000000",
         19204 => x"00000000",
         19205 => x"00000000",
         19206 => x"00000000",
         19207 => x"00000000",
         19208 => x"00000000",
         19209 => x"00000000",
         19210 => x"00000000",
         19211 => x"00000000",
         19212 => x"00000000",
         19213 => x"00000000",
         19214 => x"00000000",
         19215 => x"00000000",
         19216 => x"00000000",
         19217 => x"00000000",
         19218 => x"00000000",
         19219 => x"00000000",
         19220 => x"00000000",
         19221 => x"00000000",
         19222 => x"00000000",
         19223 => x"00000000",
         19224 => x"00000000",
         19225 => x"00000000",
         19226 => x"00000000",
         19227 => x"00000000",
         19228 => x"00000000",
         19229 => x"00000000",
         19230 => x"00000000",
         19231 => x"00000000",
         19232 => x"00000000",
         19233 => x"00000000",
         19234 => x"00000000",
         19235 => x"00000000",
         19236 => x"00000000",
         19237 => x"00000000",
         19238 => x"00000000",
         19239 => x"00000000",
         19240 => x"00000000",
         19241 => x"00000000",
         19242 => x"00000000",
         19243 => x"00000000",
         19244 => x"00000000",
         19245 => x"00000000",
         19246 => x"00000000",
         19247 => x"00000000",
         19248 => x"00000000",
         19249 => x"00000000",
         19250 => x"00000000",
         19251 => x"00000000",
         19252 => x"00000000",
         19253 => x"00000000",
         19254 => x"00000000",
         19255 => x"00000000",
         19256 => x"00000000",
         19257 => x"00000000",
         19258 => x"00000000",
         19259 => x"00000000",
         19260 => x"00000000",
         19261 => x"00000000",
         19262 => x"00000000",
         19263 => x"00000000",
         19264 => x"00000000",
         19265 => x"00000000",
         19266 => x"00000000",
         19267 => x"00000000",
         19268 => x"00000000",
         19269 => x"00000000",
         19270 => x"00000000",
         19271 => x"00000000",
         19272 => x"00000000",
         19273 => x"00000000",
         19274 => x"00000000",
         19275 => x"00000000",
         19276 => x"00000000",
         19277 => x"00000000",
         19278 => x"00000000",
         19279 => x"00000000",
         19280 => x"00000000",
         19281 => x"00000000",
         19282 => x"00000000",
         19283 => x"00000000",
         19284 => x"00000000",
         19285 => x"00000000",
         19286 => x"00000000",
         19287 => x"00000000",
         19288 => x"00000000",
         19289 => x"00000000",
         19290 => x"00000000",
         19291 => x"00000000",
         19292 => x"00000000",
         19293 => x"00000000",
         19294 => x"00000000",
         19295 => x"00000000",
         19296 => x"00000000",
         19297 => x"00000000",
         19298 => x"00000000",
         19299 => x"00000000",
         19300 => x"00000000",
         19301 => x"00000000",
         19302 => x"00000000",
         19303 => x"00000000",
         19304 => x"00000000",
         19305 => x"00000000",
         19306 => x"00000000",
         19307 => x"00000000",
         19308 => x"00000000",
         19309 => x"00000000",
         19310 => x"00000000",
         19311 => x"00000000",
         19312 => x"00000000",
         19313 => x"00000000",
         19314 => x"00000000",
         19315 => x"00000000",
         19316 => x"00000000",
         19317 => x"00000000",
         19318 => x"00000000",
         19319 => x"00000000",
         19320 => x"00000000",
         19321 => x"00000000",
         19322 => x"00000000",
         19323 => x"00000000",
         19324 => x"00000000",
         19325 => x"00000000",
         19326 => x"00000000",
         19327 => x"00000000",
         19328 => x"00000000",
         19329 => x"00000000",
         19330 => x"00000000",
         19331 => x"00000000",
         19332 => x"00000000",
         19333 => x"00000000",
         19334 => x"00000000",
         19335 => x"00000000",
         19336 => x"00000000",
         19337 => x"00000000",
         19338 => x"00000000",
         19339 => x"00000000",
         19340 => x"00000000",
         19341 => x"00000000",
         19342 => x"00000000",
         19343 => x"00000000",
         19344 => x"00000000",
         19345 => x"00000000",
         19346 => x"00000000",
         19347 => x"00000000",
         19348 => x"00000000",
         19349 => x"00000000",
         19350 => x"00000000",
         19351 => x"00000000",
         19352 => x"00000000",
         19353 => x"00000000",
         19354 => x"00000000",
         19355 => x"00000000",
         19356 => x"00000000",
         19357 => x"00000000",
         19358 => x"00000000",
         19359 => x"00000000",
         19360 => x"00000000",
         19361 => x"00000000",
         19362 => x"00000000",
         19363 => x"00000000",
         19364 => x"00000000",
         19365 => x"00000000",
         19366 => x"00000000",
         19367 => x"00000000",
         19368 => x"00000000",
         19369 => x"00000000",
         19370 => x"00000000",
         19371 => x"00000000",
         19372 => x"00000000",
         19373 => x"00000000",
         19374 => x"00000000",
         19375 => x"00000000",
         19376 => x"00000000",
         19377 => x"00000000",
         19378 => x"00000000",
         19379 => x"00000000",
         19380 => x"00000000",
         19381 => x"00000000",
         19382 => x"00000000",
         19383 => x"00000000",
         19384 => x"00000000",
         19385 => x"00000000",
         19386 => x"00000000",
         19387 => x"00000000",
         19388 => x"00000000",
         19389 => x"00000000",
         19390 => x"00000000",
         19391 => x"00000000",
         19392 => x"00000000",
         19393 => x"00000000",
         19394 => x"00000000",
         19395 => x"00000000",
         19396 => x"00000000",
         19397 => x"00000000",
         19398 => x"00000000",
         19399 => x"00000000",
         19400 => x"00000000",
         19401 => x"00000000",
         19402 => x"00000000",
         19403 => x"00000000",
         19404 => x"00000000",
         19405 => x"00000000",
         19406 => x"00000000",
         19407 => x"00000000",
         19408 => x"00000000",
         19409 => x"00000000",
         19410 => x"00000000",
         19411 => x"00000000",
         19412 => x"00000000",
         19413 => x"00000000",
         19414 => x"00000000",
         19415 => x"00000000",
         19416 => x"00000000",
         19417 => x"00000000",
         19418 => x"00000000",
         19419 => x"00000000",
         19420 => x"00000000",
         19421 => x"00000000",
         19422 => x"00000000",
         19423 => x"00000000",
         19424 => x"00000000",
         19425 => x"00000000",
         19426 => x"00000000",
         19427 => x"00000000",
         19428 => x"00000000",
         19429 => x"00000000",
         19430 => x"00000000",
         19431 => x"00000000",
         19432 => x"00000000",
         19433 => x"00000000",
         19434 => x"00000000",
         19435 => x"00000000",
         19436 => x"00000000",
         19437 => x"00000000",
         19438 => x"00000000",
         19439 => x"00000000",
         19440 => x"00000000",
         19441 => x"00000000",
         19442 => x"00000000",
         19443 => x"00000000",
         19444 => x"00000000",
         19445 => x"00000000",
         19446 => x"00000000",
         19447 => x"00000000",
         19448 => x"00000000",
         19449 => x"00000000",
         19450 => x"00000000",
         19451 => x"00000000",
         19452 => x"00000000",
         19453 => x"00000000",
         19454 => x"00000000",
         19455 => x"00000000",
         19456 => x"00000000",
         19457 => x"00000000",
         19458 => x"00000000",
         19459 => x"00000000",
         19460 => x"00000000",
         19461 => x"00000000",
         19462 => x"00000000",
         19463 => x"00000000",
         19464 => x"00000000",
         19465 => x"00000000",
         19466 => x"00000000",
         19467 => x"00000000",
         19468 => x"00000000",
         19469 => x"00000000",
         19470 => x"00000000",
         19471 => x"00000000",
         19472 => x"00000000",
         19473 => x"00000000",
         19474 => x"00000000",
         19475 => x"00000000",
         19476 => x"00000000",
         19477 => x"00000000",
         19478 => x"00000000",
         19479 => x"00000000",
         19480 => x"00000000",
         19481 => x"00000000",
         19482 => x"00000000",
         19483 => x"00000000",
         19484 => x"00000000",
         19485 => x"00000000",
         19486 => x"00000000",
         19487 => x"00000000",
         19488 => x"00000000",
         19489 => x"00000000",
         19490 => x"00000000",
         19491 => x"00000000",
         19492 => x"00000000",
         19493 => x"00000000",
         19494 => x"00000000",
         19495 => x"00000000",
         19496 => x"00000000",
         19497 => x"00000000",
         19498 => x"00000000",
         19499 => x"00000000",
         19500 => x"00000000",
         19501 => x"00000000",
         19502 => x"00000000",
         19503 => x"00000000",
         19504 => x"00000000",
         19505 => x"00000000",
         19506 => x"00000000",
         19507 => x"00000000",
         19508 => x"00000000",
         19509 => x"00000000",
         19510 => x"00000000",
         19511 => x"00000000",
         19512 => x"00000000",
         19513 => x"00000000",
         19514 => x"00000000",
         19515 => x"00000000",
         19516 => x"00000000",
         19517 => x"00000000",
         19518 => x"00000000",
         19519 => x"00000000",
         19520 => x"00000000",
         19521 => x"00000000",
         19522 => x"00000000",
         19523 => x"00000000",
         19524 => x"00000000",
         19525 => x"00000000",
         19526 => x"00000000",
         19527 => x"00000000",
         19528 => x"00000000",
         19529 => x"00000000",
         19530 => x"00000000",
         19531 => x"00000000",
         19532 => x"00000000",
         19533 => x"00000000",
         19534 => x"00000000",
         19535 => x"00000000",
         19536 => x"00000000",
         19537 => x"00000000",
         19538 => x"00000000",
         19539 => x"00000000",
         19540 => x"00000000",
         19541 => x"00000000",
         19542 => x"00000000",
         19543 => x"00000000",
         19544 => x"00000000",
         19545 => x"00000000",
         19546 => x"00000000",
         19547 => x"00000000",
         19548 => x"00000000",
         19549 => x"00000000",
         19550 => x"00000000",
         19551 => x"00000000",
         19552 => x"00000000",
         19553 => x"00000000",
         19554 => x"00000000",
         19555 => x"00000000",
         19556 => x"00000000",
         19557 => x"00000000",
         19558 => x"00000000",
         19559 => x"00000000",
         19560 => x"00000000",
         19561 => x"00000000",
         19562 => x"00000000",
         19563 => x"00000000",
         19564 => x"00000000",
         19565 => x"00000000",
         19566 => x"00000000",
         19567 => x"00000000",
         19568 => x"00000000",
         19569 => x"00000000",
         19570 => x"00000000",
         19571 => x"00000000",
         19572 => x"00000000",
         19573 => x"00000000",
         19574 => x"00000000",
         19575 => x"00000000",
         19576 => x"00000000",
         19577 => x"00000000",
         19578 => x"00000000",
         19579 => x"00000000",
         19580 => x"00000000",
         19581 => x"00000000",
         19582 => x"00000000",
         19583 => x"00000000",
         19584 => x"00000000",
         19585 => x"00000000",
         19586 => x"00000000",
         19587 => x"00000000",
         19588 => x"00000000",
         19589 => x"00000000",
         19590 => x"00000000",
         19591 => x"00000000",
         19592 => x"00000000",
         19593 => x"00000000",
         19594 => x"00000000",
         19595 => x"00000000",
         19596 => x"00000000",
         19597 => x"00000000",
         19598 => x"00000000",
         19599 => x"00000000",
         19600 => x"00000000",
         19601 => x"00000000",
         19602 => x"00000000",
         19603 => x"00000000",
         19604 => x"00000000",
         19605 => x"00000000",
         19606 => x"00000000",
         19607 => x"00000000",
         19608 => x"00000000",
         19609 => x"00000000",
         19610 => x"00000000",
         19611 => x"00000000",
         19612 => x"00000000",
         19613 => x"00000000",
         19614 => x"00000000",
         19615 => x"00000000",
         19616 => x"00000000",
         19617 => x"00000000",
         19618 => x"00000000",
         19619 => x"00000000",
         19620 => x"00000000",
         19621 => x"00000000",
         19622 => x"00000000",
         19623 => x"00000000",
         19624 => x"00000000",
         19625 => x"00000000",
         19626 => x"00000000",
         19627 => x"00000000",
         19628 => x"00000000",
         19629 => x"00000000",
         19630 => x"00000000",
         19631 => x"00000000",
         19632 => x"00000000",
         19633 => x"00000000",
         19634 => x"00000000",
         19635 => x"00000000",
         19636 => x"00000000",
         19637 => x"00000000",
         19638 => x"00000000",
         19639 => x"00000000",
         19640 => x"00000000",
         19641 => x"00000000",
         19642 => x"00000000",
         19643 => x"00000000",
         19644 => x"00000000",
         19645 => x"00000000",
         19646 => x"00000000",
         19647 => x"00000000",
         19648 => x"00000000",
         19649 => x"00000000",
         19650 => x"00000000",
         19651 => x"00000000",
         19652 => x"00000000",
         19653 => x"00000000",
         19654 => x"00000000",
         19655 => x"00000000",
         19656 => x"00000000",
         19657 => x"00000000",
         19658 => x"00000000",
         19659 => x"00000000",
         19660 => x"00000000",
         19661 => x"00000000",
         19662 => x"00000000",
         19663 => x"00000000",
         19664 => x"00000000",
         19665 => x"00000000",
         19666 => x"00000000",
         19667 => x"00000000",
         19668 => x"00000000",
         19669 => x"00000000",
         19670 => x"00000000",
         19671 => x"00000000",
         19672 => x"00000000",
         19673 => x"00000000",
         19674 => x"00000000",
         19675 => x"00000000",
         19676 => x"00000000",
         19677 => x"00000000",
         19678 => x"00000000",
         19679 => x"00000000",
         19680 => x"00000000",
         19681 => x"00000000",
         19682 => x"00000000",
         19683 => x"00000000",
         19684 => x"00000000",
         19685 => x"00000000",
         19686 => x"00000000",
         19687 => x"00000000",
         19688 => x"00000000",
         19689 => x"00000000",
         19690 => x"00000000",
         19691 => x"00000000",
         19692 => x"00000000",
         19693 => x"00000000",
         19694 => x"00000000",
         19695 => x"00000000",
         19696 => x"00000000",
         19697 => x"00000000",
         19698 => x"00000000",
         19699 => x"00000000",
         19700 => x"00000000",
         19701 => x"00000000",
         19702 => x"00000000",
         19703 => x"00000000",
         19704 => x"00000000",
         19705 => x"00000000",
         19706 => x"00000000",
         19707 => x"00000000",
         19708 => x"00000000",
         19709 => x"00000000",
         19710 => x"00000000",
         19711 => x"00000000",
         19712 => x"00000000",
         19713 => x"00000000",
         19714 => x"00000000",
         19715 => x"00000000",
         19716 => x"00000000",
         19717 => x"00000000",
         19718 => x"00000000",
         19719 => x"00000000",
         19720 => x"00000000",
         19721 => x"00000000",
         19722 => x"00000000",
         19723 => x"00000000",
         19724 => x"00000000",
         19725 => x"00000000",
         19726 => x"00000000",
         19727 => x"00000000",
         19728 => x"00000000",
         19729 => x"00000000",
         19730 => x"00000000",
         19731 => x"00000000",
         19732 => x"00000000",
         19733 => x"00000000",
         19734 => x"00000000",
         19735 => x"00000000",
         19736 => x"00000000",
         19737 => x"00000000",
         19738 => x"00000000",
         19739 => x"00000000",
         19740 => x"00000000",
         19741 => x"00000000",
         19742 => x"00000000",
         19743 => x"00000000",
         19744 => x"00000000",
         19745 => x"00000000",
         19746 => x"00000000",
         19747 => x"00000000",
         19748 => x"00000000",
         19749 => x"00000000",
         19750 => x"00000000",
         19751 => x"00000000",
         19752 => x"00000000",
         19753 => x"00000000",
         19754 => x"00000000",
         19755 => x"00000000",
         19756 => x"00000000",
         19757 => x"00000000",
         19758 => x"00000000",
         19759 => x"00000000",
         19760 => x"00000000",
         19761 => x"00000000",
         19762 => x"00000000",
         19763 => x"00000000",
         19764 => x"00000000",
         19765 => x"00000000",
         19766 => x"00000000",
         19767 => x"00000000",
         19768 => x"00000000",
         19769 => x"00000000",
         19770 => x"00000000",
         19771 => x"00000000",
         19772 => x"00000000",
         19773 => x"00000000",
         19774 => x"00000000",
         19775 => x"00000000",
         19776 => x"00000000",
         19777 => x"00000000",
         19778 => x"00000000",
         19779 => x"00000000",
         19780 => x"00000000",
         19781 => x"00000000",
         19782 => x"00000000",
         19783 => x"00000000",
         19784 => x"00000000",
         19785 => x"00000000",
         19786 => x"00000000",
         19787 => x"00000000",
         19788 => x"00000000",
         19789 => x"00000000",
         19790 => x"00000000",
         19791 => x"00000000",
         19792 => x"00000000",
         19793 => x"00000000",
         19794 => x"00000000",
         19795 => x"00000000",
         19796 => x"00000000",
         19797 => x"00000000",
         19798 => x"00000000",
         19799 => x"00000000",
         19800 => x"00000000",
         19801 => x"00000000",
         19802 => x"00000000",
         19803 => x"00000000",
         19804 => x"00000000",
         19805 => x"00000000",
         19806 => x"00000000",
         19807 => x"00000000",
         19808 => x"00000000",
         19809 => x"00000000",
         19810 => x"00000000",
         19811 => x"00000000",
         19812 => x"00000000",
         19813 => x"00000000",
         19814 => x"00000000",
         19815 => x"00000000",
         19816 => x"00000000",
         19817 => x"00000000",
         19818 => x"00000000",
         19819 => x"00000000",
         19820 => x"00000000",
         19821 => x"00000000",
         19822 => x"00000000",
         19823 => x"00000000",
         19824 => x"00000000",
         19825 => x"00000000",
         19826 => x"00000000",
         19827 => x"00000000",
         19828 => x"00000000",
         19829 => x"00000000",
         19830 => x"00000000",
         19831 => x"00000000",
         19832 => x"00000000",
         19833 => x"00000000",
         19834 => x"00000000",
         19835 => x"00000000",
         19836 => x"00000000",
         19837 => x"00000000",
         19838 => x"00000000",
         19839 => x"00000000",
         19840 => x"00000000",
         19841 => x"00000000",
         19842 => x"00000000",
         19843 => x"00000000",
         19844 => x"00000000",
         19845 => x"00000000",
         19846 => x"00000000",
         19847 => x"00000000",
         19848 => x"00000000",
         19849 => x"00000000",
         19850 => x"00000000",
         19851 => x"00000000",
         19852 => x"00000000",
         19853 => x"00000000",
         19854 => x"00000000",
         19855 => x"00000000",
         19856 => x"00000000",
         19857 => x"00000000",
         19858 => x"00000000",
         19859 => x"00000000",
         19860 => x"00000000",
         19861 => x"00000000",
         19862 => x"00000000",
         19863 => x"00000000",
         19864 => x"00000000",
         19865 => x"00000000",
         19866 => x"00000000",
         19867 => x"00000000",
         19868 => x"00000000",
         19869 => x"00000000",
         19870 => x"00000000",
         19871 => x"00000000",
         19872 => x"00000000",
         19873 => x"00000000",
         19874 => x"00000000",
         19875 => x"00000000",
         19876 => x"00000000",
         19877 => x"00000000",
         19878 => x"00000000",
         19879 => x"00000000",
         19880 => x"00000000",
         19881 => x"00000000",
         19882 => x"00000000",
         19883 => x"00000000",
         19884 => x"00000000",
         19885 => x"00000000",
         19886 => x"00000000",
         19887 => x"00000000",
         19888 => x"00000000",
         19889 => x"00000000",
         19890 => x"00000000",
         19891 => x"00000000",
         19892 => x"00000000",
         19893 => x"00000000",
         19894 => x"00000000",
         19895 => x"00000000",
         19896 => x"00000000",
         19897 => x"00000000",
         19898 => x"00000000",
         19899 => x"00000000",
         19900 => x"00000000",
         19901 => x"00000000",
         19902 => x"00000000",
         19903 => x"00000000",
         19904 => x"00000000",
         19905 => x"00000000",
         19906 => x"00000000",
         19907 => x"00000000",
         19908 => x"00000000",
         19909 => x"00000000",
         19910 => x"00000000",
         19911 => x"00000000",
         19912 => x"00000000",
         19913 => x"00000000",
         19914 => x"00000000",
         19915 => x"00000000",
         19916 => x"00000000",
         19917 => x"00000000",
         19918 => x"00000000",
         19919 => x"00000000",
         19920 => x"00000000",
         19921 => x"00000000",
         19922 => x"00000000",
         19923 => x"00000000",
         19924 => x"00000000",
         19925 => x"00000000",
         19926 => x"00000000",
         19927 => x"00000000",
         19928 => x"00000000",
         19929 => x"00000000",
         19930 => x"00000000",
         19931 => x"00000000",
         19932 => x"00000000",
         19933 => x"00000000",
         19934 => x"00000000",
         19935 => x"00000000",
         19936 => x"00000000",
         19937 => x"00000000",
         19938 => x"00000000",
         19939 => x"00000000",
         19940 => x"00000000",
         19941 => x"00000000",
         19942 => x"00000000",
         19943 => x"00000000",
         19944 => x"00000000",
         19945 => x"00000000",
         19946 => x"00000000",
         19947 => x"00000000",
         19948 => x"00000000",
         19949 => x"00000000",
         19950 => x"00000000",
         19951 => x"00000000",
         19952 => x"00000000",
         19953 => x"00000000",
         19954 => x"00000000",
         19955 => x"00000000",
         19956 => x"00000000",
         19957 => x"00000000",
         19958 => x"00000000",
         19959 => x"00000000",
         19960 => x"00000000",
         19961 => x"00000000",
         19962 => x"00000000",
         19963 => x"00000000",
         19964 => x"00000000",
         19965 => x"00000000",
         19966 => x"00000000",
         19967 => x"00000000",
         19968 => x"00000000",
         19969 => x"00000000",
         19970 => x"00000000",
         19971 => x"00000000",
         19972 => x"00000000",
         19973 => x"00000000",
         19974 => x"00000000",
         19975 => x"00000000",
         19976 => x"00000000",
         19977 => x"00000000",
         19978 => x"00000000",
         19979 => x"00000000",
         19980 => x"00000000",
         19981 => x"00000000",
         19982 => x"00000000",
         19983 => x"00000000",
         19984 => x"00000000",
         19985 => x"00000000",
         19986 => x"00000000",
         19987 => x"00000000",
         19988 => x"00000000",
         19989 => x"00000000",
         19990 => x"00000000",
         19991 => x"00000000",
         19992 => x"00000000",
         19993 => x"00000000",
         19994 => x"00000000",
         19995 => x"00000000",
         19996 => x"00000000",
         19997 => x"00000000",
         19998 => x"00000000",
         19999 => x"00000000",
         20000 => x"00000000",
         20001 => x"00000000",
         20002 => x"00000000",
         20003 => x"00000000",
         20004 => x"00000000",
         20005 => x"00000000",
         20006 => x"00000000",
         20007 => x"00000000",
         20008 => x"00000000",
         20009 => x"00000000",
         20010 => x"00000000",
         20011 => x"00000000",
         20012 => x"00000000",
         20013 => x"00000000",
         20014 => x"00000000",
         20015 => x"00000000",
         20016 => x"00000000",
         20017 => x"00000000",
         20018 => x"00000000",
         20019 => x"00000000",
         20020 => x"00000000",
         20021 => x"00000000",
         20022 => x"00000000",
         20023 => x"00000000",
         20024 => x"00000000",
         20025 => x"00000000",
         20026 => x"00000000",
         20027 => x"00000000",
         20028 => x"00000000",
         20029 => x"00000000",
         20030 => x"00000000",
         20031 => x"00000000",
         20032 => x"00000000",
         20033 => x"00000000",
         20034 => x"00000000",
         20035 => x"00000000",
         20036 => x"00000000",
         20037 => x"00000000",
         20038 => x"00000000",
         20039 => x"00000000",
         20040 => x"00000000",
         20041 => x"00000000",
         20042 => x"00000000",
         20043 => x"00000000",
         20044 => x"00000000",
         20045 => x"00000000",
         20046 => x"00000000",
         20047 => x"00000000",
         20048 => x"00000000",
         20049 => x"00000000",
         20050 => x"00000000",
         20051 => x"00000000",
         20052 => x"00000000",
         20053 => x"00000000",
         20054 => x"00000000",
         20055 => x"00000000",
         20056 => x"00000000",
         20057 => x"00000000",
         20058 => x"00000000",
         20059 => x"00000000",
         20060 => x"00000000",
         20061 => x"00000000",
         20062 => x"00000000",
         20063 => x"00000000",
         20064 => x"00000000",
         20065 => x"00000000",
         20066 => x"00000000",
         20067 => x"00000000",
         20068 => x"00000000",
         20069 => x"00000000",
         20070 => x"00000000",
         20071 => x"00000000",
         20072 => x"00000000",
         20073 => x"00000000",
         20074 => x"00000000",
         20075 => x"00000000",
         20076 => x"00000000",
         20077 => x"00000000",
         20078 => x"00000000",
         20079 => x"00000000",
         20080 => x"00000000",
         20081 => x"00000000",
         20082 => x"00000000",
         20083 => x"00000000",
         20084 => x"00000000",
         20085 => x"00000000",
         20086 => x"00000000",
         20087 => x"00000000",
         20088 => x"00000000",
         20089 => x"00000000",
         20090 => x"00000000",
         20091 => x"00000000",
         20092 => x"00000000",
         20093 => x"00000000",
         20094 => x"00000000",
         20095 => x"00000000",
         20096 => x"00000000",
         20097 => x"00000000",
         20098 => x"00000000",
         20099 => x"00000000",
         20100 => x"00000000",
         20101 => x"00000000",
         20102 => x"00000000",
         20103 => x"00000000",
         20104 => x"00000000",
         20105 => x"00000000",
         20106 => x"00000000",
         20107 => x"00000000",
         20108 => x"00000000",
         20109 => x"00000000",
         20110 => x"00000000",
         20111 => x"00000000",
         20112 => x"00000000",
         20113 => x"00000000",
         20114 => x"00000000",
         20115 => x"00000000",
         20116 => x"00000000",
         20117 => x"00000000",
         20118 => x"00000000",
         20119 => x"00000000",
         20120 => x"00000000",
         20121 => x"00000000",
         20122 => x"00000000",
         20123 => x"00000000",
         20124 => x"00000000",
         20125 => x"00000000",
         20126 => x"00000000",
         20127 => x"00000000",
         20128 => x"00000000",
         20129 => x"00000000",
         20130 => x"00000000",
         20131 => x"00000000",
         20132 => x"00000000",
         20133 => x"00000000",
         20134 => x"00000000",
         20135 => x"00000000",
         20136 => x"00000000",
         20137 => x"00000000",
         20138 => x"00000000",
         20139 => x"00000000",
         20140 => x"00000000",
         20141 => x"00000000",
         20142 => x"00000000",
         20143 => x"00000000",
         20144 => x"00000000",
         20145 => x"00000000",
         20146 => x"00000000",
         20147 => x"00000000",
         20148 => x"00000000",
         20149 => x"00000000",
         20150 => x"00000000",
         20151 => x"00000000",
         20152 => x"00000000",
         20153 => x"00000000",
         20154 => x"00000000",
         20155 => x"00000000",
         20156 => x"00000000",
         20157 => x"00000000",
         20158 => x"00000000",
         20159 => x"00000000",
         20160 => x"00000000",
         20161 => x"00000000",
         20162 => x"00000000",
         20163 => x"00000000",
         20164 => x"00000000",
         20165 => x"00000000",
         20166 => x"00000000",
         20167 => x"00000000",
         20168 => x"00000000",
         20169 => x"00000000",
         20170 => x"00000000",
         20171 => x"00000000",
         20172 => x"00000000",
         20173 => x"00000000",
         20174 => x"00000000",
         20175 => x"00000000",
         20176 => x"00000000",
         20177 => x"00000000",
         20178 => x"00000000",
         20179 => x"00000000",
         20180 => x"00000000",
         20181 => x"00000000",
         20182 => x"00000000",
         20183 => x"00000000",
         20184 => x"00000000",
         20185 => x"00000000",
         20186 => x"00000000",
         20187 => x"00000000",
         20188 => x"00000000",
         20189 => x"00000000",
         20190 => x"00000000",
         20191 => x"00000000",
         20192 => x"00000000",
         20193 => x"00000000",
         20194 => x"00000000",
         20195 => x"00000000",
         20196 => x"00000000",
         20197 => x"00000000",
         20198 => x"00000000",
         20199 => x"00000000",
         20200 => x"00000000",
         20201 => x"00000000",
         20202 => x"00000000",
         20203 => x"00000000",
         20204 => x"00000000",
         20205 => x"00000000",
         20206 => x"00003219",
         20207 => x"50000100",
         20208 => x"00000000",
         20209 => x"cce0f2f3",
         20210 => x"cecff6f7",
         20211 => x"f8f9fafb",
         20212 => x"fcfdfeff",
         20213 => x"e1c1c2c3",
         20214 => x"c4c5c6e2",
         20215 => x"e3e4e5e6",
         20216 => x"ebeeeff4",
         20217 => x"00616263",
         20218 => x"64656667",
         20219 => x"68696b6a",
         20220 => x"2f2a2e2d",
         20221 => x"20212223",
         20222 => x"24252627",
         20223 => x"28294f2c",
         20224 => x"512b5749",
         20225 => x"55010203",
         20226 => x"04050607",
         20227 => x"08090a0b",
         20228 => x"0c0d0e0f",
         20229 => x"10111213",
         20230 => x"14151617",
         20231 => x"18191a52",
         20232 => x"5954be3c",
         20233 => x"c7818283",
         20234 => x"84858687",
         20235 => x"88898a8b",
         20236 => x"8c8d8e8f",
         20237 => x"90919293",
         20238 => x"94959697",
         20239 => x"98999abc",
         20240 => x"8040a5c0",
         20241 => x"00000000",
         20242 => x"00000000",
         20243 => x"00000000",
         20244 => x"00000000",
         20245 => x"00000000",
         20246 => x"00000000",
         20247 => x"00000000",
         20248 => x"00000000",
         20249 => x"00000000",
         20250 => x"00000000",
         20251 => x"00000000",
         20252 => x"00000000",
         20253 => x"00000000",
         20254 => x"00000000",
         20255 => x"00000000",
         20256 => x"00000000",
         20257 => x"00000000",
         20258 => x"00000000",
         20259 => x"00000000",
         20260 => x"00000000",
         20261 => x"00000000",
         20262 => x"00000000",
         20263 => x"00000000",
         20264 => x"00000000",
         20265 => x"00000000",
         20266 => x"00000000",
         20267 => x"00000000",
         20268 => x"00000000",
         20269 => x"00000000",
         20270 => x"00000000",
         20271 => x"00020003",
         20272 => x"00040101",
         20273 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

