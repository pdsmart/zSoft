-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b83ff",
          2049 => x"f80d0b0b",
          2050 => x"0b93b904",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b93",
          2121 => x"9d040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b9380",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b82ac",
          2210 => x"cc738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"93850400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b80c5",
          2219 => x"9f2d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b80c7",
          2227 => x"8b2d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"95040b0b",
          2317 => x"0b8ca404",
          2318 => x"0b0b0b8c",
          2319 => x"b3040b0b",
          2320 => x"0b8cc204",
          2321 => x"0b0b0b8c",
          2322 => x"d1040b0b",
          2323 => x"0b8ce004",
          2324 => x"0b0b0b8c",
          2325 => x"f0040b0b",
          2326 => x"0b8d8004",
          2327 => x"0b0b0b8d",
          2328 => x"8f040b0b",
          2329 => x"0b8d9e04",
          2330 => x"0b0b0b8d",
          2331 => x"ad040b0b",
          2332 => x"0b8dbd04",
          2333 => x"0b0b0b8d",
          2334 => x"cd040b0b",
          2335 => x"0b8ddd04",
          2336 => x"0b0b0b8d",
          2337 => x"ed040b0b",
          2338 => x"0b8dfd04",
          2339 => x"0b0b0b8e",
          2340 => x"8d040b0b",
          2341 => x"0b8e9d04",
          2342 => x"0b0b0b8e",
          2343 => x"ad040b0b",
          2344 => x"0b8ebd04",
          2345 => x"0b0b0b8e",
          2346 => x"cd040b0b",
          2347 => x"0b8edd04",
          2348 => x"0b0b0b8e",
          2349 => x"ed040b0b",
          2350 => x"0b8efd04",
          2351 => x"0b0b0b8f",
          2352 => x"8d040b0b",
          2353 => x"0b8f9d04",
          2354 => x"0b0b0b8f",
          2355 => x"ad040b0b",
          2356 => x"0b8fbd04",
          2357 => x"0b0b0b8f",
          2358 => x"cd040b0b",
          2359 => x"0b8fdd04",
          2360 => x"0b0b0b8f",
          2361 => x"ed040b0b",
          2362 => x"0b8ffd04",
          2363 => x"0b0b0b90",
          2364 => x"8d040b0b",
          2365 => x"0b909d04",
          2366 => x"0b0b0b90",
          2367 => x"ad040b0b",
          2368 => x"0b90bd04",
          2369 => x"0b0b0b90",
          2370 => x"cd040b0b",
          2371 => x"0b90dd04",
          2372 => x"0b0b0b90",
          2373 => x"ed040b0b",
          2374 => x"0b90fd04",
          2375 => x"0b0b0b91",
          2376 => x"8d040b0b",
          2377 => x"0b919d04",
          2378 => x"0b0b0b91",
          2379 => x"ad040b0b",
          2380 => x"0b91bd04",
          2381 => x"0b0b0b91",
          2382 => x"cd040b0b",
          2383 => x"0b91dd04",
          2384 => x"0b0b0b91",
          2385 => x"ed040b0b",
          2386 => x"0b91fd04",
          2387 => x"0b0b0b92",
          2388 => x"8d040b0b",
          2389 => x"0b929d04",
          2390 => x"0b0b0b92",
          2391 => x"ad040b0b",
          2392 => x"0b92bd04",
          2393 => x"0b0b0b92",
          2394 => x"cd04ffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0482d6e4",
          2434 => x"0c80f7d4",
          2435 => x"2d82d6e4",
          2436 => x"08848090",
          2437 => x"0482d6e4",
          2438 => x"0cb3b22d",
          2439 => x"82d6e408",
          2440 => x"84809004",
          2441 => x"82d6e40c",
          2442 => x"afe32d82",
          2443 => x"d6e40884",
          2444 => x"80900482",
          2445 => x"d6e40caf",
          2446 => x"ad2d82d6",
          2447 => x"e4088480",
          2448 => x"900482d6",
          2449 => x"e40c94ad",
          2450 => x"2d82d6e4",
          2451 => x"08848090",
          2452 => x"0482d6e4",
          2453 => x"0cb1c22d",
          2454 => x"82d6e408",
          2455 => x"84809004",
          2456 => x"82d6e40c",
          2457 => x"80d0f72d",
          2458 => x"82d6e408",
          2459 => x"84809004",
          2460 => x"82d6e40c",
          2461 => x"80cba62d",
          2462 => x"82d6e408",
          2463 => x"84809004",
          2464 => x"82d6e40c",
          2465 => x"93d82d82",
          2466 => x"d6e40884",
          2467 => x"80900482",
          2468 => x"d6e40c96",
          2469 => x"c02d82d6",
          2470 => x"e4088480",
          2471 => x"900482d6",
          2472 => x"e40c97cd",
          2473 => x"2d82d6e4",
          2474 => x"08848090",
          2475 => x"0482d6e4",
          2476 => x"0c80f9fa",
          2477 => x"2d82d6e4",
          2478 => x"08848090",
          2479 => x"0482d6e4",
          2480 => x"0c80fac9",
          2481 => x"2d82d6e4",
          2482 => x"08848090",
          2483 => x"0482d6e4",
          2484 => x"0c80f399",
          2485 => x"2d82d6e4",
          2486 => x"08848090",
          2487 => x"0482d6e4",
          2488 => x"0c80f590",
          2489 => x"2d82d6e4",
          2490 => x"08848090",
          2491 => x"0482d6e4",
          2492 => x"0c80f6c3",
          2493 => x"2d82d6e4",
          2494 => x"08848090",
          2495 => x"0482d6e4",
          2496 => x"0c81ecad",
          2497 => x"2d82d6e4",
          2498 => x"08848090",
          2499 => x"0482d6e4",
          2500 => x"0c81f9ac",
          2501 => x"2d82d6e4",
          2502 => x"08848090",
          2503 => x"0482d6e4",
          2504 => x"0c81f192",
          2505 => x"2d82d6e4",
          2506 => x"08848090",
          2507 => x"0482d6e4",
          2508 => x"0c81f492",
          2509 => x"2d82d6e4",
          2510 => x"08848090",
          2511 => x"0482d6e4",
          2512 => x"0c81feea",
          2513 => x"2d82d6e4",
          2514 => x"08848090",
          2515 => x"0482d6e4",
          2516 => x"0c8287d3",
          2517 => x"2d82d6e4",
          2518 => x"08848090",
          2519 => x"0482d6e4",
          2520 => x"0c81f889",
          2521 => x"2d82d6e4",
          2522 => x"08848090",
          2523 => x"0482d6e4",
          2524 => x"0c82828d",
          2525 => x"2d82d6e4",
          2526 => x"08848090",
          2527 => x"0482d6e4",
          2528 => x"0c8283ad",
          2529 => x"2d82d6e4",
          2530 => x"08848090",
          2531 => x"0482d6e4",
          2532 => x"0c8283cc",
          2533 => x"2d82d6e4",
          2534 => x"08848090",
          2535 => x"0482d6e4",
          2536 => x"0c828bc0",
          2537 => x"2d82d6e4",
          2538 => x"08848090",
          2539 => x"0482d6e4",
          2540 => x"0c8289a2",
          2541 => x"2d82d6e4",
          2542 => x"08848090",
          2543 => x"0482d6e4",
          2544 => x"0c828e9c",
          2545 => x"2d82d6e4",
          2546 => x"08848090",
          2547 => x"0482d6e4",
          2548 => x"0c8284d2",
          2549 => x"2d82d6e4",
          2550 => x"08848090",
          2551 => x"0482d6e4",
          2552 => x"0c8291a1",
          2553 => x"2d82d6e4",
          2554 => x"08848090",
          2555 => x"0482d6e4",
          2556 => x"0c8292a2",
          2557 => x"2d82d6e4",
          2558 => x"08848090",
          2559 => x"0482d6e4",
          2560 => x"0c81fa8c",
          2561 => x"2d82d6e4",
          2562 => x"08848090",
          2563 => x"0482d6e4",
          2564 => x"0c81f9e5",
          2565 => x"2d82d6e4",
          2566 => x"08848090",
          2567 => x"0482d6e4",
          2568 => x"0c81fb90",
          2569 => x"2d82d6e4",
          2570 => x"08848090",
          2571 => x"0482d6e4",
          2572 => x"0c8285a9",
          2573 => x"2d82d6e4",
          2574 => x"08848090",
          2575 => x"0482d6e4",
          2576 => x"0c829393",
          2577 => x"2d82d6e4",
          2578 => x"08848090",
          2579 => x"0482d6e4",
          2580 => x"0c82959e",
          2581 => x"2d82d6e4",
          2582 => x"08848090",
          2583 => x"0482d6e4",
          2584 => x"0c8298a5",
          2585 => x"2d82d6e4",
          2586 => x"08848090",
          2587 => x"0482d6e4",
          2588 => x"0c81ebcc",
          2589 => x"2d82d6e4",
          2590 => x"08848090",
          2591 => x"0482d6e4",
          2592 => x"0c829b91",
          2593 => x"2d82d6e4",
          2594 => x"08848090",
          2595 => x"0482d6e4",
          2596 => x"0c82a9c6",
          2597 => x"2d82d6e4",
          2598 => x"08848090",
          2599 => x"0482d6e4",
          2600 => x"0c82a7b2",
          2601 => x"2d82d6e4",
          2602 => x"08848090",
          2603 => x"0482d6e4",
          2604 => x"0c81abd4",
          2605 => x"2d82d6e4",
          2606 => x"08848090",
          2607 => x"0482d6e4",
          2608 => x"0c81adbe",
          2609 => x"2d82d6e4",
          2610 => x"08848090",
          2611 => x"0482d6e4",
          2612 => x"0c81afa2",
          2613 => x"2d82d6e4",
          2614 => x"08848090",
          2615 => x"0482d6e4",
          2616 => x"0c80f3c2",
          2617 => x"2d82d6e4",
          2618 => x"08848090",
          2619 => x"0482d6e4",
          2620 => x"0c80f4e6",
          2621 => x"2d82d6e4",
          2622 => x"08848090",
          2623 => x"0482d6e4",
          2624 => x"0c80f8c9",
          2625 => x"2d82d6e4",
          2626 => x"08848090",
          2627 => x"0482d6e4",
          2628 => x"0c80d7bf",
          2629 => x"2d82d6e4",
          2630 => x"08848090",
          2631 => x"0482d6e4",
          2632 => x"0c81a5e8",
          2633 => x"2d82d6e4",
          2634 => x"08848090",
          2635 => x"0482d6e4",
          2636 => x"0c81a690",
          2637 => x"2d82d6e4",
          2638 => x"08848090",
          2639 => x"0482d6e4",
          2640 => x"0c81aa88",
          2641 => x"2d82d6e4",
          2642 => x"08848090",
          2643 => x"0482d6e4",
          2644 => x"0c81a2d2",
          2645 => x"2d82d6e4",
          2646 => x"08848090",
          2647 => x"043c0400",
          2648 => x"00101010",
          2649 => x"10101010",
          2650 => x"10101010",
          2651 => x"10101010",
          2652 => x"10101010",
          2653 => x"10101010",
          2654 => x"10101010",
          2655 => x"10101010",
          2656 => x"53510400",
          2657 => x"007381ff",
          2658 => x"06738306",
          2659 => x"09810583",
          2660 => x"05101010",
          2661 => x"2b0772fc",
          2662 => x"060c5151",
          2663 => x"04727280",
          2664 => x"728106ff",
          2665 => x"05097206",
          2666 => x"05711052",
          2667 => x"720a100a",
          2668 => x"5372ed38",
          2669 => x"51515351",
          2670 => x"0482d6d8",
          2671 => x"7082f2c4",
          2672 => x"278e3880",
          2673 => x"71708405",
          2674 => x"530c0b0b",
          2675 => x"0b93bc04",
          2676 => x"8c815180",
          2677 => x"f0ec0400",
          2678 => x"82d6e408",
          2679 => x"0282d6e4",
          2680 => x"0cfb3d0d",
          2681 => x"82d6e408",
          2682 => x"8c057082",
          2683 => x"d6e408fc",
          2684 => x"050c82d6",
          2685 => x"e408fc05",
          2686 => x"085482d6",
          2687 => x"e4088805",
          2688 => x"085382f2",
          2689 => x"bc085254",
          2690 => x"849a3f82",
          2691 => x"d6d80870",
          2692 => x"82d6e408",
          2693 => x"f8050c82",
          2694 => x"d6e408f8",
          2695 => x"05087082",
          2696 => x"d6d80c51",
          2697 => x"54873d0d",
          2698 => x"82d6e40c",
          2699 => x"0482d6e4",
          2700 => x"080282d6",
          2701 => x"e40cfb3d",
          2702 => x"0d82d6e4",
          2703 => x"08900508",
          2704 => x"85113370",
          2705 => x"81327081",
          2706 => x"06515151",
          2707 => x"52718f38",
          2708 => x"800b82d6",
          2709 => x"e4088c05",
          2710 => x"08258338",
          2711 => x"8d39800b",
          2712 => x"82d6e408",
          2713 => x"f4050c81",
          2714 => x"c43982d6",
          2715 => x"e4088c05",
          2716 => x"08ff0582",
          2717 => x"d6e4088c",
          2718 => x"050c800b",
          2719 => x"82d6e408",
          2720 => x"f8050c82",
          2721 => x"d6e40888",
          2722 => x"050882d6",
          2723 => x"e408fc05",
          2724 => x"0c82d6e4",
          2725 => x"08f80508",
          2726 => x"8a2e80f6",
          2727 => x"38800b82",
          2728 => x"d6e4088c",
          2729 => x"05082580",
          2730 => x"e93882d6",
          2731 => x"e4089005",
          2732 => x"0851a090",
          2733 => x"3f82d6d8",
          2734 => x"087082d6",
          2735 => x"e408f805",
          2736 => x"0c5282d6",
          2737 => x"e408f805",
          2738 => x"08ff2e09",
          2739 => x"81068d38",
          2740 => x"800b82d6",
          2741 => x"e408f405",
          2742 => x"0c80d239",
          2743 => x"82d6e408",
          2744 => x"fc050882",
          2745 => x"d6e408f8",
          2746 => x"05085353",
          2747 => x"71733482",
          2748 => x"d6e4088c",
          2749 => x"0508ff05",
          2750 => x"82d6e408",
          2751 => x"8c050c82",
          2752 => x"d6e408fc",
          2753 => x"05088105",
          2754 => x"82d6e408",
          2755 => x"fc050cff",
          2756 => x"803982d6",
          2757 => x"e408fc05",
          2758 => x"08528072",
          2759 => x"3482d6e4",
          2760 => x"08880508",
          2761 => x"7082d6e4",
          2762 => x"08f4050c",
          2763 => x"5282d6e4",
          2764 => x"08f40508",
          2765 => x"82d6d80c",
          2766 => x"873d0d82",
          2767 => x"d6e40c04",
          2768 => x"82d6e408",
          2769 => x"0282d6e4",
          2770 => x"0cf43d0d",
          2771 => x"860b82d6",
          2772 => x"e408e505",
          2773 => x"3482d6e4",
          2774 => x"08880508",
          2775 => x"82d6e408",
          2776 => x"e0050cfe",
          2777 => x"0a0b82d6",
          2778 => x"e408e805",
          2779 => x"0c82d6e4",
          2780 => x"08900570",
          2781 => x"82d6e408",
          2782 => x"fc050c82",
          2783 => x"d6e408fc",
          2784 => x"05085482",
          2785 => x"d6e4088c",
          2786 => x"05085382",
          2787 => x"d6e408e0",
          2788 => x"05705351",
          2789 => x"54818d3f",
          2790 => x"82d6d808",
          2791 => x"7082d6e4",
          2792 => x"08dc050c",
          2793 => x"82d6e408",
          2794 => x"ec050882",
          2795 => x"d6e40888",
          2796 => x"05080551",
          2797 => x"54807434",
          2798 => x"82d6e408",
          2799 => x"dc050870",
          2800 => x"82d6d80c",
          2801 => x"548e3d0d",
          2802 => x"82d6e40c",
          2803 => x"0482d6e4",
          2804 => x"080282d6",
          2805 => x"e40cfb3d",
          2806 => x"0d82d6e4",
          2807 => x"08900570",
          2808 => x"82d6e408",
          2809 => x"fc050c82",
          2810 => x"d6e408fc",
          2811 => x"05085482",
          2812 => x"d6e4088c",
          2813 => x"05085382",
          2814 => x"d6e40888",
          2815 => x"05085254",
          2816 => x"a33f82d6",
          2817 => x"d8087082",
          2818 => x"d6e408f8",
          2819 => x"050c82d6",
          2820 => x"e408f805",
          2821 => x"087082d6",
          2822 => x"d80c5154",
          2823 => x"873d0d82",
          2824 => x"d6e40c04",
          2825 => x"82d6e408",
          2826 => x"0282d6e4",
          2827 => x"0ced3d0d",
          2828 => x"800b82d6",
          2829 => x"e408e405",
          2830 => x"2382d6e4",
          2831 => x"08880508",
          2832 => x"53800b8c",
          2833 => x"140c82d6",
          2834 => x"e4088805",
          2835 => x"08851133",
          2836 => x"70812a70",
          2837 => x"81327081",
          2838 => x"06515151",
          2839 => x"51537280",
          2840 => x"2e8d38ff",
          2841 => x"0b82d6e4",
          2842 => x"08e0050c",
          2843 => x"96ac3982",
          2844 => x"d6e4088c",
          2845 => x"05085372",
          2846 => x"33537282",
          2847 => x"d6e408f8",
          2848 => x"05347281",
          2849 => x"ff065372",
          2850 => x"802e95fa",
          2851 => x"3882d6e4",
          2852 => x"088c0508",
          2853 => x"810582d6",
          2854 => x"e4088c05",
          2855 => x"0c82d6e4",
          2856 => x"08e40522",
          2857 => x"70810651",
          2858 => x"5372802e",
          2859 => x"958b3882",
          2860 => x"d6e408f8",
          2861 => x"053353af",
          2862 => x"732781fc",
          2863 => x"3882d6e4",
          2864 => x"08f80533",
          2865 => x"5372b926",
          2866 => x"81ee3882",
          2867 => x"d6e408f8",
          2868 => x"05335372",
          2869 => x"b02e0981",
          2870 => x"0680c538",
          2871 => x"82d6e408",
          2872 => x"e8053370",
          2873 => x"982b7098",
          2874 => x"2c515153",
          2875 => x"72b23882",
          2876 => x"d6e408e4",
          2877 => x"05227083",
          2878 => x"2a708132",
          2879 => x"70810651",
          2880 => x"51515372",
          2881 => x"802e9938",
          2882 => x"82d6e408",
          2883 => x"e4052270",
          2884 => x"82800751",
          2885 => x"537282d6",
          2886 => x"e408e405",
          2887 => x"23fed039",
          2888 => x"82d6e408",
          2889 => x"e8053370",
          2890 => x"982b7098",
          2891 => x"2c707083",
          2892 => x"2b721173",
          2893 => x"11515151",
          2894 => x"53515553",
          2895 => x"7282d6e4",
          2896 => x"08e80534",
          2897 => x"82d6e408",
          2898 => x"e8053354",
          2899 => x"82d6e408",
          2900 => x"f8053370",
          2901 => x"15d01151",
          2902 => x"51537282",
          2903 => x"d6e408e8",
          2904 => x"053482d6",
          2905 => x"e408e805",
          2906 => x"3370982b",
          2907 => x"70982c51",
          2908 => x"51537280",
          2909 => x"258b3880",
          2910 => x"ff0b82d6",
          2911 => x"e408e805",
          2912 => x"3482d6e4",
          2913 => x"08e40522",
          2914 => x"70832a70",
          2915 => x"81065151",
          2916 => x"5372fddb",
          2917 => x"3882d6e4",
          2918 => x"08e80533",
          2919 => x"70882b70",
          2920 => x"902b7090",
          2921 => x"2c70882c",
          2922 => x"51515151",
          2923 => x"537282d6",
          2924 => x"e408ec05",
          2925 => x"23fdb839",
          2926 => x"82d6e408",
          2927 => x"e4052270",
          2928 => x"832a7081",
          2929 => x"06515153",
          2930 => x"72802e9d",
          2931 => x"3882d6e4",
          2932 => x"08e80533",
          2933 => x"70982b70",
          2934 => x"982c5151",
          2935 => x"53728a38",
          2936 => x"810b82d6",
          2937 => x"e408e805",
          2938 => x"3482d6e4",
          2939 => x"08f80533",
          2940 => x"e01182d6",
          2941 => x"e408c405",
          2942 => x"0c5382d6",
          2943 => x"e408c405",
          2944 => x"0880d826",
          2945 => x"92943882",
          2946 => x"d6e408c4",
          2947 => x"05087082",
          2948 => x"2b82aebc",
          2949 => x"11700851",
          2950 => x"51515372",
          2951 => x"0482d6e4",
          2952 => x"08e40522",
          2953 => x"70900751",
          2954 => x"537282d6",
          2955 => x"e408e405",
          2956 => x"2382d6e4",
          2957 => x"08e40522",
          2958 => x"70a00751",
          2959 => x"537282d6",
          2960 => x"e408e405",
          2961 => x"23fca839",
          2962 => x"82d6e408",
          2963 => x"e4052270",
          2964 => x"81800751",
          2965 => x"537282d6",
          2966 => x"e408e405",
          2967 => x"23fc9039",
          2968 => x"82d6e408",
          2969 => x"e4052270",
          2970 => x"80c00751",
          2971 => x"537282d6",
          2972 => x"e408e405",
          2973 => x"23fbf839",
          2974 => x"82d6e408",
          2975 => x"e4052270",
          2976 => x"88075153",
          2977 => x"7282d6e4",
          2978 => x"08e40523",
          2979 => x"800b82d6",
          2980 => x"e408e805",
          2981 => x"34fbd839",
          2982 => x"82d6e408",
          2983 => x"e4052270",
          2984 => x"84075153",
          2985 => x"7282d6e4",
          2986 => x"08e40523",
          2987 => x"fbc139bf",
          2988 => x"0b82d6e4",
          2989 => x"08fc0534",
          2990 => x"82d6e408",
          2991 => x"ec0522ff",
          2992 => x"11515372",
          2993 => x"82d6e408",
          2994 => x"ec052380",
          2995 => x"e30b82d6",
          2996 => x"e408f805",
          2997 => x"348da839",
          2998 => x"82d6e408",
          2999 => x"90050882",
          3000 => x"d6e40890",
          3001 => x"05088405",
          3002 => x"82d6e408",
          3003 => x"90050c70",
          3004 => x"08515372",
          3005 => x"82d6e408",
          3006 => x"fc053482",
          3007 => x"d6e408ec",
          3008 => x"0522ff11",
          3009 => x"51537282",
          3010 => x"d6e408ec",
          3011 => x"05238cef",
          3012 => x"3982d6e4",
          3013 => x"08900508",
          3014 => x"82d6e408",
          3015 => x"90050884",
          3016 => x"0582d6e4",
          3017 => x"0890050c",
          3018 => x"700882d6",
          3019 => x"e408fc05",
          3020 => x"0c82d6e4",
          3021 => x"08e40522",
          3022 => x"70832a70",
          3023 => x"81065151",
          3024 => x"51537280",
          3025 => x"2eab3882",
          3026 => x"d6e408e8",
          3027 => x"05337098",
          3028 => x"2b537298",
          3029 => x"2c5382d6",
          3030 => x"e408fc05",
          3031 => x"085253a4",
          3032 => x"833f82d6",
          3033 => x"d8085372",
          3034 => x"82d6e408",
          3035 => x"f4052399",
          3036 => x"3982d6e4",
          3037 => x"08fc0508",
          3038 => x"519d8a3f",
          3039 => x"82d6d808",
          3040 => x"537282d6",
          3041 => x"e408f405",
          3042 => x"2382d6e4",
          3043 => x"08ec0522",
          3044 => x"5382d6e4",
          3045 => x"08f40522",
          3046 => x"73713154",
          3047 => x"547282d6",
          3048 => x"e408ec05",
          3049 => x"238bd839",
          3050 => x"82d6e408",
          3051 => x"90050882",
          3052 => x"d6e40890",
          3053 => x"05088405",
          3054 => x"82d6e408",
          3055 => x"90050c70",
          3056 => x"0882d6e4",
          3057 => x"08fc050c",
          3058 => x"82d6e408",
          3059 => x"e4052270",
          3060 => x"832a7081",
          3061 => x"06515151",
          3062 => x"5372802e",
          3063 => x"ab3882d6",
          3064 => x"e408e805",
          3065 => x"3370982b",
          3066 => x"5372982c",
          3067 => x"5382d6e4",
          3068 => x"08fc0508",
          3069 => x"5253a2ec",
          3070 => x"3f82d6d8",
          3071 => x"08537282",
          3072 => x"d6e408f4",
          3073 => x"05239939",
          3074 => x"82d6e408",
          3075 => x"fc050851",
          3076 => x"9bf33f82",
          3077 => x"d6d80853",
          3078 => x"7282d6e4",
          3079 => x"08f40523",
          3080 => x"82d6e408",
          3081 => x"ec052253",
          3082 => x"82d6e408",
          3083 => x"f4052273",
          3084 => x"71315454",
          3085 => x"7282d6e4",
          3086 => x"08ec0523",
          3087 => x"8ac13982",
          3088 => x"d6e408e4",
          3089 => x"05227082",
          3090 => x"2a708106",
          3091 => x"51515372",
          3092 => x"802ea438",
          3093 => x"82d6e408",
          3094 => x"90050882",
          3095 => x"d6e40890",
          3096 => x"05088405",
          3097 => x"82d6e408",
          3098 => x"90050c70",
          3099 => x"0882d6e4",
          3100 => x"08dc050c",
          3101 => x"53a23982",
          3102 => x"d6e40890",
          3103 => x"050882d6",
          3104 => x"e4089005",
          3105 => x"08840582",
          3106 => x"d6e40890",
          3107 => x"050c7008",
          3108 => x"82d6e408",
          3109 => x"dc050c53",
          3110 => x"82d6e408",
          3111 => x"dc050882",
          3112 => x"d6e408fc",
          3113 => x"050c82d6",
          3114 => x"e408fc05",
          3115 => x"088025a4",
          3116 => x"3882d6e4",
          3117 => x"08e40522",
          3118 => x"70820751",
          3119 => x"537282d6",
          3120 => x"e408e405",
          3121 => x"2382d6e4",
          3122 => x"08fc0508",
          3123 => x"3082d6e4",
          3124 => x"08fc050c",
          3125 => x"82d6e408",
          3126 => x"e4052270",
          3127 => x"ffbf0651",
          3128 => x"537282d6",
          3129 => x"e408e405",
          3130 => x"2381af39",
          3131 => x"880b82d6",
          3132 => x"e408f405",
          3133 => x"23a93982",
          3134 => x"d6e408e4",
          3135 => x"05227080",
          3136 => x"c0075153",
          3137 => x"7282d6e4",
          3138 => x"08e40523",
          3139 => x"80f80b82",
          3140 => x"d6e408f8",
          3141 => x"0534900b",
          3142 => x"82d6e408",
          3143 => x"f4052382",
          3144 => x"d6e408e4",
          3145 => x"05227082",
          3146 => x"2a708106",
          3147 => x"51515372",
          3148 => x"802ea438",
          3149 => x"82d6e408",
          3150 => x"90050882",
          3151 => x"d6e40890",
          3152 => x"05088405",
          3153 => x"82d6e408",
          3154 => x"90050c70",
          3155 => x"0882d6e4",
          3156 => x"08d8050c",
          3157 => x"53a23982",
          3158 => x"d6e40890",
          3159 => x"050882d6",
          3160 => x"e4089005",
          3161 => x"08840582",
          3162 => x"d6e40890",
          3163 => x"050c7008",
          3164 => x"82d6e408",
          3165 => x"d8050c53",
          3166 => x"82d6e408",
          3167 => x"d8050882",
          3168 => x"d6e408fc",
          3169 => x"050c82d6",
          3170 => x"e408e405",
          3171 => x"2270cf06",
          3172 => x"51537282",
          3173 => x"d6e408e4",
          3174 => x"052382d6",
          3175 => x"e80b82d6",
          3176 => x"e408f005",
          3177 => x"0c82d6e4",
          3178 => x"08f00508",
          3179 => x"82d6e408",
          3180 => x"f4052282",
          3181 => x"d6e408fc",
          3182 => x"05087155",
          3183 => x"70545654",
          3184 => x"55a59e3f",
          3185 => x"82d6d808",
          3186 => x"53727534",
          3187 => x"82d6e408",
          3188 => x"f0050882",
          3189 => x"d6e408d4",
          3190 => x"050c82d6",
          3191 => x"e408f005",
          3192 => x"08703351",
          3193 => x"53897327",
          3194 => x"a43882d6",
          3195 => x"e408f005",
          3196 => x"08537233",
          3197 => x"5482d6e4",
          3198 => x"08f80533",
          3199 => x"7015df11",
          3200 => x"51515372",
          3201 => x"82d6e408",
          3202 => x"d0053497",
          3203 => x"3982d6e4",
          3204 => x"08f00508",
          3205 => x"537233b0",
          3206 => x"11515372",
          3207 => x"82d6e408",
          3208 => x"d0053482",
          3209 => x"d6e408d4",
          3210 => x"05085382",
          3211 => x"d6e408d0",
          3212 => x"05337334",
          3213 => x"82d6e408",
          3214 => x"f0050881",
          3215 => x"0582d6e4",
          3216 => x"08f0050c",
          3217 => x"82d6e408",
          3218 => x"f4052270",
          3219 => x"5382d6e4",
          3220 => x"08fc0508",
          3221 => x"5253a3d6",
          3222 => x"3f82d6d8",
          3223 => x"087082d6",
          3224 => x"e408fc05",
          3225 => x"0c5382d6",
          3226 => x"e408fc05",
          3227 => x"08802e84",
          3228 => x"38feb239",
          3229 => x"82d6e408",
          3230 => x"f0050882",
          3231 => x"d6e85455",
          3232 => x"72547470",
          3233 => x"75315153",
          3234 => x"7282d6e4",
          3235 => x"08fc0534",
          3236 => x"82d6e408",
          3237 => x"e4052270",
          3238 => x"b2065153",
          3239 => x"72802e94",
          3240 => x"3882d6e4",
          3241 => x"08ec0522",
          3242 => x"ff115153",
          3243 => x"7282d6e4",
          3244 => x"08ec0523",
          3245 => x"82d6e408",
          3246 => x"e4052270",
          3247 => x"862a7081",
          3248 => x"06515153",
          3249 => x"72802e80",
          3250 => x"e73882d6",
          3251 => x"e408ec05",
          3252 => x"2270902b",
          3253 => x"82d6e408",
          3254 => x"cc050c82",
          3255 => x"d6e408cc",
          3256 => x"0508902c",
          3257 => x"82d6e408",
          3258 => x"cc050c82",
          3259 => x"d6e408f4",
          3260 => x"05225153",
          3261 => x"72902e09",
          3262 => x"81069538",
          3263 => x"82d6e408",
          3264 => x"cc0508fe",
          3265 => x"05537282",
          3266 => x"d6e408c8",
          3267 => x"05239339",
          3268 => x"82d6e408",
          3269 => x"cc0508ff",
          3270 => x"05537282",
          3271 => x"d6e408c8",
          3272 => x"052382d6",
          3273 => x"e408c805",
          3274 => x"2282d6e4",
          3275 => x"08ec0523",
          3276 => x"82d6e408",
          3277 => x"e4052270",
          3278 => x"832a7081",
          3279 => x"06515153",
          3280 => x"72802e80",
          3281 => x"d03882d6",
          3282 => x"e408e805",
          3283 => x"3370982b",
          3284 => x"70982c82",
          3285 => x"d6e408fc",
          3286 => x"05335751",
          3287 => x"51537274",
          3288 => x"24973882",
          3289 => x"d6e408e4",
          3290 => x"052270f7",
          3291 => x"06515372",
          3292 => x"82d6e408",
          3293 => x"e405239d",
          3294 => x"3982d6e4",
          3295 => x"08e80533",
          3296 => x"5382d6e4",
          3297 => x"08fc0533",
          3298 => x"73713154",
          3299 => x"547282d6",
          3300 => x"e408e805",
          3301 => x"3482d6e4",
          3302 => x"08e40522",
          3303 => x"70832a70",
          3304 => x"81065151",
          3305 => x"5372802e",
          3306 => x"b13882d6",
          3307 => x"e408e805",
          3308 => x"3370882b",
          3309 => x"70902b70",
          3310 => x"902c7088",
          3311 => x"2c515151",
          3312 => x"51537254",
          3313 => x"82d6e408",
          3314 => x"ec052270",
          3315 => x"75315153",
          3316 => x"7282d6e4",
          3317 => x"08ec0523",
          3318 => x"af3982d6",
          3319 => x"e408fc05",
          3320 => x"3370882b",
          3321 => x"70902b70",
          3322 => x"902c7088",
          3323 => x"2c515151",
          3324 => x"51537254",
          3325 => x"82d6e408",
          3326 => x"ec052270",
          3327 => x"75315153",
          3328 => x"7282d6e4",
          3329 => x"08ec0523",
          3330 => x"82d6e408",
          3331 => x"e4052270",
          3332 => x"83800651",
          3333 => x"5372b038",
          3334 => x"82d6e408",
          3335 => x"ec0522ff",
          3336 => x"11545472",
          3337 => x"82d6e408",
          3338 => x"ec052373",
          3339 => x"902b7090",
          3340 => x"2c515380",
          3341 => x"73259038",
          3342 => x"82d6e408",
          3343 => x"88050852",
          3344 => x"a0518aee",
          3345 => x"3fd23982",
          3346 => x"d6e408e4",
          3347 => x"05227081",
          3348 => x"2a708106",
          3349 => x"51515372",
          3350 => x"802e9138",
          3351 => x"82d6e408",
          3352 => x"88050852",
          3353 => x"ad518aca",
          3354 => x"3f80c739",
          3355 => x"82d6e408",
          3356 => x"e4052270",
          3357 => x"842a7081",
          3358 => x"06515153",
          3359 => x"72802e90",
          3360 => x"3882d6e4",
          3361 => x"08880508",
          3362 => x"52ab518a",
          3363 => x"a53fa339",
          3364 => x"82d6e408",
          3365 => x"e4052270",
          3366 => x"852a7081",
          3367 => x"06515153",
          3368 => x"72802e8e",
          3369 => x"3882d6e4",
          3370 => x"08880508",
          3371 => x"52a0518a",
          3372 => x"813f82d6",
          3373 => x"e408e405",
          3374 => x"2270862a",
          3375 => x"70810651",
          3376 => x"51537280",
          3377 => x"2eb13882",
          3378 => x"d6e40888",
          3379 => x"050852b0",
          3380 => x"5189df3f",
          3381 => x"82d6e408",
          3382 => x"f4052253",
          3383 => x"72902e09",
          3384 => x"81069438",
          3385 => x"82d6e408",
          3386 => x"88050852",
          3387 => x"82d6e408",
          3388 => x"f8053351",
          3389 => x"89bc3f82",
          3390 => x"d6e408e4",
          3391 => x"05227088",
          3392 => x"2a708106",
          3393 => x"51515372",
          3394 => x"802eb038",
          3395 => x"82d6e408",
          3396 => x"ec0522ff",
          3397 => x"11545472",
          3398 => x"82d6e408",
          3399 => x"ec052373",
          3400 => x"902b7090",
          3401 => x"2c515380",
          3402 => x"73259038",
          3403 => x"82d6e408",
          3404 => x"88050852",
          3405 => x"b05188fa",
          3406 => x"3fd23982",
          3407 => x"d6e408e4",
          3408 => x"05227083",
          3409 => x"2a708106",
          3410 => x"51515372",
          3411 => x"802eb038",
          3412 => x"82d6e408",
          3413 => x"e80533ff",
          3414 => x"11545472",
          3415 => x"82d6e408",
          3416 => x"e8053473",
          3417 => x"982b7098",
          3418 => x"2c515380",
          3419 => x"73259038",
          3420 => x"82d6e408",
          3421 => x"88050852",
          3422 => x"b05188b6",
          3423 => x"3fd23982",
          3424 => x"d6e408e4",
          3425 => x"05227087",
          3426 => x"2a708106",
          3427 => x"51515372",
          3428 => x"b03882d6",
          3429 => x"e408ec05",
          3430 => x"22ff1154",
          3431 => x"547282d6",
          3432 => x"e408ec05",
          3433 => x"2373902b",
          3434 => x"70902c51",
          3435 => x"53807325",
          3436 => x"903882d6",
          3437 => x"e4088805",
          3438 => x"0852a051",
          3439 => x"87f43fd2",
          3440 => x"3982d6e4",
          3441 => x"08f80533",
          3442 => x"537280e3",
          3443 => x"2e098106",
          3444 => x"973882d6",
          3445 => x"e4088805",
          3446 => x"085282d6",
          3447 => x"e408fc05",
          3448 => x"335187ce",
          3449 => x"3f81ee39",
          3450 => x"82d6e408",
          3451 => x"f8053353",
          3452 => x"7280f32e",
          3453 => x"09810680",
          3454 => x"cb3882d6",
          3455 => x"e408f405",
          3456 => x"22ff1151",
          3457 => x"537282d6",
          3458 => x"e408f405",
          3459 => x"237283ff",
          3460 => x"ff065372",
          3461 => x"83ffff2e",
          3462 => x"81bb3882",
          3463 => x"d6e40888",
          3464 => x"05085282",
          3465 => x"d6e408fc",
          3466 => x"05087033",
          3467 => x"5282d6e4",
          3468 => x"08fc0508",
          3469 => x"810582d6",
          3470 => x"e408fc05",
          3471 => x"0c5386f2",
          3472 => x"3fffb739",
          3473 => x"82d6e408",
          3474 => x"f8053353",
          3475 => x"7280d32e",
          3476 => x"09810680",
          3477 => x"cb3882d6",
          3478 => x"e408f405",
          3479 => x"22ff1151",
          3480 => x"537282d6",
          3481 => x"e408f405",
          3482 => x"237283ff",
          3483 => x"ff065372",
          3484 => x"83ffff2e",
          3485 => x"80df3882",
          3486 => x"d6e40888",
          3487 => x"05085282",
          3488 => x"d6e408fc",
          3489 => x"05087033",
          3490 => x"525386a6",
          3491 => x"3f82d6e4",
          3492 => x"08fc0508",
          3493 => x"810582d6",
          3494 => x"e408fc05",
          3495 => x"0cffb739",
          3496 => x"82d6e408",
          3497 => x"f0050882",
          3498 => x"d6e82ea9",
          3499 => x"3882d6e4",
          3500 => x"08880508",
          3501 => x"5282d6e4",
          3502 => x"08f00508",
          3503 => x"ff0582d6",
          3504 => x"e408f005",
          3505 => x"0c82d6e4",
          3506 => x"08f00508",
          3507 => x"70335253",
          3508 => x"85e03fcc",
          3509 => x"3982d6e4",
          3510 => x"08e40522",
          3511 => x"70872a70",
          3512 => x"81065151",
          3513 => x"5372802e",
          3514 => x"80c33882",
          3515 => x"d6e408ec",
          3516 => x"0522ff11",
          3517 => x"54547282",
          3518 => x"d6e408ec",
          3519 => x"05237390",
          3520 => x"2b70902c",
          3521 => x"51538073",
          3522 => x"25a33882",
          3523 => x"d6e40888",
          3524 => x"050852a0",
          3525 => x"51859b3f",
          3526 => x"d23982d6",
          3527 => x"e4088805",
          3528 => x"085282d6",
          3529 => x"e408f805",
          3530 => x"33518586",
          3531 => x"3f800b82",
          3532 => x"d6e408e4",
          3533 => x"0523eab7",
          3534 => x"3982d6e4",
          3535 => x"08f80533",
          3536 => x"5372a52e",
          3537 => x"098106a8",
          3538 => x"38810b82",
          3539 => x"d6e408e4",
          3540 => x"0523800b",
          3541 => x"82d6e408",
          3542 => x"ec052380",
          3543 => x"0b82d6e4",
          3544 => x"08e80534",
          3545 => x"8a0b82d6",
          3546 => x"e408f405",
          3547 => x"23ea8039",
          3548 => x"82d6e408",
          3549 => x"88050852",
          3550 => x"82d6e408",
          3551 => x"f8053351",
          3552 => x"84b03fe9",
          3553 => x"ea3982d6",
          3554 => x"e4088805",
          3555 => x"088c1108",
          3556 => x"7082d6e4",
          3557 => x"08e0050c",
          3558 => x"515382d6",
          3559 => x"e408e005",
          3560 => x"0882d6d8",
          3561 => x"0c953d0d",
          3562 => x"82d6e40c",
          3563 => x"0482d6e4",
          3564 => x"080282d6",
          3565 => x"e40cfd3d",
          3566 => x"0d82f2b8",
          3567 => x"085382d6",
          3568 => x"e4088c05",
          3569 => x"085282d6",
          3570 => x"e4088805",
          3571 => x"0851e4dd",
          3572 => x"3f82d6d8",
          3573 => x"087082d6",
          3574 => x"d80c5485",
          3575 => x"3d0d82d6",
          3576 => x"e40c0482",
          3577 => x"d6e40802",
          3578 => x"82d6e40c",
          3579 => x"fb3d0d80",
          3580 => x"0b82d6e4",
          3581 => x"08f8050c",
          3582 => x"82f2bc08",
          3583 => x"85113370",
          3584 => x"812a7081",
          3585 => x"32708106",
          3586 => x"51515151",
          3587 => x"5372802e",
          3588 => x"8d38ff0b",
          3589 => x"82d6e408",
          3590 => x"f4050c81",
          3591 => x"923982d6",
          3592 => x"e4088805",
          3593 => x"08537233",
          3594 => x"82d6e408",
          3595 => x"88050881",
          3596 => x"0582d6e4",
          3597 => x"0888050c",
          3598 => x"537282d6",
          3599 => x"e408fc05",
          3600 => x"347281ff",
          3601 => x"06537280",
          3602 => x"2eb03882",
          3603 => x"f2bc0882",
          3604 => x"f2bc0853",
          3605 => x"82d6e408",
          3606 => x"fc053352",
          3607 => x"90110851",
          3608 => x"53722d82",
          3609 => x"d6d80853",
          3610 => x"72802eff",
          3611 => x"b138ff0b",
          3612 => x"82d6e408",
          3613 => x"f8050cff",
          3614 => x"a53982f2",
          3615 => x"bc0882f2",
          3616 => x"bc085353",
          3617 => x"8a519013",
          3618 => x"0853722d",
          3619 => x"82d6d808",
          3620 => x"5372802e",
          3621 => x"8a38ff0b",
          3622 => x"82d6e408",
          3623 => x"f8050c82",
          3624 => x"d6e408f8",
          3625 => x"05087082",
          3626 => x"d6e408f4",
          3627 => x"050c5382",
          3628 => x"d6e408f4",
          3629 => x"050882d6",
          3630 => x"d80c873d",
          3631 => x"0d82d6e4",
          3632 => x"0c0482d6",
          3633 => x"e4080282",
          3634 => x"d6e40cfb",
          3635 => x"3d0d800b",
          3636 => x"82d6e408",
          3637 => x"f8050c82",
          3638 => x"d6e4088c",
          3639 => x"05088511",
          3640 => x"3370812a",
          3641 => x"70813270",
          3642 => x"81065151",
          3643 => x"51515372",
          3644 => x"802e8d38",
          3645 => x"ff0b82d6",
          3646 => x"e408f405",
          3647 => x"0c80f339",
          3648 => x"82d6e408",
          3649 => x"88050853",
          3650 => x"723382d6",
          3651 => x"e4088805",
          3652 => x"08810582",
          3653 => x"d6e40888",
          3654 => x"050c5372",
          3655 => x"82d6e408",
          3656 => x"fc053472",
          3657 => x"81ff0653",
          3658 => x"72802eb6",
          3659 => x"3882d6e4",
          3660 => x"088c0508",
          3661 => x"82d6e408",
          3662 => x"8c050853",
          3663 => x"82d6e408",
          3664 => x"fc053352",
          3665 => x"90110851",
          3666 => x"53722d82",
          3667 => x"d6d80853",
          3668 => x"72802eff",
          3669 => x"ab38ff0b",
          3670 => x"82d6e408",
          3671 => x"f8050cff",
          3672 => x"9f3982d6",
          3673 => x"e408f805",
          3674 => x"087082d6",
          3675 => x"e408f405",
          3676 => x"0c5382d6",
          3677 => x"e408f405",
          3678 => x"0882d6d8",
          3679 => x"0c873d0d",
          3680 => x"82d6e40c",
          3681 => x"0482d6e4",
          3682 => x"080282d6",
          3683 => x"e40cfe3d",
          3684 => x"0d82f2bc",
          3685 => x"085282d6",
          3686 => x"e4088805",
          3687 => x"0851933f",
          3688 => x"82d6d808",
          3689 => x"7082d6d8",
          3690 => x"0c53843d",
          3691 => x"0d82d6e4",
          3692 => x"0c0482d6",
          3693 => x"e4080282",
          3694 => x"d6e40cfb",
          3695 => x"3d0d82d6",
          3696 => x"e4088c05",
          3697 => x"08851133",
          3698 => x"70812a70",
          3699 => x"81327081",
          3700 => x"06515151",
          3701 => x"51537280",
          3702 => x"2e8d38ff",
          3703 => x"0b82d6e4",
          3704 => x"08fc050c",
          3705 => x"81cb3982",
          3706 => x"d6e4088c",
          3707 => x"05088511",
          3708 => x"3370822a",
          3709 => x"70810651",
          3710 => x"51515372",
          3711 => x"802e80db",
          3712 => x"3882d6e4",
          3713 => x"088c0508",
          3714 => x"82d6e408",
          3715 => x"8c050854",
          3716 => x"548c1408",
          3717 => x"88140825",
          3718 => x"9f3882d6",
          3719 => x"e4088c05",
          3720 => x"08700870",
          3721 => x"82d6e408",
          3722 => x"88050852",
          3723 => x"57545472",
          3724 => x"75347308",
          3725 => x"8105740c",
          3726 => x"82d6e408",
          3727 => x"8c05088c",
          3728 => x"11088105",
          3729 => x"8c120c82",
          3730 => x"d6e40888",
          3731 => x"05087082",
          3732 => x"d6e408fc",
          3733 => x"050c5153",
          3734 => x"80d73982",
          3735 => x"d6e4088c",
          3736 => x"050882d6",
          3737 => x"e4088c05",
          3738 => x"085382d6",
          3739 => x"e4088805",
          3740 => x"087081ff",
          3741 => x"06539012",
          3742 => x"08515454",
          3743 => x"722d82d6",
          3744 => x"d8085372",
          3745 => x"a33882d6",
          3746 => x"e4088c05",
          3747 => x"088c1108",
          3748 => x"81058c12",
          3749 => x"0c82d6e4",
          3750 => x"08880508",
          3751 => x"7082d6e4",
          3752 => x"08fc050c",
          3753 => x"51538a39",
          3754 => x"ff0b82d6",
          3755 => x"e408fc05",
          3756 => x"0c82d6e4",
          3757 => x"08fc0508",
          3758 => x"82d6d80c",
          3759 => x"873d0d82",
          3760 => x"d6e40c04",
          3761 => x"82d6e408",
          3762 => x"0282d6e4",
          3763 => x"0cf93d0d",
          3764 => x"82d6e408",
          3765 => x"88050885",
          3766 => x"11337081",
          3767 => x"32708106",
          3768 => x"51515152",
          3769 => x"71802e8d",
          3770 => x"38ff0b82",
          3771 => x"d6e408f8",
          3772 => x"050c8394",
          3773 => x"3982d6e4",
          3774 => x"08880508",
          3775 => x"85113370",
          3776 => x"862a7081",
          3777 => x"06515151",
          3778 => x"5271802e",
          3779 => x"80c53882",
          3780 => x"d6e40888",
          3781 => x"050882d6",
          3782 => x"e4088805",
          3783 => x"08535385",
          3784 => x"123370ff",
          3785 => x"bf065152",
          3786 => x"71851434",
          3787 => x"82d6e408",
          3788 => x"8805088c",
          3789 => x"11088105",
          3790 => x"8c120c82",
          3791 => x"d6e40888",
          3792 => x"05088411",
          3793 => x"337082d6",
          3794 => x"e408f805",
          3795 => x"0c515152",
          3796 => x"82b63982",
          3797 => x"d6e40888",
          3798 => x"05088511",
          3799 => x"3370822a",
          3800 => x"70810651",
          3801 => x"51515271",
          3802 => x"802e80d7",
          3803 => x"3882d6e4",
          3804 => x"08880508",
          3805 => x"70087033",
          3806 => x"82d6e408",
          3807 => x"fc050c51",
          3808 => x"5282d6e4",
          3809 => x"08fc0508",
          3810 => x"a93882d6",
          3811 => x"e4088805",
          3812 => x"0882d6e4",
          3813 => x"08880508",
          3814 => x"53538512",
          3815 => x"3370a007",
          3816 => x"51527185",
          3817 => x"1434ff0b",
          3818 => x"82d6e408",
          3819 => x"f8050c81",
          3820 => x"d73982d6",
          3821 => x"e4088805",
          3822 => x"08700881",
          3823 => x"05710c52",
          3824 => x"81a13982",
          3825 => x"d6e40888",
          3826 => x"050882d6",
          3827 => x"e4088805",
          3828 => x"08529411",
          3829 => x"08515271",
          3830 => x"2d82d6d8",
          3831 => x"087082d6",
          3832 => x"e408fc05",
          3833 => x"0c5282d6",
          3834 => x"e408fc05",
          3835 => x"08802580",
          3836 => x"f23882d6",
          3837 => x"e4088805",
          3838 => x"0882d6e4",
          3839 => x"08f4050c",
          3840 => x"82d6e408",
          3841 => x"88050885",
          3842 => x"113382d6",
          3843 => x"e408f005",
          3844 => x"0c5282d6",
          3845 => x"e408fc05",
          3846 => x"08ff2e09",
          3847 => x"81069538",
          3848 => x"82d6e408",
          3849 => x"f0050890",
          3850 => x"07527182",
          3851 => x"d6e408ec",
          3852 => x"05349339",
          3853 => x"82d6e408",
          3854 => x"f00508a0",
          3855 => x"07527182",
          3856 => x"d6e408ec",
          3857 => x"053482d6",
          3858 => x"e408f405",
          3859 => x"085282d6",
          3860 => x"e408ec05",
          3861 => x"33851334",
          3862 => x"ff0b82d6",
          3863 => x"e408f805",
          3864 => x"0ca63982",
          3865 => x"d6e40888",
          3866 => x"05088c11",
          3867 => x"0881058c",
          3868 => x"120c82d6",
          3869 => x"e408fc05",
          3870 => x"087081ff",
          3871 => x"067082d6",
          3872 => x"e408f805",
          3873 => x"0c515152",
          3874 => x"82d6e408",
          3875 => x"f8050882",
          3876 => x"d6d80c89",
          3877 => x"3d0d82d6",
          3878 => x"e40c0482",
          3879 => x"d6e40802",
          3880 => x"82d6e40c",
          3881 => x"fd3d0d82",
          3882 => x"d6e40888",
          3883 => x"050882d6",
          3884 => x"e408fc05",
          3885 => x"0c82d6e4",
          3886 => x"088c0508",
          3887 => x"82d6e408",
          3888 => x"f8050c82",
          3889 => x"d6e40890",
          3890 => x"0508802e",
          3891 => x"82a23882",
          3892 => x"d6e408f8",
          3893 => x"050882d6",
          3894 => x"e408fc05",
          3895 => x"082681ac",
          3896 => x"3882d6e4",
          3897 => x"08f80508",
          3898 => x"82d6e408",
          3899 => x"90050805",
          3900 => x"5182d6e4",
          3901 => x"08fc0508",
          3902 => x"71278190",
          3903 => x"3882d6e4",
          3904 => x"08fc0508",
          3905 => x"82d6e408",
          3906 => x"90050805",
          3907 => x"82d6e408",
          3908 => x"fc050c82",
          3909 => x"d6e408f8",
          3910 => x"050882d6",
          3911 => x"e4089005",
          3912 => x"080582d6",
          3913 => x"e408f805",
          3914 => x"0c82d6e4",
          3915 => x"08900508",
          3916 => x"810582d6",
          3917 => x"e4089005",
          3918 => x"0c82d6e4",
          3919 => x"08900508",
          3920 => x"ff0582d6",
          3921 => x"e4089005",
          3922 => x"0c82d6e4",
          3923 => x"08900508",
          3924 => x"802e819c",
          3925 => x"3882d6e4",
          3926 => x"08fc0508",
          3927 => x"ff0582d6",
          3928 => x"e408fc05",
          3929 => x"0c82d6e4",
          3930 => x"08f80508",
          3931 => x"ff0582d6",
          3932 => x"e408f805",
          3933 => x"0c82d6e4",
          3934 => x"08fc0508",
          3935 => x"82d6e408",
          3936 => x"f8050853",
          3937 => x"51713371",
          3938 => x"34ffae39",
          3939 => x"82d6e408",
          3940 => x"90050881",
          3941 => x"0582d6e4",
          3942 => x"0890050c",
          3943 => x"82d6e408",
          3944 => x"900508ff",
          3945 => x"0582d6e4",
          3946 => x"0890050c",
          3947 => x"82d6e408",
          3948 => x"90050880",
          3949 => x"2eba3882",
          3950 => x"d6e408f8",
          3951 => x"05085170",
          3952 => x"3382d6e4",
          3953 => x"08f80508",
          3954 => x"810582d6",
          3955 => x"e408f805",
          3956 => x"0c82d6e4",
          3957 => x"08fc0508",
          3958 => x"52527171",
          3959 => x"3482d6e4",
          3960 => x"08fc0508",
          3961 => x"810582d6",
          3962 => x"e408fc05",
          3963 => x"0cffad39",
          3964 => x"82d6e408",
          3965 => x"88050870",
          3966 => x"82d6d80c",
          3967 => x"51853d0d",
          3968 => x"82d6e40c",
          3969 => x"0482d6e4",
          3970 => x"080282d6",
          3971 => x"e40cfe3d",
          3972 => x"0d82d6e4",
          3973 => x"08880508",
          3974 => x"82d6e408",
          3975 => x"fc050c82",
          3976 => x"d6e408fc",
          3977 => x"05085271",
          3978 => x"3382d6e4",
          3979 => x"08fc0508",
          3980 => x"810582d6",
          3981 => x"e408fc05",
          3982 => x"0c7081ff",
          3983 => x"06515170",
          3984 => x"802e8338",
          3985 => x"da3982d6",
          3986 => x"e408fc05",
          3987 => x"08ff0582",
          3988 => x"d6e408fc",
          3989 => x"050c82d6",
          3990 => x"e408fc05",
          3991 => x"0882d6e4",
          3992 => x"08880508",
          3993 => x"317082d6",
          3994 => x"d80c5184",
          3995 => x"3d0d82d6",
          3996 => x"e40c0482",
          3997 => x"d6e40802",
          3998 => x"82d6e40c",
          3999 => x"fe3d0d82",
          4000 => x"d6e40888",
          4001 => x"050882d6",
          4002 => x"e408fc05",
          4003 => x"0c82d6e4",
          4004 => x"088c0508",
          4005 => x"52713382",
          4006 => x"d6e4088c",
          4007 => x"05088105",
          4008 => x"82d6e408",
          4009 => x"8c050c82",
          4010 => x"d6e408fc",
          4011 => x"05085351",
          4012 => x"70723482",
          4013 => x"d6e408fc",
          4014 => x"05088105",
          4015 => x"82d6e408",
          4016 => x"fc050c70",
          4017 => x"81ff0651",
          4018 => x"70802e84",
          4019 => x"38ffbe39",
          4020 => x"82d6e408",
          4021 => x"88050870",
          4022 => x"82d6d80c",
          4023 => x"51843d0d",
          4024 => x"82d6e40c",
          4025 => x"0482d6e4",
          4026 => x"080282d6",
          4027 => x"e40cfd3d",
          4028 => x"0d82d6e4",
          4029 => x"08880508",
          4030 => x"82d6e408",
          4031 => x"fc050c82",
          4032 => x"d6e4088c",
          4033 => x"050882d6",
          4034 => x"e408f805",
          4035 => x"0c82d6e4",
          4036 => x"08900508",
          4037 => x"802e80e5",
          4038 => x"3882d6e4",
          4039 => x"08900508",
          4040 => x"810582d6",
          4041 => x"e4089005",
          4042 => x"0c82d6e4",
          4043 => x"08900508",
          4044 => x"ff0582d6",
          4045 => x"e4089005",
          4046 => x"0c82d6e4",
          4047 => x"08900508",
          4048 => x"802eba38",
          4049 => x"82d6e408",
          4050 => x"f8050851",
          4051 => x"703382d6",
          4052 => x"e408f805",
          4053 => x"08810582",
          4054 => x"d6e408f8",
          4055 => x"050c82d6",
          4056 => x"e408fc05",
          4057 => x"08525271",
          4058 => x"713482d6",
          4059 => x"e408fc05",
          4060 => x"08810582",
          4061 => x"d6e408fc",
          4062 => x"050cffad",
          4063 => x"3982d6e4",
          4064 => x"08880508",
          4065 => x"7082d6d8",
          4066 => x"0c51853d",
          4067 => x"0d82d6e4",
          4068 => x"0c0482d6",
          4069 => x"e4080282",
          4070 => x"d6e40cfd",
          4071 => x"3d0d82d6",
          4072 => x"e4089005",
          4073 => x"08802e81",
          4074 => x"f43882d6",
          4075 => x"e4088c05",
          4076 => x"08527133",
          4077 => x"82d6e408",
          4078 => x"8c050881",
          4079 => x"0582d6e4",
          4080 => x"088c050c",
          4081 => x"82d6e408",
          4082 => x"88050870",
          4083 => x"337281ff",
          4084 => x"06535454",
          4085 => x"5171712e",
          4086 => x"843880ce",
          4087 => x"3982d6e4",
          4088 => x"08880508",
          4089 => x"52713382",
          4090 => x"d6e40888",
          4091 => x"05088105",
          4092 => x"82d6e408",
          4093 => x"88050c70",
          4094 => x"81ff0651",
          4095 => x"51708d38",
          4096 => x"800b82d6",
          4097 => x"e408fc05",
          4098 => x"0c819b39",
          4099 => x"82d6e408",
          4100 => x"900508ff",
          4101 => x"0582d6e4",
          4102 => x"0890050c",
          4103 => x"82d6e408",
          4104 => x"90050880",
          4105 => x"2e8438ff",
          4106 => x"813982d6",
          4107 => x"e4089005",
          4108 => x"08802e80",
          4109 => x"e83882d6",
          4110 => x"e4088805",
          4111 => x"08703352",
          4112 => x"53708d38",
          4113 => x"ff0b82d6",
          4114 => x"e408fc05",
          4115 => x"0c80d739",
          4116 => x"82d6e408",
          4117 => x"8c0508ff",
          4118 => x"0582d6e4",
          4119 => x"088c050c",
          4120 => x"82d6e408",
          4121 => x"8c050870",
          4122 => x"33525270",
          4123 => x"8c38810b",
          4124 => x"82d6e408",
          4125 => x"fc050cae",
          4126 => x"3982d6e4",
          4127 => x"08880508",
          4128 => x"703382d6",
          4129 => x"e4088c05",
          4130 => x"08703372",
          4131 => x"71317082",
          4132 => x"d6e408fc",
          4133 => x"050c5355",
          4134 => x"5252538a",
          4135 => x"39800b82",
          4136 => x"d6e408fc",
          4137 => x"050c82d6",
          4138 => x"e408fc05",
          4139 => x"0882d6d8",
          4140 => x"0c853d0d",
          4141 => x"82d6e40c",
          4142 => x"0482d6e4",
          4143 => x"080282d6",
          4144 => x"e40cfa3d",
          4145 => x"0d82d6e4",
          4146 => x"088c0508",
          4147 => x"5282d6e4",
          4148 => x"08880508",
          4149 => x"51818d3f",
          4150 => x"82d6d808",
          4151 => x"7082d6e4",
          4152 => x"08f8050c",
          4153 => x"82d6e408",
          4154 => x"f8050881",
          4155 => x"05705351",
          4156 => x"5480e3f4",
          4157 => x"3f82d6d8",
          4158 => x"087082d6",
          4159 => x"e408fc05",
          4160 => x"0c5482d6",
          4161 => x"e408fc05",
          4162 => x"088c3880",
          4163 => x"0b82d6e4",
          4164 => x"08f4050c",
          4165 => x"bc3982d6",
          4166 => x"e408fc05",
          4167 => x"0882d6e4",
          4168 => x"08f80508",
          4169 => x"05548074",
          4170 => x"3482d6e4",
          4171 => x"08f80508",
          4172 => x"5382d6e4",
          4173 => x"08880508",
          4174 => x"5282d6e4",
          4175 => x"08fc0508",
          4176 => x"51fba23f",
          4177 => x"82d6d808",
          4178 => x"7082d6e4",
          4179 => x"08f4050c",
          4180 => x"5482d6e4",
          4181 => x"08f40508",
          4182 => x"82d6d80c",
          4183 => x"883d0d82",
          4184 => x"d6e40c04",
          4185 => x"82d6e408",
          4186 => x"0282d6e4",
          4187 => x"0cfd3d0d",
          4188 => x"82d6e408",
          4189 => x"88050882",
          4190 => x"d6e408f8",
          4191 => x"050c82d6",
          4192 => x"e4088c05",
          4193 => x"088d3880",
          4194 => x"0b82d6e4",
          4195 => x"08fc050c",
          4196 => x"80ec3982",
          4197 => x"d6e408f8",
          4198 => x"05085271",
          4199 => x"3382d6e4",
          4200 => x"08f80508",
          4201 => x"810582d6",
          4202 => x"e408f805",
          4203 => x"0c7081ff",
          4204 => x"06515170",
          4205 => x"802e9f38",
          4206 => x"82d6e408",
          4207 => x"8c0508ff",
          4208 => x"0582d6e4",
          4209 => x"088c050c",
          4210 => x"82d6e408",
          4211 => x"8c0508ff",
          4212 => x"2e8438ff",
          4213 => x"be3982d6",
          4214 => x"e408f805",
          4215 => x"08ff0582",
          4216 => x"d6e408f8",
          4217 => x"050c82d6",
          4218 => x"e408f805",
          4219 => x"0882d6e4",
          4220 => x"08880508",
          4221 => x"317082d6",
          4222 => x"e408fc05",
          4223 => x"0c5182d6",
          4224 => x"e408fc05",
          4225 => x"0882d6d8",
          4226 => x"0c853d0d",
          4227 => x"82d6e40c",
          4228 => x"0482d6e4",
          4229 => x"080282d6",
          4230 => x"e40cfe3d",
          4231 => x"0d82d6e4",
          4232 => x"08880508",
          4233 => x"82d6e408",
          4234 => x"fc050c82",
          4235 => x"d6e40890",
          4236 => x"0508802e",
          4237 => x"80d43882",
          4238 => x"d6e40890",
          4239 => x"05088105",
          4240 => x"82d6e408",
          4241 => x"90050c82",
          4242 => x"d6e40890",
          4243 => x"0508ff05",
          4244 => x"82d6e408",
          4245 => x"90050c82",
          4246 => x"d6e40890",
          4247 => x"0508802e",
          4248 => x"a93882d6",
          4249 => x"e4088c05",
          4250 => x"08517082",
          4251 => x"d6e408fc",
          4252 => x"05085252",
          4253 => x"71713482",
          4254 => x"d6e408fc",
          4255 => x"05088105",
          4256 => x"82d6e408",
          4257 => x"fc050cff",
          4258 => x"be3982d6",
          4259 => x"e4088805",
          4260 => x"087082d6",
          4261 => x"d80c5184",
          4262 => x"3d0d82d6",
          4263 => x"e40c0482",
          4264 => x"d6e40802",
          4265 => x"82d6e40c",
          4266 => x"f93d0d80",
          4267 => x"0b82d6e4",
          4268 => x"08fc050c",
          4269 => x"82d6e408",
          4270 => x"88050880",
          4271 => x"25b93882",
          4272 => x"d6e40888",
          4273 => x"05083082",
          4274 => x"d6e40888",
          4275 => x"050c800b",
          4276 => x"82d6e408",
          4277 => x"f4050c82",
          4278 => x"d6e408fc",
          4279 => x"05088a38",
          4280 => x"810b82d6",
          4281 => x"e408f405",
          4282 => x"0c82d6e4",
          4283 => x"08f40508",
          4284 => x"82d6e408",
          4285 => x"fc050c82",
          4286 => x"d6e4088c",
          4287 => x"05088025",
          4288 => x"b93882d6",
          4289 => x"e4088c05",
          4290 => x"083082d6",
          4291 => x"e4088c05",
          4292 => x"0c800b82",
          4293 => x"d6e408f0",
          4294 => x"050c82d6",
          4295 => x"e408fc05",
          4296 => x"088a3881",
          4297 => x"0b82d6e4",
          4298 => x"08f0050c",
          4299 => x"82d6e408",
          4300 => x"f0050882",
          4301 => x"d6e408fc",
          4302 => x"050c8053",
          4303 => x"82d6e408",
          4304 => x"8c050852",
          4305 => x"82d6e408",
          4306 => x"88050851",
          4307 => x"82c53f82",
          4308 => x"d6d80870",
          4309 => x"82d6e408",
          4310 => x"f8050c54",
          4311 => x"82d6e408",
          4312 => x"fc050880",
          4313 => x"2e903882",
          4314 => x"d6e408f8",
          4315 => x"05083082",
          4316 => x"d6e408f8",
          4317 => x"050c82d6",
          4318 => x"e408f805",
          4319 => x"087082d6",
          4320 => x"d80c5489",
          4321 => x"3d0d82d6",
          4322 => x"e40c0482",
          4323 => x"d6e40802",
          4324 => x"82d6e40c",
          4325 => x"fb3d0d80",
          4326 => x"0b82d6e4",
          4327 => x"08fc050c",
          4328 => x"82d6e408",
          4329 => x"88050880",
          4330 => x"25993882",
          4331 => x"d6e40888",
          4332 => x"05083082",
          4333 => x"d6e40888",
          4334 => x"050c810b",
          4335 => x"82d6e408",
          4336 => x"fc050c82",
          4337 => x"d6e4088c",
          4338 => x"05088025",
          4339 => x"903882d6",
          4340 => x"e4088c05",
          4341 => x"083082d6",
          4342 => x"e4088c05",
          4343 => x"0c815382",
          4344 => x"d6e4088c",
          4345 => x"05085282",
          4346 => x"d6e40888",
          4347 => x"05085181",
          4348 => x"a23f82d6",
          4349 => x"d8087082",
          4350 => x"d6e408f8",
          4351 => x"050c5482",
          4352 => x"d6e408fc",
          4353 => x"0508802e",
          4354 => x"903882d6",
          4355 => x"e408f805",
          4356 => x"083082d6",
          4357 => x"e408f805",
          4358 => x"0c82d6e4",
          4359 => x"08f80508",
          4360 => x"7082d6d8",
          4361 => x"0c54873d",
          4362 => x"0d82d6e4",
          4363 => x"0c0482d6",
          4364 => x"e4080282",
          4365 => x"d6e40cfd",
          4366 => x"3d0d8053",
          4367 => x"82d6e408",
          4368 => x"8c050852",
          4369 => x"82d6e408",
          4370 => x"88050851",
          4371 => x"80c53f82",
          4372 => x"d6d80870",
          4373 => x"82d6d80c",
          4374 => x"54853d0d",
          4375 => x"82d6e40c",
          4376 => x"0482d6e4",
          4377 => x"080282d6",
          4378 => x"e40cfd3d",
          4379 => x"0d815382",
          4380 => x"d6e4088c",
          4381 => x"05085282",
          4382 => x"d6e40888",
          4383 => x"05085193",
          4384 => x"3f82d6d8",
          4385 => x"087082d6",
          4386 => x"d80c5485",
          4387 => x"3d0d82d6",
          4388 => x"e40c0482",
          4389 => x"d6e40802",
          4390 => x"82d6e40c",
          4391 => x"fd3d0d81",
          4392 => x"0b82d6e4",
          4393 => x"08fc050c",
          4394 => x"800b82d6",
          4395 => x"e408f805",
          4396 => x"0c82d6e4",
          4397 => x"088c0508",
          4398 => x"82d6e408",
          4399 => x"88050827",
          4400 => x"b93882d6",
          4401 => x"e408fc05",
          4402 => x"08802eae",
          4403 => x"38800b82",
          4404 => x"d6e4088c",
          4405 => x"050824a2",
          4406 => x"3882d6e4",
          4407 => x"088c0508",
          4408 => x"1082d6e4",
          4409 => x"088c050c",
          4410 => x"82d6e408",
          4411 => x"fc050810",
          4412 => x"82d6e408",
          4413 => x"fc050cff",
          4414 => x"b83982d6",
          4415 => x"e408fc05",
          4416 => x"08802e80",
          4417 => x"e13882d6",
          4418 => x"e4088c05",
          4419 => x"0882d6e4",
          4420 => x"08880508",
          4421 => x"26ad3882",
          4422 => x"d6e40888",
          4423 => x"050882d6",
          4424 => x"e4088c05",
          4425 => x"083182d6",
          4426 => x"e4088805",
          4427 => x"0c82d6e4",
          4428 => x"08f80508",
          4429 => x"82d6e408",
          4430 => x"fc050807",
          4431 => x"82d6e408",
          4432 => x"f8050c82",
          4433 => x"d6e408fc",
          4434 => x"0508812a",
          4435 => x"82d6e408",
          4436 => x"fc050c82",
          4437 => x"d6e4088c",
          4438 => x"0508812a",
          4439 => x"82d6e408",
          4440 => x"8c050cff",
          4441 => x"953982d6",
          4442 => x"e4089005",
          4443 => x"08802e93",
          4444 => x"3882d6e4",
          4445 => x"08880508",
          4446 => x"7082d6e4",
          4447 => x"08f4050c",
          4448 => x"51913982",
          4449 => x"d6e408f8",
          4450 => x"05087082",
          4451 => x"d6e408f4",
          4452 => x"050c5182",
          4453 => x"d6e408f4",
          4454 => x"050882d6",
          4455 => x"d80c853d",
          4456 => x"0d82d6e4",
          4457 => x"0c0482d6",
          4458 => x"e4080282",
          4459 => x"d6e40cf7",
          4460 => x"3d0d800b",
          4461 => x"82d6e408",
          4462 => x"f0053482",
          4463 => x"d6e4088c",
          4464 => x"05085380",
          4465 => x"730c82d6",
          4466 => x"e4088805",
          4467 => x"08700851",
          4468 => x"53723353",
          4469 => x"7282d6e4",
          4470 => x"08f80534",
          4471 => x"7281ff06",
          4472 => x"5372a02e",
          4473 => x"09810691",
          4474 => x"3882d6e4",
          4475 => x"08880508",
          4476 => x"70088105",
          4477 => x"710c53ce",
          4478 => x"3982d6e4",
          4479 => x"08f80533",
          4480 => x"5372ad2e",
          4481 => x"098106a4",
          4482 => x"38810b82",
          4483 => x"d6e408f0",
          4484 => x"053482d6",
          4485 => x"e4088805",
          4486 => x"08700881",
          4487 => x"05710c70",
          4488 => x"08515372",
          4489 => x"3382d6e4",
          4490 => x"08f80534",
          4491 => x"82d6e408",
          4492 => x"f8053353",
          4493 => x"72b02e09",
          4494 => x"810681dc",
          4495 => x"3882d6e4",
          4496 => x"08880508",
          4497 => x"70088105",
          4498 => x"710c7008",
          4499 => x"51537233",
          4500 => x"82d6e408",
          4501 => x"f8053482",
          4502 => x"d6e408f8",
          4503 => x"053382d6",
          4504 => x"e408e805",
          4505 => x"0c82d6e4",
          4506 => x"08e80508",
          4507 => x"80e22eb6",
          4508 => x"3882d6e4",
          4509 => x"08e80508",
          4510 => x"80f82e84",
          4511 => x"3880cd39",
          4512 => x"900b82d6",
          4513 => x"e408f405",
          4514 => x"3482d6e4",
          4515 => x"08880508",
          4516 => x"70088105",
          4517 => x"710c7008",
          4518 => x"51537233",
          4519 => x"82d6e408",
          4520 => x"f8053481",
          4521 => x"a439820b",
          4522 => x"82d6e408",
          4523 => x"f4053482",
          4524 => x"d6e40888",
          4525 => x"05087008",
          4526 => x"8105710c",
          4527 => x"70085153",
          4528 => x"723382d6",
          4529 => x"e408f805",
          4530 => x"3480fe39",
          4531 => x"82d6e408",
          4532 => x"f8053353",
          4533 => x"72a0268d",
          4534 => x"38810b82",
          4535 => x"d6e408ec",
          4536 => x"050c8380",
          4537 => x"3982d6e4",
          4538 => x"08f80533",
          4539 => x"53af7327",
          4540 => x"903882d6",
          4541 => x"e408f805",
          4542 => x"335372b9",
          4543 => x"2683388d",
          4544 => x"39800b82",
          4545 => x"d6e408ec",
          4546 => x"050c82d8",
          4547 => x"39880b82",
          4548 => x"d6e408f4",
          4549 => x"0534b239",
          4550 => x"82d6e408",
          4551 => x"f8053353",
          4552 => x"af732790",
          4553 => x"3882d6e4",
          4554 => x"08f80533",
          4555 => x"5372b926",
          4556 => x"83388d39",
          4557 => x"800b82d6",
          4558 => x"e408ec05",
          4559 => x"0c82a539",
          4560 => x"8a0b82d6",
          4561 => x"e408f405",
          4562 => x"34800b82",
          4563 => x"d6e408fc",
          4564 => x"050c82d6",
          4565 => x"e408f805",
          4566 => x"3353a073",
          4567 => x"2781cf38",
          4568 => x"82d6e408",
          4569 => x"f8053353",
          4570 => x"80e07327",
          4571 => x"943882d6",
          4572 => x"e408f805",
          4573 => x"33e01151",
          4574 => x"537282d6",
          4575 => x"e408f805",
          4576 => x"3482d6e4",
          4577 => x"08f80533",
          4578 => x"d0115153",
          4579 => x"7282d6e4",
          4580 => x"08f80534",
          4581 => x"82d6e408",
          4582 => x"f8053353",
          4583 => x"907327ad",
          4584 => x"3882d6e4",
          4585 => x"08f80533",
          4586 => x"f9115153",
          4587 => x"7282d6e4",
          4588 => x"08f80534",
          4589 => x"82d6e408",
          4590 => x"f8053353",
          4591 => x"7289268d",
          4592 => x"38800b82",
          4593 => x"d6e408ec",
          4594 => x"050c8198",
          4595 => x"3982d6e4",
          4596 => x"08f80533",
          4597 => x"82d6e408",
          4598 => x"f4053354",
          4599 => x"54727426",
          4600 => x"8d38800b",
          4601 => x"82d6e408",
          4602 => x"ec050c80",
          4603 => x"f73982d6",
          4604 => x"e408f405",
          4605 => x"337082d6",
          4606 => x"e408fc05",
          4607 => x"082982d6",
          4608 => x"e408f805",
          4609 => x"33701282",
          4610 => x"d6e408fc",
          4611 => x"050c82d6",
          4612 => x"e4088805",
          4613 => x"08700881",
          4614 => x"05710c70",
          4615 => x"08515152",
          4616 => x"55537233",
          4617 => x"82d6e408",
          4618 => x"f80534fe",
          4619 => x"a53982d6",
          4620 => x"e408f005",
          4621 => x"33537280",
          4622 => x"2e903882",
          4623 => x"d6e408fc",
          4624 => x"05083082",
          4625 => x"d6e408fc",
          4626 => x"050c82d6",
          4627 => x"e4088c05",
          4628 => x"0882d6e4",
          4629 => x"08fc0508",
          4630 => x"710c5381",
          4631 => x"0b82d6e4",
          4632 => x"08ec050c",
          4633 => x"82d6e408",
          4634 => x"ec050882",
          4635 => x"d6d80c8b",
          4636 => x"3d0d82d6",
          4637 => x"e40c0482",
          4638 => x"d6e40802",
          4639 => x"82d6e40c",
          4640 => x"f73d0d80",
          4641 => x"0b82d6e4",
          4642 => x"08f00534",
          4643 => x"82d6e408",
          4644 => x"8c050853",
          4645 => x"80730c82",
          4646 => x"d6e40888",
          4647 => x"05087008",
          4648 => x"51537233",
          4649 => x"537282d6",
          4650 => x"e408f805",
          4651 => x"347281ff",
          4652 => x"065372a0",
          4653 => x"2e098106",
          4654 => x"913882d6",
          4655 => x"e4088805",
          4656 => x"08700881",
          4657 => x"05710c53",
          4658 => x"ce3982d6",
          4659 => x"e408f805",
          4660 => x"335372ad",
          4661 => x"2e098106",
          4662 => x"a438810b",
          4663 => x"82d6e408",
          4664 => x"f0053482",
          4665 => x"d6e40888",
          4666 => x"05087008",
          4667 => x"8105710c",
          4668 => x"70085153",
          4669 => x"723382d6",
          4670 => x"e408f805",
          4671 => x"3482d6e4",
          4672 => x"08f80533",
          4673 => x"5372b02e",
          4674 => x"09810681",
          4675 => x"dc3882d6",
          4676 => x"e4088805",
          4677 => x"08700881",
          4678 => x"05710c70",
          4679 => x"08515372",
          4680 => x"3382d6e4",
          4681 => x"08f80534",
          4682 => x"82d6e408",
          4683 => x"f8053382",
          4684 => x"d6e408e8",
          4685 => x"050c82d6",
          4686 => x"e408e805",
          4687 => x"0880e22e",
          4688 => x"b63882d6",
          4689 => x"e408e805",
          4690 => x"0880f82e",
          4691 => x"843880cd",
          4692 => x"39900b82",
          4693 => x"d6e408f4",
          4694 => x"053482d6",
          4695 => x"e4088805",
          4696 => x"08700881",
          4697 => x"05710c70",
          4698 => x"08515372",
          4699 => x"3382d6e4",
          4700 => x"08f80534",
          4701 => x"81a43982",
          4702 => x"0b82d6e4",
          4703 => x"08f40534",
          4704 => x"82d6e408",
          4705 => x"88050870",
          4706 => x"08810571",
          4707 => x"0c700851",
          4708 => x"53723382",
          4709 => x"d6e408f8",
          4710 => x"053480fe",
          4711 => x"3982d6e4",
          4712 => x"08f80533",
          4713 => x"5372a026",
          4714 => x"8d38810b",
          4715 => x"82d6e408",
          4716 => x"ec050c83",
          4717 => x"803982d6",
          4718 => x"e408f805",
          4719 => x"3353af73",
          4720 => x"27903882",
          4721 => x"d6e408f8",
          4722 => x"05335372",
          4723 => x"b9268338",
          4724 => x"8d39800b",
          4725 => x"82d6e408",
          4726 => x"ec050c82",
          4727 => x"d839880b",
          4728 => x"82d6e408",
          4729 => x"f40534b2",
          4730 => x"3982d6e4",
          4731 => x"08f80533",
          4732 => x"53af7327",
          4733 => x"903882d6",
          4734 => x"e408f805",
          4735 => x"335372b9",
          4736 => x"2683388d",
          4737 => x"39800b82",
          4738 => x"d6e408ec",
          4739 => x"050c82a5",
          4740 => x"398a0b82",
          4741 => x"d6e408f4",
          4742 => x"0534800b",
          4743 => x"82d6e408",
          4744 => x"fc050c82",
          4745 => x"d6e408f8",
          4746 => x"053353a0",
          4747 => x"732781cf",
          4748 => x"3882d6e4",
          4749 => x"08f80533",
          4750 => x"5380e073",
          4751 => x"27943882",
          4752 => x"d6e408f8",
          4753 => x"0533e011",
          4754 => x"51537282",
          4755 => x"d6e408f8",
          4756 => x"053482d6",
          4757 => x"e408f805",
          4758 => x"33d01151",
          4759 => x"537282d6",
          4760 => x"e408f805",
          4761 => x"3482d6e4",
          4762 => x"08f80533",
          4763 => x"53907327",
          4764 => x"ad3882d6",
          4765 => x"e408f805",
          4766 => x"33f91151",
          4767 => x"537282d6",
          4768 => x"e408f805",
          4769 => x"3482d6e4",
          4770 => x"08f80533",
          4771 => x"53728926",
          4772 => x"8d38800b",
          4773 => x"82d6e408",
          4774 => x"ec050c81",
          4775 => x"983982d6",
          4776 => x"e408f805",
          4777 => x"3382d6e4",
          4778 => x"08f40533",
          4779 => x"54547274",
          4780 => x"268d3880",
          4781 => x"0b82d6e4",
          4782 => x"08ec050c",
          4783 => x"80f73982",
          4784 => x"d6e408f4",
          4785 => x"05337082",
          4786 => x"d6e408fc",
          4787 => x"05082982",
          4788 => x"d6e408f8",
          4789 => x"05337012",
          4790 => x"82d6e408",
          4791 => x"fc050c82",
          4792 => x"d6e40888",
          4793 => x"05087008",
          4794 => x"8105710c",
          4795 => x"70085151",
          4796 => x"52555372",
          4797 => x"3382d6e4",
          4798 => x"08f80534",
          4799 => x"fea53982",
          4800 => x"d6e408f0",
          4801 => x"05335372",
          4802 => x"802e9038",
          4803 => x"82d6e408",
          4804 => x"fc050830",
          4805 => x"82d6e408",
          4806 => x"fc050c82",
          4807 => x"d6e4088c",
          4808 => x"050882d6",
          4809 => x"e408fc05",
          4810 => x"08710c53",
          4811 => x"810b82d6",
          4812 => x"e408ec05",
          4813 => x"0c82d6e4",
          4814 => x"08ec0508",
          4815 => x"82d6d80c",
          4816 => x"8b3d0d82",
          4817 => x"d6e40c04",
          4818 => x"f83d0d7a",
          4819 => x"70087056",
          4820 => x"56597480",
          4821 => x"2e80df38",
          4822 => x"8c397715",
          4823 => x"790c8516",
          4824 => x"335480d2",
          4825 => x"39743354",
          4826 => x"73a02e09",
          4827 => x"81068638",
          4828 => x"811555f1",
          4829 => x"39805776",
          4830 => x"902982d0",
          4831 => x"cc057008",
          4832 => x"5256e581",
          4833 => x"3f82d6d8",
          4834 => x"0882d6d8",
          4835 => x"08547553",
          4836 => x"76085258",
          4837 => x"e7fc3f82",
          4838 => x"d6d8088b",
          4839 => x"38841633",
          4840 => x"5473812e",
          4841 => x"ffb43881",
          4842 => x"177081ff",
          4843 => x"06585499",
          4844 => x"7727c438",
          4845 => x"ff547382",
          4846 => x"d6d80c8a",
          4847 => x"3d0d04ff",
          4848 => x"3d0d7352",
          4849 => x"71932681",
          4850 => x"8e387184",
          4851 => x"2982acdc",
          4852 => x"05527108",
          4853 => x"0482b2cc",
          4854 => x"51818039",
          4855 => x"82b2d851",
          4856 => x"80f93982",
          4857 => x"b2e85180",
          4858 => x"f23982b2",
          4859 => x"f85180eb",
          4860 => x"3982b388",
          4861 => x"5180e439",
          4862 => x"82b39851",
          4863 => x"80dd3982",
          4864 => x"b3ac5180",
          4865 => x"d63982b3",
          4866 => x"bc5180cf",
          4867 => x"3982b3d4",
          4868 => x"5180c839",
          4869 => x"82b3ec51",
          4870 => x"80c13982",
          4871 => x"b48451bb",
          4872 => x"3982b4a0",
          4873 => x"51b53982",
          4874 => x"b4b451af",
          4875 => x"3982b4dc",
          4876 => x"51a93982",
          4877 => x"b4ec51a3",
          4878 => x"3982b58c",
          4879 => x"519d3982",
          4880 => x"b59c5197",
          4881 => x"3982b5b4",
          4882 => x"51913982",
          4883 => x"b5cc518b",
          4884 => x"3982b5e4",
          4885 => x"51853982",
          4886 => x"b5f051d7",
          4887 => x"863f833d",
          4888 => x"0d04fb3d",
          4889 => x"0d777956",
          4890 => x"567487e7",
          4891 => x"268a3874",
          4892 => x"527587e8",
          4893 => x"29519039",
          4894 => x"87e85274",
          4895 => x"51efaf3f",
          4896 => x"82d6d808",
          4897 => x"527551ef",
          4898 => x"a53f82d6",
          4899 => x"d8085479",
          4900 => x"53755282",
          4901 => x"b68051ff",
          4902 => x"babe3f87",
          4903 => x"3d0d04ec",
          4904 => x"3d0d6602",
          4905 => x"840580e3",
          4906 => x"05335b57",
          4907 => x"80687830",
          4908 => x"707a0773",
          4909 => x"25515759",
          4910 => x"59785677",
          4911 => x"87ff2683",
          4912 => x"38815674",
          4913 => x"76077081",
          4914 => x"ff065155",
          4915 => x"93567481",
          4916 => x"82388153",
          4917 => x"76528c3d",
          4918 => x"70525681",
          4919 => x"92cf3f82",
          4920 => x"d6d80857",
          4921 => x"82d6d808",
          4922 => x"b93882d6",
          4923 => x"d80887c0",
          4924 => x"98880c82",
          4925 => x"d6d80859",
          4926 => x"963dd405",
          4927 => x"54848053",
          4928 => x"77527551",
          4929 => x"81978b3f",
          4930 => x"82d6d808",
          4931 => x"5782d6d8",
          4932 => x"0890387a",
          4933 => x"5574802e",
          4934 => x"89387419",
          4935 => x"75195959",
          4936 => x"d739963d",
          4937 => x"d8055181",
          4938 => x"9f823f76",
          4939 => x"30707807",
          4940 => x"80257b30",
          4941 => x"709f2a72",
          4942 => x"06515751",
          4943 => x"5674802e",
          4944 => x"903882b6",
          4945 => x"a45387c0",
          4946 => x"98880852",
          4947 => x"7851fe92",
          4948 => x"3f765675",
          4949 => x"82d6d80c",
          4950 => x"963d0d04",
          4951 => x"f73d0d7d",
          4952 => x"028405bb",
          4953 => x"0533595a",
          4954 => x"ff598053",
          4955 => x"7c527b51",
          4956 => x"fead3f82",
          4957 => x"d6d80880",
          4958 => x"cb387780",
          4959 => x"2e883877",
          4960 => x"812ebf38",
          4961 => x"bf3982f2",
          4962 => x"b85782f2",
          4963 => x"b85682f2",
          4964 => x"b85582f2",
          4965 => x"c0085482",
          4966 => x"f2bc0853",
          4967 => x"82f2b808",
          4968 => x"5282b6ac",
          4969 => x"51ffb8b0",
          4970 => x"3f82f2b8",
          4971 => x"56625561",
          4972 => x"5482d6d8",
          4973 => x"5360527f",
          4974 => x"51792d82",
          4975 => x"d6d80859",
          4976 => x"83397904",
          4977 => x"7882d6d8",
          4978 => x"0c8b3d0d",
          4979 => x"04f33d0d",
          4980 => x"7f616302",
          4981 => x"8c0580cf",
          4982 => x"05337373",
          4983 => x"1568415f",
          4984 => x"5c5c5e5e",
          4985 => x"5e7a5282",
          4986 => x"b6e051ff",
          4987 => x"b7ea3f82",
          4988 => x"b6e851ff",
          4989 => x"b7e23f80",
          4990 => x"55747927",
          4991 => x"8180387b",
          4992 => x"902e8938",
          4993 => x"7ba02ea7",
          4994 => x"3880c639",
          4995 => x"74185372",
          4996 => x"7a278e38",
          4997 => x"72225282",
          4998 => x"b6ec51ff",
          4999 => x"b7ba3f89",
          5000 => x"3982b6f8",
          5001 => x"51ffb7b0",
          5002 => x"3f821555",
          5003 => x"80c33974",
          5004 => x"1853727a",
          5005 => x"278e3872",
          5006 => x"085282b6",
          5007 => x"e051ffb7",
          5008 => x"973f8939",
          5009 => x"82b6f451",
          5010 => x"ffb78d3f",
          5011 => x"841555a1",
          5012 => x"39741853",
          5013 => x"727a278e",
          5014 => x"38723352",
          5015 => x"82b78051",
          5016 => x"ffb6f53f",
          5017 => x"893982b7",
          5018 => x"8851ffb6",
          5019 => x"eb3f8115",
          5020 => x"5582f2bc",
          5021 => x"0852a051",
          5022 => x"d6b83ffe",
          5023 => x"fc3982b7",
          5024 => x"8c51ffb6",
          5025 => x"d33f8055",
          5026 => x"74792780",
          5027 => x"c6387418",
          5028 => x"70335553",
          5029 => x"8056727a",
          5030 => x"27833881",
          5031 => x"5680539f",
          5032 => x"74278338",
          5033 => x"81537573",
          5034 => x"067081ff",
          5035 => x"06515372",
          5036 => x"802e9038",
          5037 => x"7380fe26",
          5038 => x"8a3882f2",
          5039 => x"bc085273",
          5040 => x"51883982",
          5041 => x"f2bc0852",
          5042 => x"a051d5e6",
          5043 => x"3f811555",
          5044 => x"ffb63982",
          5045 => x"b79051d2",
          5046 => x"8a3f7818",
          5047 => x"791c5c58",
          5048 => x"9ce73f82",
          5049 => x"d6d80898",
          5050 => x"2b70982c",
          5051 => x"515776a0",
          5052 => x"2e098106",
          5053 => x"aa389cd1",
          5054 => x"3f82d6d8",
          5055 => x"08982b70",
          5056 => x"982c70a0",
          5057 => x"32703072",
          5058 => x"9b327030",
          5059 => x"70720773",
          5060 => x"75070651",
          5061 => x"58585957",
          5062 => x"51578073",
          5063 => x"24d83876",
          5064 => x"9b2e0981",
          5065 => x"06853880",
          5066 => x"538c397c",
          5067 => x"1e537278",
          5068 => x"26fdb238",
          5069 => x"ff537282",
          5070 => x"d6d80c8f",
          5071 => x"3d0d04fc",
          5072 => x"3d0d029b",
          5073 => x"053382b7",
          5074 => x"945382b7",
          5075 => x"985255ff",
          5076 => x"b5863f82",
          5077 => x"d4a42251",
          5078 => x"a5c03f82",
          5079 => x"b7a45482",
          5080 => x"b7b05382",
          5081 => x"d4a53352",
          5082 => x"82b7b851",
          5083 => x"ffb4e93f",
          5084 => x"74802e84",
          5085 => x"38a0f43f",
          5086 => x"863d0d04",
          5087 => x"fe3d0d87",
          5088 => x"c0968008",
          5089 => x"53a5dc3f",
          5090 => x"815199bd",
          5091 => x"3f82b7d4",
          5092 => x"5199ce3f",
          5093 => x"805199b1",
          5094 => x"3f72812a",
          5095 => x"70810651",
          5096 => x"5271802e",
          5097 => x"92388151",
          5098 => x"999f3f82",
          5099 => x"b7ec5199",
          5100 => x"b03f8051",
          5101 => x"99933f72",
          5102 => x"822a7081",
          5103 => x"06515271",
          5104 => x"802e9238",
          5105 => x"81519981",
          5106 => x"3f82b7fc",
          5107 => x"5199923f",
          5108 => x"805198f5",
          5109 => x"3f72832a",
          5110 => x"70810651",
          5111 => x"5271802e",
          5112 => x"92388151",
          5113 => x"98e33f82",
          5114 => x"b88c5198",
          5115 => x"f43f8051",
          5116 => x"98d73f72",
          5117 => x"842a7081",
          5118 => x"06515271",
          5119 => x"802e9238",
          5120 => x"815198c5",
          5121 => x"3f82b8a0",
          5122 => x"5198d63f",
          5123 => x"805198b9",
          5124 => x"3f72852a",
          5125 => x"70810651",
          5126 => x"5271802e",
          5127 => x"92388151",
          5128 => x"98a73f82",
          5129 => x"b8b45198",
          5130 => x"b83f8051",
          5131 => x"989b3f72",
          5132 => x"862a7081",
          5133 => x"06515271",
          5134 => x"802e9238",
          5135 => x"81519889",
          5136 => x"3f82b8c8",
          5137 => x"51989a3f",
          5138 => x"805197fd",
          5139 => x"3f72872a",
          5140 => x"70810651",
          5141 => x"5271802e",
          5142 => x"92388151",
          5143 => x"97eb3f82",
          5144 => x"b8dc5197",
          5145 => x"fc3f8051",
          5146 => x"97df3f72",
          5147 => x"882a7081",
          5148 => x"06515271",
          5149 => x"802e9238",
          5150 => x"815197cd",
          5151 => x"3f82b8f0",
          5152 => x"5197de3f",
          5153 => x"805197c1",
          5154 => x"3fa3e03f",
          5155 => x"843d0d04",
          5156 => x"fb3d0d77",
          5157 => x"028405a3",
          5158 => x"05337055",
          5159 => x"56568052",
          5160 => x"7551e2ed",
          5161 => x"3f0b0b82",
          5162 => x"d0c83354",
          5163 => x"73a93881",
          5164 => x"5382b9ac",
          5165 => x"5282ede8",
          5166 => x"51818af1",
          5167 => x"3f82d6d8",
          5168 => x"08307082",
          5169 => x"d6d80807",
          5170 => x"80258271",
          5171 => x"31515154",
          5172 => x"730b0b82",
          5173 => x"d0c8340b",
          5174 => x"0b82d0c8",
          5175 => x"33547381",
          5176 => x"2e098106",
          5177 => x"af3882ed",
          5178 => x"e8537452",
          5179 => x"755181c5",
          5180 => x"c13f82d6",
          5181 => x"d808802e",
          5182 => x"8b3882d6",
          5183 => x"d80851cd",
          5184 => x"e23f9139",
          5185 => x"82ede851",
          5186 => x"8197a13f",
          5187 => x"820b0b0b",
          5188 => x"82d0c834",
          5189 => x"0b0b82d0",
          5190 => x"c8335473",
          5191 => x"822e0981",
          5192 => x"068c3882",
          5193 => x"b9bc5374",
          5194 => x"527551a9",
          5195 => x"d83f800b",
          5196 => x"82d6d80c",
          5197 => x"873d0d04",
          5198 => x"cd3d0d80",
          5199 => x"70415eff",
          5200 => x"7e82ede4",
          5201 => x"0c5f8152",
          5202 => x"7d5180c8",
          5203 => x"883f82d6",
          5204 => x"d80881ff",
          5205 => x"0659787e",
          5206 => x"2e098106",
          5207 => x"a338973d",
          5208 => x"59835382",
          5209 => x"b9c45278",
          5210 => x"51dafa3f",
          5211 => x"7d537852",
          5212 => x"82d88451",
          5213 => x"8188d53f",
          5214 => x"82d6d808",
          5215 => x"7e2e8838",
          5216 => x"82b9c851",
          5217 => x"8ddf3981",
          5218 => x"70415e82",
          5219 => x"ba8051ff",
          5220 => x"b0c63f97",
          5221 => x"3d70475a",
          5222 => x"80f85279",
          5223 => x"51fdf13f",
          5224 => x"b53dff84",
          5225 => x"0551f3a0",
          5226 => x"3f82d6d8",
          5227 => x"08902b70",
          5228 => x"902c5159",
          5229 => x"7880c22e",
          5230 => x"87a33878",
          5231 => x"80c224b2",
          5232 => x"3878bd2e",
          5233 => x"81d23878",
          5234 => x"bd249038",
          5235 => x"78802eff",
          5236 => x"ba3878bc",
          5237 => x"2e80da38",
          5238 => x"8ad63978",
          5239 => x"80c02e83",
          5240 => x"99387880",
          5241 => x"c02485cd",
          5242 => x"3878bf2e",
          5243 => x"828c388a",
          5244 => x"bf397880",
          5245 => x"f92e89db",
          5246 => x"387880f9",
          5247 => x"24923878",
          5248 => x"80c32e88",
          5249 => x"8a387880",
          5250 => x"f82e89a3",
          5251 => x"388aa139",
          5252 => x"7881832e",
          5253 => x"8a883878",
          5254 => x"8183248b",
          5255 => x"38788182",
          5256 => x"2e89ed38",
          5257 => x"8a8a3978",
          5258 => x"81852e89",
          5259 => x"fd388a80",
          5260 => x"39b53dff",
          5261 => x"801153ff",
          5262 => x"840551ec",
          5263 => x"ba3f82d6",
          5264 => x"d808802e",
          5265 => x"fec538b5",
          5266 => x"3dfefc11",
          5267 => x"53ff8405",
          5268 => x"51eca43f",
          5269 => x"82d6d808",
          5270 => x"802efeaf",
          5271 => x"38b53dfe",
          5272 => x"f81153ff",
          5273 => x"840551ec",
          5274 => x"8e3f82d6",
          5275 => x"d8088638",
          5276 => x"82d6d808",
          5277 => x"4382ba84",
          5278 => x"51ffaedc",
          5279 => x"3f64645c",
          5280 => x"5a797b27",
          5281 => x"81ec3862",
          5282 => x"59787a70",
          5283 => x"84055c0c",
          5284 => x"7a7a26f5",
          5285 => x"3881db39",
          5286 => x"b53dff80",
          5287 => x"1153ff84",
          5288 => x"0551ebd3",
          5289 => x"3f82d6d8",
          5290 => x"08802efd",
          5291 => x"de38b53d",
          5292 => x"fefc1153",
          5293 => x"ff840551",
          5294 => x"ebbd3f82",
          5295 => x"d6d80880",
          5296 => x"2efdc838",
          5297 => x"b53dfef8",
          5298 => x"1153ff84",
          5299 => x"0551eba7",
          5300 => x"3f82d6d8",
          5301 => x"08802efd",
          5302 => x"b23882ba",
          5303 => x"9451ffad",
          5304 => x"f73f645a",
          5305 => x"79642781",
          5306 => x"89386259",
          5307 => x"79708105",
          5308 => x"5b337934",
          5309 => x"62810543",
          5310 => x"eb39b53d",
          5311 => x"ff801153",
          5312 => x"ff840551",
          5313 => x"eaf13f82",
          5314 => x"d6d80880",
          5315 => x"2efcfc38",
          5316 => x"b53dfefc",
          5317 => x"1153ff84",
          5318 => x"0551eadb",
          5319 => x"3f82d6d8",
          5320 => x"08802efc",
          5321 => x"e638b53d",
          5322 => x"fef81153",
          5323 => x"ff840551",
          5324 => x"eac53f82",
          5325 => x"d6d80880",
          5326 => x"2efcd038",
          5327 => x"82baa051",
          5328 => x"ffad953f",
          5329 => x"645a7964",
          5330 => x"27a83862",
          5331 => x"70337b33",
          5332 => x"5e5a5b78",
          5333 => x"7c2e9238",
          5334 => x"78557a54",
          5335 => x"79335379",
          5336 => x"5282bab0",
          5337 => x"51ffacf0",
          5338 => x"3f811a63",
          5339 => x"8105445a",
          5340 => x"d5398a51",
          5341 => x"cc8f3ffc",
          5342 => x"9239b53d",
          5343 => x"ff801153",
          5344 => x"ff840551",
          5345 => x"e9f13f82",
          5346 => x"d6d80880",
          5347 => x"df3882d4",
          5348 => x"b8335978",
          5349 => x"802e8938",
          5350 => x"82d3f008",
          5351 => x"4580cd39",
          5352 => x"82d4b933",
          5353 => x"5978802e",
          5354 => x"883882d3",
          5355 => x"f80845bc",
          5356 => x"3982d4ba",
          5357 => x"33597880",
          5358 => x"2e883882",
          5359 => x"d4800845",
          5360 => x"ab3982d4",
          5361 => x"bb335978",
          5362 => x"802e8838",
          5363 => x"82d48808",
          5364 => x"459a3982",
          5365 => x"d4b63359",
          5366 => x"78802e88",
          5367 => x"3882d490",
          5368 => x"08458939",
          5369 => x"82d4a008",
          5370 => x"fc800545",
          5371 => x"b53dfefc",
          5372 => x"1153ff84",
          5373 => x"0551e8ff",
          5374 => x"3f82d6d8",
          5375 => x"0880de38",
          5376 => x"82d4b833",
          5377 => x"5978802e",
          5378 => x"893882d3",
          5379 => x"f4084480",
          5380 => x"cc3982d4",
          5381 => x"b9335978",
          5382 => x"802e8838",
          5383 => x"82d3fc08",
          5384 => x"44bb3982",
          5385 => x"d4ba3359",
          5386 => x"78802e88",
          5387 => x"3882d484",
          5388 => x"0844aa39",
          5389 => x"82d4bb33",
          5390 => x"5978802e",
          5391 => x"883882d4",
          5392 => x"8c084499",
          5393 => x"3982d4b6",
          5394 => x"33597880",
          5395 => x"2e883882",
          5396 => x"d4940844",
          5397 => x"883982d4",
          5398 => x"a0088805",
          5399 => x"44b53dfe",
          5400 => x"f81153ff",
          5401 => x"840551e8",
          5402 => x"8e3f82d6",
          5403 => x"d808802e",
          5404 => x"a7388063",
          5405 => x"5c5c7a88",
          5406 => x"2e833881",
          5407 => x"5c7a9032",
          5408 => x"70307072",
          5409 => x"079f2a70",
          5410 => x"7f065151",
          5411 => x"5a5a7880",
          5412 => x"2e88387a",
          5413 => x"a02e8338",
          5414 => x"884382ba",
          5415 => x"cc51c6c3",
          5416 => x"3fa05564",
          5417 => x"54625363",
          5418 => x"526451f2",
          5419 => x"a03f82ba",
          5420 => x"d85187b1",
          5421 => x"39b53dff",
          5422 => x"801153ff",
          5423 => x"840551e7",
          5424 => x"b63f82d6",
          5425 => x"d808802e",
          5426 => x"f9c138b5",
          5427 => x"3dfefc11",
          5428 => x"53ff8405",
          5429 => x"51e7a03f",
          5430 => x"82d6d808",
          5431 => x"802ea438",
          5432 => x"64590280",
          5433 => x"cf053379",
          5434 => x"34648105",
          5435 => x"45b53dfe",
          5436 => x"fc1153ff",
          5437 => x"840551e6",
          5438 => x"fe3f82d6",
          5439 => x"d808e138",
          5440 => x"f9893964",
          5441 => x"70335452",
          5442 => x"82bae451",
          5443 => x"ffa9c93f",
          5444 => x"82f2b808",
          5445 => x"5380f852",
          5446 => x"7951ffaa",
          5447 => x"903f7946",
          5448 => x"79335978",
          5449 => x"ae2ef8e3",
          5450 => x"389f7927",
          5451 => x"9f38b53d",
          5452 => x"fefc1153",
          5453 => x"ff840551",
          5454 => x"e6bd3f82",
          5455 => x"d6d80880",
          5456 => x"2e913864",
          5457 => x"590280cf",
          5458 => x"05337934",
          5459 => x"64810545",
          5460 => x"ffb13982",
          5461 => x"baf051c5",
          5462 => x"8a3fffa7",
          5463 => x"39b53dfe",
          5464 => x"f41153ff",
          5465 => x"840551e0",
          5466 => x"bd3f82d6",
          5467 => x"d808802e",
          5468 => x"f89938b5",
          5469 => x"3dfef011",
          5470 => x"53ff8405",
          5471 => x"51e0a73f",
          5472 => x"82d6d808",
          5473 => x"802ea638",
          5474 => x"61590280",
          5475 => x"c2052279",
          5476 => x"7082055b",
          5477 => x"237842b5",
          5478 => x"3dfef011",
          5479 => x"53ff8405",
          5480 => x"51e0833f",
          5481 => x"82d6d808",
          5482 => x"df38f7df",
          5483 => x"39617022",
          5484 => x"545282ba",
          5485 => x"f451ffa8",
          5486 => x"9f3f82f2",
          5487 => x"b8085380",
          5488 => x"f8527951",
          5489 => x"ffa8e63f",
          5490 => x"79467933",
          5491 => x"5978ae2e",
          5492 => x"f7b93878",
          5493 => x"9f268738",
          5494 => x"61820542",
          5495 => x"d039b53d",
          5496 => x"fef01153",
          5497 => x"ff840551",
          5498 => x"dfbc3f82",
          5499 => x"d6d80880",
          5500 => x"2e933861",
          5501 => x"590280c2",
          5502 => x"05227970",
          5503 => x"82055b23",
          5504 => x"7842ffa9",
          5505 => x"3982baf0",
          5506 => x"51c3d83f",
          5507 => x"ff9f39b5",
          5508 => x"3dfef411",
          5509 => x"53ff8405",
          5510 => x"51df8b3f",
          5511 => x"82d6d808",
          5512 => x"802ef6e7",
          5513 => x"38b53dfe",
          5514 => x"f01153ff",
          5515 => x"840551de",
          5516 => x"f53f82d6",
          5517 => x"d808802e",
          5518 => x"a0386161",
          5519 => x"710c5961",
          5520 => x"840542b5",
          5521 => x"3dfef011",
          5522 => x"53ff8405",
          5523 => x"51ded73f",
          5524 => x"82d6d808",
          5525 => x"e538f6b3",
          5526 => x"39617008",
          5527 => x"545282bb",
          5528 => x"8051ffa6",
          5529 => x"f33f82f2",
          5530 => x"b8085380",
          5531 => x"f8527951",
          5532 => x"ffa7ba3f",
          5533 => x"79467933",
          5534 => x"5978ae2e",
          5535 => x"f68d389f",
          5536 => x"79279b38",
          5537 => x"b53dfef0",
          5538 => x"1153ff84",
          5539 => x"0551de96",
          5540 => x"3f82d6d8",
          5541 => x"08802e8d",
          5542 => x"38616171",
          5543 => x"0c596184",
          5544 => x"0542ffb5",
          5545 => x"3982baf0",
          5546 => x"51c2b83f",
          5547 => x"ffab39b5",
          5548 => x"3dff8011",
          5549 => x"53ff8405",
          5550 => x"51e3bc3f",
          5551 => x"82d6d808",
          5552 => x"802ef5c7",
          5553 => x"38645282",
          5554 => x"bb9051ff",
          5555 => x"a68a3f64",
          5556 => x"597804b5",
          5557 => x"3dff8011",
          5558 => x"53ff8405",
          5559 => x"51e3983f",
          5560 => x"82d6d808",
          5561 => x"802ef5a3",
          5562 => x"38645282",
          5563 => x"bbac51ff",
          5564 => x"a5e63f64",
          5565 => x"59782d82",
          5566 => x"d6d80880",
          5567 => x"2ef58c38",
          5568 => x"82d6d808",
          5569 => x"5282bbc8",
          5570 => x"51ffa5cc",
          5571 => x"3ff4fc39",
          5572 => x"82bbe451",
          5573 => x"c1cd3fff",
          5574 => x"a59f3ff4",
          5575 => x"ee3982bc",
          5576 => x"8051c1bf",
          5577 => x"3f8059ff",
          5578 => x"a83991bf",
          5579 => x"3ff4dc39",
          5580 => x"973d3359",
          5581 => x"78802ef4",
          5582 => x"d23880f8",
          5583 => x"527951d2",
          5584 => x"f83f82d6",
          5585 => x"d8085d82",
          5586 => x"d6d80880",
          5587 => x"2e829238",
          5588 => x"82d6d808",
          5589 => x"46b53dff",
          5590 => x"84055184",
          5591 => x"e53f82d6",
          5592 => x"d808607f",
          5593 => x"065a5c78",
          5594 => x"802e81d2",
          5595 => x"3882d6d8",
          5596 => x"0851cd91",
          5597 => x"3f82d6d8",
          5598 => x"088f2681",
          5599 => x"c138815b",
          5600 => x"7a822eb2",
          5601 => x"387a8224",
          5602 => x"89387a81",
          5603 => x"2e8c3880",
          5604 => x"ca397a83",
          5605 => x"2ead3880",
          5606 => x"c23982bc",
          5607 => x"94567b55",
          5608 => x"82bc9854",
          5609 => x"805382bc",
          5610 => x"9c52b53d",
          5611 => x"ffb00551",
          5612 => x"ffa78d3f",
          5613 => x"b8397b52",
          5614 => x"b53dffb0",
          5615 => x"0551cdb3",
          5616 => x"3fab397b",
          5617 => x"5582bc98",
          5618 => x"54805382",
          5619 => x"bcac52b5",
          5620 => x"3dffb005",
          5621 => x"51ffa6e8",
          5622 => x"3f93397b",
          5623 => x"54805382",
          5624 => x"bcb852b5",
          5625 => x"3dffb005",
          5626 => x"51ffa6d4",
          5627 => x"3f82d3f0",
          5628 => x"5882d788",
          5629 => x"577c5665",
          5630 => x"55805484",
          5631 => x"80805384",
          5632 => x"808052b5",
          5633 => x"3dffb005",
          5634 => x"51ead13f",
          5635 => x"82d6d808",
          5636 => x"82d6d808",
          5637 => x"09703070",
          5638 => x"72078025",
          5639 => x"515b5b5f",
          5640 => x"805a7a83",
          5641 => x"26833881",
          5642 => x"5a787a06",
          5643 => x"5978802e",
          5644 => x"8d38811b",
          5645 => x"7081ff06",
          5646 => x"5c597afe",
          5647 => x"c3387f81",
          5648 => x"327e8132",
          5649 => x"07597889",
          5650 => x"387eff2e",
          5651 => x"09810689",
          5652 => x"3882bcc0",
          5653 => x"51ffbf8b",
          5654 => x"3f7c51b1",
          5655 => x"f53ff2ab",
          5656 => x"3982bcd0",
          5657 => x"51ffbefb",
          5658 => x"3ff2a039",
          5659 => x"f63d0d80",
          5660 => x"0b82d788",
          5661 => x"3487c094",
          5662 => x"8c085387",
          5663 => x"84805272",
          5664 => x"51d7ab3f",
          5665 => x"82d6d808",
          5666 => x"902b87c0",
          5667 => x"948c0855",
          5668 => x"53878480",
          5669 => x"527351d7",
          5670 => x"953f7282",
          5671 => x"d6d80807",
          5672 => x"87c0948c",
          5673 => x"0c87c094",
          5674 => x"9c085387",
          5675 => x"84805272",
          5676 => x"51d6fb3f",
          5677 => x"82d6d808",
          5678 => x"902b87c0",
          5679 => x"949c0855",
          5680 => x"53878480",
          5681 => x"527351d6",
          5682 => x"e53f7282",
          5683 => x"d6d80807",
          5684 => x"87c0949c",
          5685 => x"0c8c8083",
          5686 => x"0b87c094",
          5687 => x"840c8c80",
          5688 => x"830b87c0",
          5689 => x"94940c87",
          5690 => x"a0a08053",
          5691 => x"80737084",
          5692 => x"05550c87",
          5693 => x"a0affe73",
          5694 => x"27f23887",
          5695 => x"a0b08053",
          5696 => x"878bc5e2",
          5697 => x"f1737084",
          5698 => x"05550c87",
          5699 => x"a0bffe73",
          5700 => x"27ee3880",
          5701 => x"5280c851",
          5702 => x"a79e3f80",
          5703 => x"5280c551",
          5704 => x"a7963f80",
          5705 => x"5280cc51",
          5706 => x"a78e3f80",
          5707 => x"5280cc51",
          5708 => x"a7863f80",
          5709 => x"5280cf51",
          5710 => x"a6fe3f80",
          5711 => x"528a51a6",
          5712 => x"f73f8052",
          5713 => x"be51a6f0",
          5714 => x"3f8199b8",
          5715 => x"59819aca",
          5716 => x"5a830284",
          5717 => x"05950534",
          5718 => x"805b853d",
          5719 => x"7082f2c0",
          5720 => x"0c7082f2",
          5721 => x"b80c82f2",
          5722 => x"bc0c82bc",
          5723 => x"fc51ffbc",
          5724 => x"f23f88ab",
          5725 => x"3f91ec3f",
          5726 => x"82bd8c51",
          5727 => x"ffbce43f",
          5728 => x"82bd9851",
          5729 => x"ffbcdc3f",
          5730 => x"80defc51",
          5731 => x"91d03f81",
          5732 => x"51ebac3f",
          5733 => x"efa23f80",
          5734 => x"04fe3d0d",
          5735 => x"80528353",
          5736 => x"71882b52",
          5737 => x"86d43f82",
          5738 => x"d6d80881",
          5739 => x"ff067207",
          5740 => x"ff145452",
          5741 => x"728025e8",
          5742 => x"387182d6",
          5743 => x"d80c843d",
          5744 => x"0d04fc3d",
          5745 => x"0d767008",
          5746 => x"54558073",
          5747 => x"52547274",
          5748 => x"2e818a38",
          5749 => x"72335170",
          5750 => x"a02e0981",
          5751 => x"06863881",
          5752 => x"1353f139",
          5753 => x"72335170",
          5754 => x"a22e0981",
          5755 => x"06863881",
          5756 => x"13538154",
          5757 => x"72527381",
          5758 => x"2e098106",
          5759 => x"9f388439",
          5760 => x"81125280",
          5761 => x"72335254",
          5762 => x"70a22e83",
          5763 => x"38815470",
          5764 => x"802e9d38",
          5765 => x"73ea3898",
          5766 => x"39811252",
          5767 => x"80723352",
          5768 => x"5470a02e",
          5769 => x"83388154",
          5770 => x"70802e84",
          5771 => x"3873ea38",
          5772 => x"80723352",
          5773 => x"5470a02e",
          5774 => x"09810683",
          5775 => x"38815470",
          5776 => x"a2327030",
          5777 => x"70802576",
          5778 => x"07515151",
          5779 => x"70802e88",
          5780 => x"38807270",
          5781 => x"81055434",
          5782 => x"71750c72",
          5783 => x"517082d6",
          5784 => x"d80c863d",
          5785 => x"0d04fc3d",
          5786 => x"0d765372",
          5787 => x"08802e91",
          5788 => x"38863dfc",
          5789 => x"05527251",
          5790 => x"d6ac3f82",
          5791 => x"d6d80885",
          5792 => x"38805383",
          5793 => x"39745372",
          5794 => x"82d6d80c",
          5795 => x"863d0d04",
          5796 => x"fc3d0d76",
          5797 => x"821133ff",
          5798 => x"05525381",
          5799 => x"52708b26",
          5800 => x"81983883",
          5801 => x"1333ff05",
          5802 => x"51825270",
          5803 => x"9e26818a",
          5804 => x"38841333",
          5805 => x"51835270",
          5806 => x"972680fe",
          5807 => x"38851333",
          5808 => x"51845270",
          5809 => x"bb2680f2",
          5810 => x"38861333",
          5811 => x"51855270",
          5812 => x"bb2680e6",
          5813 => x"38881322",
          5814 => x"55865274",
          5815 => x"87e72680",
          5816 => x"d9388a13",
          5817 => x"22548752",
          5818 => x"7387e726",
          5819 => x"80cc3881",
          5820 => x"0b87c098",
          5821 => x"9c0c7222",
          5822 => x"87c098bc",
          5823 => x"0c821333",
          5824 => x"87c098b8",
          5825 => x"0c831333",
          5826 => x"87c098b4",
          5827 => x"0c841333",
          5828 => x"87c098b0",
          5829 => x"0c851333",
          5830 => x"87c098ac",
          5831 => x"0c861333",
          5832 => x"87c098a8",
          5833 => x"0c7487c0",
          5834 => x"98a40c73",
          5835 => x"87c098a0",
          5836 => x"0c800b87",
          5837 => x"c0989c0c",
          5838 => x"80527182",
          5839 => x"d6d80c86",
          5840 => x"3d0d04f3",
          5841 => x"3d0d7f5b",
          5842 => x"87c0989c",
          5843 => x"5d817d0c",
          5844 => x"87c098bc",
          5845 => x"085e7d7b",
          5846 => x"2387c098",
          5847 => x"b8085a79",
          5848 => x"821c3487",
          5849 => x"c098b408",
          5850 => x"5a79831c",
          5851 => x"3487c098",
          5852 => x"b0085a79",
          5853 => x"841c3487",
          5854 => x"c098ac08",
          5855 => x"5a79851c",
          5856 => x"3487c098",
          5857 => x"a8085a79",
          5858 => x"861c3487",
          5859 => x"c098a408",
          5860 => x"5c7b881c",
          5861 => x"2387c098",
          5862 => x"a0085a79",
          5863 => x"8a1c2380",
          5864 => x"7d0c7983",
          5865 => x"ffff0659",
          5866 => x"7b83ffff",
          5867 => x"0658861b",
          5868 => x"3357851b",
          5869 => x"3356841b",
          5870 => x"3355831b",
          5871 => x"3354821b",
          5872 => x"33537d83",
          5873 => x"ffff0652",
          5874 => x"82bdb051",
          5875 => x"ff9c893f",
          5876 => x"8f3d0d04",
          5877 => x"fb3d0d02",
          5878 => x"9f053382",
          5879 => x"d3ec3370",
          5880 => x"81ff0658",
          5881 => x"555587c0",
          5882 => x"94845175",
          5883 => x"802e8638",
          5884 => x"87c09494",
          5885 => x"51700870",
          5886 => x"962a7081",
          5887 => x"06535452",
          5888 => x"70802e8c",
          5889 => x"3871912a",
          5890 => x"70810651",
          5891 => x"5170d738",
          5892 => x"72813270",
          5893 => x"81065151",
          5894 => x"70802e8d",
          5895 => x"3871932a",
          5896 => x"70810651",
          5897 => x"5170ffbe",
          5898 => x"387381ff",
          5899 => x"065187c0",
          5900 => x"94805270",
          5901 => x"802e8638",
          5902 => x"87c09490",
          5903 => x"5274720c",
          5904 => x"7482d6d8",
          5905 => x"0c873d0d",
          5906 => x"04ff3d0d",
          5907 => x"028f0533",
          5908 => x"7030709f",
          5909 => x"2a515252",
          5910 => x"7082d3ec",
          5911 => x"34833d0d",
          5912 => x"04f93d0d",
          5913 => x"79548074",
          5914 => x"337081ff",
          5915 => x"06535357",
          5916 => x"70772e80",
          5917 => x"fc387181",
          5918 => x"ff068115",
          5919 => x"82d3ec33",
          5920 => x"7081ff06",
          5921 => x"59575558",
          5922 => x"87c09484",
          5923 => x"5175802e",
          5924 => x"863887c0",
          5925 => x"94945170",
          5926 => x"0870962a",
          5927 => x"70810653",
          5928 => x"54527080",
          5929 => x"2e8c3871",
          5930 => x"912a7081",
          5931 => x"06515170",
          5932 => x"d7387281",
          5933 => x"32708106",
          5934 => x"51517080",
          5935 => x"2e8d3871",
          5936 => x"932a7081",
          5937 => x"06515170",
          5938 => x"ffbe3874",
          5939 => x"81ff0651",
          5940 => x"87c09480",
          5941 => x"5270802e",
          5942 => x"863887c0",
          5943 => x"94905277",
          5944 => x"720c8117",
          5945 => x"74337081",
          5946 => x"ff065353",
          5947 => x"5770ff86",
          5948 => x"387682d6",
          5949 => x"d80c893d",
          5950 => x"0d04fe3d",
          5951 => x"0d82d3ec",
          5952 => x"337081ff",
          5953 => x"06545287",
          5954 => x"c0948451",
          5955 => x"72802e86",
          5956 => x"3887c094",
          5957 => x"94517008",
          5958 => x"70822a70",
          5959 => x"81065151",
          5960 => x"5170802e",
          5961 => x"e2387181",
          5962 => x"ff065187",
          5963 => x"c0948052",
          5964 => x"70802e86",
          5965 => x"3887c094",
          5966 => x"90527108",
          5967 => x"7081ff06",
          5968 => x"82d6d80c",
          5969 => x"51843d0d",
          5970 => x"04fe3d0d",
          5971 => x"82d3ec33",
          5972 => x"7081ff06",
          5973 => x"525387c0",
          5974 => x"94845270",
          5975 => x"802e8638",
          5976 => x"87c09494",
          5977 => x"52710870",
          5978 => x"822a7081",
          5979 => x"06515151",
          5980 => x"ff527080",
          5981 => x"2ea03872",
          5982 => x"81ff0651",
          5983 => x"87c09480",
          5984 => x"5270802e",
          5985 => x"863887c0",
          5986 => x"94905271",
          5987 => x"0870982b",
          5988 => x"70982c51",
          5989 => x"53517182",
          5990 => x"d6d80c84",
          5991 => x"3d0d04ff",
          5992 => x"3d0d87c0",
          5993 => x"9e800870",
          5994 => x"9c2a8a06",
          5995 => x"51517080",
          5996 => x"2e84b438",
          5997 => x"87c09ea4",
          5998 => x"0882d3f0",
          5999 => x"0c87c09e",
          6000 => x"a80882d3",
          6001 => x"f40c87c0",
          6002 => x"9e940882",
          6003 => x"d3f80c87",
          6004 => x"c09e9808",
          6005 => x"82d3fc0c",
          6006 => x"87c09e9c",
          6007 => x"0882d480",
          6008 => x"0c87c09e",
          6009 => x"a00882d4",
          6010 => x"840c87c0",
          6011 => x"9eac0882",
          6012 => x"d4880c87",
          6013 => x"c09eb008",
          6014 => x"82d48c0c",
          6015 => x"87c09eb4",
          6016 => x"0882d490",
          6017 => x"0c87c09e",
          6018 => x"b80882d4",
          6019 => x"940c87c0",
          6020 => x"9ebc0882",
          6021 => x"d4980c87",
          6022 => x"c09ec008",
          6023 => x"82d49c0c",
          6024 => x"87c09ec4",
          6025 => x"0882d4a0",
          6026 => x"0c87c09e",
          6027 => x"80085170",
          6028 => x"82d4a423",
          6029 => x"87c09e84",
          6030 => x"0882d4a8",
          6031 => x"0c87c09e",
          6032 => x"880882d4",
          6033 => x"ac0c87c0",
          6034 => x"9e8c0882",
          6035 => x"d4b00c81",
          6036 => x"0b82d4b4",
          6037 => x"34800b87",
          6038 => x"c09e9008",
          6039 => x"7084800a",
          6040 => x"06515252",
          6041 => x"70802e83",
          6042 => x"38815271",
          6043 => x"82d4b534",
          6044 => x"800b87c0",
          6045 => x"9e900870",
          6046 => x"88800a06",
          6047 => x"51525270",
          6048 => x"802e8338",
          6049 => x"81527182",
          6050 => x"d4b63480",
          6051 => x"0b87c09e",
          6052 => x"90087090",
          6053 => x"800a0651",
          6054 => x"52527080",
          6055 => x"2e833881",
          6056 => x"527182d4",
          6057 => x"b734800b",
          6058 => x"87c09e90",
          6059 => x"08708880",
          6060 => x"80065152",
          6061 => x"5270802e",
          6062 => x"83388152",
          6063 => x"7182d4b8",
          6064 => x"34800b87",
          6065 => x"c09e9008",
          6066 => x"70a08080",
          6067 => x"06515252",
          6068 => x"70802e83",
          6069 => x"38815271",
          6070 => x"82d4b934",
          6071 => x"800b87c0",
          6072 => x"9e900870",
          6073 => x"90808006",
          6074 => x"51525270",
          6075 => x"802e8338",
          6076 => x"81527182",
          6077 => x"d4ba3480",
          6078 => x"0b87c09e",
          6079 => x"90087084",
          6080 => x"80800651",
          6081 => x"52527080",
          6082 => x"2e833881",
          6083 => x"527182d4",
          6084 => x"bb34800b",
          6085 => x"87c09e90",
          6086 => x"08708280",
          6087 => x"80065152",
          6088 => x"5270802e",
          6089 => x"83388152",
          6090 => x"7182d4bc",
          6091 => x"34800b87",
          6092 => x"c09e9008",
          6093 => x"70818080",
          6094 => x"06515252",
          6095 => x"70802e83",
          6096 => x"38815271",
          6097 => x"82d4bd34",
          6098 => x"800b87c0",
          6099 => x"9e900870",
          6100 => x"80c08006",
          6101 => x"51525270",
          6102 => x"802e8338",
          6103 => x"81527182",
          6104 => x"d4be3480",
          6105 => x"0b87c09e",
          6106 => x"900870a0",
          6107 => x"80065152",
          6108 => x"5270802e",
          6109 => x"83388152",
          6110 => x"7182d4bf",
          6111 => x"3487c09e",
          6112 => x"90087098",
          6113 => x"8006708a",
          6114 => x"2a515151",
          6115 => x"7082d4c0",
          6116 => x"34800b87",
          6117 => x"c09e9008",
          6118 => x"70848006",
          6119 => x"51525270",
          6120 => x"802e8338",
          6121 => x"81527182",
          6122 => x"d4c13487",
          6123 => x"c09e9008",
          6124 => x"7083f006",
          6125 => x"70842a51",
          6126 => x"51517082",
          6127 => x"d4c23480",
          6128 => x"0b87c09e",
          6129 => x"90087088",
          6130 => x"06515252",
          6131 => x"70802e83",
          6132 => x"38815271",
          6133 => x"82d4c334",
          6134 => x"87c09e90",
          6135 => x"08708706",
          6136 => x"51517082",
          6137 => x"d4c43483",
          6138 => x"3d0d04fb",
          6139 => x"3d0d82bd",
          6140 => x"c851ff93",
          6141 => x"e33f82d4",
          6142 => x"b4335473",
          6143 => x"802e8938",
          6144 => x"82bddc51",
          6145 => x"ff93d13f",
          6146 => x"82bdf051",
          6147 => x"ffafd43f",
          6148 => x"82d4b633",
          6149 => x"5473802e",
          6150 => x"943882d4",
          6151 => x"900882d4",
          6152 => x"94081154",
          6153 => x"5282be88",
          6154 => x"51ff93ac",
          6155 => x"3f82d4bb",
          6156 => x"33547380",
          6157 => x"2e943882",
          6158 => x"d4880882",
          6159 => x"d48c0811",
          6160 => x"545282be",
          6161 => x"a451ff93",
          6162 => x"8f3f82d4",
          6163 => x"b8335473",
          6164 => x"802e9438",
          6165 => x"82d3f008",
          6166 => x"82d3f408",
          6167 => x"11545282",
          6168 => x"bec051ff",
          6169 => x"92f23f82",
          6170 => x"d4b93354",
          6171 => x"73802e94",
          6172 => x"3882d3f8",
          6173 => x"0882d3fc",
          6174 => x"08115452",
          6175 => x"82bedc51",
          6176 => x"ff92d53f",
          6177 => x"82d4ba33",
          6178 => x"5473802e",
          6179 => x"943882d4",
          6180 => x"800882d4",
          6181 => x"84081154",
          6182 => x"5282bef8",
          6183 => x"51ff92b8",
          6184 => x"3f82d4bf",
          6185 => x"33547380",
          6186 => x"2e8e3882",
          6187 => x"d4c03352",
          6188 => x"82bf9451",
          6189 => x"ff92a13f",
          6190 => x"82d4c333",
          6191 => x"5473802e",
          6192 => x"8e3882d4",
          6193 => x"c4335282",
          6194 => x"bfb451ff",
          6195 => x"928a3f82",
          6196 => x"d4c13354",
          6197 => x"73802e8e",
          6198 => x"3882d4c2",
          6199 => x"335282bf",
          6200 => x"d451ff91",
          6201 => x"f33f82d4",
          6202 => x"b5335473",
          6203 => x"802e8938",
          6204 => x"82bff451",
          6205 => x"ffadec3f",
          6206 => x"82d4b733",
          6207 => x"5473802e",
          6208 => x"893882c0",
          6209 => x"8851ffad",
          6210 => x"da3f82d4",
          6211 => x"bc335473",
          6212 => x"802e8938",
          6213 => x"82c09451",
          6214 => x"ffadc83f",
          6215 => x"82d4bd33",
          6216 => x"5473802e",
          6217 => x"893882c0",
          6218 => x"a051ffad",
          6219 => x"b63f82d4",
          6220 => x"be335473",
          6221 => x"802e8938",
          6222 => x"82c0a851",
          6223 => x"ffada43f",
          6224 => x"82c0b051",
          6225 => x"ffad9c3f",
          6226 => x"82d49808",
          6227 => x"5282c0bc",
          6228 => x"51ff9184",
          6229 => x"3f82d49c",
          6230 => x"085282c0",
          6231 => x"e451ff90",
          6232 => x"f73f82d4",
          6233 => x"a0085282",
          6234 => x"c18c51ff",
          6235 => x"90ea3f82",
          6236 => x"c1b451ff",
          6237 => x"aced3f82",
          6238 => x"d4a42252",
          6239 => x"82c1bc51",
          6240 => x"ff90d53f",
          6241 => x"82d4a808",
          6242 => x"56bd84c0",
          6243 => x"527551c5",
          6244 => x"9d3f82d6",
          6245 => x"d808bd84",
          6246 => x"c0297671",
          6247 => x"31545482",
          6248 => x"d6d80852",
          6249 => x"82c1e451",
          6250 => x"ff90ad3f",
          6251 => x"82d4bb33",
          6252 => x"5473802e",
          6253 => x"a93882d4",
          6254 => x"ac0856bd",
          6255 => x"84c05275",
          6256 => x"51c4eb3f",
          6257 => x"82d6d808",
          6258 => x"bd84c029",
          6259 => x"76713154",
          6260 => x"5482d6d8",
          6261 => x"085282c2",
          6262 => x"9051ff8f",
          6263 => x"fb3f82d4",
          6264 => x"b6335473",
          6265 => x"802ea938",
          6266 => x"82d4b008",
          6267 => x"56bd84c0",
          6268 => x"527551c4",
          6269 => x"b93f82d6",
          6270 => x"d808bd84",
          6271 => x"c0297671",
          6272 => x"31545482",
          6273 => x"d6d80852",
          6274 => x"82c2bc51",
          6275 => x"ff8fc93f",
          6276 => x"8a51ffae",
          6277 => x"f03f873d",
          6278 => x"0d04fe3d",
          6279 => x"0d029205",
          6280 => x"33ff0552",
          6281 => x"718426aa",
          6282 => x"38718429",
          6283 => x"82adac05",
          6284 => x"52710804",
          6285 => x"82c2e851",
          6286 => x"9d3982c2",
          6287 => x"f0519739",
          6288 => x"82c2f851",
          6289 => x"913982c3",
          6290 => x"80518b39",
          6291 => x"82c38451",
          6292 => x"853982c3",
          6293 => x"8c51ff8e",
          6294 => x"ff3f843d",
          6295 => x"0d047188",
          6296 => x"800c0480",
          6297 => x"0b87c096",
          6298 => x"840c0482",
          6299 => x"d4c80887",
          6300 => x"c096840c",
          6301 => x"04fd3d0d",
          6302 => x"76982b70",
          6303 => x"982c7998",
          6304 => x"2b70982c",
          6305 => x"72101370",
          6306 => x"822b5153",
          6307 => x"51545151",
          6308 => x"800b82c3",
          6309 => x"98123355",
          6310 => x"53717425",
          6311 => x"9c3882c3",
          6312 => x"94110812",
          6313 => x"02840597",
          6314 => x"05337133",
          6315 => x"52525270",
          6316 => x"722e0981",
          6317 => x"06833881",
          6318 => x"537282d6",
          6319 => x"d80c853d",
          6320 => x"0d04fb3d",
          6321 => x"0d790284",
          6322 => x"05a30533",
          6323 => x"71335556",
          6324 => x"5472802e",
          6325 => x"b13882f2",
          6326 => x"bc085288",
          6327 => x"51ffadd2",
          6328 => x"3f82f2bc",
          6329 => x"0852a051",
          6330 => x"ffadc73f",
          6331 => x"82f2bc08",
          6332 => x"528851ff",
          6333 => x"adbc3f73",
          6334 => x"33ff0553",
          6335 => x"72743472",
          6336 => x"81ff0653",
          6337 => x"cc397751",
          6338 => x"ff8dcd3f",
          6339 => x"74743487",
          6340 => x"3d0d04f6",
          6341 => x"3d0d7c02",
          6342 => x"8405b705",
          6343 => x"33028805",
          6344 => x"bb053382",
          6345 => x"d5a43370",
          6346 => x"842982d4",
          6347 => x"cc057008",
          6348 => x"5159595a",
          6349 => x"58597480",
          6350 => x"2e863874",
          6351 => x"519c933f",
          6352 => x"82d5a433",
          6353 => x"70842982",
          6354 => x"d4cc0581",
          6355 => x"19705458",
          6356 => x"565a9f94",
          6357 => x"3f82d6d8",
          6358 => x"08750c82",
          6359 => x"d5a43370",
          6360 => x"842982d4",
          6361 => x"cc057008",
          6362 => x"51565a74",
          6363 => x"802ea738",
          6364 => x"75537852",
          6365 => x"7451ffb6",
          6366 => x"ec3f82d5",
          6367 => x"a4338105",
          6368 => x"557482d5",
          6369 => x"a4347481",
          6370 => x"ff065593",
          6371 => x"75278738",
          6372 => x"800b82d5",
          6373 => x"a4347780",
          6374 => x"2eb63882",
          6375 => x"d5a00856",
          6376 => x"75802eac",
          6377 => x"3882d59c",
          6378 => x"335574a4",
          6379 => x"388c3dfc",
          6380 => x"05547653",
          6381 => x"78527551",
          6382 => x"80ecd73f",
          6383 => x"82d5a008",
          6384 => x"528a5181",
          6385 => x"a2803f82",
          6386 => x"d5a00851",
          6387 => x"80f0ba3f",
          6388 => x"8c3d0d04",
          6389 => x"fd3d0d82",
          6390 => x"d4cc5393",
          6391 => x"54720852",
          6392 => x"71802e89",
          6393 => x"3871519a",
          6394 => x"e93f8073",
          6395 => x"0cff1484",
          6396 => x"14545473",
          6397 => x"8025e638",
          6398 => x"800b82d5",
          6399 => x"a43482d5",
          6400 => x"a0085271",
          6401 => x"802e9538",
          6402 => x"715180f1",
          6403 => x"9f3f82d5",
          6404 => x"a008519a",
          6405 => x"bd3f800b",
          6406 => x"82d5a00c",
          6407 => x"853d0d04",
          6408 => x"dc3d0d81",
          6409 => x"57805282",
          6410 => x"d5a00851",
          6411 => x"80f6bb3f",
          6412 => x"82d6d808",
          6413 => x"80d33882",
          6414 => x"d5a00853",
          6415 => x"80f85288",
          6416 => x"3d705256",
          6417 => x"819eeb3f",
          6418 => x"82d6d808",
          6419 => x"802eba38",
          6420 => x"7551ffb3",
          6421 => x"b03f82d6",
          6422 => x"d8085580",
          6423 => x"0b82d6d8",
          6424 => x"08259d38",
          6425 => x"82d6d808",
          6426 => x"ff057017",
          6427 => x"55558074",
          6428 => x"34755376",
          6429 => x"52811782",
          6430 => x"c6885257",
          6431 => x"ff8ad93f",
          6432 => x"74ff2e09",
          6433 => x"8106ffaf",
          6434 => x"38a63d0d",
          6435 => x"04d93d0d",
          6436 => x"aa3d08ad",
          6437 => x"3d085a5a",
          6438 => x"81705858",
          6439 => x"805282d5",
          6440 => x"a0085180",
          6441 => x"f5c43f82",
          6442 => x"d6d80881",
          6443 => x"9538ff0b",
          6444 => x"82d5a008",
          6445 => x"545580f8",
          6446 => x"528b3d70",
          6447 => x"5256819d",
          6448 => x"f13f82d6",
          6449 => x"d808802e",
          6450 => x"a5387551",
          6451 => x"ffb2b63f",
          6452 => x"82d6d808",
          6453 => x"81185855",
          6454 => x"800b82d6",
          6455 => x"d808258e",
          6456 => x"3882d6d8",
          6457 => x"08ff0570",
          6458 => x"17555580",
          6459 => x"74347409",
          6460 => x"70307072",
          6461 => x"079f2a51",
          6462 => x"55557877",
          6463 => x"2e853873",
          6464 => x"ffac3882",
          6465 => x"d5a0088c",
          6466 => x"11085351",
          6467 => x"80f4db3f",
          6468 => x"82d6d808",
          6469 => x"802e8938",
          6470 => x"82c69451",
          6471 => x"ff89b93f",
          6472 => x"78772e09",
          6473 => x"81069b38",
          6474 => x"75527951",
          6475 => x"ffb2c43f",
          6476 => x"7951ffb1",
          6477 => x"d03fab3d",
          6478 => x"085482d6",
          6479 => x"d8087434",
          6480 => x"80587782",
          6481 => x"d6d80ca9",
          6482 => x"3d0d04f6",
          6483 => x"3d0d7c7e",
          6484 => x"715c7172",
          6485 => x"3357595a",
          6486 => x"5873a02e",
          6487 => x"098106a2",
          6488 => x"38783378",
          6489 => x"05567776",
          6490 => x"27983881",
          6491 => x"17705b70",
          6492 => x"71335658",
          6493 => x"5573a02e",
          6494 => x"09810686",
          6495 => x"38757526",
          6496 => x"ea388054",
          6497 => x"73882982",
          6498 => x"d5a80570",
          6499 => x"085255ff",
          6500 => x"b0f33f82",
          6501 => x"d6d80853",
          6502 => x"79527408",
          6503 => x"51ffb3f2",
          6504 => x"3f82d6d8",
          6505 => x"0880c538",
          6506 => x"84153355",
          6507 => x"74812e88",
          6508 => x"3874822e",
          6509 => x"8838b539",
          6510 => x"fce63fac",
          6511 => x"39811a5a",
          6512 => x"8c3dfc11",
          6513 => x"53f80551",
          6514 => x"c5ad3f82",
          6515 => x"d6d80880",
          6516 => x"2e9a38ff",
          6517 => x"1b537852",
          6518 => x"7751fdb1",
          6519 => x"3f82d6d8",
          6520 => x"0881ff06",
          6521 => x"55748538",
          6522 => x"74549139",
          6523 => x"81147081",
          6524 => x"ff065154",
          6525 => x"827427ff",
          6526 => x"8b388054",
          6527 => x"7382d6d8",
          6528 => x"0c8c3d0d",
          6529 => x"04d33d0d",
          6530 => x"b03d08b2",
          6531 => x"3d08b43d",
          6532 => x"08595f5a",
          6533 => x"800baf3d",
          6534 => x"3482d5a4",
          6535 => x"3382d5a0",
          6536 => x"08555b73",
          6537 => x"81cb3873",
          6538 => x"82d59c33",
          6539 => x"55557383",
          6540 => x"38815576",
          6541 => x"802e81bc",
          6542 => x"38817076",
          6543 => x"06555673",
          6544 => x"802e81ad",
          6545 => x"38a85199",
          6546 => x"9f3f82d6",
          6547 => x"d80882d5",
          6548 => x"a00c82d6",
          6549 => x"d808802e",
          6550 => x"81923893",
          6551 => x"53765282",
          6552 => x"d6d80851",
          6553 => x"80dfc63f",
          6554 => x"82d6d808",
          6555 => x"802e8c38",
          6556 => x"82c6c051",
          6557 => x"ffa2ec3f",
          6558 => x"80f73982",
          6559 => x"d6d8085b",
          6560 => x"82d5a008",
          6561 => x"5380f852",
          6562 => x"903d7052",
          6563 => x"54819aa2",
          6564 => x"3f82d6d8",
          6565 => x"085682d6",
          6566 => x"d808742e",
          6567 => x"09810680",
          6568 => x"d03882d6",
          6569 => x"d80851ff",
          6570 => x"aedb3f82",
          6571 => x"d6d80855",
          6572 => x"800b82d6",
          6573 => x"d80825a9",
          6574 => x"3882d6d8",
          6575 => x"08ff0570",
          6576 => x"17555580",
          6577 => x"74348053",
          6578 => x"7481ff06",
          6579 => x"527551f8",
          6580 => x"c23f811b",
          6581 => x"7081ff06",
          6582 => x"5c54937b",
          6583 => x"27833880",
          6584 => x"5b74ff2e",
          6585 => x"098106ff",
          6586 => x"97388639",
          6587 => x"7582d59c",
          6588 => x"34768c38",
          6589 => x"82d5a008",
          6590 => x"802e8438",
          6591 => x"f9d63f8f",
          6592 => x"3d5decc5",
          6593 => x"3f82d6d8",
          6594 => x"08982b70",
          6595 => x"982c5159",
          6596 => x"78ff2eee",
          6597 => x"387881ff",
          6598 => x"0682ee94",
          6599 => x"3370982b",
          6600 => x"70982c82",
          6601 => x"ee903370",
          6602 => x"982b7097",
          6603 => x"2c71982c",
          6604 => x"05708429",
          6605 => x"82c39405",
          6606 => x"70081570",
          6607 => x"33515151",
          6608 => x"51595951",
          6609 => x"595d5881",
          6610 => x"5673782e",
          6611 => x"80e93877",
          6612 => x"7427b438",
          6613 => x"7481800a",
          6614 => x"2981ff0a",
          6615 => x"0570982c",
          6616 => x"51558075",
          6617 => x"2480ce38",
          6618 => x"76537452",
          6619 => x"7751f685",
          6620 => x"3f82d6d8",
          6621 => x"0881ff06",
          6622 => x"5473802e",
          6623 => x"d7387482",
          6624 => x"ee903481",
          6625 => x"56b13974",
          6626 => x"81800a29",
          6627 => x"81800a05",
          6628 => x"70982c70",
          6629 => x"81ff0656",
          6630 => x"51557395",
          6631 => x"26973876",
          6632 => x"53745277",
          6633 => x"51f5ce3f",
          6634 => x"82d6d808",
          6635 => x"81ff0654",
          6636 => x"73cc38d3",
          6637 => x"39805675",
          6638 => x"802e80ca",
          6639 => x"38811c55",
          6640 => x"7482ee94",
          6641 => x"3474982b",
          6642 => x"70982c82",
          6643 => x"ee903370",
          6644 => x"982b7098",
          6645 => x"2c701011",
          6646 => x"70822b82",
          6647 => x"c3981133",
          6648 => x"5e515151",
          6649 => x"57585155",
          6650 => x"74772e09",
          6651 => x"8106fe92",
          6652 => x"3882c39c",
          6653 => x"14087d0c",
          6654 => x"800b82ee",
          6655 => x"9434800b",
          6656 => x"82ee9034",
          6657 => x"92397582",
          6658 => x"ee943475",
          6659 => x"82ee9034",
          6660 => x"78af3d34",
          6661 => x"757d0c7e",
          6662 => x"54739526",
          6663 => x"fde13873",
          6664 => x"842982ad",
          6665 => x"c0055473",
          6666 => x"080482ee",
          6667 => x"9c335473",
          6668 => x"7e2efdcb",
          6669 => x"3882ee98",
          6670 => x"33557375",
          6671 => x"27ab3874",
          6672 => x"982b7098",
          6673 => x"2c515573",
          6674 => x"75249e38",
          6675 => x"741a5473",
          6676 => x"33811534",
          6677 => x"7481800a",
          6678 => x"2981ff0a",
          6679 => x"0570982c",
          6680 => x"82ee9c33",
          6681 => x"565155df",
          6682 => x"3982ee9c",
          6683 => x"33811156",
          6684 => x"547482ee",
          6685 => x"9c34731a",
          6686 => x"54ae3d33",
          6687 => x"743482ee",
          6688 => x"98335473",
          6689 => x"7e258938",
          6690 => x"81145473",
          6691 => x"82ee9834",
          6692 => x"82ee9c33",
          6693 => x"7081800a",
          6694 => x"2981ff0a",
          6695 => x"0570982c",
          6696 => x"82ee9833",
          6697 => x"5a515656",
          6698 => x"747725a8",
          6699 => x"3882f2bc",
          6700 => x"0852741a",
          6701 => x"70335254",
          6702 => x"ffa1f73f",
          6703 => x"7481800a",
          6704 => x"2981800a",
          6705 => x"0570982c",
          6706 => x"82ee9833",
          6707 => x"56515573",
          6708 => x"7524da38",
          6709 => x"82ee9c33",
          6710 => x"70982b70",
          6711 => x"982c82ee",
          6712 => x"98335a51",
          6713 => x"56567477",
          6714 => x"25fc9438",
          6715 => x"82f2bc08",
          6716 => x"528851ff",
          6717 => x"a1bc3f74",
          6718 => x"81800a29",
          6719 => x"81800a05",
          6720 => x"70982c82",
          6721 => x"ee983356",
          6722 => x"51557375",
          6723 => x"24de38fb",
          6724 => x"ee39837a",
          6725 => x"34800b81",
          6726 => x"1b3482ee",
          6727 => x"9c538052",
          6728 => x"82b6a051",
          6729 => x"f39c3f81",
          6730 => x"fd3982ee",
          6731 => x"9c337081",
          6732 => x"ff065555",
          6733 => x"73802efb",
          6734 => x"c63882ee",
          6735 => x"9833ff05",
          6736 => x"547382ee",
          6737 => x"9834ff15",
          6738 => x"547382ee",
          6739 => x"9c3482f2",
          6740 => x"bc085288",
          6741 => x"51ffa0da",
          6742 => x"3f82ee9c",
          6743 => x"3370982b",
          6744 => x"70982c82",
          6745 => x"ee983357",
          6746 => x"51565774",
          6747 => x"7425ad38",
          6748 => x"741a5481",
          6749 => x"14337434",
          6750 => x"82f2bc08",
          6751 => x"52733351",
          6752 => x"ffa0af3f",
          6753 => x"7481800a",
          6754 => x"2981800a",
          6755 => x"0570982c",
          6756 => x"82ee9833",
          6757 => x"58515575",
          6758 => x"7524d538",
          6759 => x"82f2bc08",
          6760 => x"52a051ff",
          6761 => x"a08c3f82",
          6762 => x"ee9c3370",
          6763 => x"982b7098",
          6764 => x"2c82ee98",
          6765 => x"33575156",
          6766 => x"57747424",
          6767 => x"fac13882",
          6768 => x"f2bc0852",
          6769 => x"8851ff9f",
          6770 => x"e93f7481",
          6771 => x"800a2981",
          6772 => x"800a0570",
          6773 => x"982c82ee",
          6774 => x"98335851",
          6775 => x"55757525",
          6776 => x"de38fa9b",
          6777 => x"3982ee98",
          6778 => x"337a0554",
          6779 => x"80743482",
          6780 => x"f2bc0852",
          6781 => x"8a51ff9f",
          6782 => x"b93f82ee",
          6783 => x"98527951",
          6784 => x"f6c93f82",
          6785 => x"d6d80881",
          6786 => x"ff065473",
          6787 => x"963882ee",
          6788 => x"98335473",
          6789 => x"802e8f38",
          6790 => x"81537352",
          6791 => x"7951f1f3",
          6792 => x"3f843980",
          6793 => x"7a34800b",
          6794 => x"82ee9c34",
          6795 => x"800b82ee",
          6796 => x"98347982",
          6797 => x"d6d80caf",
          6798 => x"3d0d0482",
          6799 => x"ee9c3354",
          6800 => x"73802ef9",
          6801 => x"ba3882f2",
          6802 => x"bc085288",
          6803 => x"51ff9ee2",
          6804 => x"3f82ee9c",
          6805 => x"33ff0554",
          6806 => x"7382ee9c",
          6807 => x"347381ff",
          6808 => x"0654dd39",
          6809 => x"82ee9c33",
          6810 => x"82ee9833",
          6811 => x"55557375",
          6812 => x"2ef98c38",
          6813 => x"ff145473",
          6814 => x"82ee9834",
          6815 => x"74982b70",
          6816 => x"982c7581",
          6817 => x"ff065651",
          6818 => x"55747425",
          6819 => x"ad38741a",
          6820 => x"54811433",
          6821 => x"743482f2",
          6822 => x"bc085273",
          6823 => x"3351ff9e",
          6824 => x"913f7481",
          6825 => x"800a2981",
          6826 => x"800a0570",
          6827 => x"982c82ee",
          6828 => x"98335851",
          6829 => x"55757524",
          6830 => x"d53882f2",
          6831 => x"bc0852a0",
          6832 => x"51ff9dee",
          6833 => x"3f82ee9c",
          6834 => x"3370982b",
          6835 => x"70982c82",
          6836 => x"ee983357",
          6837 => x"51565774",
          6838 => x"7424f8a3",
          6839 => x"3882f2bc",
          6840 => x"08528851",
          6841 => x"ff9dcb3f",
          6842 => x"7481800a",
          6843 => x"2981800a",
          6844 => x"0570982c",
          6845 => x"82ee9833",
          6846 => x"58515575",
          6847 => x"7525de38",
          6848 => x"f7fd3982",
          6849 => x"ee9c3370",
          6850 => x"81ff0682",
          6851 => x"ee983359",
          6852 => x"56547477",
          6853 => x"27f7e838",
          6854 => x"82f2bc08",
          6855 => x"52811454",
          6856 => x"7382ee9c",
          6857 => x"34741a70",
          6858 => x"335254ff",
          6859 => x"9d843f82",
          6860 => x"ee9c3370",
          6861 => x"81ff0682",
          6862 => x"ee983358",
          6863 => x"56547575",
          6864 => x"26d638f7",
          6865 => x"ba3982ee",
          6866 => x"9c538052",
          6867 => x"82b6a051",
          6868 => x"eef03f80",
          6869 => x"0b82ee9c",
          6870 => x"34800b82",
          6871 => x"ee9834f7",
          6872 => x"9e397ab0",
          6873 => x"3882d598",
          6874 => x"08557480",
          6875 => x"2ea63874",
          6876 => x"51ffa591",
          6877 => x"3f82d6d8",
          6878 => x"0882ee98",
          6879 => x"3482d6d8",
          6880 => x"0881ff06",
          6881 => x"81055374",
          6882 => x"527951ff",
          6883 => x"a6d73f93",
          6884 => x"5b81c039",
          6885 => x"7a842982",
          6886 => x"d4cc05fc",
          6887 => x"11085654",
          6888 => x"74802ea7",
          6889 => x"387451ff",
          6890 => x"a4db3f82",
          6891 => x"d6d80882",
          6892 => x"ee983482",
          6893 => x"d6d80881",
          6894 => x"ff068105",
          6895 => x"53745279",
          6896 => x"51ffa6a1",
          6897 => x"3fff1b54",
          6898 => x"80fa3973",
          6899 => x"08557480",
          6900 => x"2ef6ac38",
          6901 => x"7451ffa4",
          6902 => x"ac3f9939",
          6903 => x"7a932e09",
          6904 => x"8106ae38",
          6905 => x"82d4cc08",
          6906 => x"5574802e",
          6907 => x"a4387451",
          6908 => x"ffa4923f",
          6909 => x"82d6d808",
          6910 => x"82ee9834",
          6911 => x"82d6d808",
          6912 => x"81ff0681",
          6913 => x"05537452",
          6914 => x"7951ffa5",
          6915 => x"d83f80c3",
          6916 => x"397a8429",
          6917 => x"82d4d005",
          6918 => x"70085654",
          6919 => x"74802eab",
          6920 => x"387451ff",
          6921 => x"a3df3f82",
          6922 => x"d6d80882",
          6923 => x"ee983482",
          6924 => x"d6d80881",
          6925 => x"ff068105",
          6926 => x"53745279",
          6927 => x"51ffa5a5",
          6928 => x"3f811b54",
          6929 => x"7381ff06",
          6930 => x"5b893974",
          6931 => x"82ee9834",
          6932 => x"747a3482",
          6933 => x"ee9c5382",
          6934 => x"ee983352",
          6935 => x"7951ece2",
          6936 => x"3ff59c39",
          6937 => x"82ee9c33",
          6938 => x"7081ff06",
          6939 => x"82ee9833",
          6940 => x"59565474",
          6941 => x"7727f587",
          6942 => x"3882f2bc",
          6943 => x"08528114",
          6944 => x"547382ee",
          6945 => x"9c34741a",
          6946 => x"70335254",
          6947 => x"ff9aa33f",
          6948 => x"f4ed3982",
          6949 => x"ee9c3354",
          6950 => x"73802ef4",
          6951 => x"e23882f2",
          6952 => x"bc085288",
          6953 => x"51ff9a8a",
          6954 => x"3f82ee9c",
          6955 => x"33ff0554",
          6956 => x"7382ee9c",
          6957 => x"34f4c839",
          6958 => x"ff3d0d02",
          6959 => x"8f053352",
          6960 => x"718a2e09",
          6961 => x"8106a038",
          6962 => x"82d6c408",
          6963 => x"810582d6",
          6964 => x"c40c980b",
          6965 => x"82d6c408",
          6966 => x"25873898",
          6967 => x"0b82d6c4",
          6968 => x"0c800b82",
          6969 => x"d6c80c82",
          6970 => x"d6c40884",
          6971 => x"2982d6c4",
          6972 => x"08057088",
          6973 => x"2982d6c8",
          6974 => x"080587a0",
          6975 => x"a0801170",
          6976 => x"82d6c00c",
          6977 => x"51515182",
          6978 => x"d5c01233",
          6979 => x"713482d6",
          6980 => x"c8088105",
          6981 => x"82d6c80c",
          6982 => x"a70b82d6",
          6983 => x"c80825a0",
          6984 => x"3882d6c4",
          6985 => x"08810582",
          6986 => x"d6c40c98",
          6987 => x"0b82d6c4",
          6988 => x"08258738",
          6989 => x"980b82d6",
          6990 => x"c40c800b",
          6991 => x"82d6c80c",
          6992 => x"800b82d6",
          6993 => x"d80c833d",
          6994 => x"0d04ff0b",
          6995 => x"82d6d80c",
          6996 => x"04f93d0d",
          6997 => x"83bff40b",
          6998 => x"82d6d00c",
          6999 => x"84800b82",
          7000 => x"d6cc23a0",
          7001 => x"80538052",
          7002 => x"83bff451",
          7003 => x"ffa9a23f",
          7004 => x"82d6d008",
          7005 => x"54805877",
          7006 => x"74348157",
          7007 => x"76811534",
          7008 => x"82d6d008",
          7009 => x"54778415",
          7010 => x"34768515",
          7011 => x"3482d6d0",
          7012 => x"08547786",
          7013 => x"15347687",
          7014 => x"153482d6",
          7015 => x"d00882d6",
          7016 => x"cc22ff05",
          7017 => x"fe808007",
          7018 => x"7083ffff",
          7019 => x"0670882a",
          7020 => x"58515556",
          7021 => x"74881734",
          7022 => x"73891734",
          7023 => x"82d6cc22",
          7024 => x"70882982",
          7025 => x"d6d00805",
          7026 => x"f8115155",
          7027 => x"55778215",
          7028 => x"34768315",
          7029 => x"34893d0d",
          7030 => x"04ff3d0d",
          7031 => x"73528151",
          7032 => x"8472278f",
          7033 => x"38fb1283",
          7034 => x"2a821170",
          7035 => x"83ffff06",
          7036 => x"51515170",
          7037 => x"82d6d80c",
          7038 => x"833d0d04",
          7039 => x"f93d0d02",
          7040 => x"a6052202",
          7041 => x"8405aa05",
          7042 => x"22710582",
          7043 => x"d6d00871",
          7044 => x"832b7111",
          7045 => x"74832b73",
          7046 => x"11703381",
          7047 => x"12337188",
          7048 => x"2b0702a4",
          7049 => x"05ae0522",
          7050 => x"7181ffff",
          7051 => x"06077088",
          7052 => x"2a535152",
          7053 => x"59545b5b",
          7054 => x"57535455",
          7055 => x"71773470",
          7056 => x"81183482",
          7057 => x"d6d00814",
          7058 => x"75882a52",
          7059 => x"54708215",
          7060 => x"34748315",
          7061 => x"3482d6d0",
          7062 => x"08701770",
          7063 => x"33811233",
          7064 => x"71882b07",
          7065 => x"70832b8f",
          7066 => x"fff80651",
          7067 => x"52565271",
          7068 => x"057383ff",
          7069 => x"ff067088",
          7070 => x"2a545451",
          7071 => x"71821234",
          7072 => x"7281ff06",
          7073 => x"53728312",
          7074 => x"3482d6d0",
          7075 => x"08165671",
          7076 => x"76347281",
          7077 => x"1734893d",
          7078 => x"0d04fb3d",
          7079 => x"0d82d6d0",
          7080 => x"08028405",
          7081 => x"9e052270",
          7082 => x"832b7211",
          7083 => x"86113387",
          7084 => x"1233718b",
          7085 => x"2b71832b",
          7086 => x"07585b59",
          7087 => x"52555272",
          7088 => x"05841233",
          7089 => x"85133371",
          7090 => x"882b0770",
          7091 => x"882a5456",
          7092 => x"56527084",
          7093 => x"13347385",
          7094 => x"133482d6",
          7095 => x"d0087014",
          7096 => x"84113385",
          7097 => x"1233718b",
          7098 => x"2b71832b",
          7099 => x"07565957",
          7100 => x"52720586",
          7101 => x"12338713",
          7102 => x"3371882b",
          7103 => x"0770882a",
          7104 => x"54565652",
          7105 => x"70861334",
          7106 => x"73871334",
          7107 => x"82d6d008",
          7108 => x"13703381",
          7109 => x"12337188",
          7110 => x"2b077081",
          7111 => x"ffff0670",
          7112 => x"882a5351",
          7113 => x"53535371",
          7114 => x"73347081",
          7115 => x"1434873d",
          7116 => x"0d04fa3d",
          7117 => x"0d02a205",
          7118 => x"2282d6d0",
          7119 => x"0871832b",
          7120 => x"71117033",
          7121 => x"81123371",
          7122 => x"882b0770",
          7123 => x"88291570",
          7124 => x"33811233",
          7125 => x"71982b71",
          7126 => x"902b0753",
          7127 => x"5f535552",
          7128 => x"5a565753",
          7129 => x"54718025",
          7130 => x"80f63872",
          7131 => x"51feab3f",
          7132 => x"82d6d008",
          7133 => x"70167033",
          7134 => x"81123371",
          7135 => x"8b2b7183",
          7136 => x"2b077411",
          7137 => x"70338112",
          7138 => x"3371882b",
          7139 => x"0770832b",
          7140 => x"8ffff806",
          7141 => x"51525451",
          7142 => x"535a5853",
          7143 => x"72057488",
          7144 => x"2a545272",
          7145 => x"82133473",
          7146 => x"83133482",
          7147 => x"d6d00870",
          7148 => x"16703381",
          7149 => x"1233718b",
          7150 => x"2b71832b",
          7151 => x"07565957",
          7152 => x"55720570",
          7153 => x"33811233",
          7154 => x"71882b07",
          7155 => x"7081ffff",
          7156 => x"0670882a",
          7157 => x"57515258",
          7158 => x"52727434",
          7159 => x"71811534",
          7160 => x"883d0d04",
          7161 => x"fb3d0d82",
          7162 => x"d6d00802",
          7163 => x"84059e05",
          7164 => x"2270832b",
          7165 => x"72118211",
          7166 => x"33831233",
          7167 => x"718b2b71",
          7168 => x"832b0759",
          7169 => x"5b595256",
          7170 => x"52730571",
          7171 => x"33811333",
          7172 => x"71882b07",
          7173 => x"028c05a2",
          7174 => x"05227107",
          7175 => x"70882a53",
          7176 => x"51535353",
          7177 => x"71733470",
          7178 => x"81143482",
          7179 => x"d6d00870",
          7180 => x"15703381",
          7181 => x"1233718b",
          7182 => x"2b71832b",
          7183 => x"07565957",
          7184 => x"52720582",
          7185 => x"12338313",
          7186 => x"3371882b",
          7187 => x"0770882a",
          7188 => x"54555652",
          7189 => x"70821334",
          7190 => x"72831334",
          7191 => x"82d6d008",
          7192 => x"14821133",
          7193 => x"83123371",
          7194 => x"882b0782",
          7195 => x"d6d80c52",
          7196 => x"54873d0d",
          7197 => x"04f73d0d",
          7198 => x"7b82d6d0",
          7199 => x"0831832a",
          7200 => x"7083ffff",
          7201 => x"06705357",
          7202 => x"53fda73f",
          7203 => x"82d6d008",
          7204 => x"76832b71",
          7205 => x"11821133",
          7206 => x"83123371",
          7207 => x"8b2b7183",
          7208 => x"2b077511",
          7209 => x"70338112",
          7210 => x"3371982b",
          7211 => x"71902b07",
          7212 => x"53424051",
          7213 => x"535b5855",
          7214 => x"59547280",
          7215 => x"258d3882",
          7216 => x"80805275",
          7217 => x"51fe9d3f",
          7218 => x"81843984",
          7219 => x"14338515",
          7220 => x"33718b2b",
          7221 => x"71832b07",
          7222 => x"76117988",
          7223 => x"2a535155",
          7224 => x"58557686",
          7225 => x"14347581",
          7226 => x"ff065675",
          7227 => x"87143482",
          7228 => x"d6d00870",
          7229 => x"19841233",
          7230 => x"85133371",
          7231 => x"882b0770",
          7232 => x"882a5457",
          7233 => x"5b565372",
          7234 => x"84163473",
          7235 => x"85163482",
          7236 => x"d6d00818",
          7237 => x"53800b86",
          7238 => x"1434800b",
          7239 => x"87143482",
          7240 => x"d6d00853",
          7241 => x"76841434",
          7242 => x"75851434",
          7243 => x"82d6d008",
          7244 => x"18703381",
          7245 => x"12337188",
          7246 => x"2b077082",
          7247 => x"80800770",
          7248 => x"882a5351",
          7249 => x"55565474",
          7250 => x"74347281",
          7251 => x"15348b3d",
          7252 => x"0d04ff3d",
          7253 => x"0d735282",
          7254 => x"d6d00884",
          7255 => x"38f7f23f",
          7256 => x"71802e86",
          7257 => x"387151fe",
          7258 => x"8c3f833d",
          7259 => x"0d04f53d",
          7260 => x"0d807e52",
          7261 => x"58f8e23f",
          7262 => x"82d6d808",
          7263 => x"83ffff06",
          7264 => x"82d6d008",
          7265 => x"84113385",
          7266 => x"12337188",
          7267 => x"2b07705f",
          7268 => x"5956585a",
          7269 => x"81ffff59",
          7270 => x"75782e80",
          7271 => x"cb387588",
          7272 => x"29177033",
          7273 => x"81123371",
          7274 => x"882b0770",
          7275 => x"81ffff06",
          7276 => x"79317083",
          7277 => x"ffff0670",
          7278 => x"7f275253",
          7279 => x"51565955",
          7280 => x"7779278a",
          7281 => x"3873802e",
          7282 => x"85387578",
          7283 => x"5a5b8415",
          7284 => x"33851633",
          7285 => x"71882b07",
          7286 => x"575475c2",
          7287 => x"387881ff",
          7288 => x"ff2e8538",
          7289 => x"7a795956",
          7290 => x"8076832b",
          7291 => x"82d6d008",
          7292 => x"11703381",
          7293 => x"12337188",
          7294 => x"2b077081",
          7295 => x"ffff0651",
          7296 => x"525a565c",
          7297 => x"5573752e",
          7298 => x"83388155",
          7299 => x"80547978",
          7300 => x"2681cc38",
          7301 => x"74547480",
          7302 => x"2e81c438",
          7303 => x"777a2e09",
          7304 => x"81068938",
          7305 => x"7551f8f2",
          7306 => x"3f81ac39",
          7307 => x"82808053",
          7308 => x"79527551",
          7309 => x"f7c63f82",
          7310 => x"d6d00870",
          7311 => x"1c861133",
          7312 => x"87123371",
          7313 => x"8b2b7183",
          7314 => x"2b07535a",
          7315 => x"5e557405",
          7316 => x"7a177083",
          7317 => x"ffff0670",
          7318 => x"882a5c59",
          7319 => x"56547884",
          7320 => x"15347681",
          7321 => x"ff065776",
          7322 => x"85153482",
          7323 => x"d6d00875",
          7324 => x"832b7111",
          7325 => x"721e8611",
          7326 => x"33871233",
          7327 => x"71882b07",
          7328 => x"70882a53",
          7329 => x"5b5e535a",
          7330 => x"56547386",
          7331 => x"19347587",
          7332 => x"193482d6",
          7333 => x"d008701c",
          7334 => x"84113385",
          7335 => x"1233718b",
          7336 => x"2b71832b",
          7337 => x"07535d5a",
          7338 => x"55740554",
          7339 => x"78861534",
          7340 => x"76871534",
          7341 => x"82d6d008",
          7342 => x"7016711d",
          7343 => x"84113385",
          7344 => x"12337188",
          7345 => x"2b077088",
          7346 => x"2a535a5f",
          7347 => x"52565473",
          7348 => x"84163475",
          7349 => x"85163482",
          7350 => x"d6d0081b",
          7351 => x"84055473",
          7352 => x"82d6d80c",
          7353 => x"8d3d0d04",
          7354 => x"fe3d0d74",
          7355 => x"5282d6d0",
          7356 => x"088438f4",
          7357 => x"dc3f7153",
          7358 => x"71802e8b",
          7359 => x"387151fc",
          7360 => x"ed3f82d6",
          7361 => x"d8085372",
          7362 => x"82d6d80c",
          7363 => x"843d0d04",
          7364 => x"ee3d0d64",
          7365 => x"66405c80",
          7366 => x"70424082",
          7367 => x"d6d00860",
          7368 => x"2e098106",
          7369 => x"8438f4a9",
          7370 => x"3f7b8e38",
          7371 => x"7e51ffb8",
          7372 => x"3f82d6d8",
          7373 => x"085483c7",
          7374 => x"397e8b38",
          7375 => x"7b51fc92",
          7376 => x"3f7e5483",
          7377 => x"ba397e51",
          7378 => x"f58f3f82",
          7379 => x"d6d80883",
          7380 => x"ffff0682",
          7381 => x"d6d0087d",
          7382 => x"7131832a",
          7383 => x"7083ffff",
          7384 => x"0670832b",
          7385 => x"73117033",
          7386 => x"81123371",
          7387 => x"882b0770",
          7388 => x"75317083",
          7389 => x"ffff0670",
          7390 => x"8829fc05",
          7391 => x"7388291a",
          7392 => x"70338112",
          7393 => x"3371882b",
          7394 => x"0770902b",
          7395 => x"53444e53",
          7396 => x"4841525c",
          7397 => x"545b415c",
          7398 => x"565b5b73",
          7399 => x"80258f38",
          7400 => x"7681ffff",
          7401 => x"06753170",
          7402 => x"83ffff06",
          7403 => x"42548216",
          7404 => x"33831733",
          7405 => x"71882b07",
          7406 => x"7088291c",
          7407 => x"70338112",
          7408 => x"3371982b",
          7409 => x"71902b07",
          7410 => x"53474552",
          7411 => x"56547380",
          7412 => x"258b3878",
          7413 => x"75317083",
          7414 => x"ffff0641",
          7415 => x"54777b27",
          7416 => x"81fe3860",
          7417 => x"1854737b",
          7418 => x"2e098106",
          7419 => x"8f387851",
          7420 => x"f6c03f7a",
          7421 => x"83ffff06",
          7422 => x"5881e539",
          7423 => x"7f8e387a",
          7424 => x"74248938",
          7425 => x"7851f6aa",
          7426 => x"3f81a539",
          7427 => x"7f18557a",
          7428 => x"752480c8",
          7429 => x"38791d82",
          7430 => x"11338312",
          7431 => x"3371882b",
          7432 => x"07535754",
          7433 => x"f4f43f80",
          7434 => x"527851f7",
          7435 => x"b73f82d6",
          7436 => x"d80883ff",
          7437 => x"ff067e54",
          7438 => x"7c537083",
          7439 => x"2b82d6d0",
          7440 => x"08118405",
          7441 => x"535559ff",
          7442 => x"90d13f82",
          7443 => x"d6d00814",
          7444 => x"84057583",
          7445 => x"ffff0659",
          7446 => x"5c818539",
          7447 => x"6015547a",
          7448 => x"742480d4",
          7449 => x"387851f5",
          7450 => x"c93f82d6",
          7451 => x"d0081d82",
          7452 => x"11338312",
          7453 => x"3371882b",
          7454 => x"07534354",
          7455 => x"f49c3f80",
          7456 => x"527851f6",
          7457 => x"df3f82d6",
          7458 => x"d80883ff",
          7459 => x"ff067e54",
          7460 => x"7c537083",
          7461 => x"2b82d6d0",
          7462 => x"08118405",
          7463 => x"535559ff",
          7464 => x"8ff93f82",
          7465 => x"d6d00814",
          7466 => x"84056062",
          7467 => x"0519555c",
          7468 => x"7383ffff",
          7469 => x"0658a939",
          7470 => x"7b7f5254",
          7471 => x"f9b03f82",
          7472 => x"d6d8085c",
          7473 => x"82d6d808",
          7474 => x"802e9338",
          7475 => x"7d537352",
          7476 => x"82d6d808",
          7477 => x"51ff948d",
          7478 => x"3f7351f7",
          7479 => x"983f7a58",
          7480 => x"7a782799",
          7481 => x"3880537a",
          7482 => x"527851f2",
          7483 => x"8f3f7a19",
          7484 => x"832b82d6",
          7485 => x"d0080584",
          7486 => x"0551f6f9",
          7487 => x"3f7b5473",
          7488 => x"82d6d80c",
          7489 => x"943d0d04",
          7490 => x"fc3d0d77",
          7491 => x"77297052",
          7492 => x"54fbd53f",
          7493 => x"82d6d808",
          7494 => x"5582d6d8",
          7495 => x"08802e8e",
          7496 => x"38735380",
          7497 => x"5282d6d8",
          7498 => x"0851ff99",
          7499 => x"e43f7482",
          7500 => x"d6d80c86",
          7501 => x"3d0d04ff",
          7502 => x"3d0d028f",
          7503 => x"05335181",
          7504 => x"52707226",
          7505 => x"873882d6",
          7506 => x"d4113352",
          7507 => x"7182d6d8",
          7508 => x"0c833d0d",
          7509 => x"04fc3d0d",
          7510 => x"029b0533",
          7511 => x"0284059f",
          7512 => x"05335653",
          7513 => x"83517281",
          7514 => x"2680e038",
          7515 => x"72842b87",
          7516 => x"c0928c11",
          7517 => x"53518854",
          7518 => x"74802e84",
          7519 => x"38818854",
          7520 => x"73720c87",
          7521 => x"c0928c11",
          7522 => x"5181710c",
          7523 => x"850b87c0",
          7524 => x"988c0c70",
          7525 => x"52710870",
          7526 => x"82065151",
          7527 => x"70802e8a",
          7528 => x"3887c098",
          7529 => x"8c085170",
          7530 => x"ec387108",
          7531 => x"fc808006",
          7532 => x"52719238",
          7533 => x"87c0988c",
          7534 => x"08517080",
          7535 => x"2e873871",
          7536 => x"82d6d414",
          7537 => x"3482d6d4",
          7538 => x"13335170",
          7539 => x"82d6d80c",
          7540 => x"863d0d04",
          7541 => x"f33d0d60",
          7542 => x"6264028c",
          7543 => x"05bf0533",
          7544 => x"5740585b",
          7545 => x"8374525a",
          7546 => x"fecd3f82",
          7547 => x"d6d80881",
          7548 => x"067a5452",
          7549 => x"7181be38",
          7550 => x"71727584",
          7551 => x"2b87c092",
          7552 => x"801187c0",
          7553 => x"928c1287",
          7554 => x"c0928413",
          7555 => x"415a4057",
          7556 => x"5a58850b",
          7557 => x"87c0988c",
          7558 => x"0c767d0c",
          7559 => x"84760c75",
          7560 => x"0870852a",
          7561 => x"70810651",
          7562 => x"53547180",
          7563 => x"2e8e387b",
          7564 => x"0852717b",
          7565 => x"7081055d",
          7566 => x"34811959",
          7567 => x"8074a206",
          7568 => x"53537173",
          7569 => x"2e833881",
          7570 => x"537883ff",
          7571 => x"268f3872",
          7572 => x"802e8a38",
          7573 => x"87c0988c",
          7574 => x"085271c3",
          7575 => x"3887c098",
          7576 => x"8c085271",
          7577 => x"802e8738",
          7578 => x"7884802e",
          7579 => x"99388176",
          7580 => x"0c87c092",
          7581 => x"8c155372",
          7582 => x"08708206",
          7583 => x"515271f7",
          7584 => x"38ff1a5a",
          7585 => x"8d398480",
          7586 => x"17811970",
          7587 => x"81ff065a",
          7588 => x"53577980",
          7589 => x"2e903873",
          7590 => x"fc808006",
          7591 => x"52718738",
          7592 => x"7d7826fe",
          7593 => x"ed3873fc",
          7594 => x"80800652",
          7595 => x"71802e83",
          7596 => x"38815271",
          7597 => x"537282d6",
          7598 => x"d80c8f3d",
          7599 => x"0d04f33d",
          7600 => x"0d606264",
          7601 => x"028c05bf",
          7602 => x"05335740",
          7603 => x"585b8359",
          7604 => x"80745258",
          7605 => x"fce13f82",
          7606 => x"d6d80881",
          7607 => x"06795452",
          7608 => x"71782e09",
          7609 => x"810681b1",
          7610 => x"38777484",
          7611 => x"2b87c092",
          7612 => x"801187c0",
          7613 => x"928c1287",
          7614 => x"c0928413",
          7615 => x"40595f56",
          7616 => x"5a850b87",
          7617 => x"c0988c0c",
          7618 => x"767d0c82",
          7619 => x"760c8058",
          7620 => x"75087084",
          7621 => x"2a708106",
          7622 => x"51535471",
          7623 => x"802e8c38",
          7624 => x"7a708105",
          7625 => x"5c337c0c",
          7626 => x"81185873",
          7627 => x"812a7081",
          7628 => x"06515271",
          7629 => x"802e8a38",
          7630 => x"87c0988c",
          7631 => x"085271d0",
          7632 => x"3887c098",
          7633 => x"8c085271",
          7634 => x"802e8738",
          7635 => x"7784802e",
          7636 => x"99388176",
          7637 => x"0c87c092",
          7638 => x"8c155372",
          7639 => x"08708206",
          7640 => x"515271f7",
          7641 => x"38ff1959",
          7642 => x"8d39811a",
          7643 => x"7081ff06",
          7644 => x"84801959",
          7645 => x"5b527880",
          7646 => x"2e903873",
          7647 => x"fc808006",
          7648 => x"52718738",
          7649 => x"7d7a26fe",
          7650 => x"f83873fc",
          7651 => x"80800652",
          7652 => x"71802e83",
          7653 => x"38815271",
          7654 => x"537282d6",
          7655 => x"d80c8f3d",
          7656 => x"0d04fa3d",
          7657 => x"0d7a0284",
          7658 => x"05a30533",
          7659 => x"028805a7",
          7660 => x"05337154",
          7661 => x"545657fa",
          7662 => x"fe3f82d6",
          7663 => x"d8088106",
          7664 => x"53835472",
          7665 => x"80fe3885",
          7666 => x"0b87c098",
          7667 => x"8c0c8156",
          7668 => x"71762e80",
          7669 => x"dc387176",
          7670 => x"24933874",
          7671 => x"842b87c0",
          7672 => x"928c1154",
          7673 => x"5471802e",
          7674 => x"8d3880d4",
          7675 => x"3971832e",
          7676 => x"80c63880",
          7677 => x"cb397208",
          7678 => x"70812a70",
          7679 => x"81065151",
          7680 => x"5271802e",
          7681 => x"8a3887c0",
          7682 => x"988c0852",
          7683 => x"71e83887",
          7684 => x"c0988c08",
          7685 => x"52719638",
          7686 => x"81730c87",
          7687 => x"c0928c14",
          7688 => x"53720870",
          7689 => x"82065152",
          7690 => x"71f73896",
          7691 => x"39805692",
          7692 => x"3988800a",
          7693 => x"770c8539",
          7694 => x"8180770c",
          7695 => x"72568339",
          7696 => x"84567554",
          7697 => x"7382d6d8",
          7698 => x"0c883d0d",
          7699 => x"04fe3d0d",
          7700 => x"74811133",
          7701 => x"71337188",
          7702 => x"2b0782d6",
          7703 => x"d80c5351",
          7704 => x"843d0d04",
          7705 => x"fd3d0d75",
          7706 => x"83113382",
          7707 => x"12337190",
          7708 => x"2b71882b",
          7709 => x"07811433",
          7710 => x"70720788",
          7711 => x"2b753371",
          7712 => x"0782d6d8",
          7713 => x"0c525354",
          7714 => x"56545285",
          7715 => x"3d0d04ff",
          7716 => x"3d0d7302",
          7717 => x"84059205",
          7718 => x"22525270",
          7719 => x"72708105",
          7720 => x"54347088",
          7721 => x"2a517072",
          7722 => x"34833d0d",
          7723 => x"04ff3d0d",
          7724 => x"73755252",
          7725 => x"70727081",
          7726 => x"05543470",
          7727 => x"882a5170",
          7728 => x"72708105",
          7729 => x"54347088",
          7730 => x"2a517072",
          7731 => x"70810554",
          7732 => x"3470882a",
          7733 => x"51707234",
          7734 => x"833d0d04",
          7735 => x"fe3d0d76",
          7736 => x"75775454",
          7737 => x"5170802e",
          7738 => x"92387170",
          7739 => x"81055333",
          7740 => x"73708105",
          7741 => x"5534ff11",
          7742 => x"51eb3984",
          7743 => x"3d0d04fe",
          7744 => x"3d0d7577",
          7745 => x"76545253",
          7746 => x"72727081",
          7747 => x"055434ff",
          7748 => x"115170f4",
          7749 => x"38843d0d",
          7750 => x"04fc3d0d",
          7751 => x"78777956",
          7752 => x"56537470",
          7753 => x"81055633",
          7754 => x"74708105",
          7755 => x"56337171",
          7756 => x"31ff1656",
          7757 => x"52525272",
          7758 => x"802e8638",
          7759 => x"71802ee2",
          7760 => x"387182d6",
          7761 => x"d80c863d",
          7762 => x"0d04fe3d",
          7763 => x"0d747654",
          7764 => x"51893971",
          7765 => x"732e8a38",
          7766 => x"81115170",
          7767 => x"335271f3",
          7768 => x"38703382",
          7769 => x"d6d80c84",
          7770 => x"3d0d0480",
          7771 => x"0b82d6d8",
          7772 => x"0c04fb3d",
          7773 => x"0d777008",
          7774 => x"70708105",
          7775 => x"52337054",
          7776 => x"555556e7",
          7777 => x"3fff5582",
          7778 => x"d6d808a2",
          7779 => x"3872802e",
          7780 => x"983883b5",
          7781 => x"52725180",
          7782 => x"f7b63f82",
          7783 => x"d6d80883",
          7784 => x"ffff0653",
          7785 => x"72802e86",
          7786 => x"3873760c",
          7787 => x"72557482",
          7788 => x"d6d80c87",
          7789 => x"3d0d04f7",
          7790 => x"3d0d7b56",
          7791 => x"800b8317",
          7792 => x"33565a74",
          7793 => x"7a2e80d6",
          7794 => x"388154b4",
          7795 => x"160853b8",
          7796 => x"16705381",
          7797 => x"17335259",
          7798 => x"f9e43f82",
          7799 => x"d6d8087a",
          7800 => x"2e098106",
          7801 => x"b73882d6",
          7802 => x"d8088317",
          7803 => x"34b41608",
          7804 => x"70a81808",
          7805 => x"31a01808",
          7806 => x"59565874",
          7807 => x"77279f38",
          7808 => x"82163355",
          7809 => x"74822e09",
          7810 => x"81069338",
          7811 => x"81547618",
          7812 => x"53785281",
          7813 => x"163351f9",
          7814 => x"a53f8339",
          7815 => x"815a7982",
          7816 => x"d6d80c8b",
          7817 => x"3d0d04fa",
          7818 => x"3d0d787a",
          7819 => x"56568057",
          7820 => x"74b41708",
          7821 => x"2eaf3875",
          7822 => x"51fefc3f",
          7823 => x"82d6d808",
          7824 => x"5782d6d8",
          7825 => x"089f3881",
          7826 => x"547453b8",
          7827 => x"16528116",
          7828 => x"3351f780",
          7829 => x"3f82d6d8",
          7830 => x"08802e85",
          7831 => x"38ff5581",
          7832 => x"5774b417",
          7833 => x"0c7682d6",
          7834 => x"d80c883d",
          7835 => x"0d04f83d",
          7836 => x"0d7a7052",
          7837 => x"57fec03f",
          7838 => x"82d6d808",
          7839 => x"5882d6d8",
          7840 => x"08819138",
          7841 => x"76335574",
          7842 => x"832e0981",
          7843 => x"0680f038",
          7844 => x"84173359",
          7845 => x"78812e09",
          7846 => x"810680e3",
          7847 => x"38848053",
          7848 => x"82d6d808",
          7849 => x"52b81770",
          7850 => x"5256fcd3",
          7851 => x"3f82d4d5",
          7852 => x"5284b617",
          7853 => x"51fbd83f",
          7854 => x"848b85a4",
          7855 => x"d2527551",
          7856 => x"fbeb3f86",
          7857 => x"8a85e4f2",
          7858 => x"52849c17",
          7859 => x"51fbde3f",
          7860 => x"94170852",
          7861 => x"84a01751",
          7862 => x"fbd33f90",
          7863 => x"17085284",
          7864 => x"a41751fb",
          7865 => x"c83fa417",
          7866 => x"08810570",
          7867 => x"b4190c79",
          7868 => x"55537552",
          7869 => x"81173351",
          7870 => x"f7c43f77",
          7871 => x"84183480",
          7872 => x"53805281",
          7873 => x"173351f9",
          7874 => x"993f82d6",
          7875 => x"d808802e",
          7876 => x"83388158",
          7877 => x"7782d6d8",
          7878 => x"0c8a3d0d",
          7879 => x"04fb3d0d",
          7880 => x"77fe1a9c",
          7881 => x"1208fe05",
          7882 => x"55565480",
          7883 => x"56747327",
          7884 => x"8d388a14",
          7885 => x"22757129",
          7886 => x"b0160805",
          7887 => x"57537582",
          7888 => x"d6d80c87",
          7889 => x"3d0d04f9",
          7890 => x"3d0d7a7a",
          7891 => x"70085654",
          7892 => x"57817727",
          7893 => x"81df3876",
          7894 => x"9c150827",
          7895 => x"81d738ff",
          7896 => x"74335458",
          7897 => x"72822e80",
          7898 => x"f5387282",
          7899 => x"24893872",
          7900 => x"812e8d38",
          7901 => x"81bf3972",
          7902 => x"832e818e",
          7903 => x"3881b639",
          7904 => x"76812a17",
          7905 => x"70892aa8",
          7906 => x"16080553",
          7907 => x"745255fd",
          7908 => x"963f82d6",
          7909 => x"d808819f",
          7910 => x"387483ff",
          7911 => x"0614b811",
          7912 => x"33811770",
          7913 => x"892aa818",
          7914 => x"08055576",
          7915 => x"54575753",
          7916 => x"fcf53f82",
          7917 => x"d6d80880",
          7918 => x"fe387483",
          7919 => x"ff0614b8",
          7920 => x"11337088",
          7921 => x"2b780779",
          7922 => x"81067184",
          7923 => x"2a5c5258",
          7924 => x"51537280",
          7925 => x"e238759f",
          7926 => x"ff065880",
          7927 => x"da397688",
          7928 => x"2aa81508",
          7929 => x"05527351",
          7930 => x"fcbd3f82",
          7931 => x"d6d80880",
          7932 => x"c6387610",
          7933 => x"83fe0674",
          7934 => x"05b80551",
          7935 => x"f8cf3f82",
          7936 => x"d6d80883",
          7937 => x"ffff0658",
          7938 => x"ae397687",
          7939 => x"2aa81508",
          7940 => x"05527351",
          7941 => x"fc913f82",
          7942 => x"d6d8089b",
          7943 => x"3876822b",
          7944 => x"83fc0674",
          7945 => x"05b80551",
          7946 => x"f8ba3f82",
          7947 => x"d6d808f0",
          7948 => x"0a065883",
          7949 => x"39815877",
          7950 => x"82d6d80c",
          7951 => x"893d0d04",
          7952 => x"f83d0d7a",
          7953 => x"7c7e5a58",
          7954 => x"56825981",
          7955 => x"7727829e",
          7956 => x"38769c17",
          7957 => x"08278296",
          7958 => x"38753353",
          7959 => x"72792e81",
          7960 => x"9d387279",
          7961 => x"24893872",
          7962 => x"812e8d38",
          7963 => x"82803972",
          7964 => x"832e81b8",
          7965 => x"3881f739",
          7966 => x"76812a17",
          7967 => x"70892aa8",
          7968 => x"18080553",
          7969 => x"765255fb",
          7970 => x"9e3f82d6",
          7971 => x"d8085982",
          7972 => x"d6d80881",
          7973 => x"d9387483",
          7974 => x"ff0616b8",
          7975 => x"05811678",
          7976 => x"81065956",
          7977 => x"54775376",
          7978 => x"802e8f38",
          7979 => x"77842b9f",
          7980 => x"f0067433",
          7981 => x"8f067107",
          7982 => x"51537274",
          7983 => x"34810b83",
          7984 => x"17347489",
          7985 => x"2aa81708",
          7986 => x"05527551",
          7987 => x"fad93f82",
          7988 => x"d6d80859",
          7989 => x"82d6d808",
          7990 => x"81943874",
          7991 => x"83ff0616",
          7992 => x"b8057884",
          7993 => x"2a545476",
          7994 => x"8f387788",
          7995 => x"2a743381",
          7996 => x"f006718f",
          7997 => x"06075153",
          7998 => x"72743480",
          7999 => x"ec397688",
          8000 => x"2aa81708",
          8001 => x"05527551",
          8002 => x"fa9d3f82",
          8003 => x"d6d80859",
          8004 => x"82d6d808",
          8005 => x"80d83877",
          8006 => x"83ffff06",
          8007 => x"52761083",
          8008 => x"fe067605",
          8009 => x"b80551f6",
          8010 => x"e63fbe39",
          8011 => x"76872aa8",
          8012 => x"17080552",
          8013 => x"7551f9ef",
          8014 => x"3f82d6d8",
          8015 => x"085982d6",
          8016 => x"d808ab38",
          8017 => x"77f00a06",
          8018 => x"77822b83",
          8019 => x"fc067018",
          8020 => x"b8057054",
          8021 => x"515454f6",
          8022 => x"8b3f82d6",
          8023 => x"d8088f0a",
          8024 => x"06740752",
          8025 => x"7251f6c5",
          8026 => x"3f810b83",
          8027 => x"17347882",
          8028 => x"d6d80c8a",
          8029 => x"3d0d04f8",
          8030 => x"3d0d7a7c",
          8031 => x"7e720859",
          8032 => x"56565981",
          8033 => x"7527a438",
          8034 => x"749c1708",
          8035 => x"279d3873",
          8036 => x"802eaa38",
          8037 => x"ff537352",
          8038 => x"7551fda4",
          8039 => x"3f82d6d8",
          8040 => x"085482d6",
          8041 => x"d80880f2",
          8042 => x"38933982",
          8043 => x"5480eb39",
          8044 => x"815480e6",
          8045 => x"3982d6d8",
          8046 => x"085480de",
          8047 => x"39745278",
          8048 => x"51fb843f",
          8049 => x"82d6d808",
          8050 => x"5882d6d8",
          8051 => x"08802e80",
          8052 => x"c73882d6",
          8053 => x"d808812e",
          8054 => x"d23882d6",
          8055 => x"d808ff2e",
          8056 => x"cf388053",
          8057 => x"74527551",
          8058 => x"fcd63f82",
          8059 => x"d6d808c5",
          8060 => x"389c1608",
          8061 => x"fe119418",
          8062 => x"08575557",
          8063 => x"74742790",
          8064 => x"38811594",
          8065 => x"170c8416",
          8066 => x"33810754",
          8067 => x"73841734",
          8068 => x"77557678",
          8069 => x"26ffa638",
          8070 => x"80547382",
          8071 => x"d6d80c8a",
          8072 => x"3d0d04f6",
          8073 => x"3d0d7c7e",
          8074 => x"7108595b",
          8075 => x"5b799538",
          8076 => x"90170858",
          8077 => x"77802e88",
          8078 => x"389c1708",
          8079 => x"7826b238",
          8080 => x"8158ae39",
          8081 => x"79527a51",
          8082 => x"f9fd3f81",
          8083 => x"557482d6",
          8084 => x"d8082782",
          8085 => x"e03882d6",
          8086 => x"d8085582",
          8087 => x"d6d808ff",
          8088 => x"2e82d238",
          8089 => x"9c170882",
          8090 => x"d6d80826",
          8091 => x"82c73879",
          8092 => x"58941708",
          8093 => x"70565473",
          8094 => x"802e82b9",
          8095 => x"38777a2e",
          8096 => x"09810680",
          8097 => x"e238811a",
          8098 => x"569c1708",
          8099 => x"76268338",
          8100 => x"82567552",
          8101 => x"7a51f9af",
          8102 => x"3f805982",
          8103 => x"d6d80881",
          8104 => x"2e098106",
          8105 => x"863882d6",
          8106 => x"d8085982",
          8107 => x"d6d80809",
          8108 => x"70307072",
          8109 => x"07802570",
          8110 => x"7c0782d6",
          8111 => x"d8085451",
          8112 => x"51555573",
          8113 => x"81ef3882",
          8114 => x"d6d80880",
          8115 => x"2e953890",
          8116 => x"17085481",
          8117 => x"74279038",
          8118 => x"739c1808",
          8119 => x"27893873",
          8120 => x"58853975",
          8121 => x"80db3877",
          8122 => x"56811656",
          8123 => x"9c170876",
          8124 => x"26893882",
          8125 => x"56757826",
          8126 => x"81ac3875",
          8127 => x"527a51f8",
          8128 => x"c63f82d6",
          8129 => x"d808802e",
          8130 => x"b8388059",
          8131 => x"82d6d808",
          8132 => x"812e0981",
          8133 => x"06863882",
          8134 => x"d6d80859",
          8135 => x"82d6d808",
          8136 => x"09703070",
          8137 => x"72078025",
          8138 => x"707c0751",
          8139 => x"51555573",
          8140 => x"80f83875",
          8141 => x"782e0981",
          8142 => x"06ffae38",
          8143 => x"735580f5",
          8144 => x"39ff5375",
          8145 => x"527651f9",
          8146 => x"f73f82d6",
          8147 => x"d80882d6",
          8148 => x"d8083070",
          8149 => x"82d6d808",
          8150 => x"07802551",
          8151 => x"55557980",
          8152 => x"2e943873",
          8153 => x"802e8f38",
          8154 => x"75537952",
          8155 => x"7651f9d0",
          8156 => x"3f82d6d8",
          8157 => x"085574a5",
          8158 => x"38759018",
          8159 => x"0c9c1708",
          8160 => x"fe059418",
          8161 => x"08565474",
          8162 => x"74268638",
          8163 => x"ff159418",
          8164 => x"0c841733",
          8165 => x"81075473",
          8166 => x"84183497",
          8167 => x"39ff5674",
          8168 => x"812e9038",
          8169 => x"8c398055",
          8170 => x"8c3982d6",
          8171 => x"d8085585",
          8172 => x"39815675",
          8173 => x"557482d6",
          8174 => x"d80c8c3d",
          8175 => x"0d04f83d",
          8176 => x"0d7a7052",
          8177 => x"55f3f03f",
          8178 => x"82d6d808",
          8179 => x"58815682",
          8180 => x"d6d80880",
          8181 => x"d8387b52",
          8182 => x"7451f6c1",
          8183 => x"3f82d6d8",
          8184 => x"0882d6d8",
          8185 => x"08b4170c",
          8186 => x"59848053",
          8187 => x"7752b815",
          8188 => x"705257f2",
          8189 => x"8a3f7756",
          8190 => x"84398116",
          8191 => x"568a1522",
          8192 => x"58757827",
          8193 => x"97388154",
          8194 => x"75195376",
          8195 => x"52811533",
          8196 => x"51edab3f",
          8197 => x"82d6d808",
          8198 => x"802edf38",
          8199 => x"8a152276",
          8200 => x"32703070",
          8201 => x"7207709f",
          8202 => x"2a535156",
          8203 => x"567582d6",
          8204 => x"d80c8a3d",
          8205 => x"0d04f83d",
          8206 => x"0d7a7c71",
          8207 => x"08585657",
          8208 => x"74f0800a",
          8209 => x"2680f138",
          8210 => x"749f0653",
          8211 => x"7280e938",
          8212 => x"7490180c",
          8213 => x"88170854",
          8214 => x"73aa3875",
          8215 => x"33538273",
          8216 => x"278838ac",
          8217 => x"16085473",
          8218 => x"9b387485",
          8219 => x"2a53820b",
          8220 => x"8817225a",
          8221 => x"58727927",
          8222 => x"80fe38ac",
          8223 => x"16089818",
          8224 => x"0c80cd39",
          8225 => x"8a162270",
          8226 => x"892b5458",
          8227 => x"727526b2",
          8228 => x"38735276",
          8229 => x"51f5b03f",
          8230 => x"82d6d808",
          8231 => x"5482d6d8",
          8232 => x"08ff2ebd",
          8233 => x"38810b82",
          8234 => x"d6d80827",
          8235 => x"8b389c16",
          8236 => x"0882d6d8",
          8237 => x"08268538",
          8238 => x"8258bd39",
          8239 => x"74733155",
          8240 => x"cb397352",
          8241 => x"7551f4d5",
          8242 => x"3f82d6d8",
          8243 => x"0898180c",
          8244 => x"7394180c",
          8245 => x"98170853",
          8246 => x"82587280",
          8247 => x"2e9a3885",
          8248 => x"39815894",
          8249 => x"3974892a",
          8250 => x"1398180c",
          8251 => x"7483ff06",
          8252 => x"16b8059c",
          8253 => x"180c8058",
          8254 => x"7782d6d8",
          8255 => x"0c8a3d0d",
          8256 => x"04f83d0d",
          8257 => x"7a700890",
          8258 => x"1208a005",
          8259 => x"595754f0",
          8260 => x"800a7727",
          8261 => x"8638800b",
          8262 => x"98150c98",
          8263 => x"14085384",
          8264 => x"5572802e",
          8265 => x"81cb3876",
          8266 => x"83ff0658",
          8267 => x"7781b538",
          8268 => x"81139815",
          8269 => x"0c941408",
          8270 => x"55749238",
          8271 => x"76852a88",
          8272 => x"17225653",
          8273 => x"74732681",
          8274 => x"9b3880c0",
          8275 => x"398a1622",
          8276 => x"ff057789",
          8277 => x"2a065372",
          8278 => x"818a3874",
          8279 => x"527351f3",
          8280 => x"e63f82d6",
          8281 => x"d8085382",
          8282 => x"55810b82",
          8283 => x"d6d80827",
          8284 => x"80ff3881",
          8285 => x"5582d6d8",
          8286 => x"08ff2e80",
          8287 => x"f4389c16",
          8288 => x"0882d6d8",
          8289 => x"082680ca",
          8290 => x"387b8a38",
          8291 => x"7798150c",
          8292 => x"845580dd",
          8293 => x"39941408",
          8294 => x"527351f9",
          8295 => x"863f82d6",
          8296 => x"d8085387",
          8297 => x"5582d6d8",
          8298 => x"08802e80",
          8299 => x"c4388255",
          8300 => x"82d6d808",
          8301 => x"812eba38",
          8302 => x"815582d6",
          8303 => x"d808ff2e",
          8304 => x"b03882d6",
          8305 => x"d8085275",
          8306 => x"51fbf33f",
          8307 => x"82d6d808",
          8308 => x"a0387294",
          8309 => x"150c7252",
          8310 => x"7551f2c1",
          8311 => x"3f82d6d8",
          8312 => x"0898150c",
          8313 => x"7690150c",
          8314 => x"7716b805",
          8315 => x"9c150c80",
          8316 => x"557482d6",
          8317 => x"d80c8a3d",
          8318 => x"0d04f73d",
          8319 => x"0d7b7d71",
          8320 => x"085b5b57",
          8321 => x"80527651",
          8322 => x"fcac3f82",
          8323 => x"d6d80854",
          8324 => x"82d6d808",
          8325 => x"80ec3882",
          8326 => x"d6d80856",
          8327 => x"98170852",
          8328 => x"7851f083",
          8329 => x"3f82d6d8",
          8330 => x"085482d6",
          8331 => x"d80880d2",
          8332 => x"3882d6d8",
          8333 => x"089c1808",
          8334 => x"70335154",
          8335 => x"587281e5",
          8336 => x"2e098106",
          8337 => x"83388158",
          8338 => x"82d6d808",
          8339 => x"55728338",
          8340 => x"81557775",
          8341 => x"07537280",
          8342 => x"2e8e3881",
          8343 => x"1656757a",
          8344 => x"2e098106",
          8345 => x"8838a539",
          8346 => x"82d6d808",
          8347 => x"56815276",
          8348 => x"51fd8e3f",
          8349 => x"82d6d808",
          8350 => x"5482d6d8",
          8351 => x"08802eff",
          8352 => x"9b387384",
          8353 => x"2e098106",
          8354 => x"83388754",
          8355 => x"7382d6d8",
          8356 => x"0c8b3d0d",
          8357 => x"04fd3d0d",
          8358 => x"769a1152",
          8359 => x"54ebae3f",
          8360 => x"82d6d808",
          8361 => x"83ffff06",
          8362 => x"76703351",
          8363 => x"53537183",
          8364 => x"2e098106",
          8365 => x"90389414",
          8366 => x"51eb923f",
          8367 => x"82d6d808",
          8368 => x"902b7307",
          8369 => x"537282d6",
          8370 => x"d80c853d",
          8371 => x"0d04fc3d",
          8372 => x"0d777970",
          8373 => x"83ffff06",
          8374 => x"549a1253",
          8375 => x"5555ebaf",
          8376 => x"3f767033",
          8377 => x"51537283",
          8378 => x"2e098106",
          8379 => x"8b387390",
          8380 => x"2a529415",
          8381 => x"51eb983f",
          8382 => x"863d0d04",
          8383 => x"fd3d0d75",
          8384 => x"5480518b",
          8385 => x"5370812a",
          8386 => x"71818029",
          8387 => x"05747081",
          8388 => x"05563371",
          8389 => x"057081ff",
          8390 => x"06ff1656",
          8391 => x"51515172",
          8392 => x"e4387082",
          8393 => x"d6d80c85",
          8394 => x"3d0d04f2",
          8395 => x"3d0d6062",
          8396 => x"40598479",
          8397 => x"085f5b81",
          8398 => x"ff705d5d",
          8399 => x"98190880",
          8400 => x"2e838038",
          8401 => x"98190852",
          8402 => x"7d51eddb",
          8403 => x"3f82d6d8",
          8404 => x"085b82d6",
          8405 => x"d80882eb",
          8406 => x"389c1908",
          8407 => x"70335555",
          8408 => x"73863884",
          8409 => x"5b82dc39",
          8410 => x"8b1533bf",
          8411 => x"067081ff",
          8412 => x"06585372",
          8413 => x"861a3482",
          8414 => x"d6d80856",
          8415 => x"7381e52e",
          8416 => x"09810683",
          8417 => x"38815682",
          8418 => x"d6d80853",
          8419 => x"73ae2e09",
          8420 => x"81068338",
          8421 => x"81537573",
          8422 => x"07537299",
          8423 => x"3882d6d8",
          8424 => x"0877df06",
          8425 => x"54567288",
          8426 => x"2e098106",
          8427 => x"83388156",
          8428 => x"757f2e87",
          8429 => x"3881ff5c",
          8430 => x"81ef3976",
          8431 => x"8f2e0981",
          8432 => x"0681ca38",
          8433 => x"73862a70",
          8434 => x"81065153",
          8435 => x"72802e92",
          8436 => x"388d1533",
          8437 => x"7481bf06",
          8438 => x"70901c08",
          8439 => x"ac1d0c56",
          8440 => x"5d5d737c",
          8441 => x"2e098106",
          8442 => x"819c388d",
          8443 => x"1533537c",
          8444 => x"732e0981",
          8445 => x"06818f38",
          8446 => x"8c1e089a",
          8447 => x"16525ae8",
          8448 => x"cc3f82d6",
          8449 => x"d80883ff",
          8450 => x"ff065372",
          8451 => x"80f83874",
          8452 => x"337081bf",
          8453 => x"068d29f3",
          8454 => x"05515481",
          8455 => x"7b585882",
          8456 => x"c7d41733",
          8457 => x"750551e8",
          8458 => x"a43f82d6",
          8459 => x"d80883ff",
          8460 => x"ff065677",
          8461 => x"802e9638",
          8462 => x"7381fe26",
          8463 => x"80c83873",
          8464 => x"101a7659",
          8465 => x"53757323",
          8466 => x"8114548b",
          8467 => x"397583ff",
          8468 => x"ff2e0981",
          8469 => x"06b03881",
          8470 => x"17578c77",
          8471 => x"27c13874",
          8472 => x"3370862a",
          8473 => x"70810651",
          8474 => x"54557280",
          8475 => x"2e8e3873",
          8476 => x"81fe2692",
          8477 => x"3873101a",
          8478 => x"53807323",
          8479 => x"ff1c7081",
          8480 => x"ff065153",
          8481 => x"843981ff",
          8482 => x"53725c9d",
          8483 => x"397b9338",
          8484 => x"7451fce8",
          8485 => x"3f82d6d8",
          8486 => x"0881ff06",
          8487 => x"53727d2e",
          8488 => x"a738ff0b",
          8489 => x"ac1a0ca0",
          8490 => x"39805278",
          8491 => x"51f8d23f",
          8492 => x"82d6d808",
          8493 => x"5b82d6d8",
          8494 => x"08893898",
          8495 => x"1908fd84",
          8496 => x"38863980",
          8497 => x"0b981a0c",
          8498 => x"7a82d6d8",
          8499 => x"0c903d0d",
          8500 => x"04f23d0d",
          8501 => x"60700840",
          8502 => x"59805278",
          8503 => x"51f6d73f",
          8504 => x"82d6d808",
          8505 => x"5882d6d8",
          8506 => x"0883a438",
          8507 => x"81ff705f",
          8508 => x"5cff0bac",
          8509 => x"1a0c9819",
          8510 => x"08527e51",
          8511 => x"eaa93f82",
          8512 => x"d6d80858",
          8513 => x"82d6d808",
          8514 => x"8385389c",
          8515 => x"19087033",
          8516 => x"57577586",
          8517 => x"38845882",
          8518 => x"f6398b17",
          8519 => x"33bf0670",
          8520 => x"81ff0656",
          8521 => x"5473861a",
          8522 => x"347581e5",
          8523 => x"2e82c338",
          8524 => x"74832a70",
          8525 => x"81065154",
          8526 => x"748f2e8e",
          8527 => x"387382b2",
          8528 => x"38748f2e",
          8529 => x"09810681",
          8530 => x"f738ab19",
          8531 => x"3370862a",
          8532 => x"70810651",
          8533 => x"55557382",
          8534 => x"a1387586",
          8535 => x"2a708106",
          8536 => x"51547380",
          8537 => x"2e92388d",
          8538 => x"17337681",
          8539 => x"bf067090",
          8540 => x"1c08ac1d",
          8541 => x"0c585d5e",
          8542 => x"757c2e09",
          8543 => x"810681b9",
          8544 => x"388d1733",
          8545 => x"567d762e",
          8546 => x"09810681",
          8547 => x"ac388c1f",
          8548 => x"089a1852",
          8549 => x"5de5b63f",
          8550 => x"82d6d808",
          8551 => x"83ffff06",
          8552 => x"55748195",
          8553 => x"38763370",
          8554 => x"bf068d29",
          8555 => x"f3055956",
          8556 => x"81755c5a",
          8557 => x"82c7d41b",
          8558 => x"33770551",
          8559 => x"e58f3f82",
          8560 => x"d6d80883",
          8561 => x"ffff0656",
          8562 => x"79802eb1",
          8563 => x"387781fe",
          8564 => x"2680e638",
          8565 => x"755180df",
          8566 => x"b43f82d6",
          8567 => x"d8087810",
          8568 => x"1e702253",
          8569 => x"55811959",
          8570 => x"5580dfa1",
          8571 => x"3f7482d6",
          8572 => x"d8082e09",
          8573 => x"810680c1",
          8574 => x"38755a8b",
          8575 => x"397583ff",
          8576 => x"ff2e0981",
          8577 => x"06b33881",
          8578 => x"1b5b8c7b",
          8579 => x"27ffa538",
          8580 => x"76337086",
          8581 => x"2a708106",
          8582 => x"51555779",
          8583 => x"802e9038",
          8584 => x"73802e8b",
          8585 => x"3877101d",
          8586 => x"70225154",
          8587 => x"738b38ff",
          8588 => x"1c7081ff",
          8589 => x"06515484",
          8590 => x"3981ff54",
          8591 => x"735cbb39",
          8592 => x"7b933876",
          8593 => x"51f9b53f",
          8594 => x"82d6d808",
          8595 => x"81ff0654",
          8596 => x"737e2ebb",
          8597 => x"38ab1933",
          8598 => x"81065473",
          8599 => x"95388b53",
          8600 => x"a019529c",
          8601 => x"190851e5",
          8602 => x"b03f82d6",
          8603 => x"d808802e",
          8604 => x"9e3881ff",
          8605 => x"5cff0bac",
          8606 => x"1a0c8052",
          8607 => x"7851f581",
          8608 => x"3f82d6d8",
          8609 => x"085882d6",
          8610 => x"d808802e",
          8611 => x"fce83877",
          8612 => x"82d6d80c",
          8613 => x"903d0d04",
          8614 => x"ee3d0d64",
          8615 => x"7008ab12",
          8616 => x"3381a006",
          8617 => x"565d5a86",
          8618 => x"557385b5",
          8619 => x"38738c1d",
          8620 => x"08702256",
          8621 => x"565d7380",
          8622 => x"2e8d3881",
          8623 => x"1d701016",
          8624 => x"70225155",
          8625 => x"5df0398c",
          8626 => x"53a01a70",
          8627 => x"53923d70",
          8628 => x"535f59e4",
          8629 => x"873f0280",
          8630 => x"cb053381",
          8631 => x"06547380",
          8632 => x"2e82a838",
          8633 => x"80c00bab",
          8634 => x"1b34815b",
          8635 => x"8c1c087b",
          8636 => x"56588b53",
          8637 => x"7d527851",
          8638 => x"e3e23f85",
          8639 => x"7b2780c6",
          8640 => x"387a5677",
          8641 => x"227083ff",
          8642 => x"ff065555",
          8643 => x"73802eb4",
          8644 => x"387483ff",
          8645 => x"ff068219",
          8646 => x"59558f57",
          8647 => x"74810676",
          8648 => x"10077581",
          8649 => x"2a71902a",
          8650 => x"70810651",
          8651 => x"56565673",
          8652 => x"802e8738",
          8653 => x"7584a0a1",
          8654 => x"3256ff17",
          8655 => x"57768025",
          8656 => x"db38c039",
          8657 => x"75558702",
          8658 => x"8405bf05",
          8659 => x"575774b0",
          8660 => x"07bf0654",
          8661 => x"b9742784",
          8662 => x"38871454",
          8663 => x"737634ff",
          8664 => x"16ff1876",
          8665 => x"842a5758",
          8666 => x"5674e338",
          8667 => x"943dec05",
          8668 => x"175480fe",
          8669 => x"74348077",
          8670 => x"27b53878",
          8671 => x"335473a0",
          8672 => x"2ead3874",
          8673 => x"19703352",
          8674 => x"54e3e03f",
          8675 => x"82d6d808",
          8676 => x"802e8c38",
          8677 => x"ff175474",
          8678 => x"742e9438",
          8679 => x"81155581",
          8680 => x"15557477",
          8681 => x"27893874",
          8682 => x"19703351",
          8683 => x"54d03994",
          8684 => x"3d7705eb",
          8685 => x"05547815",
          8686 => x"81165658",
          8687 => x"a0567687",
          8688 => x"268a3881",
          8689 => x"17811570",
          8690 => x"33585557",
          8691 => x"75783487",
          8692 => x"7527e338",
          8693 => x"7951f9f9",
          8694 => x"3f82d6d8",
          8695 => x"088b3881",
          8696 => x"1b5b80e3",
          8697 => x"7b27fe84",
          8698 => x"3887557a",
          8699 => x"80e42e82",
          8700 => x"f03882d6",
          8701 => x"d8085582",
          8702 => x"d6d80884",
          8703 => x"2e098106",
          8704 => x"82df3802",
          8705 => x"80cb0533",
          8706 => x"ab1b3402",
          8707 => x"80cb0533",
          8708 => x"70812a70",
          8709 => x"81065155",
          8710 => x"5e815973",
          8711 => x"802e9038",
          8712 => x"8d528c1d",
          8713 => x"51fef886",
          8714 => x"3f82d6d8",
          8715 => x"08195978",
          8716 => x"527951f3",
          8717 => x"c53f82d6",
          8718 => x"d8085782",
          8719 => x"d6d80882",
          8720 => x"9e38ff19",
          8721 => x"5978802e",
          8722 => x"81d43878",
          8723 => x"852b901b",
          8724 => x"08713153",
          8725 => x"547951ef",
          8726 => x"dd3f82d6",
          8727 => x"d8085782",
          8728 => x"d6d80881",
          8729 => x"fa38a01a",
          8730 => x"51f5913f",
          8731 => x"82d6d808",
          8732 => x"81ff065d",
          8733 => x"981a0852",
          8734 => x"7b51e3ab",
          8735 => x"3f82d6d8",
          8736 => x"085782d6",
          8737 => x"d80881d7",
          8738 => x"388c1c08",
          8739 => x"9c1b087a",
          8740 => x"81ff065a",
          8741 => x"575b7c8d",
          8742 => x"17348f0b",
          8743 => x"8b173482",
          8744 => x"d6d8088c",
          8745 => x"173482d6",
          8746 => x"d808529a",
          8747 => x"1651dfdf",
          8748 => x"3f778d29",
          8749 => x"f3057755",
          8750 => x"557383ff",
          8751 => x"ff2e8b38",
          8752 => x"74101b70",
          8753 => x"22811757",
          8754 => x"51547352",
          8755 => x"82c7d417",
          8756 => x"33760551",
          8757 => x"dfb93f73",
          8758 => x"853883ff",
          8759 => x"ff548117",
          8760 => x"578c7727",
          8761 => x"d4387383",
          8762 => x"ffff2e8b",
          8763 => x"3874101b",
          8764 => x"70225154",
          8765 => x"73863877",
          8766 => x"80c00758",
          8767 => x"77763481",
          8768 => x"0b831d34",
          8769 => x"80527951",
          8770 => x"eff73f82",
          8771 => x"d6d80857",
          8772 => x"82d6d808",
          8773 => x"80c938ff",
          8774 => x"195978fe",
          8775 => x"d738981a",
          8776 => x"08527b51",
          8777 => x"e2813f82",
          8778 => x"d6d80857",
          8779 => x"82d6d808",
          8780 => x"ae38a053",
          8781 => x"82d6d808",
          8782 => x"529c1a08",
          8783 => x"51dfc03f",
          8784 => x"8b53a01a",
          8785 => x"529c1a08",
          8786 => x"51df913f",
          8787 => x"9c1a08ab",
          8788 => x"1b339806",
          8789 => x"5555738c",
          8790 => x"1634810b",
          8791 => x"831d3476",
          8792 => x"557482d6",
          8793 => x"d80c943d",
          8794 => x"0d04fa3d",
          8795 => x"0d787008",
          8796 => x"901208ac",
          8797 => x"13085659",
          8798 => x"575572ff",
          8799 => x"2e943872",
          8800 => x"527451ed",
          8801 => x"b13f82d6",
          8802 => x"d8085482",
          8803 => x"d6d80880",
          8804 => x"c9389815",
          8805 => x"08527551",
          8806 => x"e18d3f82",
          8807 => x"d6d80854",
          8808 => x"82d6d808",
          8809 => x"ab389c15",
          8810 => x"0853e573",
          8811 => x"34810b83",
          8812 => x"17349015",
          8813 => x"087727a2",
          8814 => x"3882d6d8",
          8815 => x"08527451",
          8816 => x"eebf3f82",
          8817 => x"d6d80854",
          8818 => x"82d6d808",
          8819 => x"802ec338",
          8820 => x"73842e09",
          8821 => x"81068338",
          8822 => x"82547382",
          8823 => x"d6d80c88",
          8824 => x"3d0d04f4",
          8825 => x"3d0d7e60",
          8826 => x"71085f59",
          8827 => x"5c800b96",
          8828 => x"1934981c",
          8829 => x"08802e83",
          8830 => x"e238ac1c",
          8831 => x"08ff2e81",
          8832 => x"bb388070",
          8833 => x"717f8c05",
          8834 => x"08702257",
          8835 => x"575b5c57",
          8836 => x"72772e81",
          8837 => x"9d387810",
          8838 => x"14702281",
          8839 => x"1b5b5653",
          8840 => x"7a973880",
          8841 => x"d0801570",
          8842 => x"83ffff06",
          8843 => x"5153728f",
          8844 => x"ff268638",
          8845 => x"745b80df",
          8846 => x"39761896",
          8847 => x"1181ff79",
          8848 => x"31585b54",
          8849 => x"83b5527a",
          8850 => x"902b7507",
          8851 => x"5180d598",
          8852 => x"3f82d6d8",
          8853 => x"0883ffff",
          8854 => x"065581ff",
          8855 => x"75279538",
          8856 => x"817627a5",
          8857 => x"3874882a",
          8858 => x"53727a34",
          8859 => x"74971534",
          8860 => x"82559f39",
          8861 => x"74307630",
          8862 => x"70780780",
          8863 => x"25728025",
          8864 => x"07525454",
          8865 => x"73802e85",
          8866 => x"3880579a",
          8867 => x"39747a34",
          8868 => x"81557417",
          8869 => x"57805b8c",
          8870 => x"1d087910",
          8871 => x"11702251",
          8872 => x"545472fe",
          8873 => x"f1387a30",
          8874 => x"70802570",
          8875 => x"30790659",
          8876 => x"51537717",
          8877 => x"94055380",
          8878 => x"0b821434",
          8879 => x"8070891a",
          8880 => x"585a579c",
          8881 => x"1c081970",
          8882 => x"33811b5b",
          8883 => x"565374a0",
          8884 => x"2eb73874",
          8885 => x"852e0981",
          8886 => x"06843881",
          8887 => x"e5557889",
          8888 => x"32703070",
          8889 => x"72078025",
          8890 => x"51545476",
          8891 => x"8b269038",
          8892 => x"72802e8b",
          8893 => x"38ae7670",
          8894 => x"81055834",
          8895 => x"81175774",
          8896 => x"76708105",
          8897 => x"58348117",
          8898 => x"578a7927",
          8899 => x"ffb53877",
          8900 => x"17880553",
          8901 => x"800b8114",
          8902 => x"34961833",
          8903 => x"53728187",
          8904 => x"38768b38",
          8905 => x"bf0b9619",
          8906 => x"34815780",
          8907 => x"e1397273",
          8908 => x"891a3355",
          8909 => x"5a577280",
          8910 => x"2e80d338",
          8911 => x"96188919",
          8912 => x"55567333",
          8913 => x"ffbf1154",
          8914 => x"55729926",
          8915 => x"aa389c1c",
          8916 => x"088c1133",
          8917 => x"51538879",
          8918 => x"27873872",
          8919 => x"842a5385",
          8920 => x"3972832a",
          8921 => x"53728106",
          8922 => x"5372802e",
          8923 => x"8a38a015",
          8924 => x"7083ffff",
          8925 => x"06565374",
          8926 => x"76708105",
          8927 => x"58348119",
          8928 => x"81158119",
          8929 => x"71335659",
          8930 => x"555972ff",
          8931 => x"b5387717",
          8932 => x"94055380",
          8933 => x"0b821434",
          8934 => x"9c1c088c",
          8935 => x"11335153",
          8936 => x"72853872",
          8937 => x"8919349c",
          8938 => x"1c08538b",
          8939 => x"13338819",
          8940 => x"349c1c08",
          8941 => x"9c115253",
          8942 => x"d9aa3f82",
          8943 => x"d6d80878",
          8944 => x"0c961351",
          8945 => x"d9873f82",
          8946 => x"d6d80886",
          8947 => x"19239813",
          8948 => x"51d8fa3f",
          8949 => x"82d6d808",
          8950 => x"8419238e",
          8951 => x"3d0d04f0",
          8952 => x"3d0d6270",
          8953 => x"08415e80",
          8954 => x"64703351",
          8955 => x"555573af",
          8956 => x"2e833881",
          8957 => x"557380dc",
          8958 => x"2e923874",
          8959 => x"802e8d38",
          8960 => x"7f980508",
          8961 => x"881f0caa",
          8962 => x"39811544",
          8963 => x"80647033",
          8964 => x"56565673",
          8965 => x"af2e0981",
          8966 => x"06833881",
          8967 => x"567380dc",
          8968 => x"32703070",
          8969 => x"80257807",
          8970 => x"51515473",
          8971 => x"dc387388",
          8972 => x"1f0c6370",
          8973 => x"33515473",
          8974 => x"9f269638",
          8975 => x"ff800bab",
          8976 => x"1f348052",
          8977 => x"7d51e7ee",
          8978 => x"3f82d6d8",
          8979 => x"085687e1",
          8980 => x"3963417d",
          8981 => x"088c1108",
          8982 => x"5b548059",
          8983 => x"923dfc05",
          8984 => x"51da8f3f",
          8985 => x"82d6d808",
          8986 => x"ff2e82b1",
          8987 => x"3883ffff",
          8988 => x"0b82d6d8",
          8989 => x"08279238",
          8990 => x"78101a82",
          8991 => x"d6d80890",
          8992 => x"2a555573",
          8993 => x"75238119",
          8994 => x"5982d6d8",
          8995 => x"0883ffff",
          8996 => x"0670af32",
          8997 => x"70309f73",
          8998 => x"27718025",
          8999 => x"07515155",
          9000 => x"5673b438",
          9001 => x"7580dc2e",
          9002 => x"ae387580",
          9003 => x"ff269138",
          9004 => x"755282c6",
          9005 => x"f051d992",
          9006 => x"3f82d6d8",
          9007 => x"0881de38",
          9008 => x"7881fe26",
          9009 => x"81d73878",
          9010 => x"101a5475",
          9011 => x"74238119",
          9012 => x"59ff8939",
          9013 => x"81154180",
          9014 => x"61703356",
          9015 => x"565773af",
          9016 => x"2e098106",
          9017 => x"83388157",
          9018 => x"7380dc32",
          9019 => x"70307080",
          9020 => x"25790751",
          9021 => x"515473dc",
          9022 => x"3874449f",
          9023 => x"7627822b",
          9024 => x"5778812e",
          9025 => x"0981068c",
          9026 => x"38792254",
          9027 => x"73ae2ea5",
          9028 => x"3880d239",
          9029 => x"78822e09",
          9030 => x"810680c9",
          9031 => x"38821a22",
          9032 => x"5473ae2e",
          9033 => x"09810680",
          9034 => x"c1387922",
          9035 => x"5473ae2e",
          9036 => x"098106b6",
          9037 => x"3878101a",
          9038 => x"54807423",
          9039 => x"800ba01f",
          9040 => x"5658ae54",
          9041 => x"78782683",
          9042 => x"38a05473",
          9043 => x"75708105",
          9044 => x"57348118",
          9045 => x"588a7827",
          9046 => x"e93876a0",
          9047 => x"075473ab",
          9048 => x"1f3484c4",
          9049 => x"3978802e",
          9050 => x"a8387810",
          9051 => x"1afe0555",
          9052 => x"7422fe16",
          9053 => x"7172a032",
          9054 => x"7030709f",
          9055 => x"2a515153",
          9056 => x"58565475",
          9057 => x"ae2e8438",
          9058 => x"738738ff",
          9059 => x"195978e0",
          9060 => x"3878197a",
          9061 => x"11555680",
          9062 => x"7423788d",
          9063 => x"38865685",
          9064 => x"90397683",
          9065 => x"07578399",
          9066 => x"39807a22",
          9067 => x"7083ffff",
          9068 => x"0656565d",
          9069 => x"73a02e09",
          9070 => x"81069338",
          9071 => x"811d7010",
          9072 => x"1b702251",
          9073 => x"555d73a0",
          9074 => x"2ef2387c",
          9075 => x"8f387483",
          9076 => x"ffff0654",
          9077 => x"73ae2e09",
          9078 => x"81068538",
          9079 => x"76830757",
          9080 => x"78802eaa",
          9081 => x"387916fe",
          9082 => x"05702251",
          9083 => x"5473ae2e",
          9084 => x"9d387810",
          9085 => x"1afe0555",
          9086 => x"ff195978",
          9087 => x"802e8f38",
          9088 => x"fe157022",
          9089 => x"555573ae",
          9090 => x"2e098106",
          9091 => x"eb388b53",
          9092 => x"a052a01e",
          9093 => x"51d5e83f",
          9094 => x"8070595c",
          9095 => x"885f7c10",
          9096 => x"1a702281",
          9097 => x"1f5f5754",
          9098 => x"75802e82",
          9099 => x"943875a0",
          9100 => x"2e963875",
          9101 => x"ae327030",
          9102 => x"70802551",
          9103 => x"51547c79",
          9104 => x"2e8c3873",
          9105 => x"802e8938",
          9106 => x"76830757",
          9107 => x"d1398054",
          9108 => x"735b7e78",
          9109 => x"26833881",
          9110 => x"5b7c7932",
          9111 => x"70307072",
          9112 => x"07802570",
          9113 => x"7e075151",
          9114 => x"55557380",
          9115 => x"2ea6387e",
          9116 => x"8b2efeae",
          9117 => x"387c792e",
          9118 => x"8b387683",
          9119 => x"07577c79",
          9120 => x"2681be38",
          9121 => x"785d8858",
          9122 => x"8b7c822b",
          9123 => x"81fc065d",
          9124 => x"5fff8b39",
          9125 => x"80ff7627",
          9126 => x"af387682",
          9127 => x"075783b5",
          9128 => x"52755180",
          9129 => x"ccc23f82",
          9130 => x"d6d80883",
          9131 => x"ffff0670",
          9132 => x"872a7081",
          9133 => x"06515556",
          9134 => x"73802e8c",
          9135 => x"387580ff",
          9136 => x"0682c7e4",
          9137 => x"11335754",
          9138 => x"81ff7627",
          9139 => x"a438ff1f",
          9140 => x"54737826",
          9141 => x"8a387683",
          9142 => x"077f5957",
          9143 => x"fec0397d",
          9144 => x"18a00576",
          9145 => x"882a5555",
          9146 => x"73753481",
          9147 => x"185880c3",
          9148 => x"3975802e",
          9149 => x"92387552",
          9150 => x"82c6fc51",
          9151 => x"d4cc3f82",
          9152 => x"d6d80880",
          9153 => x"2e8a3880",
          9154 => x"df778307",
          9155 => x"5856a439",
          9156 => x"ffbf1654",
          9157 => x"73992685",
          9158 => x"387b8207",
          9159 => x"5cff9f16",
          9160 => x"54739926",
          9161 => x"8e387b81",
          9162 => x"07e01770",
          9163 => x"83ffff06",
          9164 => x"58555c7d",
          9165 => x"18a00554",
          9166 => x"75743481",
          9167 => x"1858fdde",
          9168 => x"39a01e33",
          9169 => x"547381e5",
          9170 => x"2e098106",
          9171 => x"8638850b",
          9172 => x"a01f347e",
          9173 => x"882e0981",
          9174 => x"0688387b",
          9175 => x"822b81fc",
          9176 => x"065c7b8c",
          9177 => x"0654738c",
          9178 => x"2e8d387b",
          9179 => x"83065473",
          9180 => x"832e0981",
          9181 => x"06853876",
          9182 => x"82075776",
          9183 => x"812a7081",
          9184 => x"06515473",
          9185 => x"9f387b81",
          9186 => x"06547380",
          9187 => x"2e853876",
          9188 => x"9007577b",
          9189 => x"822a7081",
          9190 => x"06515473",
          9191 => x"802e8538",
          9192 => x"76880757",
          9193 => x"76ab1f34",
          9194 => x"7d51eaa5",
          9195 => x"3f82d6d8",
          9196 => x"08ab1f33",
          9197 => x"565682d6",
          9198 => x"d808802e",
          9199 => x"be3882d6",
          9200 => x"d808842e",
          9201 => x"09810680",
          9202 => x"e8387485",
          9203 => x"2a708106",
          9204 => x"76822a57",
          9205 => x"51547380",
          9206 => x"2e963874",
          9207 => x"81065473",
          9208 => x"802ef8ed",
          9209 => x"38ff800b",
          9210 => x"ab1f3480",
          9211 => x"5680c239",
          9212 => x"74810654",
          9213 => x"73bb3885",
          9214 => x"56b73974",
          9215 => x"822a7081",
          9216 => x"06515473",
          9217 => x"ac38861e",
          9218 => x"3370842a",
          9219 => x"70810651",
          9220 => x"55557380",
          9221 => x"2ee13890",
          9222 => x"1e0883ff",
          9223 => x"066005b8",
          9224 => x"05527f51",
          9225 => x"e4ef3f82",
          9226 => x"d6d80888",
          9227 => x"1f0cf8a1",
          9228 => x"397582d6",
          9229 => x"d80c923d",
          9230 => x"0d04f63d",
          9231 => x"0d7c5bff",
          9232 => x"7b087071",
          9233 => x"7355595c",
          9234 => x"55597380",
          9235 => x"2e81c638",
          9236 => x"75708105",
          9237 => x"5733709f",
          9238 => x"26525271",
          9239 => x"ba2e8d38",
          9240 => x"70ee3871",
          9241 => x"ba2e0981",
          9242 => x"0681a538",
          9243 => x"7333d011",
          9244 => x"7081ff06",
          9245 => x"51525370",
          9246 => x"89269138",
          9247 => x"82147381",
          9248 => x"ff06d005",
          9249 => x"56527176",
          9250 => x"2e80f738",
          9251 => x"800b82c7",
          9252 => x"c4595577",
          9253 => x"087a5557",
          9254 => x"76708105",
          9255 => x"58337470",
          9256 => x"81055633",
          9257 => x"ff9f1253",
          9258 => x"53537099",
          9259 => x"268938e0",
          9260 => x"137081ff",
          9261 => x"065451ff",
          9262 => x"9f125170",
          9263 => x"99268938",
          9264 => x"e0127081",
          9265 => x"ff065351",
          9266 => x"7230709f",
          9267 => x"2a515172",
          9268 => x"722e0981",
          9269 => x"06853870",
          9270 => x"ffbe3872",
          9271 => x"30747732",
          9272 => x"70307072",
          9273 => x"079f2a73",
          9274 => x"9f2a0753",
          9275 => x"54545170",
          9276 => x"802e8f38",
          9277 => x"81158419",
          9278 => x"59558375",
          9279 => x"25ff9438",
          9280 => x"8b397483",
          9281 => x"24863874",
          9282 => x"767c0c59",
          9283 => x"78518639",
          9284 => x"82eeb433",
          9285 => x"517082d6",
          9286 => x"d80c8c3d",
          9287 => x"0d04fa3d",
          9288 => x"0d785680",
          9289 => x"0b831734",
          9290 => x"ff0bb417",
          9291 => x"0c795275",
          9292 => x"51d1f43f",
          9293 => x"845582d6",
          9294 => x"d8088180",
          9295 => x"3884b616",
          9296 => x"51ce8a3f",
          9297 => x"82d6d808",
          9298 => x"83ffff06",
          9299 => x"54835573",
          9300 => x"82d4d52e",
          9301 => x"09810680",
          9302 => x"e338800b",
          9303 => x"b8173356",
          9304 => x"577481e9",
          9305 => x"2e098106",
          9306 => x"83388157",
          9307 => x"7481eb32",
          9308 => x"70307080",
          9309 => x"25790751",
          9310 => x"5154738a",
          9311 => x"387481e8",
          9312 => x"2e098106",
          9313 => x"b5388353",
          9314 => x"82c78452",
          9315 => x"80ee1651",
          9316 => x"cf873f82",
          9317 => x"d6d80855",
          9318 => x"82d6d808",
          9319 => x"802e9d38",
          9320 => x"855382c7",
          9321 => x"8852818a",
          9322 => x"1651ceed",
          9323 => x"3f82d6d8",
          9324 => x"085582d6",
          9325 => x"d808802e",
          9326 => x"83388255",
          9327 => x"7482d6d8",
          9328 => x"0c883d0d",
          9329 => x"04f23d0d",
          9330 => x"61028405",
          9331 => x"80cb0533",
          9332 => x"58558075",
          9333 => x"0c6051fc",
          9334 => x"e13f82d6",
          9335 => x"d808588b",
          9336 => x"56800b82",
          9337 => x"d6d80824",
          9338 => x"87843882",
          9339 => x"d6d80884",
          9340 => x"2982eea0",
          9341 => x"05700855",
          9342 => x"538c5673",
          9343 => x"802e86ee",
          9344 => x"3873750c",
          9345 => x"7681fe06",
          9346 => x"74335457",
          9347 => x"72802eae",
          9348 => x"38811433",
          9349 => x"51c6a03f",
          9350 => x"82d6d808",
          9351 => x"81ff0670",
          9352 => x"81065455",
          9353 => x"72983876",
          9354 => x"802e86c0",
          9355 => x"3874822a",
          9356 => x"70810651",
          9357 => x"538a5672",
          9358 => x"86b43886",
          9359 => x"af398074",
          9360 => x"34778115",
          9361 => x"34815281",
          9362 => x"143351c6",
          9363 => x"883f82d6",
          9364 => x"d80881ff",
          9365 => x"06708106",
          9366 => x"54558356",
          9367 => x"72868f38",
          9368 => x"76802e8f",
          9369 => x"3874822a",
          9370 => x"70810651",
          9371 => x"538a5672",
          9372 => x"85fc3880",
          9373 => x"70537452",
          9374 => x"5bfda33f",
          9375 => x"82d6d808",
          9376 => x"81ff0657",
          9377 => x"76822e09",
          9378 => x"810680e2",
          9379 => x"388c3d74",
          9380 => x"56588356",
          9381 => x"83fa1533",
          9382 => x"70585372",
          9383 => x"802e8d38",
          9384 => x"83fe1551",
          9385 => x"cbbe3f82",
          9386 => x"d6d80857",
          9387 => x"76787084",
          9388 => x"055a0cff",
          9389 => x"16901656",
          9390 => x"56758025",
          9391 => x"d738800b",
          9392 => x"8d3d5456",
          9393 => x"72708405",
          9394 => x"54085b83",
          9395 => x"577a802e",
          9396 => x"95387a52",
          9397 => x"7351fcc6",
          9398 => x"3f82d6d8",
          9399 => x"0881ff06",
          9400 => x"57817727",
          9401 => x"89388116",
          9402 => x"56837627",
          9403 => x"d7388156",
          9404 => x"76842e84",
          9405 => x"f9388d56",
          9406 => x"76812684",
          9407 => x"f13880c3",
          9408 => x"1451cac9",
          9409 => x"3f82d6d8",
          9410 => x"0883ffff",
          9411 => x"06537284",
          9412 => x"802e0981",
          9413 => x"0684d738",
          9414 => x"80ce1451",
          9415 => x"caaf3f82",
          9416 => x"d6d80883",
          9417 => x"ffff0658",
          9418 => x"778d3880",
          9419 => x"dc1451ca",
          9420 => x"b33f82d6",
          9421 => x"d8085877",
          9422 => x"a0150c80",
          9423 => x"c8143382",
          9424 => x"153480c8",
          9425 => x"1433ff11",
          9426 => x"7081ff06",
          9427 => x"5154558d",
          9428 => x"56728126",
          9429 => x"84983874",
          9430 => x"81ff0678",
          9431 => x"712980c5",
          9432 => x"16335259",
          9433 => x"53728a15",
          9434 => x"2372802e",
          9435 => x"8b38ff13",
          9436 => x"73065372",
          9437 => x"802e8638",
          9438 => x"8d5683f2",
          9439 => x"3980c914",
          9440 => x"51c9ca3f",
          9441 => x"82d6d808",
          9442 => x"5382d6d8",
          9443 => x"08881523",
          9444 => x"728f0657",
          9445 => x"8d567683",
          9446 => x"d53880cb",
          9447 => x"1451c9ad",
          9448 => x"3f82d6d8",
          9449 => x"0883ffff",
          9450 => x"0655748d",
          9451 => x"3880d814",
          9452 => x"51c9b13f",
          9453 => x"82d6d808",
          9454 => x"5580c614",
          9455 => x"51c98e3f",
          9456 => x"82d6d808",
          9457 => x"83ffff06",
          9458 => x"538d5672",
          9459 => x"802e839e",
          9460 => x"38881422",
          9461 => x"78147184",
          9462 => x"2a055a5a",
          9463 => x"78752683",
          9464 => x"8d388a14",
          9465 => x"22527479",
          9466 => x"3151fee0",
          9467 => x"c13f82d6",
          9468 => x"d8085582",
          9469 => x"d6d80880",
          9470 => x"2e82f338",
          9471 => x"82d6d808",
          9472 => x"80ffffff",
          9473 => x"f5268338",
          9474 => x"83577483",
          9475 => x"fff52683",
          9476 => x"38825774",
          9477 => x"9ff52685",
          9478 => x"38815789",
          9479 => x"398d5676",
          9480 => x"802e82ca",
          9481 => x"38821570",
          9482 => x"9c160c7b",
          9483 => x"a4160c73",
          9484 => x"1c70a817",
          9485 => x"0c7a1db0",
          9486 => x"170c5455",
          9487 => x"76832e09",
          9488 => x"8106af38",
          9489 => x"80e21451",
          9490 => x"c8833f82",
          9491 => x"d6d80883",
          9492 => x"ffff0653",
          9493 => x"8d567282",
          9494 => x"95387982",
          9495 => x"913880e4",
          9496 => x"1451c880",
          9497 => x"3f82d6d8",
          9498 => x"08ac150c",
          9499 => x"74822b53",
          9500 => x"a2398d56",
          9501 => x"79802e81",
          9502 => x"f5387713",
          9503 => x"ac150c74",
          9504 => x"15537682",
          9505 => x"2e8d3874",
          9506 => x"10157081",
          9507 => x"2a768106",
          9508 => x"05515383",
          9509 => x"ff13892a",
          9510 => x"538d5672",
          9511 => x"a0150826",
          9512 => x"81cc38ff",
          9513 => x"0b94150c",
          9514 => x"ff0b9015",
          9515 => x"0cff800b",
          9516 => x"84153476",
          9517 => x"832e0981",
          9518 => x"06819238",
          9519 => x"80e81451",
          9520 => x"c78b3f82",
          9521 => x"d6d80883",
          9522 => x"ffff0653",
          9523 => x"72812e09",
          9524 => x"810680f9",
          9525 => x"38811b52",
          9526 => x"7351cacb",
          9527 => x"3f82d6d8",
          9528 => x"0880ea38",
          9529 => x"82d6d808",
          9530 => x"84153484",
          9531 => x"b61451c6",
          9532 => x"dc3f82d6",
          9533 => x"d80883ff",
          9534 => x"ff065372",
          9535 => x"82d4d52e",
          9536 => x"09810680",
          9537 => x"c838b814",
          9538 => x"51c6d93f",
          9539 => x"82d6d808",
          9540 => x"848b85a4",
          9541 => x"d22e0981",
          9542 => x"06b33884",
          9543 => x"9c1451c6",
          9544 => x"c33f82d6",
          9545 => x"d808868a",
          9546 => x"85e4f22e",
          9547 => x"0981069d",
          9548 => x"3884a014",
          9549 => x"51c6ad3f",
          9550 => x"82d6d808",
          9551 => x"94150c84",
          9552 => x"a41451c6",
          9553 => x"9f3f82d6",
          9554 => x"d8089015",
          9555 => x"0c767434",
          9556 => x"82eeb022",
          9557 => x"81055372",
          9558 => x"82eeb023",
          9559 => x"72861523",
          9560 => x"82eeb80b",
          9561 => x"8c150c80",
          9562 => x"0b98150c",
          9563 => x"80567582",
          9564 => x"d6d80c90",
          9565 => x"3d0d04fb",
          9566 => x"3d0d7754",
          9567 => x"89557380",
          9568 => x"2eba3873",
          9569 => x"08537280",
          9570 => x"2eb23872",
          9571 => x"33527180",
          9572 => x"2eaa3886",
          9573 => x"13228415",
          9574 => x"22575271",
          9575 => x"762e0981",
          9576 => x"069a3881",
          9577 => x"133351ff",
          9578 => x"bf8d3f82",
          9579 => x"d6d80881",
          9580 => x"06527188",
          9581 => x"38717408",
          9582 => x"54558339",
          9583 => x"80537873",
          9584 => x"710c5274",
          9585 => x"82d6d80c",
          9586 => x"873d0d04",
          9587 => x"fa3d0d02",
          9588 => x"ab05337a",
          9589 => x"58893dfc",
          9590 => x"055256f4",
          9591 => x"dd3f8b54",
          9592 => x"800b82d6",
          9593 => x"d80824bc",
          9594 => x"3882d6d8",
          9595 => x"08842982",
          9596 => x"eea00570",
          9597 => x"08555573",
          9598 => x"802e8438",
          9599 => x"80743478",
          9600 => x"5473802e",
          9601 => x"84388074",
          9602 => x"3478750c",
          9603 => x"75547580",
          9604 => x"2e923880",
          9605 => x"53893d70",
          9606 => x"53840551",
          9607 => x"f7a73f82",
          9608 => x"d6d80854",
          9609 => x"7382d6d8",
          9610 => x"0c883d0d",
          9611 => x"04ea3d0d",
          9612 => x"68028405",
          9613 => x"80eb0533",
          9614 => x"59598954",
          9615 => x"78802e84",
          9616 => x"c83877bf",
          9617 => x"06705499",
          9618 => x"3dcc0553",
          9619 => x"9a3d8405",
          9620 => x"5258f6f1",
          9621 => x"3f82d6d8",
          9622 => x"085582d6",
          9623 => x"d80884a4",
          9624 => x"387a5c69",
          9625 => x"528c3d70",
          9626 => x"5256eaf3",
          9627 => x"3f82d6d8",
          9628 => x"085582d6",
          9629 => x"d8089238",
          9630 => x"0280d705",
          9631 => x"3370982b",
          9632 => x"55577380",
          9633 => x"25833886",
          9634 => x"55779c06",
          9635 => x"5473802e",
          9636 => x"81ab3874",
          9637 => x"802e9538",
          9638 => x"74842e09",
          9639 => x"8106aa38",
          9640 => x"7551dff4",
          9641 => x"3f82d6d8",
          9642 => x"08559e39",
          9643 => x"02b20533",
          9644 => x"91065473",
          9645 => x"81b83877",
          9646 => x"822a7081",
          9647 => x"06515473",
          9648 => x"802e8e38",
          9649 => x"885583bc",
          9650 => x"39778807",
          9651 => x"587483b4",
          9652 => x"3877832a",
          9653 => x"70810651",
          9654 => x"5473802e",
          9655 => x"81af3862",
          9656 => x"527a51d7",
          9657 => x"b03f82d6",
          9658 => x"d8085682",
          9659 => x"88b20a52",
          9660 => x"628e0551",
          9661 => x"c3b73f62",
          9662 => x"54a00b8b",
          9663 => x"15348053",
          9664 => x"62527a51",
          9665 => x"d7c83f80",
          9666 => x"52629c05",
          9667 => x"51c39e3f",
          9668 => x"7a54810b",
          9669 => x"83153475",
          9670 => x"802e80f1",
          9671 => x"387ab411",
          9672 => x"08515480",
          9673 => x"53755298",
          9674 => x"3dd00551",
          9675 => x"ccc93f82",
          9676 => x"d6d80855",
          9677 => x"82d6d808",
          9678 => x"82ca38b7",
          9679 => x"397482c4",
          9680 => x"3802b205",
          9681 => x"3370842a",
          9682 => x"70810651",
          9683 => x"55567380",
          9684 => x"2e863884",
          9685 => x"5582ad39",
          9686 => x"77812a70",
          9687 => x"81065154",
          9688 => x"73802ea9",
          9689 => x"38758106",
          9690 => x"5473802e",
          9691 => x"a0388755",
          9692 => x"82923973",
          9693 => x"527a51c5",
          9694 => x"ae3f82d6",
          9695 => x"d8087bff",
          9696 => x"1890120c",
          9697 => x"555582d6",
          9698 => x"d80881f8",
          9699 => x"3877832a",
          9700 => x"70810651",
          9701 => x"5473802e",
          9702 => x"86387780",
          9703 => x"c007587a",
          9704 => x"b41108a0",
          9705 => x"1b0c63a4",
          9706 => x"1b0c6353",
          9707 => x"705257d5",
          9708 => x"e43f82d6",
          9709 => x"d80882d6",
          9710 => x"d808881b",
          9711 => x"0c639c05",
          9712 => x"525ac1a0",
          9713 => x"3f82d6d8",
          9714 => x"0882d6d8",
          9715 => x"088c1b0c",
          9716 => x"777a0c56",
          9717 => x"86172284",
          9718 => x"1a237790",
          9719 => x"1a34800b",
          9720 => x"911a3480",
          9721 => x"0b9c1a0c",
          9722 => x"800b941a",
          9723 => x"0c77852a",
          9724 => x"70810651",
          9725 => x"5473802e",
          9726 => x"818d3882",
          9727 => x"d6d80880",
          9728 => x"2e818438",
          9729 => x"82d6d808",
          9730 => x"941a0c8a",
          9731 => x"17227089",
          9732 => x"2b7b5259",
          9733 => x"57a83976",
          9734 => x"527851c6",
          9735 => x"aa3f82d6",
          9736 => x"d8085782",
          9737 => x"d6d80881",
          9738 => x"26833882",
          9739 => x"5582d6d8",
          9740 => x"08ff2e09",
          9741 => x"81068338",
          9742 => x"79557578",
          9743 => x"31567430",
          9744 => x"70760780",
          9745 => x"25515477",
          9746 => x"76278a38",
          9747 => x"81707506",
          9748 => x"555a73c3",
          9749 => x"3876981a",
          9750 => x"0c74a938",
          9751 => x"7583ff06",
          9752 => x"5473802e",
          9753 => x"a2387652",
          9754 => x"7a51c5b1",
          9755 => x"3f82d6d8",
          9756 => x"08853882",
          9757 => x"558e3975",
          9758 => x"892a82d6",
          9759 => x"d808059c",
          9760 => x"1a0c8439",
          9761 => x"80790c74",
          9762 => x"547382d6",
          9763 => x"d80c983d",
          9764 => x"0d04f23d",
          9765 => x"0d606365",
          9766 => x"6440405d",
          9767 => x"59807e0c",
          9768 => x"903dfc05",
          9769 => x"527851f9",
          9770 => x"ce3f82d6",
          9771 => x"d8085582",
          9772 => x"d6d8088a",
          9773 => x"38911933",
          9774 => x"5574802e",
          9775 => x"86387456",
          9776 => x"82c73990",
          9777 => x"19338106",
          9778 => x"55875674",
          9779 => x"802e82b9",
          9780 => x"38953982",
          9781 => x"0b911a34",
          9782 => x"825682ad",
          9783 => x"39810b91",
          9784 => x"1a348156",
          9785 => x"82a3398c",
          9786 => x"1908941a",
          9787 => x"08315574",
          9788 => x"7c278338",
          9789 => x"745c7b80",
          9790 => x"2e828c38",
          9791 => x"94190870",
          9792 => x"83ff0656",
          9793 => x"567481b4",
          9794 => x"387e8a11",
          9795 => x"22ff0577",
          9796 => x"892a065b",
          9797 => x"5579a838",
          9798 => x"75873888",
          9799 => x"1908558f",
          9800 => x"39981908",
          9801 => x"527851c4",
          9802 => x"9e3f82d6",
          9803 => x"d8085581",
          9804 => x"7527ff9f",
          9805 => x"3874ff2e",
          9806 => x"ffa33874",
          9807 => x"981a0c98",
          9808 => x"1908527e",
          9809 => x"51c3d63f",
          9810 => x"82d6d808",
          9811 => x"802eff83",
          9812 => x"3882d6d8",
          9813 => x"081a7c89",
          9814 => x"2a595777",
          9815 => x"802e80d8",
          9816 => x"38771a7f",
          9817 => x"8a112258",
          9818 => x"5c557575",
          9819 => x"27853875",
          9820 => x"7a315877",
          9821 => x"5476537c",
          9822 => x"52811b33",
          9823 => x"51ffb8d4",
          9824 => x"3f82d6d8",
          9825 => x"08fed638",
          9826 => x"7e831133",
          9827 => x"56567480",
          9828 => x"2ea038b4",
          9829 => x"16087731",
          9830 => x"55747827",
          9831 => x"95388480",
          9832 => x"53b81652",
          9833 => x"b4160877",
          9834 => x"31892b7d",
          9835 => x"0551ffbe",
          9836 => x"ab3f7789",
          9837 => x"2b56ba39",
          9838 => x"769c1a0c",
          9839 => x"94190883",
          9840 => x"ff068480",
          9841 => x"71315755",
          9842 => x"7b762783",
          9843 => x"387b569c",
          9844 => x"1908527e",
          9845 => x"51c0d03f",
          9846 => x"82d6d808",
          9847 => x"fdff3875",
          9848 => x"53941908",
          9849 => x"83ff061f",
          9850 => x"b805527c",
          9851 => x"51ffbdec",
          9852 => x"3f7b7631",
          9853 => x"7e08177f",
          9854 => x"0c761e94",
          9855 => x"1b081894",
          9856 => x"1c0c5e5c",
          9857 => x"fdf03980",
          9858 => x"567582d6",
          9859 => x"d80c903d",
          9860 => x"0d04f23d",
          9861 => x"0d606365",
          9862 => x"6440405d",
          9863 => x"58807e0c",
          9864 => x"903dfc05",
          9865 => x"527751f6",
          9866 => x"ce3f82d6",
          9867 => x"d8085582",
          9868 => x"d6d8088a",
          9869 => x"38911833",
          9870 => x"5574802e",
          9871 => x"86387456",
          9872 => x"83be3990",
          9873 => x"18337081",
          9874 => x"2a708106",
          9875 => x"51565687",
          9876 => x"5674802e",
          9877 => x"83aa3895",
          9878 => x"39820b91",
          9879 => x"19348256",
          9880 => x"839e3981",
          9881 => x"0b911934",
          9882 => x"81568394",
          9883 => x"39941808",
          9884 => x"7c115656",
          9885 => x"74762784",
          9886 => x"3875095c",
          9887 => x"7b802e82",
          9888 => x"f2389418",
          9889 => x"087083ff",
          9890 => x"06565674",
          9891 => x"8281387e",
          9892 => x"8a1122ff",
          9893 => x"0577892a",
          9894 => x"065c557a",
          9895 => x"bf38758c",
          9896 => x"38881808",
          9897 => x"55749c38",
          9898 => x"7a528539",
          9899 => x"98180852",
          9900 => x"7751c6ef",
          9901 => x"3f82d6d8",
          9902 => x"085582d6",
          9903 => x"d808802e",
          9904 => x"82b13874",
          9905 => x"812eff91",
          9906 => x"3874ff2e",
          9907 => x"ff953874",
          9908 => x"98190c88",
          9909 => x"18088538",
          9910 => x"7488190c",
          9911 => x"7e55b415",
          9912 => x"089c1908",
          9913 => x"2e098106",
          9914 => x"8e387451",
          9915 => x"ffbdc83f",
          9916 => x"82d6d808",
          9917 => x"feed3898",
          9918 => x"1808527e",
          9919 => x"51c09e3f",
          9920 => x"82d6d808",
          9921 => x"802efed1",
          9922 => x"3882d6d8",
          9923 => x"081b7c89",
          9924 => x"2a5a5778",
          9925 => x"802e80d7",
          9926 => x"38781b7f",
          9927 => x"8a112258",
          9928 => x"5b557575",
          9929 => x"27853875",
          9930 => x"7b315978",
          9931 => x"5476537c",
          9932 => x"52811a33",
          9933 => x"51ffb786",
          9934 => x"3f82d6d8",
          9935 => x"08fea438",
          9936 => x"7eb41108",
          9937 => x"78315656",
          9938 => x"7479279c",
          9939 => x"38848053",
          9940 => x"b4160877",
          9941 => x"31892b7d",
          9942 => x"0552b816",
          9943 => x"51ffbafc",
          9944 => x"3f7e5580",
          9945 => x"0b831634",
          9946 => x"78892b56",
          9947 => x"80de398c",
          9948 => x"18089419",
          9949 => x"08269438",
          9950 => x"7e51ffbc",
          9951 => x"ba3f82d6",
          9952 => x"d808fddf",
          9953 => x"387e77b4",
          9954 => x"120c5576",
          9955 => x"9c190c94",
          9956 => x"180883ff",
          9957 => x"06848071",
          9958 => x"3157557b",
          9959 => x"76278338",
          9960 => x"7b569c18",
          9961 => x"08527e51",
          9962 => x"ffbcfc3f",
          9963 => x"82d6d808",
          9964 => x"fdb13875",
          9965 => x"537c5294",
          9966 => x"180883ff",
          9967 => x"061fb805",
          9968 => x"51ffba98",
          9969 => x"3f7e5581",
          9970 => x"0b831634",
          9971 => x"7b76317e",
          9972 => x"08177f0c",
          9973 => x"761e941a",
          9974 => x"08187094",
          9975 => x"1c0c8c1b",
          9976 => x"0858585e",
          9977 => x"5c747627",
          9978 => x"83387555",
          9979 => x"748c190c",
          9980 => x"fd8a3990",
          9981 => x"183380c0",
          9982 => x"07557490",
          9983 => x"19348056",
          9984 => x"7582d6d8",
          9985 => x"0c903d0d",
          9986 => x"04f83d0d",
          9987 => x"7a8b3dfc",
          9988 => x"05537052",
          9989 => x"56f2e03f",
          9990 => x"82d6d808",
          9991 => x"5782d6d8",
          9992 => x"08818038",
          9993 => x"90163370",
          9994 => x"862a7081",
          9995 => x"06515555",
          9996 => x"73802e80",
          9997 => x"ee38a016",
          9998 => x"08527851",
          9999 => x"ffbbe83f",
         10000 => x"82d6d808",
         10001 => x"5782d6d8",
         10002 => x"0880d838",
         10003 => x"a416088b",
         10004 => x"1133a007",
         10005 => x"5555738b",
         10006 => x"16348816",
         10007 => x"08537452",
         10008 => x"750851cc",
         10009 => x"e93f8c16",
         10010 => x"08529c15",
         10011 => x"51ffb8bd",
         10012 => x"3f8288b2",
         10013 => x"0a529615",
         10014 => x"51ffb8b1",
         10015 => x"3f765292",
         10016 => x"1551ffb8",
         10017 => x"8a3f7854",
         10018 => x"810b8315",
         10019 => x"347851ff",
         10020 => x"bbdc3f82",
         10021 => x"d6d80890",
         10022 => x"173381bf",
         10023 => x"06555773",
         10024 => x"90173476",
         10025 => x"82d6d80c",
         10026 => x"8a3d0d04",
         10027 => x"fc3d0d76",
         10028 => x"705254fe",
         10029 => x"d43f82d6",
         10030 => x"d8085382",
         10031 => x"d6d8089c",
         10032 => x"38863dfc",
         10033 => x"05527351",
         10034 => x"f1ad3f82",
         10035 => x"d6d80853",
         10036 => x"82d6d808",
         10037 => x"873882d6",
         10038 => x"d808740c",
         10039 => x"7282d6d8",
         10040 => x"0c863d0d",
         10041 => x"04ff3d0d",
         10042 => x"843d51e6",
         10043 => x"cd3f8b52",
         10044 => x"800b82d6",
         10045 => x"d808248b",
         10046 => x"3882d6d8",
         10047 => x"0882eeb4",
         10048 => x"34805271",
         10049 => x"82d6d80c",
         10050 => x"833d0d04",
         10051 => x"ee3d0d80",
         10052 => x"53943dcc",
         10053 => x"0552953d",
         10054 => x"51e9aa3f",
         10055 => x"82d6d808",
         10056 => x"5582d6d8",
         10057 => x"0880e038",
         10058 => x"76586452",
         10059 => x"943dd005",
         10060 => x"51ddac3f",
         10061 => x"82d6d808",
         10062 => x"5582d6d8",
         10063 => x"08bc3802",
         10064 => x"80c70533",
         10065 => x"70982b55",
         10066 => x"56738025",
         10067 => x"8938767a",
         10068 => x"98120c54",
         10069 => x"b23902a2",
         10070 => x"05337084",
         10071 => x"2a708106",
         10072 => x"51555673",
         10073 => x"802e9e38",
         10074 => x"767f5370",
         10075 => x"5254caa5",
         10076 => x"3f82d6d8",
         10077 => x"0898150c",
         10078 => x"8e3982d6",
         10079 => x"d808842e",
         10080 => x"09810683",
         10081 => x"38855574",
         10082 => x"82d6d80c",
         10083 => x"943d0d04",
         10084 => x"ffa33d0d",
         10085 => x"80e13d08",
         10086 => x"80e13d08",
         10087 => x"5b5b807a",
         10088 => x"34805380",
         10089 => x"df3dfdb4",
         10090 => x"055280e0",
         10091 => x"3d51e895",
         10092 => x"3f82d6d8",
         10093 => x"085782d6",
         10094 => x"d80883a1",
         10095 => x"387b80d4",
         10096 => x"3d0c7a7c",
         10097 => x"98110880",
         10098 => x"d83d0c55",
         10099 => x"5880d53d",
         10100 => x"08547380",
         10101 => x"2e828338",
         10102 => x"a05280d3",
         10103 => x"3d705255",
         10104 => x"c4d43f82",
         10105 => x"d6d80857",
         10106 => x"82d6d808",
         10107 => x"82ef3880",
         10108 => x"d93d0852",
         10109 => x"7b51ffb8",
         10110 => x"ae3f82d6",
         10111 => x"d8085782",
         10112 => x"d6d80882",
         10113 => x"d83880da",
         10114 => x"3d08527b",
         10115 => x"51c9863f",
         10116 => x"82d6d808",
         10117 => x"80d63d0c",
         10118 => x"76527451",
         10119 => x"c4983f82",
         10120 => x"d6d80857",
         10121 => x"82d6d808",
         10122 => x"82b33880",
         10123 => x"527451c9",
         10124 => x"fa3f82d6",
         10125 => x"d8085782",
         10126 => x"d6d808a7",
         10127 => x"3880da3d",
         10128 => x"08527b51",
         10129 => x"c8cf3f73",
         10130 => x"82d6d808",
         10131 => x"2ea63876",
         10132 => x"527451c5",
         10133 => x"ac3f82d6",
         10134 => x"d8085782",
         10135 => x"d6d80880",
         10136 => x"2ec93876",
         10137 => x"842e0981",
         10138 => x"06863882",
         10139 => x"5781ee39",
         10140 => x"7681ea38",
         10141 => x"80df3dfd",
         10142 => x"b8055274",
         10143 => x"51d6e43f",
         10144 => x"76933d78",
         10145 => x"11821133",
         10146 => x"51565a56",
         10147 => x"73802e92",
         10148 => x"380280c6",
         10149 => x"05558116",
         10150 => x"81167033",
         10151 => x"56565673",
         10152 => x"f5388116",
         10153 => x"54737826",
         10154 => x"81993875",
         10155 => x"802e9c38",
         10156 => x"78168205",
         10157 => x"55ff1880",
         10158 => x"e13d0811",
         10159 => x"ff18ff18",
         10160 => x"58585558",
         10161 => x"74337434",
         10162 => x"75eb38ff",
         10163 => x"1880e13d",
         10164 => x"08115558",
         10165 => x"af7434fd",
         10166 => x"f439777b",
         10167 => x"2e098106",
         10168 => x"8d38ff18",
         10169 => x"80e13d08",
         10170 => x"115558af",
         10171 => x"7434800b",
         10172 => x"82eeb433",
         10173 => x"70842982",
         10174 => x"c7c40570",
         10175 => x"08703352",
         10176 => x"5c565656",
         10177 => x"73762e8d",
         10178 => x"38811670",
         10179 => x"1a703351",
         10180 => x"555673f5",
         10181 => x"38821654",
         10182 => x"737826a7",
         10183 => x"38805574",
         10184 => x"76279138",
         10185 => x"74195473",
         10186 => x"337a7081",
         10187 => x"055c3481",
         10188 => x"1555ec39",
         10189 => x"ba7a7081",
         10190 => x"055c3474",
         10191 => x"ff2e0981",
         10192 => x"06853891",
         10193 => x"57973980",
         10194 => x"e03d0818",
         10195 => x"81195954",
         10196 => x"73337a70",
         10197 => x"81055c34",
         10198 => x"7a7826eb",
         10199 => x"38807a34",
         10200 => x"7682d6d8",
         10201 => x"0c80df3d",
         10202 => x"0d04f73d",
         10203 => x"0d7b7d8d",
         10204 => x"3dfc0554",
         10205 => x"71535755",
         10206 => x"ebfd3f82",
         10207 => x"d6d80853",
         10208 => x"82d6d808",
         10209 => x"82fe3891",
         10210 => x"15335372",
         10211 => x"82f6388c",
         10212 => x"15085473",
         10213 => x"76279238",
         10214 => x"90153370",
         10215 => x"812a7081",
         10216 => x"06515457",
         10217 => x"72833873",
         10218 => x"56941508",
         10219 => x"54807094",
         10220 => x"170c5875",
         10221 => x"782e829b",
         10222 => x"38798a11",
         10223 => x"2270892b",
         10224 => x"59515373",
         10225 => x"782eb738",
         10226 => x"7652ff16",
         10227 => x"51fec8de",
         10228 => x"3f82d6d8",
         10229 => x"08ff1578",
         10230 => x"54705355",
         10231 => x"53fec8ce",
         10232 => x"3f82d6d8",
         10233 => x"08732696",
         10234 => x"38763070",
         10235 => x"75067094",
         10236 => x"180c7771",
         10237 => x"31981808",
         10238 => x"57585153",
         10239 => x"b2398815",
         10240 => x"085473a7",
         10241 => x"38735274",
         10242 => x"51ffbc97",
         10243 => x"3f82d6d8",
         10244 => x"085482d6",
         10245 => x"d808812e",
         10246 => x"819d3882",
         10247 => x"d6d808ff",
         10248 => x"2e819e38",
         10249 => x"82d6d808",
         10250 => x"88160c73",
         10251 => x"98160c73",
         10252 => x"802e819f",
         10253 => x"38767627",
         10254 => x"80de3875",
         10255 => x"77319416",
         10256 => x"08189417",
         10257 => x"0c901633",
         10258 => x"70812a70",
         10259 => x"81065155",
         10260 => x"5a567280",
         10261 => x"2e9b3873",
         10262 => x"527451ff",
         10263 => x"bbc53f82",
         10264 => x"d6d80854",
         10265 => x"82d6d808",
         10266 => x"953882d6",
         10267 => x"d80856a8",
         10268 => x"39735274",
         10269 => x"51ffb5cf",
         10270 => x"3f82d6d8",
         10271 => x"085473ff",
         10272 => x"2ebf3881",
         10273 => x"7427b038",
         10274 => x"7953739c",
         10275 => x"140827a7",
         10276 => x"38739816",
         10277 => x"0cff9e39",
         10278 => x"94150816",
         10279 => x"94160c75",
         10280 => x"83ff0653",
         10281 => x"72802eab",
         10282 => x"38735279",
         10283 => x"51ffb4ed",
         10284 => x"3f82d6d8",
         10285 => x"08943882",
         10286 => x"0b911634",
         10287 => x"825380c4",
         10288 => x"39810b91",
         10289 => x"16348153",
         10290 => x"bb397589",
         10291 => x"2a82d6d8",
         10292 => x"08055894",
         10293 => x"1508548c",
         10294 => x"15087427",
         10295 => x"9038738c",
         10296 => x"160c9015",
         10297 => x"3380c007",
         10298 => x"53729016",
         10299 => x"347383ff",
         10300 => x"06537280",
         10301 => x"2e8c3877",
         10302 => x"9c16082e",
         10303 => x"8538779c",
         10304 => x"160c8053",
         10305 => x"7282d6d8",
         10306 => x"0c8b3d0d",
         10307 => x"04f93d0d",
         10308 => x"79568954",
         10309 => x"75802e81",
         10310 => x"8b388053",
         10311 => x"893dfc05",
         10312 => x"528a3d84",
         10313 => x"0551e19d",
         10314 => x"3f82d6d8",
         10315 => x"085582d6",
         10316 => x"d80880eb",
         10317 => x"3877760c",
         10318 => x"7a527551",
         10319 => x"d5a13f82",
         10320 => x"d6d80855",
         10321 => x"82d6d808",
         10322 => x"80c438ab",
         10323 => x"16337098",
         10324 => x"2b555780",
         10325 => x"7424a238",
         10326 => x"86163370",
         10327 => x"842a7081",
         10328 => x"06515557",
         10329 => x"73802eae",
         10330 => x"389c1608",
         10331 => x"527751c2",
         10332 => x"a43f82d6",
         10333 => x"d8088817",
         10334 => x"0c775486",
         10335 => x"14228417",
         10336 => x"23745275",
         10337 => x"51ffbdae",
         10338 => x"3f82d6d8",
         10339 => x"08557484",
         10340 => x"2e098106",
         10341 => x"85388555",
         10342 => x"86397480",
         10343 => x"2e843880",
         10344 => x"760c7454",
         10345 => x"7382d6d8",
         10346 => x"0c893d0d",
         10347 => x"04fc3d0d",
         10348 => x"76873dfc",
         10349 => x"05537052",
         10350 => x"53e7bc3f",
         10351 => x"82d6d808",
         10352 => x"873882d6",
         10353 => x"d808730c",
         10354 => x"863d0d04",
         10355 => x"fb3d0d77",
         10356 => x"79893dfc",
         10357 => x"05547153",
         10358 => x"5654e79b",
         10359 => x"3f82d6d8",
         10360 => x"085382d6",
         10361 => x"d80880e1",
         10362 => x"38749438",
         10363 => x"82d6d808",
         10364 => x"527351ff",
         10365 => x"bcc03f82",
         10366 => x"d6d80853",
         10367 => x"80cb3982",
         10368 => x"d6d80852",
         10369 => x"7351c2a3",
         10370 => x"3f82d6d8",
         10371 => x"085382d6",
         10372 => x"d808842e",
         10373 => x"09810685",
         10374 => x"38805387",
         10375 => x"3982d6d8",
         10376 => x"08a73874",
         10377 => x"527351cf",
         10378 => x"ba3f7252",
         10379 => x"7351ffbd",
         10380 => x"d03f82d6",
         10381 => x"d8088432",
         10382 => x"70307072",
         10383 => x"079f2c70",
         10384 => x"82d6d808",
         10385 => x"06515154",
         10386 => x"547282d6",
         10387 => x"d80c873d",
         10388 => x"0d04ed3d",
         10389 => x"0d665780",
         10390 => x"53893d70",
         10391 => x"53973d52",
         10392 => x"56dee23f",
         10393 => x"82d6d808",
         10394 => x"5582d6d8",
         10395 => x"08b23865",
         10396 => x"527551d2",
         10397 => x"ea3f82d6",
         10398 => x"d8085582",
         10399 => x"d6d808a0",
         10400 => x"380280cb",
         10401 => x"05337098",
         10402 => x"2b555873",
         10403 => x"80258538",
         10404 => x"86558d39",
         10405 => x"76802e88",
         10406 => x"38765275",
         10407 => x"51cec43f",
         10408 => x"7482d6d8",
         10409 => x"0c953d0d",
         10410 => x"04f03d0d",
         10411 => x"6365555c",
         10412 => x"8053923d",
         10413 => x"ec055293",
         10414 => x"3d51de89",
         10415 => x"3f82d6d8",
         10416 => x"085b82d6",
         10417 => x"d8088282",
         10418 => x"387c740c",
         10419 => x"73089c11",
         10420 => x"08fe1194",
         10421 => x"13085956",
         10422 => x"58557574",
         10423 => x"26913875",
         10424 => x"7c0c81e6",
         10425 => x"39815b81",
         10426 => x"ce39825b",
         10427 => x"81c93982",
         10428 => x"d6d80875",
         10429 => x"33555973",
         10430 => x"812e0981",
         10431 => x"0680c038",
         10432 => x"82755f57",
         10433 => x"7652923d",
         10434 => x"f00551ff",
         10435 => x"b0b93f82",
         10436 => x"d6d808ff",
         10437 => x"2ecf3882",
         10438 => x"d6d80881",
         10439 => x"2ecc3882",
         10440 => x"d6d80830",
         10441 => x"7082d6d8",
         10442 => x"08078025",
         10443 => x"7a058119",
         10444 => x"7f53595a",
         10445 => x"549c1408",
         10446 => x"7726c938",
         10447 => x"80f939a8",
         10448 => x"150882d6",
         10449 => x"d8085758",
         10450 => x"75983877",
         10451 => x"5281187d",
         10452 => x"5258ffad",
         10453 => x"d23f82d6",
         10454 => x"d8085b82",
         10455 => x"d6d80880",
         10456 => x"d6387c70",
         10457 => x"337712ff",
         10458 => x"1a5d5256",
         10459 => x"5474822e",
         10460 => x"0981069e",
         10461 => x"38b81451",
         10462 => x"ffa9d23f",
         10463 => x"82d6d808",
         10464 => x"83ffff06",
         10465 => x"70307080",
         10466 => x"251b8219",
         10467 => x"595b5154",
         10468 => x"9b39b814",
         10469 => x"51ffa9cc",
         10470 => x"3f82d6d8",
         10471 => x"08f00a06",
         10472 => x"70307080",
         10473 => x"251b8419",
         10474 => x"595b5154",
         10475 => x"7583ff06",
         10476 => x"7a585679",
         10477 => x"ff923878",
         10478 => x"7c0c7c79",
         10479 => x"94120c84",
         10480 => x"11338107",
         10481 => x"56547484",
         10482 => x"15347a82",
         10483 => x"d6d80c92",
         10484 => x"3d0d04f9",
         10485 => x"3d0d798a",
         10486 => x"3dfc0553",
         10487 => x"705257e3",
         10488 => x"963f82d6",
         10489 => x"d8085682",
         10490 => x"d6d80881",
         10491 => x"aa389117",
         10492 => x"33567581",
         10493 => x"a2389017",
         10494 => x"3370812a",
         10495 => x"70810651",
         10496 => x"55558755",
         10497 => x"73802e81",
         10498 => x"90389417",
         10499 => x"0854738c",
         10500 => x"18082781",
         10501 => x"8238739c",
         10502 => x"3882d6d8",
         10503 => x"08538817",
         10504 => x"08527651",
         10505 => x"ffb2d03f",
         10506 => x"82d6d808",
         10507 => x"7488190c",
         10508 => x"5680ca39",
         10509 => x"98170852",
         10510 => x"7651ffae",
         10511 => x"8a3f82d6",
         10512 => x"d808ff2e",
         10513 => x"09810683",
         10514 => x"38815682",
         10515 => x"d6d80881",
         10516 => x"2e098106",
         10517 => x"85388256",
         10518 => x"a43975a1",
         10519 => x"38775482",
         10520 => x"d6d8089c",
         10521 => x"15082795",
         10522 => x"38981708",
         10523 => x"5382d6d8",
         10524 => x"08527651",
         10525 => x"ffb2803f",
         10526 => x"82d6d808",
         10527 => x"56941708",
         10528 => x"8c180c90",
         10529 => x"173380c0",
         10530 => x"07547390",
         10531 => x"18347580",
         10532 => x"2e853875",
         10533 => x"91183475",
         10534 => x"557482d6",
         10535 => x"d80c893d",
         10536 => x"0d04e03d",
         10537 => x"0d8253a2",
         10538 => x"3dff9c05",
         10539 => x"52a33d51",
         10540 => x"da933f82",
         10541 => x"d6d80855",
         10542 => x"82d6d808",
         10543 => x"81f93878",
         10544 => x"46a33d08",
         10545 => x"52963d70",
         10546 => x"5258ce93",
         10547 => x"3f82d6d8",
         10548 => x"085582d6",
         10549 => x"d80881df",
         10550 => x"380280ff",
         10551 => x"05337085",
         10552 => x"2a708106",
         10553 => x"51555686",
         10554 => x"557381cb",
         10555 => x"3875982b",
         10556 => x"54807424",
         10557 => x"81c13802",
         10558 => x"80da0533",
         10559 => x"70810658",
         10560 => x"54875576",
         10561 => x"81b1386c",
         10562 => x"527851ff",
         10563 => x"bb873f82",
         10564 => x"d6d80874",
         10565 => x"842a7081",
         10566 => x"06515556",
         10567 => x"73802e80",
         10568 => x"d6387854",
         10569 => x"82d6d808",
         10570 => x"9815082e",
         10571 => x"81893873",
         10572 => x"5a82d6d8",
         10573 => x"085c7652",
         10574 => x"8a3d7052",
         10575 => x"54ffb5f6",
         10576 => x"3f82d6d8",
         10577 => x"085582d6",
         10578 => x"d80880eb",
         10579 => x"3882d6d8",
         10580 => x"08527351",
         10581 => x"ffbbd43f",
         10582 => x"82d6d808",
         10583 => x"5582d6d8",
         10584 => x"08863887",
         10585 => x"5580d039",
         10586 => x"82d6d808",
         10587 => x"842e8838",
         10588 => x"82d6d808",
         10589 => x"80c13877",
         10590 => x"51c7ef3f",
         10591 => x"82d6d808",
         10592 => x"82d6d808",
         10593 => x"307082d6",
         10594 => x"d8080780",
         10595 => x"25515555",
         10596 => x"75802e95",
         10597 => x"3873802e",
         10598 => x"90388053",
         10599 => x"75527751",
         10600 => x"ffafd43f",
         10601 => x"82d6d808",
         10602 => x"55748c38",
         10603 => x"7851ffa9",
         10604 => x"bd3f82d6",
         10605 => x"d8085574",
         10606 => x"82d6d80c",
         10607 => x"a23d0d04",
         10608 => x"e83d0d82",
         10609 => x"539a3dff",
         10610 => x"bc05529b",
         10611 => x"3d51d7f5",
         10612 => x"3f82d6d8",
         10613 => x"085482d6",
         10614 => x"d80882b7",
         10615 => x"38785e6a",
         10616 => x"528e3d70",
         10617 => x"5258cbf7",
         10618 => x"3f82d6d8",
         10619 => x"085482d6",
         10620 => x"d8088638",
         10621 => x"8854829b",
         10622 => x"3982d6d8",
         10623 => x"08842e09",
         10624 => x"8106828f",
         10625 => x"380280df",
         10626 => x"05337085",
         10627 => x"2a810651",
         10628 => x"55865474",
         10629 => x"81fd3878",
         10630 => x"5a74528a",
         10631 => x"3d705257",
         10632 => x"ffb0803f",
         10633 => x"82d6d808",
         10634 => x"75555682",
         10635 => x"d6d80883",
         10636 => x"38875482",
         10637 => x"d6d80881",
         10638 => x"2e098106",
         10639 => x"83388254",
         10640 => x"82d6d808",
         10641 => x"ff2e0981",
         10642 => x"06863881",
         10643 => x"5481ba39",
         10644 => x"7381b638",
         10645 => x"82d6d808",
         10646 => x"527851ff",
         10647 => x"b2e03f82",
         10648 => x"d6d80854",
         10649 => x"82d6d808",
         10650 => x"819f388b",
         10651 => x"53a052b8",
         10652 => x"1951ffa5",
         10653 => x"8a3f7854",
         10654 => x"ae0bb815",
         10655 => x"34785490",
         10656 => x"0b80c315",
         10657 => x"348288b2",
         10658 => x"0a5280ce",
         10659 => x"1951ffa4",
         10660 => x"9c3f7553",
         10661 => x"78b81153",
         10662 => x"51ffb8b2",
         10663 => x"3fa05378",
         10664 => x"b8115380",
         10665 => x"d80551ff",
         10666 => x"a4b23f78",
         10667 => x"54ae0b80",
         10668 => x"d915347f",
         10669 => x"537880d8",
         10670 => x"115351ff",
         10671 => x"b8903f78",
         10672 => x"54810b83",
         10673 => x"15347751",
         10674 => x"ffbfcd3f",
         10675 => x"82d6d808",
         10676 => x"5482d6d8",
         10677 => x"08b33882",
         10678 => x"88b20a52",
         10679 => x"64960551",
         10680 => x"ffa3ca3f",
         10681 => x"75536452",
         10682 => x"7851ffb7",
         10683 => x"e13f6454",
         10684 => x"900b8b15",
         10685 => x"34785481",
         10686 => x"0b831534",
         10687 => x"7851ffa6",
         10688 => x"ed3f82d6",
         10689 => x"d808548b",
         10690 => x"39805375",
         10691 => x"527651ff",
         10692 => x"ace53f73",
         10693 => x"82d6d80c",
         10694 => x"9a3d0d04",
         10695 => x"d83d0dab",
         10696 => x"3d840551",
         10697 => x"d2943f82",
         10698 => x"53aa3dfe",
         10699 => x"fc0552ab",
         10700 => x"3d51d591",
         10701 => x"3f82d6d8",
         10702 => x"085582d6",
         10703 => x"d80882d8",
         10704 => x"38784eab",
         10705 => x"3d08529e",
         10706 => x"3d705258",
         10707 => x"c9913f82",
         10708 => x"d6d80855",
         10709 => x"82d6d808",
         10710 => x"82be3802",
         10711 => x"819f0533",
         10712 => x"81a00654",
         10713 => x"86557382",
         10714 => x"af38a053",
         10715 => x"a53d0852",
         10716 => x"aa3dff80",
         10717 => x"0551ffa2",
         10718 => x"e33fb053",
         10719 => x"7752923d",
         10720 => x"705254ff",
         10721 => x"a2d63fac",
         10722 => x"3d085273",
         10723 => x"51c8d03f",
         10724 => x"82d6d808",
         10725 => x"5582d6d8",
         10726 => x"08973863",
         10727 => x"a13d082e",
         10728 => x"09810688",
         10729 => x"3865a33d",
         10730 => x"082e9238",
         10731 => x"885581e8",
         10732 => x"3982d6d8",
         10733 => x"08842e09",
         10734 => x"810681bb",
         10735 => x"387351ff",
         10736 => x"bdd63f82",
         10737 => x"d6d80855",
         10738 => x"82d6d808",
         10739 => x"81ca3868",
         10740 => x"569353aa",
         10741 => x"3dff8d05",
         10742 => x"528d1651",
         10743 => x"ffa1fd3f",
         10744 => x"02af0533",
         10745 => x"8b17348b",
         10746 => x"16337084",
         10747 => x"2a708106",
         10748 => x"51555573",
         10749 => x"893874a0",
         10750 => x"0754738b",
         10751 => x"17347854",
         10752 => x"810b8315",
         10753 => x"348b1633",
         10754 => x"70842a70",
         10755 => x"81065155",
         10756 => x"5573802e",
         10757 => x"80e7386f",
         10758 => x"642e80e1",
         10759 => x"38755278",
         10760 => x"51ffb4f1",
         10761 => x"3f82d6d8",
         10762 => x"08527851",
         10763 => x"ffa5ee3f",
         10764 => x"825582d6",
         10765 => x"d808802e",
         10766 => x"80de3882",
         10767 => x"d6d80852",
         10768 => x"7851ffa3",
         10769 => x"e23f82d6",
         10770 => x"d8087980",
         10771 => x"d8115858",
         10772 => x"5582d6d8",
         10773 => x"0880c138",
         10774 => x"81163354",
         10775 => x"73ae2e09",
         10776 => x"81069a38",
         10777 => x"63537552",
         10778 => x"7651ffb4",
         10779 => x"e13f7854",
         10780 => x"810b8315",
         10781 => x"34873982",
         10782 => x"d6d8089c",
         10783 => x"387751c1",
         10784 => x"e93f82d6",
         10785 => x"d8085582",
         10786 => x"d6d8088c",
         10787 => x"387851ff",
         10788 => x"a3dc3f82",
         10789 => x"d6d80855",
         10790 => x"7482d6d8",
         10791 => x"0caa3d0d",
         10792 => x"04ec3d0d",
         10793 => x"0280df05",
         10794 => x"33028405",
         10795 => x"80e30533",
         10796 => x"57578253",
         10797 => x"963dcc05",
         10798 => x"52973d51",
         10799 => x"d2873f82",
         10800 => x"d6d80855",
         10801 => x"82d6d808",
         10802 => x"80cf3878",
         10803 => x"5a665296",
         10804 => x"3dd00551",
         10805 => x"c6893f82",
         10806 => x"d6d80855",
         10807 => x"82d6d808",
         10808 => x"b8380280",
         10809 => x"cf053381",
         10810 => x"a0065486",
         10811 => x"5573aa38",
         10812 => x"75a70661",
         10813 => x"71098b12",
         10814 => x"3371067a",
         10815 => x"74060751",
         10816 => x"57555674",
         10817 => x"8b153478",
         10818 => x"54810b83",
         10819 => x"15347851",
         10820 => x"ffa2db3f",
         10821 => x"82d6d808",
         10822 => x"557482d6",
         10823 => x"d80c963d",
         10824 => x"0d04ee3d",
         10825 => x"0d655682",
         10826 => x"53943dcc",
         10827 => x"0552953d",
         10828 => x"51d1923f",
         10829 => x"82d6d808",
         10830 => x"5582d6d8",
         10831 => x"0880cb38",
         10832 => x"76586452",
         10833 => x"943dd005",
         10834 => x"51c5943f",
         10835 => x"82d6d808",
         10836 => x"5582d6d8",
         10837 => x"08b43802",
         10838 => x"80c70533",
         10839 => x"81a00654",
         10840 => x"865573a6",
         10841 => x"38841622",
         10842 => x"86172271",
         10843 => x"902b0753",
         10844 => x"54961f51",
         10845 => x"ff9eb63f",
         10846 => x"7654810b",
         10847 => x"83153476",
         10848 => x"51ffa1ea",
         10849 => x"3f82d6d8",
         10850 => x"08557482",
         10851 => x"d6d80c94",
         10852 => x"3d0d04e9",
         10853 => x"3d0d6a6c",
         10854 => x"5c5a8053",
         10855 => x"993dcc05",
         10856 => x"529a3d51",
         10857 => x"d09f3f82",
         10858 => x"d6d80882",
         10859 => x"d6d80830",
         10860 => x"7082d6d8",
         10861 => x"08078025",
         10862 => x"51555779",
         10863 => x"802e8186",
         10864 => x"38817075",
         10865 => x"06555573",
         10866 => x"802e80fa",
         10867 => x"387b5d80",
         10868 => x"5f80528d",
         10869 => x"3d705254",
         10870 => x"ffacdb3f",
         10871 => x"82d6d808",
         10872 => x"5782d6d8",
         10873 => x"0880d238",
         10874 => x"74527351",
         10875 => x"ffb2bc3f",
         10876 => x"82d6d808",
         10877 => x"5782d6d8",
         10878 => x"08bf3882",
         10879 => x"d6d80882",
         10880 => x"d6d80865",
         10881 => x"5b595678",
         10882 => x"1881197b",
         10883 => x"18565955",
         10884 => x"74337434",
         10885 => x"8116568a",
         10886 => x"7827ec38",
         10887 => x"8b56751a",
         10888 => x"54807434",
         10889 => x"75802e9e",
         10890 => x"38ff1670",
         10891 => x"1b703351",
         10892 => x"555673a0",
         10893 => x"2ee8388e",
         10894 => x"3976842e",
         10895 => x"09810686",
         10896 => x"38807a34",
         10897 => x"80577630",
         10898 => x"70780780",
         10899 => x"2551547a",
         10900 => x"802e80c1",
         10901 => x"3873802e",
         10902 => x"bc387ba4",
         10903 => x"11085351",
         10904 => x"ff9fc43f",
         10905 => x"82d6d808",
         10906 => x"5782d6d8",
         10907 => x"08a7387b",
         10908 => x"70335555",
         10909 => x"80c35673",
         10910 => x"832e8b38",
         10911 => x"80e45673",
         10912 => x"842e8338",
         10913 => x"a7567515",
         10914 => x"b80551ff",
         10915 => x"9bd63f82",
         10916 => x"d6d8087b",
         10917 => x"0c7682d6",
         10918 => x"d80c993d",
         10919 => x"0d04e63d",
         10920 => x"0d82539c",
         10921 => x"3dffb405",
         10922 => x"529d3d51",
         10923 => x"ce973f82",
         10924 => x"d6d80882",
         10925 => x"d6d80856",
         10926 => x"5482d6d8",
         10927 => x"0882dd38",
         10928 => x"8b53a052",
         10929 => x"8a3d7052",
         10930 => x"58ff9cb3",
         10931 => x"3f736d70",
         10932 => x"33515556",
         10933 => x"9f742781",
         10934 => x"86387757",
         10935 => x"9d3d51ff",
         10936 => x"9d903f82",
         10937 => x"d6d80883",
         10938 => x"ffff2680",
         10939 => x"c43882d6",
         10940 => x"d8085195",
         10941 => x"983f83b5",
         10942 => x"5282d6d8",
         10943 => x"085193e8",
         10944 => x"3f82d6d8",
         10945 => x"0883ffff",
         10946 => x"06557480",
         10947 => x"2ea33874",
         10948 => x"5282c8e4",
         10949 => x"51ff9cb2",
         10950 => x"3f82d6d8",
         10951 => x"08933881",
         10952 => x"ff752788",
         10953 => x"38758926",
         10954 => x"88388b39",
         10955 => x"8a762786",
         10956 => x"38865581",
         10957 => x"e73981ff",
         10958 => x"75278f38",
         10959 => x"74882a54",
         10960 => x"73777081",
         10961 => x"05593481",
         10962 => x"16567477",
         10963 => x"70810559",
         10964 => x"3481166d",
         10965 => x"70335155",
         10966 => x"56739f26",
         10967 => x"fefe388a",
         10968 => x"3d335486",
         10969 => x"557381e5",
         10970 => x"2e81b138",
         10971 => x"75802e99",
         10972 => x"3802a305",
         10973 => x"55751570",
         10974 => x"33515473",
         10975 => x"a02e0981",
         10976 => x"068738ff",
         10977 => x"165675ed",
         10978 => x"38784080",
         10979 => x"42805290",
         10980 => x"3d705255",
         10981 => x"ffa99f3f",
         10982 => x"82d6d808",
         10983 => x"5482d6d8",
         10984 => x"0880f738",
         10985 => x"81527451",
         10986 => x"ffaf803f",
         10987 => x"82d6d808",
         10988 => x"5482d6d8",
         10989 => x"088d3875",
         10990 => x"80c43866",
         10991 => x"54e57434",
         10992 => x"80c63982",
         10993 => x"d6d80884",
         10994 => x"2e098106",
         10995 => x"80cc3880",
         10996 => x"5475742e",
         10997 => x"80c43881",
         10998 => x"527451ff",
         10999 => x"ac9c3f82",
         11000 => x"d6d80854",
         11001 => x"82d6d808",
         11002 => x"b138a053",
         11003 => x"82d6d808",
         11004 => x"526651ff",
         11005 => x"9a893f66",
         11006 => x"54880b8b",
         11007 => x"15348b53",
         11008 => x"77526651",
         11009 => x"ff99d53f",
         11010 => x"7854810b",
         11011 => x"83153478",
         11012 => x"51ff9cda",
         11013 => x"3f82d6d8",
         11014 => x"08547355",
         11015 => x"7482d6d8",
         11016 => x"0c9c3d0d",
         11017 => x"04f23d0d",
         11018 => x"60620288",
         11019 => x"0580cb05",
         11020 => x"33933dfc",
         11021 => x"05557254",
         11022 => x"405e5ad2",
         11023 => x"ba3f82d6",
         11024 => x"d8085882",
         11025 => x"d6d80882",
         11026 => x"bd38911a",
         11027 => x"33587782",
         11028 => x"b5387c80",
         11029 => x"2e97388c",
         11030 => x"1a085978",
         11031 => x"9038901a",
         11032 => x"3370812a",
         11033 => x"70810651",
         11034 => x"55557390",
         11035 => x"38875482",
         11036 => x"97398258",
         11037 => x"82903981",
         11038 => x"58828b39",
         11039 => x"7e8a1122",
         11040 => x"70892b70",
         11041 => x"557f5456",
         11042 => x"5656feaf",
         11043 => x"a13fff14",
         11044 => x"7d067030",
         11045 => x"7072079f",
         11046 => x"2a82d6d8",
         11047 => x"08059019",
         11048 => x"087c405a",
         11049 => x"5d555581",
         11050 => x"77278838",
         11051 => x"9c160877",
         11052 => x"26833882",
         11053 => x"57767756",
         11054 => x"59805674",
         11055 => x"527951ff",
         11056 => x"9d853f81",
         11057 => x"157f5555",
         11058 => x"9c140875",
         11059 => x"26833882",
         11060 => x"5582d6d8",
         11061 => x"08812eff",
         11062 => x"993882d6",
         11063 => x"d808ff2e",
         11064 => x"ff953882",
         11065 => x"d6d8088e",
         11066 => x"38811656",
         11067 => x"757b2e09",
         11068 => x"81068738",
         11069 => x"93397459",
         11070 => x"80567477",
         11071 => x"2e098106",
         11072 => x"ffb93887",
         11073 => x"5880ff39",
         11074 => x"7d802eba",
         11075 => x"38787b55",
         11076 => x"557a802e",
         11077 => x"b4388115",
         11078 => x"5673812e",
         11079 => x"09810683",
         11080 => x"38ff5675",
         11081 => x"5374527e",
         11082 => x"51ff9e94",
         11083 => x"3f82d6d8",
         11084 => x"085882d6",
         11085 => x"d80880ce",
         11086 => x"38748116",
         11087 => x"ff165656",
         11088 => x"5c73d338",
         11089 => x"8439ff19",
         11090 => x"5c7e7c90",
         11091 => x"120c557d",
         11092 => x"802eb338",
         11093 => x"78881b0c",
         11094 => x"7c8c1b0c",
         11095 => x"901a3380",
         11096 => x"c0075473",
         11097 => x"901b349c",
         11098 => x"1508fe05",
         11099 => x"94160857",
         11100 => x"54757426",
         11101 => x"9138757b",
         11102 => x"3194160c",
         11103 => x"84153381",
         11104 => x"07547384",
         11105 => x"16347754",
         11106 => x"7382d6d8",
         11107 => x"0c903d0d",
         11108 => x"04e93d0d",
         11109 => x"6b6d0288",
         11110 => x"0580eb05",
         11111 => x"339d3d54",
         11112 => x"5a5c59c5",
         11113 => x"953f8b56",
         11114 => x"800b82d6",
         11115 => x"d808248b",
         11116 => x"f83882d6",
         11117 => x"d8088429",
         11118 => x"82eea005",
         11119 => x"70085155",
         11120 => x"74802e84",
         11121 => x"38807534",
         11122 => x"82d6d808",
         11123 => x"81ff065f",
         11124 => x"81527e51",
         11125 => x"ff8efe3f",
         11126 => x"82d6d808",
         11127 => x"81ff0670",
         11128 => x"81065657",
         11129 => x"8356748b",
         11130 => x"c0387682",
         11131 => x"2a708106",
         11132 => x"51558a56",
         11133 => x"748bb238",
         11134 => x"993dfc05",
         11135 => x"5383527e",
         11136 => x"51ff939e",
         11137 => x"3f82d6d8",
         11138 => x"08993867",
         11139 => x"5574802e",
         11140 => x"92387482",
         11141 => x"8080268b",
         11142 => x"38ff1575",
         11143 => x"06557480",
         11144 => x"2e833881",
         11145 => x"4878802e",
         11146 => x"87388480",
         11147 => x"79269238",
         11148 => x"7881800a",
         11149 => x"268b38ff",
         11150 => x"19790655",
         11151 => x"74802e86",
         11152 => x"3893568a",
         11153 => x"e4397889",
         11154 => x"2a6e892a",
         11155 => x"70892b77",
         11156 => x"59484359",
         11157 => x"7a833881",
         11158 => x"56613070",
         11159 => x"80257707",
         11160 => x"51559156",
         11161 => x"748ac238",
         11162 => x"993df805",
         11163 => x"5381527e",
         11164 => x"51ff92ae",
         11165 => x"3f815682",
         11166 => x"d6d8088a",
         11167 => x"ac387783",
         11168 => x"2a707706",
         11169 => x"82d6d808",
         11170 => x"43564574",
         11171 => x"8338bf41",
         11172 => x"66558e56",
         11173 => x"6075268a",
         11174 => x"90387461",
         11175 => x"31704855",
         11176 => x"80ff7527",
         11177 => x"8a833893",
         11178 => x"56788180",
         11179 => x"2689fa38",
         11180 => x"77812a70",
         11181 => x"81065643",
         11182 => x"74802e95",
         11183 => x"38778706",
         11184 => x"5574822e",
         11185 => x"838d3877",
         11186 => x"81065574",
         11187 => x"802e8383",
         11188 => x"38778106",
         11189 => x"55935682",
         11190 => x"5e74802e",
         11191 => x"89cb3878",
         11192 => x"5a7d832e",
         11193 => x"09810680",
         11194 => x"e13878ae",
         11195 => x"3866912a",
         11196 => x"57810b82",
         11197 => x"c9882256",
         11198 => x"5a74802e",
         11199 => x"9d387477",
         11200 => x"26983882",
         11201 => x"c9885679",
         11202 => x"10821770",
         11203 => x"2257575a",
         11204 => x"74802e86",
         11205 => x"38767527",
         11206 => x"ee387952",
         11207 => x"6651feaa",
         11208 => x"8d3f82d6",
         11209 => x"d8088429",
         11210 => x"84870570",
         11211 => x"892a5e55",
         11212 => x"a05c800b",
         11213 => x"82d6d808",
         11214 => x"fc808a05",
         11215 => x"5644fdff",
         11216 => x"f00a7527",
         11217 => x"80ec3888",
         11218 => x"d33978ae",
         11219 => x"38668c2a",
         11220 => x"57810b82",
         11221 => x"c8f82256",
         11222 => x"5a74802e",
         11223 => x"9d387477",
         11224 => x"26983882",
         11225 => x"c8f85679",
         11226 => x"10821770",
         11227 => x"2257575a",
         11228 => x"74802e86",
         11229 => x"38767527",
         11230 => x"ee387952",
         11231 => x"6651fea9",
         11232 => x"ad3f82d6",
         11233 => x"d8081084",
         11234 => x"055782d6",
         11235 => x"d8089ff5",
         11236 => x"26963881",
         11237 => x"0b82d6d8",
         11238 => x"081082d6",
         11239 => x"d8080571",
         11240 => x"11722a83",
         11241 => x"0559565e",
         11242 => x"83ff1789",
         11243 => x"2a5d815c",
         11244 => x"a044601c",
         11245 => x"7d116505",
         11246 => x"697012ff",
         11247 => x"05713070",
         11248 => x"72067431",
         11249 => x"5c525957",
         11250 => x"59407d83",
         11251 => x"2e098106",
         11252 => x"8938761c",
         11253 => x"6018415c",
         11254 => x"8439761d",
         11255 => x"5d799029",
         11256 => x"18706231",
         11257 => x"68585155",
         11258 => x"74762687",
         11259 => x"af38757c",
         11260 => x"317d317a",
         11261 => x"53706531",
         11262 => x"5255fea8",
         11263 => x"b13f82d6",
         11264 => x"d808587d",
         11265 => x"832e0981",
         11266 => x"069b3882",
         11267 => x"d6d80883",
         11268 => x"fff52680",
         11269 => x"dd387887",
         11270 => x"83387981",
         11271 => x"2a5978fd",
         11272 => x"be3886f8",
         11273 => x"397d822e",
         11274 => x"09810680",
         11275 => x"c53883ff",
         11276 => x"f50b82d6",
         11277 => x"d80827a0",
         11278 => x"38788f38",
         11279 => x"791a5574",
         11280 => x"80c02686",
         11281 => x"387459fd",
         11282 => x"96396281",
         11283 => x"06557480",
         11284 => x"2e8f3883",
         11285 => x"5efd8839",
         11286 => x"82d6d808",
         11287 => x"9ff52692",
         11288 => x"387886b8",
         11289 => x"38791a59",
         11290 => x"81807927",
         11291 => x"fcf13886",
         11292 => x"ab398055",
         11293 => x"7d812e09",
         11294 => x"81068338",
         11295 => x"7d559ff5",
         11296 => x"78278b38",
         11297 => x"74810655",
         11298 => x"8e567486",
         11299 => x"9c388480",
         11300 => x"5380527a",
         11301 => x"51ff90e7",
         11302 => x"3f8b5382",
         11303 => x"c790527a",
         11304 => x"51ff90b8",
         11305 => x"3f848052",
         11306 => x"8b1b51ff",
         11307 => x"8fe13f79",
         11308 => x"8d1c347b",
         11309 => x"83ffff06",
         11310 => x"528e1b51",
         11311 => x"ff8fd03f",
         11312 => x"810b901c",
         11313 => x"347d8332",
         11314 => x"70307096",
         11315 => x"2a848006",
         11316 => x"54515591",
         11317 => x"1b51ff8f",
         11318 => x"b63f6655",
         11319 => x"7483ffff",
         11320 => x"26903874",
         11321 => x"83ffff06",
         11322 => x"52931b51",
         11323 => x"ff8fa03f",
         11324 => x"8a397452",
         11325 => x"a01b51ff",
         11326 => x"8fb33ff8",
         11327 => x"0b951c34",
         11328 => x"bf52981b",
         11329 => x"51ff8f87",
         11330 => x"3f81ff52",
         11331 => x"9a1b51ff",
         11332 => x"8efd3f60",
         11333 => x"529c1b51",
         11334 => x"ff8f923f",
         11335 => x"7d832e09",
         11336 => x"810680cb",
         11337 => x"388288b2",
         11338 => x"0a5280c3",
         11339 => x"1b51ff8e",
         11340 => x"fc3f7c52",
         11341 => x"a41b51ff",
         11342 => x"8ef33f82",
         11343 => x"52ac1b51",
         11344 => x"ff8eea3f",
         11345 => x"8152b01b",
         11346 => x"51ff8ec3",
         11347 => x"3f8652b2",
         11348 => x"1b51ff8e",
         11349 => x"ba3fff80",
         11350 => x"0b80c01c",
         11351 => x"34a90b80",
         11352 => x"c21c3493",
         11353 => x"5382c79c",
         11354 => x"5280c71b",
         11355 => x"51ae3982",
         11356 => x"88b20a52",
         11357 => x"a71b51ff",
         11358 => x"8eb33f7c",
         11359 => x"83ffff06",
         11360 => x"52961b51",
         11361 => x"ff8e883f",
         11362 => x"ff800ba4",
         11363 => x"1c34a90b",
         11364 => x"a61c3493",
         11365 => x"5382c7b0",
         11366 => x"52ab1b51",
         11367 => x"ff8ebd3f",
         11368 => x"82d4d552",
         11369 => x"83fe1b70",
         11370 => x"5259ff8d",
         11371 => x"e23f8154",
         11372 => x"60537a52",
         11373 => x"7e51ff8a",
         11374 => x"853f8156",
         11375 => x"82d6d808",
         11376 => x"83e7387d",
         11377 => x"832e0981",
         11378 => x"0680ee38",
         11379 => x"75546086",
         11380 => x"05537a52",
         11381 => x"7e51ff89",
         11382 => x"e53f8480",
         11383 => x"5380527a",
         11384 => x"51ff8e9b",
         11385 => x"3f848b85",
         11386 => x"a4d2527a",
         11387 => x"51ff8dbd",
         11388 => x"3f868a85",
         11389 => x"e4f25283",
         11390 => x"e41b51ff",
         11391 => x"8daf3fff",
         11392 => x"185283e8",
         11393 => x"1b51ff8d",
         11394 => x"a43f8252",
         11395 => x"83ec1b51",
         11396 => x"ff8d9a3f",
         11397 => x"82d4d552",
         11398 => x"7851ff8c",
         11399 => x"f23f7554",
         11400 => x"60870553",
         11401 => x"7a527e51",
         11402 => x"ff89933f",
         11403 => x"75546016",
         11404 => x"537a527e",
         11405 => x"51ff8986",
         11406 => x"3f655380",
         11407 => x"527a51ff",
         11408 => x"8dbd3f7f",
         11409 => x"5680587d",
         11410 => x"832e0981",
         11411 => x"069a38f8",
         11412 => x"527a51ff",
         11413 => x"8cd73fff",
         11414 => x"52841b51",
         11415 => x"ff8cce3f",
         11416 => x"f00a5288",
         11417 => x"1b519139",
         11418 => x"87fffff8",
         11419 => x"557d812e",
         11420 => x"8338f855",
         11421 => x"74527a51",
         11422 => x"ff8cb23f",
         11423 => x"7c556157",
         11424 => x"74622683",
         11425 => x"38745776",
         11426 => x"5475537a",
         11427 => x"527e51ff",
         11428 => x"88ac3f82",
         11429 => x"d6d80882",
         11430 => x"87388480",
         11431 => x"5382d6d8",
         11432 => x"08527a51",
         11433 => x"ff8cd83f",
         11434 => x"76167578",
         11435 => x"31565674",
         11436 => x"cd388118",
         11437 => x"5877802e",
         11438 => x"ff8d3879",
         11439 => x"557d832e",
         11440 => x"83386355",
         11441 => x"61577462",
         11442 => x"26833874",
         11443 => x"57765475",
         11444 => x"537a527e",
         11445 => x"51ff87e6",
         11446 => x"3f82d6d8",
         11447 => x"0881c138",
         11448 => x"76167578",
         11449 => x"31565674",
         11450 => x"db388c56",
         11451 => x"7d832e93",
         11452 => x"38865666",
         11453 => x"83ffff26",
         11454 => x"8a388456",
         11455 => x"7d822e83",
         11456 => x"38815664",
         11457 => x"81065877",
         11458 => x"80fe3884",
         11459 => x"80537752",
         11460 => x"7a51ff8b",
         11461 => x"ea3f82d4",
         11462 => x"d5527851",
         11463 => x"ff8af03f",
         11464 => x"83be1b55",
         11465 => x"77753481",
         11466 => x"0b811634",
         11467 => x"810b8216",
         11468 => x"34778316",
         11469 => x"34758416",
         11470 => x"34606705",
         11471 => x"5680fdc1",
         11472 => x"527551fe",
         11473 => x"a1e83ffe",
         11474 => x"0b851634",
         11475 => x"82d6d808",
         11476 => x"822abf07",
         11477 => x"56758616",
         11478 => x"3482d6d8",
         11479 => x"08871634",
         11480 => x"605283c6",
         11481 => x"1b51ff8a",
         11482 => x"c43f6652",
         11483 => x"83ca1b51",
         11484 => x"ff8aba3f",
         11485 => x"81547753",
         11486 => x"7a527e51",
         11487 => x"ff86bf3f",
         11488 => x"815682d6",
         11489 => x"d808a238",
         11490 => x"80538052",
         11491 => x"7e51ff88",
         11492 => x"913f8156",
         11493 => x"82d6d808",
         11494 => x"90388939",
         11495 => x"8e568a39",
         11496 => x"81568639",
         11497 => x"82d6d808",
         11498 => x"567582d6",
         11499 => x"d80c993d",
         11500 => x"0d04f53d",
         11501 => x"0d7d605b",
         11502 => x"59807960",
         11503 => x"ff055a57",
         11504 => x"57767825",
         11505 => x"b4388d3d",
         11506 => x"f8115555",
         11507 => x"8153fc15",
         11508 => x"527951c9",
         11509 => x"bd3f7a81",
         11510 => x"2e098106",
         11511 => x"9c388c3d",
         11512 => x"3355748d",
         11513 => x"2edb3874",
         11514 => x"76708105",
         11515 => x"58348117",
         11516 => x"57748a2e",
         11517 => x"098106c9",
         11518 => x"38807634",
         11519 => x"78557683",
         11520 => x"38765574",
         11521 => x"82d6d80c",
         11522 => x"8d3d0d04",
         11523 => x"f73d0d7b",
         11524 => x"028405b3",
         11525 => x"05335957",
         11526 => x"778a2e09",
         11527 => x"81068738",
         11528 => x"8d527651",
         11529 => x"e73f8417",
         11530 => x"08568076",
         11531 => x"24be3888",
         11532 => x"17087717",
         11533 => x"8c055659",
         11534 => x"77753481",
         11535 => x"1656bb76",
         11536 => x"25a1388b",
         11537 => x"3dfc0554",
         11538 => x"75538c17",
         11539 => x"52760851",
         11540 => x"cbc03f79",
         11541 => x"76327030",
         11542 => x"7072079f",
         11543 => x"2a703053",
         11544 => x"51565675",
         11545 => x"84180c81",
         11546 => x"1988180c",
         11547 => x"8b3d0d04",
         11548 => x"f93d0d79",
         11549 => x"84110856",
         11550 => x"56807524",
         11551 => x"a738893d",
         11552 => x"fc055474",
         11553 => x"538c1652",
         11554 => x"750851cb",
         11555 => x"853f82d6",
         11556 => x"d8089138",
         11557 => x"84160878",
         11558 => x"2e098106",
         11559 => x"87388816",
         11560 => x"08558339",
         11561 => x"ff557482",
         11562 => x"d6d80c89",
         11563 => x"3d0d04fd",
         11564 => x"3d0d7554",
         11565 => x"80cc5380",
         11566 => x"527351ff",
         11567 => x"88c13f76",
         11568 => x"740c853d",
         11569 => x"0d04ea3d",
         11570 => x"0d0280e3",
         11571 => x"05336a53",
         11572 => x"863d7053",
         11573 => x"5454d83f",
         11574 => x"73527251",
         11575 => x"feae3f72",
         11576 => x"51ff8d3f",
         11577 => x"983d0d04",
         11578 => x"fd3d0d75",
         11579 => x"0284059a",
         11580 => x"05225553",
         11581 => x"80527280",
         11582 => x"ff268a38",
         11583 => x"7283ffff",
         11584 => x"065280c3",
         11585 => x"3983ffff",
         11586 => x"73275173",
         11587 => x"83b52e09",
         11588 => x"8106b438",
         11589 => x"70802eaf",
         11590 => x"3882c998",
         11591 => x"22517271",
         11592 => x"2e9c3881",
         11593 => x"127083ff",
         11594 => x"ff065351",
         11595 => x"7180ff26",
         11596 => x"8d387110",
         11597 => x"82c99805",
         11598 => x"70225151",
         11599 => x"e1398180",
         11600 => x"127081ff",
         11601 => x"06535171",
         11602 => x"82d6d80c",
         11603 => x"853d0d04",
         11604 => x"fe3d0d02",
         11605 => x"92052202",
         11606 => x"84059605",
         11607 => x"22535180",
         11608 => x"537080ff",
         11609 => x"26853870",
         11610 => x"539a3971",
         11611 => x"83b52e09",
         11612 => x"81069138",
         11613 => x"7081ff26",
         11614 => x"8b387010",
         11615 => x"82c79805",
         11616 => x"70225451",
         11617 => x"7282d6d8",
         11618 => x"0c843d0d",
         11619 => x"04fb3d0d",
         11620 => x"77517083",
         11621 => x"ffff2681",
         11622 => x"a7387083",
         11623 => x"ffff0682",
         11624 => x"cb985752",
         11625 => x"9fff7227",
         11626 => x"853882cf",
         11627 => x"8c567570",
         11628 => x"82055722",
         11629 => x"70307080",
         11630 => x"25727526",
         11631 => x"07515255",
         11632 => x"7080fb38",
         11633 => x"75708205",
         11634 => x"57227088",
         11635 => x"2a7181ff",
         11636 => x"06701854",
         11637 => x"52555371",
         11638 => x"712580d7",
         11639 => x"38738826",
         11640 => x"80dc3873",
         11641 => x"842982ae",
         11642 => x"98055170",
         11643 => x"08047175",
         11644 => x"31107611",
         11645 => x"70225451",
         11646 => x"5180c339",
         11647 => x"71753181",
         11648 => x"06727131",
         11649 => x"5151a439",
         11650 => x"f012519f",
         11651 => x"39e01251",
         11652 => x"9a39d012",
         11653 => x"519539e6",
         11654 => x"12519039",
         11655 => x"8812518b",
         11656 => x"39ffb012",
         11657 => x"518539c7",
         11658 => x"a0125170",
         11659 => x"83ffff06",
         11660 => x"528c3973",
         11661 => x"fef83872",
         11662 => x"101656fe",
         11663 => x"f1397151",
         11664 => x"7082d6d8",
         11665 => x"0c873d0d",
         11666 => x"04000000",
         11667 => x"00ffffff",
         11668 => x"ff00ffff",
         11669 => x"ffff00ff",
         11670 => x"ffffff00",
         11671 => x"00002c51",
         11672 => x"00002bd5",
         11673 => x"00002bdc",
         11674 => x"00002be3",
         11675 => x"00002bea",
         11676 => x"00002bf1",
         11677 => x"00002bf8",
         11678 => x"00002bff",
         11679 => x"00002c06",
         11680 => x"00002c0d",
         11681 => x"00002c14",
         11682 => x"00002c1b",
         11683 => x"00002c21",
         11684 => x"00002c27",
         11685 => x"00002c2d",
         11686 => x"00002c33",
         11687 => x"00002c39",
         11688 => x"00002c3f",
         11689 => x"00002c45",
         11690 => x"00002c4b",
         11691 => x"00004234",
         11692 => x"0000423a",
         11693 => x"00004240",
         11694 => x"00004246",
         11695 => x"0000424c",
         11696 => x"0000482a",
         11697 => x"0000492a",
         11698 => x"00004a3b",
         11699 => x"00004c93",
         11700 => x"00004912",
         11701 => x"000046ff",
         11702 => x"00004b03",
         11703 => x"00004c64",
         11704 => x"00004b46",
         11705 => x"00004bdc",
         11706 => x"00004b62",
         11707 => x"000049e5",
         11708 => x"000046ff",
         11709 => x"00004a3b",
         11710 => x"00004a64",
         11711 => x"00004b03",
         11712 => x"000046ff",
         11713 => x"000046ff",
         11714 => x"00004b62",
         11715 => x"00004bdc",
         11716 => x"00004c64",
         11717 => x"00004c93",
         11718 => x"000095ee",
         11719 => x"000095fc",
         11720 => x"00009608",
         11721 => x"0000960d",
         11722 => x"00009612",
         11723 => x"00009617",
         11724 => x"0000961c",
         11725 => x"00009621",
         11726 => x"00009627",
         11727 => x"00000e31",
         11728 => x"0000171a",
         11729 => x"0000171a",
         11730 => x"00000e60",
         11731 => x"0000171a",
         11732 => x"0000171a",
         11733 => x"0000171a",
         11734 => x"0000171a",
         11735 => x"0000171a",
         11736 => x"0000171a",
         11737 => x"0000171a",
         11738 => x"00000e1d",
         11739 => x"0000171a",
         11740 => x"00000e48",
         11741 => x"00000e78",
         11742 => x"0000171a",
         11743 => x"0000171a",
         11744 => x"0000171a",
         11745 => x"0000171a",
         11746 => x"0000171a",
         11747 => x"0000171a",
         11748 => x"0000171a",
         11749 => x"0000171a",
         11750 => x"0000171a",
         11751 => x"0000171a",
         11752 => x"0000171a",
         11753 => x"0000171a",
         11754 => x"0000171a",
         11755 => x"0000171a",
         11756 => x"0000171a",
         11757 => x"0000171a",
         11758 => x"0000171a",
         11759 => x"0000171a",
         11760 => x"0000171a",
         11761 => x"0000171a",
         11762 => x"0000171a",
         11763 => x"0000171a",
         11764 => x"0000171a",
         11765 => x"0000171a",
         11766 => x"0000171a",
         11767 => x"0000171a",
         11768 => x"0000171a",
         11769 => x"0000171a",
         11770 => x"0000171a",
         11771 => x"0000171a",
         11772 => x"0000171a",
         11773 => x"0000171a",
         11774 => x"0000171a",
         11775 => x"0000171a",
         11776 => x"0000171a",
         11777 => x"0000171a",
         11778 => x"00000fa8",
         11779 => x"0000171a",
         11780 => x"0000171a",
         11781 => x"0000171a",
         11782 => x"0000171a",
         11783 => x"00001116",
         11784 => x"0000171a",
         11785 => x"0000171a",
         11786 => x"0000171a",
         11787 => x"0000171a",
         11788 => x"0000171a",
         11789 => x"0000171a",
         11790 => x"0000171a",
         11791 => x"0000171a",
         11792 => x"0000171a",
         11793 => x"0000171a",
         11794 => x"00000ed8",
         11795 => x"0000103f",
         11796 => x"00000eaf",
         11797 => x"00000eaf",
         11798 => x"00000eaf",
         11799 => x"0000171a",
         11800 => x"0000103f",
         11801 => x"0000171a",
         11802 => x"0000171a",
         11803 => x"00000e98",
         11804 => x"0000171a",
         11805 => x"0000171a",
         11806 => x"000010ec",
         11807 => x"000010f7",
         11808 => x"0000171a",
         11809 => x"0000171a",
         11810 => x"00000f11",
         11811 => x"0000171a",
         11812 => x"0000111f",
         11813 => x"0000171a",
         11814 => x"0000171a",
         11815 => x"00001116",
         11816 => x"64696e69",
         11817 => x"74000000",
         11818 => x"64696f63",
         11819 => x"746c0000",
         11820 => x"66696e69",
         11821 => x"74000000",
         11822 => x"666c6f61",
         11823 => x"64000000",
         11824 => x"66657865",
         11825 => x"63000000",
         11826 => x"6d636c65",
         11827 => x"61720000",
         11828 => x"6d636f70",
         11829 => x"79000000",
         11830 => x"6d646966",
         11831 => x"66000000",
         11832 => x"6d64756d",
         11833 => x"70000000",
         11834 => x"6d656200",
         11835 => x"6d656800",
         11836 => x"6d657700",
         11837 => x"68696400",
         11838 => x"68696500",
         11839 => x"68666400",
         11840 => x"68666500",
         11841 => x"63616c6c",
         11842 => x"00000000",
         11843 => x"6a6d7000",
         11844 => x"72657374",
         11845 => x"61727400",
         11846 => x"72657365",
         11847 => x"74000000",
         11848 => x"696e666f",
         11849 => x"00000000",
         11850 => x"74657374",
         11851 => x"00000000",
         11852 => x"74626173",
         11853 => x"69630000",
         11854 => x"6d626173",
         11855 => x"69630000",
         11856 => x"6b696c6f",
         11857 => x"00000000",
         11858 => x"65640000",
         11859 => x"4469736b",
         11860 => x"20457272",
         11861 => x"6f720000",
         11862 => x"496e7465",
         11863 => x"726e616c",
         11864 => x"20657272",
         11865 => x"6f722e00",
         11866 => x"4469736b",
         11867 => x"206e6f74",
         11868 => x"20726561",
         11869 => x"64792e00",
         11870 => x"4e6f2066",
         11871 => x"696c6520",
         11872 => x"666f756e",
         11873 => x"642e0000",
         11874 => x"4e6f2070",
         11875 => x"61746820",
         11876 => x"666f756e",
         11877 => x"642e0000",
         11878 => x"496e7661",
         11879 => x"6c696420",
         11880 => x"66696c65",
         11881 => x"6e616d65",
         11882 => x"2e000000",
         11883 => x"41636365",
         11884 => x"73732064",
         11885 => x"656e6965",
         11886 => x"642e0000",
         11887 => x"46696c65",
         11888 => x"20616c72",
         11889 => x"65616479",
         11890 => x"20657869",
         11891 => x"7374732e",
         11892 => x"00000000",
         11893 => x"46696c65",
         11894 => x"2068616e",
         11895 => x"646c6520",
         11896 => x"696e7661",
         11897 => x"6c69642e",
         11898 => x"00000000",
         11899 => x"53442069",
         11900 => x"73207772",
         11901 => x"69746520",
         11902 => x"70726f74",
         11903 => x"65637465",
         11904 => x"642e0000",
         11905 => x"44726976",
         11906 => x"65206e75",
         11907 => x"6d626572",
         11908 => x"20697320",
         11909 => x"696e7661",
         11910 => x"6c69642e",
         11911 => x"00000000",
         11912 => x"4469736b",
         11913 => x"206e6f74",
         11914 => x"20656e61",
         11915 => x"626c6564",
         11916 => x"2e000000",
         11917 => x"4e6f2063",
         11918 => x"6f6d7061",
         11919 => x"7469626c",
         11920 => x"65206669",
         11921 => x"6c657379",
         11922 => x"7374656d",
         11923 => x"20666f75",
         11924 => x"6e64206f",
         11925 => x"6e206469",
         11926 => x"736b2e00",
         11927 => x"466f726d",
         11928 => x"61742061",
         11929 => x"626f7274",
         11930 => x"65642e00",
         11931 => x"54696d65",
         11932 => x"6f75742c",
         11933 => x"206f7065",
         11934 => x"72617469",
         11935 => x"6f6e2063",
         11936 => x"616e6365",
         11937 => x"6c6c6564",
         11938 => x"2e000000",
         11939 => x"46696c65",
         11940 => x"20697320",
         11941 => x"6c6f636b",
         11942 => x"65642e00",
         11943 => x"496e7375",
         11944 => x"66666963",
         11945 => x"69656e74",
         11946 => x"206d656d",
         11947 => x"6f72792e",
         11948 => x"00000000",
         11949 => x"546f6f20",
         11950 => x"6d616e79",
         11951 => x"206f7065",
         11952 => x"6e206669",
         11953 => x"6c65732e",
         11954 => x"00000000",
         11955 => x"50617261",
         11956 => x"6d657465",
         11957 => x"72732069",
         11958 => x"6e636f72",
         11959 => x"72656374",
         11960 => x"2e000000",
         11961 => x"53756363",
         11962 => x"6573732e",
         11963 => x"00000000",
         11964 => x"556e6b6e",
         11965 => x"6f776e20",
         11966 => x"6572726f",
         11967 => x"722e0000",
         11968 => x"0a256c75",
         11969 => x"20627974",
         11970 => x"65732025",
         11971 => x"73206174",
         11972 => x"20256c75",
         11973 => x"20627974",
         11974 => x"65732f73",
         11975 => x"65632e0a",
         11976 => x"00000000",
         11977 => x"72656164",
         11978 => x"00000000",
         11979 => x"303d2530",
         11980 => x"386c782c",
         11981 => x"20313d25",
         11982 => x"30386c78",
         11983 => x"2c20323d",
         11984 => x"2530386c",
         11985 => x"782c205f",
         11986 => x"494f423d",
         11987 => x"2530386c",
         11988 => x"78202530",
         11989 => x"386c7820",
         11990 => x"2530386c",
         11991 => x"780a0000",
         11992 => x"2530386c",
         11993 => x"58000000",
         11994 => x"3a202000",
         11995 => x"25303458",
         11996 => x"00000000",
         11997 => x"20202020",
         11998 => x"20202020",
         11999 => x"00000000",
         12000 => x"25303258",
         12001 => x"00000000",
         12002 => x"20200000",
         12003 => x"207c0000",
         12004 => x"7c000000",
         12005 => x"7a4f5300",
         12006 => x"0a2a2a20",
         12007 => x"25732028",
         12008 => x"00000000",
         12009 => x"30352f31",
         12010 => x"322f3230",
         12011 => x"32300000",
         12012 => x"76312e30",
         12013 => x"34660000",
         12014 => x"205a5055",
         12015 => x"2c207265",
         12016 => x"76202530",
         12017 => x"32782920",
         12018 => x"25732025",
         12019 => x"73202a2a",
         12020 => x"0a0a0000",
         12021 => x"5a505520",
         12022 => x"496e7465",
         12023 => x"72727570",
         12024 => x"74204861",
         12025 => x"6e646c65",
         12026 => x"72000000",
         12027 => x"54696d65",
         12028 => x"7220696e",
         12029 => x"74657272",
         12030 => x"75707400",
         12031 => x"50533220",
         12032 => x"696e7465",
         12033 => x"72727570",
         12034 => x"74000000",
         12035 => x"494f4354",
         12036 => x"4c205244",
         12037 => x"20696e74",
         12038 => x"65727275",
         12039 => x"70740000",
         12040 => x"494f4354",
         12041 => x"4c205752",
         12042 => x"20696e74",
         12043 => x"65727275",
         12044 => x"70740000",
         12045 => x"55415254",
         12046 => x"30205258",
         12047 => x"20696e74",
         12048 => x"65727275",
         12049 => x"70740000",
         12050 => x"55415254",
         12051 => x"30205458",
         12052 => x"20696e74",
         12053 => x"65727275",
         12054 => x"70740000",
         12055 => x"55415254",
         12056 => x"31205258",
         12057 => x"20696e74",
         12058 => x"65727275",
         12059 => x"70740000",
         12060 => x"55415254",
         12061 => x"31205458",
         12062 => x"20696e74",
         12063 => x"65727275",
         12064 => x"70740000",
         12065 => x"53657474",
         12066 => x"696e6720",
         12067 => x"75702074",
         12068 => x"696d6572",
         12069 => x"2e2e2e00",
         12070 => x"456e6162",
         12071 => x"6c696e67",
         12072 => x"2074696d",
         12073 => x"65722e2e",
         12074 => x"2e000000",
         12075 => x"6175746f",
         12076 => x"65786563",
         12077 => x"2e626174",
         12078 => x"00000000",
         12079 => x"7a4f532e",
         12080 => x"68737400",
         12081 => x"303a0000",
         12082 => x"4661696c",
         12083 => x"65642074",
         12084 => x"6f20696e",
         12085 => x"69746961",
         12086 => x"6c697365",
         12087 => x"20736420",
         12088 => x"63617264",
         12089 => x"20302c20",
         12090 => x"706c6561",
         12091 => x"73652069",
         12092 => x"6e697420",
         12093 => x"6d616e75",
         12094 => x"616c6c79",
         12095 => x"2e000000",
         12096 => x"2a200000",
         12097 => x"436c6561",
         12098 => x"72696e67",
         12099 => x"2e2e2e2e",
         12100 => x"00000000",
         12101 => x"436f7079",
         12102 => x"696e672e",
         12103 => x"2e2e0000",
         12104 => x"436f6d70",
         12105 => x"6172696e",
         12106 => x"672e2e2e",
         12107 => x"00000000",
         12108 => x"2530386c",
         12109 => x"78282530",
         12110 => x"3878292d",
         12111 => x"3e253038",
         12112 => x"6c782825",
         12113 => x"30387829",
         12114 => x"0a000000",
         12115 => x"44756d70",
         12116 => x"204d656d",
         12117 => x"6f727900",
         12118 => x"0a436f6d",
         12119 => x"706c6574",
         12120 => x"652e0000",
         12121 => x"2530386c",
         12122 => x"58202530",
         12123 => x"32582d00",
         12124 => x"3f3f3f00",
         12125 => x"2530386c",
         12126 => x"58202530",
         12127 => x"34582d00",
         12128 => x"2530386c",
         12129 => x"58202530",
         12130 => x"386c582d",
         12131 => x"00000000",
         12132 => x"45786563",
         12133 => x"7574696e",
         12134 => x"6720636f",
         12135 => x"64652040",
         12136 => x"20253038",
         12137 => x"6c78202e",
         12138 => x"2e2e0a00",
         12139 => x"43616c6c",
         12140 => x"696e6720",
         12141 => x"636f6465",
         12142 => x"20402025",
         12143 => x"30386c78",
         12144 => x"202e2e2e",
         12145 => x"0a000000",
         12146 => x"43616c6c",
         12147 => x"20726574",
         12148 => x"75726e65",
         12149 => x"6420636f",
         12150 => x"64652028",
         12151 => x"2564292e",
         12152 => x"0a000000",
         12153 => x"52657374",
         12154 => x"61727469",
         12155 => x"6e672061",
         12156 => x"70706c69",
         12157 => x"63617469",
         12158 => x"6f6e2e2e",
         12159 => x"2e000000",
         12160 => x"436f6c64",
         12161 => x"20726562",
         12162 => x"6f6f7469",
         12163 => x"6e672e2e",
         12164 => x"2e000000",
         12165 => x"5a505500",
         12166 => x"62696e00",
         12167 => x"25643a5c",
         12168 => x"25735c25",
         12169 => x"732e2573",
         12170 => x"00000000",
         12171 => x"25643a5c",
         12172 => x"25735c25",
         12173 => x"73000000",
         12174 => x"25643a5c",
         12175 => x"25730000",
         12176 => x"42616420",
         12177 => x"636f6d6d",
         12178 => x"616e642e",
         12179 => x"00000000",
         12180 => x"4d656d6f",
         12181 => x"72792065",
         12182 => x"78686175",
         12183 => x"73746564",
         12184 => x"2c206361",
         12185 => x"6e6e6f74",
         12186 => x"2070726f",
         12187 => x"63657373",
         12188 => x"20636f6d",
         12189 => x"6d616e64",
         12190 => x"2e000000",
         12191 => x"54657374",
         12192 => x"696e6720",
         12193 => x"7072696e",
         12194 => x"74660000",
         12195 => x"52756e6e",
         12196 => x"696e672e",
         12197 => x"2e2e0000",
         12198 => x"456e6162",
         12199 => x"6c696e67",
         12200 => x"20696e74",
         12201 => x"65727275",
         12202 => x"7074732e",
         12203 => x"2e2e0000",
         12204 => x"25642f25",
         12205 => x"642f2564",
         12206 => x"2025643a",
         12207 => x"25643a25",
         12208 => x"642e2564",
         12209 => x"25640a00",
         12210 => x"536f4320",
         12211 => x"436f6e66",
         12212 => x"69677572",
         12213 => x"6174696f",
         12214 => x"6e000000",
         12215 => x"20286672",
         12216 => x"6f6d2053",
         12217 => x"6f432063",
         12218 => x"6f6e6669",
         12219 => x"67290000",
         12220 => x"3a0a4465",
         12221 => x"76696365",
         12222 => x"7320696d",
         12223 => x"706c656d",
         12224 => x"656e7465",
         12225 => x"643a0000",
         12226 => x"20202020",
         12227 => x"57422053",
         12228 => x"4452414d",
         12229 => x"20202825",
         12230 => x"3038583a",
         12231 => x"25303858",
         12232 => x"292e0a00",
         12233 => x"20202020",
         12234 => x"53445241",
         12235 => x"4d202020",
         12236 => x"20202825",
         12237 => x"3038583a",
         12238 => x"25303858",
         12239 => x"292e0a00",
         12240 => x"20202020",
         12241 => x"494e534e",
         12242 => x"20425241",
         12243 => x"4d202825",
         12244 => x"3038583a",
         12245 => x"25303858",
         12246 => x"292e0a00",
         12247 => x"20202020",
         12248 => x"4252414d",
         12249 => x"20202020",
         12250 => x"20202825",
         12251 => x"3038583a",
         12252 => x"25303858",
         12253 => x"292e0a00",
         12254 => x"20202020",
         12255 => x"52414d20",
         12256 => x"20202020",
         12257 => x"20202825",
         12258 => x"3038583a",
         12259 => x"25303858",
         12260 => x"292e0a00",
         12261 => x"20202020",
         12262 => x"53442043",
         12263 => x"41524420",
         12264 => x"20202844",
         12265 => x"65766963",
         12266 => x"6573203d",
         12267 => x"25303264",
         12268 => x"292e0a00",
         12269 => x"20202020",
         12270 => x"54494d45",
         12271 => x"52312020",
         12272 => x"20202854",
         12273 => x"696d6572",
         12274 => x"7320203d",
         12275 => x"25303264",
         12276 => x"292e0a00",
         12277 => x"20202020",
         12278 => x"494e5452",
         12279 => x"20435452",
         12280 => x"4c202843",
         12281 => x"68616e6e",
         12282 => x"656c733d",
         12283 => x"25303264",
         12284 => x"292e0a00",
         12285 => x"20202020",
         12286 => x"57495348",
         12287 => x"424f4e45",
         12288 => x"20425553",
         12289 => x"00000000",
         12290 => x"20202020",
         12291 => x"57422049",
         12292 => x"32430000",
         12293 => x"20202020",
         12294 => x"494f4354",
         12295 => x"4c000000",
         12296 => x"20202020",
         12297 => x"50533200",
         12298 => x"20202020",
         12299 => x"53504900",
         12300 => x"41646472",
         12301 => x"65737365",
         12302 => x"733a0000",
         12303 => x"20202020",
         12304 => x"43505520",
         12305 => x"52657365",
         12306 => x"74205665",
         12307 => x"63746f72",
         12308 => x"20416464",
         12309 => x"72657373",
         12310 => x"203d2025",
         12311 => x"3038580a",
         12312 => x"00000000",
         12313 => x"20202020",
         12314 => x"43505520",
         12315 => x"4d656d6f",
         12316 => x"72792053",
         12317 => x"74617274",
         12318 => x"20416464",
         12319 => x"72657373",
         12320 => x"203d2025",
         12321 => x"3038580a",
         12322 => x"00000000",
         12323 => x"20202020",
         12324 => x"53746163",
         12325 => x"6b205374",
         12326 => x"61727420",
         12327 => x"41646472",
         12328 => x"65737320",
         12329 => x"20202020",
         12330 => x"203d2025",
         12331 => x"3038580a",
         12332 => x"00000000",
         12333 => x"4d697363",
         12334 => x"3a000000",
         12335 => x"20202020",
         12336 => x"5a505520",
         12337 => x"49642020",
         12338 => x"20202020",
         12339 => x"20202020",
         12340 => x"20202020",
         12341 => x"20202020",
         12342 => x"203d2025",
         12343 => x"3034580a",
         12344 => x"00000000",
         12345 => x"20202020",
         12346 => x"53797374",
         12347 => x"656d2043",
         12348 => x"6c6f636b",
         12349 => x"20467265",
         12350 => x"71202020",
         12351 => x"20202020",
         12352 => x"203d2025",
         12353 => x"642e2530",
         12354 => x"34644d48",
         12355 => x"7a0a0000",
         12356 => x"20202020",
         12357 => x"53445241",
         12358 => x"4d20436c",
         12359 => x"6f636b20",
         12360 => x"46726571",
         12361 => x"20202020",
         12362 => x"20202020",
         12363 => x"203d2025",
         12364 => x"642e2530",
         12365 => x"34644d48",
         12366 => x"7a0a0000",
         12367 => x"20202020",
         12368 => x"57697368",
         12369 => x"626f6e65",
         12370 => x"20534452",
         12371 => x"414d2043",
         12372 => x"6c6f636b",
         12373 => x"20467265",
         12374 => x"713d2025",
         12375 => x"642e2530",
         12376 => x"34644d48",
         12377 => x"7a0a0000",
         12378 => x"536d616c",
         12379 => x"6c000000",
         12380 => x"4d656469",
         12381 => x"756d0000",
         12382 => x"466c6578",
         12383 => x"00000000",
         12384 => x"45564f00",
         12385 => x"45564f6d",
         12386 => x"00000000",
         12387 => x"556e6b6e",
         12388 => x"6f776e00",
         12389 => x"0000a2f0",
         12390 => x"01000000",
         12391 => x"00000002",
         12392 => x"0000a2ec",
         12393 => x"01000000",
         12394 => x"00000003",
         12395 => x"0000a2e8",
         12396 => x"01000000",
         12397 => x"00000004",
         12398 => x"0000a2e4",
         12399 => x"01000000",
         12400 => x"00000005",
         12401 => x"0000a2e0",
         12402 => x"01000000",
         12403 => x"00000006",
         12404 => x"0000a2dc",
         12405 => x"01000000",
         12406 => x"00000007",
         12407 => x"0000a2d8",
         12408 => x"01000000",
         12409 => x"00000001",
         12410 => x"0000a2d4",
         12411 => x"01000000",
         12412 => x"00000008",
         12413 => x"0000a2d0",
         12414 => x"01000000",
         12415 => x"0000000b",
         12416 => x"0000a2cc",
         12417 => x"01000000",
         12418 => x"00000009",
         12419 => x"0000a2c8",
         12420 => x"01000000",
         12421 => x"0000000a",
         12422 => x"0000a2c4",
         12423 => x"04000000",
         12424 => x"0000000d",
         12425 => x"0000a2c0",
         12426 => x"04000000",
         12427 => x"0000000c",
         12428 => x"0000a2bc",
         12429 => x"04000000",
         12430 => x"0000000e",
         12431 => x"0000a2b8",
         12432 => x"03000000",
         12433 => x"0000000f",
         12434 => x"0000a2b4",
         12435 => x"04000000",
         12436 => x"0000000f",
         12437 => x"0000a2b0",
         12438 => x"04000000",
         12439 => x"00000010",
         12440 => x"0000a2ac",
         12441 => x"04000000",
         12442 => x"00000011",
         12443 => x"0000a2a8",
         12444 => x"03000000",
         12445 => x"00000012",
         12446 => x"0000a2a4",
         12447 => x"03000000",
         12448 => x"00000013",
         12449 => x"0000a2a0",
         12450 => x"03000000",
         12451 => x"00000014",
         12452 => x"0000a29c",
         12453 => x"03000000",
         12454 => x"00000015",
         12455 => x"1b5b4400",
         12456 => x"1b5b4300",
         12457 => x"1b5b4200",
         12458 => x"1b5b4100",
         12459 => x"1b5b367e",
         12460 => x"1b5b357e",
         12461 => x"1b5b347e",
         12462 => x"1b304600",
         12463 => x"1b5b337e",
         12464 => x"1b5b327e",
         12465 => x"1b5b317e",
         12466 => x"10000000",
         12467 => x"0e000000",
         12468 => x"0d000000",
         12469 => x"0b000000",
         12470 => x"08000000",
         12471 => x"06000000",
         12472 => x"05000000",
         12473 => x"04000000",
         12474 => x"03000000",
         12475 => x"02000000",
         12476 => x"01000000",
         12477 => x"68697374",
         12478 => x"6f727900",
         12479 => x"68697374",
         12480 => x"00000000",
         12481 => x"21000000",
         12482 => x"2530346c",
         12483 => x"75202025",
         12484 => x"730a0000",
         12485 => x"4661696c",
         12486 => x"65642074",
         12487 => x"6f207265",
         12488 => x"73657420",
         12489 => x"74686520",
         12490 => x"68697374",
         12491 => x"6f727920",
         12492 => x"66696c65",
         12493 => x"20746f20",
         12494 => x"454f462e",
         12495 => x"00000000",
         12496 => x"43616e6e",
         12497 => x"6f74206f",
         12498 => x"70656e2f",
         12499 => x"63726561",
         12500 => x"74652068",
         12501 => x"6973746f",
         12502 => x"72792066",
         12503 => x"696c652c",
         12504 => x"20646973",
         12505 => x"61626c69",
         12506 => x"6e672e00",
         12507 => x"53440000",
         12508 => x"222a3a3c",
         12509 => x"3e3f7c7f",
         12510 => x"00000000",
         12511 => x"2b2c3b3d",
         12512 => x"5b5d0000",
         12513 => x"46415400",
         12514 => x"46415433",
         12515 => x"32000000",
         12516 => x"ebfe904d",
         12517 => x"53444f53",
         12518 => x"352e3000",
         12519 => x"4e4f204e",
         12520 => x"414d4520",
         12521 => x"20202046",
         12522 => x"41543332",
         12523 => x"20202000",
         12524 => x"4e4f204e",
         12525 => x"414d4520",
         12526 => x"20202046",
         12527 => x"41542020",
         12528 => x"20202000",
         12529 => x"0000a36c",
         12530 => x"00000000",
         12531 => x"00000000",
         12532 => x"00000000",
         12533 => x"01030507",
         12534 => x"090e1012",
         12535 => x"1416181c",
         12536 => x"1e000000",
         12537 => x"809a4541",
         12538 => x"8e418f80",
         12539 => x"45454549",
         12540 => x"49498e8f",
         12541 => x"9092924f",
         12542 => x"994f5555",
         12543 => x"59999a9b",
         12544 => x"9c9d9e9f",
         12545 => x"41494f55",
         12546 => x"a5a5a6a7",
         12547 => x"a8a9aaab",
         12548 => x"acadaeaf",
         12549 => x"b0b1b2b3",
         12550 => x"b4b5b6b7",
         12551 => x"b8b9babb",
         12552 => x"bcbdbebf",
         12553 => x"c0c1c2c3",
         12554 => x"c4c5c6c7",
         12555 => x"c8c9cacb",
         12556 => x"cccdcecf",
         12557 => x"d0d1d2d3",
         12558 => x"d4d5d6d7",
         12559 => x"d8d9dadb",
         12560 => x"dcdddedf",
         12561 => x"e0e1e2e3",
         12562 => x"e4e5e6e7",
         12563 => x"e8e9eaeb",
         12564 => x"ecedeeef",
         12565 => x"f0f1f2f3",
         12566 => x"f4f5f6f7",
         12567 => x"f8f9fafb",
         12568 => x"fcfdfeff",
         12569 => x"2b2e2c3b",
         12570 => x"3d5b5d2f",
         12571 => x"5c222a3a",
         12572 => x"3c3e3f7c",
         12573 => x"7f000000",
         12574 => x"00010004",
         12575 => x"00100040",
         12576 => x"01000200",
         12577 => x"00000000",
         12578 => x"00010002",
         12579 => x"00040008",
         12580 => x"00100020",
         12581 => x"00000000",
         12582 => x"00c700fc",
         12583 => x"00e900e2",
         12584 => x"00e400e0",
         12585 => x"00e500e7",
         12586 => x"00ea00eb",
         12587 => x"00e800ef",
         12588 => x"00ee00ec",
         12589 => x"00c400c5",
         12590 => x"00c900e6",
         12591 => x"00c600f4",
         12592 => x"00f600f2",
         12593 => x"00fb00f9",
         12594 => x"00ff00d6",
         12595 => x"00dc00a2",
         12596 => x"00a300a5",
         12597 => x"20a70192",
         12598 => x"00e100ed",
         12599 => x"00f300fa",
         12600 => x"00f100d1",
         12601 => x"00aa00ba",
         12602 => x"00bf2310",
         12603 => x"00ac00bd",
         12604 => x"00bc00a1",
         12605 => x"00ab00bb",
         12606 => x"25912592",
         12607 => x"25932502",
         12608 => x"25242561",
         12609 => x"25622556",
         12610 => x"25552563",
         12611 => x"25512557",
         12612 => x"255d255c",
         12613 => x"255b2510",
         12614 => x"25142534",
         12615 => x"252c251c",
         12616 => x"2500253c",
         12617 => x"255e255f",
         12618 => x"255a2554",
         12619 => x"25692566",
         12620 => x"25602550",
         12621 => x"256c2567",
         12622 => x"25682564",
         12623 => x"25652559",
         12624 => x"25582552",
         12625 => x"2553256b",
         12626 => x"256a2518",
         12627 => x"250c2588",
         12628 => x"2584258c",
         12629 => x"25902580",
         12630 => x"03b100df",
         12631 => x"039303c0",
         12632 => x"03a303c3",
         12633 => x"00b503c4",
         12634 => x"03a60398",
         12635 => x"03a903b4",
         12636 => x"221e03c6",
         12637 => x"03b52229",
         12638 => x"226100b1",
         12639 => x"22652264",
         12640 => x"23202321",
         12641 => x"00f72248",
         12642 => x"00b02219",
         12643 => x"00b7221a",
         12644 => x"207f00b2",
         12645 => x"25a000a0",
         12646 => x"0061031a",
         12647 => x"00e00317",
         12648 => x"00f80307",
         12649 => x"00ff0001",
         12650 => x"01780100",
         12651 => x"01300132",
         12652 => x"01060139",
         12653 => x"0110014a",
         12654 => x"012e0179",
         12655 => x"01060180",
         12656 => x"004d0243",
         12657 => x"01810182",
         12658 => x"01820184",
         12659 => x"01840186",
         12660 => x"01870187",
         12661 => x"0189018a",
         12662 => x"018b018b",
         12663 => x"018d018e",
         12664 => x"018f0190",
         12665 => x"01910191",
         12666 => x"01930194",
         12667 => x"01f60196",
         12668 => x"01970198",
         12669 => x"0198023d",
         12670 => x"019b019c",
         12671 => x"019d0220",
         12672 => x"019f01a0",
         12673 => x"01a001a2",
         12674 => x"01a201a4",
         12675 => x"01a401a6",
         12676 => x"01a701a7",
         12677 => x"01a901aa",
         12678 => x"01ab01ac",
         12679 => x"01ac01ae",
         12680 => x"01af01af",
         12681 => x"01b101b2",
         12682 => x"01b301b3",
         12683 => x"01b501b5",
         12684 => x"01b701b8",
         12685 => x"01b801ba",
         12686 => x"01bb01bc",
         12687 => x"01bc01be",
         12688 => x"01f701c0",
         12689 => x"01c101c2",
         12690 => x"01c301c4",
         12691 => x"01c501c4",
         12692 => x"01c701c8",
         12693 => x"01c701ca",
         12694 => x"01cb01ca",
         12695 => x"01cd0110",
         12696 => x"01dd0001",
         12697 => x"018e01de",
         12698 => x"011201f3",
         12699 => x"000301f1",
         12700 => x"01f401f4",
         12701 => x"01f80128",
         12702 => x"02220112",
         12703 => x"023a0009",
         12704 => x"2c65023b",
         12705 => x"023b023d",
         12706 => x"2c66023f",
         12707 => x"02400241",
         12708 => x"02410246",
         12709 => x"010a0253",
         12710 => x"00400181",
         12711 => x"01860255",
         12712 => x"0189018a",
         12713 => x"0258018f",
         12714 => x"025a0190",
         12715 => x"025c025d",
         12716 => x"025e025f",
         12717 => x"01930261",
         12718 => x"02620194",
         12719 => x"02640265",
         12720 => x"02660267",
         12721 => x"01970196",
         12722 => x"026a2c62",
         12723 => x"026c026d",
         12724 => x"026e019c",
         12725 => x"02700271",
         12726 => x"019d0273",
         12727 => x"0274019f",
         12728 => x"02760277",
         12729 => x"02780279",
         12730 => x"027a027b",
         12731 => x"027c2c64",
         12732 => x"027e027f",
         12733 => x"01a60281",
         12734 => x"028201a9",
         12735 => x"02840285",
         12736 => x"02860287",
         12737 => x"01ae0244",
         12738 => x"01b101b2",
         12739 => x"0245028d",
         12740 => x"028e028f",
         12741 => x"02900291",
         12742 => x"01b7037b",
         12743 => x"000303fd",
         12744 => x"03fe03ff",
         12745 => x"03ac0004",
         12746 => x"03860388",
         12747 => x"0389038a",
         12748 => x"03b10311",
         12749 => x"03c20002",
         12750 => x"03a303a3",
         12751 => x"03c40308",
         12752 => x"03cc0003",
         12753 => x"038c038e",
         12754 => x"038f03d8",
         12755 => x"011803f2",
         12756 => x"000a03f9",
         12757 => x"03f303f4",
         12758 => x"03f503f6",
         12759 => x"03f703f7",
         12760 => x"03f903fa",
         12761 => x"03fa0430",
         12762 => x"03200450",
         12763 => x"07100460",
         12764 => x"0122048a",
         12765 => x"013604c1",
         12766 => x"010e04cf",
         12767 => x"000104c0",
         12768 => x"04d00144",
         12769 => x"05610426",
         12770 => x"00000000",
         12771 => x"1d7d0001",
         12772 => x"2c631e00",
         12773 => x"01961ea0",
         12774 => x"015a1f00",
         12775 => x"06081f10",
         12776 => x"06061f20",
         12777 => x"06081f30",
         12778 => x"06081f40",
         12779 => x"06061f51",
         12780 => x"00071f59",
         12781 => x"1f521f5b",
         12782 => x"1f541f5d",
         12783 => x"1f561f5f",
         12784 => x"1f600608",
         12785 => x"1f70000e",
         12786 => x"1fba1fbb",
         12787 => x"1fc81fc9",
         12788 => x"1fca1fcb",
         12789 => x"1fda1fdb",
         12790 => x"1ff81ff9",
         12791 => x"1fea1feb",
         12792 => x"1ffa1ffb",
         12793 => x"1f800608",
         12794 => x"1f900608",
         12795 => x"1fa00608",
         12796 => x"1fb00004",
         12797 => x"1fb81fb9",
         12798 => x"1fb21fbc",
         12799 => x"1fcc0001",
         12800 => x"1fc31fd0",
         12801 => x"06021fe0",
         12802 => x"06021fe5",
         12803 => x"00011fec",
         12804 => x"1ff30001",
         12805 => x"1ffc214e",
         12806 => x"00012132",
         12807 => x"21700210",
         12808 => x"21840001",
         12809 => x"218324d0",
         12810 => x"051a2c30",
         12811 => x"042f2c60",
         12812 => x"01022c67",
         12813 => x"01062c75",
         12814 => x"01022c80",
         12815 => x"01642d00",
         12816 => x"0826ff41",
         12817 => x"031a0000",
         12818 => x"00000000",
         12819 => x"000098a0",
         12820 => x"01020100",
         12821 => x"00000000",
         12822 => x"00000000",
         12823 => x"000098a8",
         12824 => x"01040100",
         12825 => x"00000000",
         12826 => x"00000000",
         12827 => x"000098b0",
         12828 => x"01140300",
         12829 => x"00000000",
         12830 => x"00000000",
         12831 => x"000098b8",
         12832 => x"012b0300",
         12833 => x"00000000",
         12834 => x"00000000",
         12835 => x"000098c0",
         12836 => x"01300300",
         12837 => x"00000000",
         12838 => x"00000000",
         12839 => x"000098c8",
         12840 => x"013c0400",
         12841 => x"00000000",
         12842 => x"00000000",
         12843 => x"000098d0",
         12844 => x"013d0400",
         12845 => x"00000000",
         12846 => x"00000000",
         12847 => x"000098d8",
         12848 => x"013f0400",
         12849 => x"00000000",
         12850 => x"00000000",
         12851 => x"000098e0",
         12852 => x"01400400",
         12853 => x"00000000",
         12854 => x"00000000",
         12855 => x"000098e8",
         12856 => x"01410400",
         12857 => x"00000000",
         12858 => x"00000000",
         12859 => x"000098ec",
         12860 => x"01420400",
         12861 => x"00000000",
         12862 => x"00000000",
         12863 => x"000098f0",
         12864 => x"01430400",
         12865 => x"00000000",
         12866 => x"00000000",
         12867 => x"000098f4",
         12868 => x"01500500",
         12869 => x"00000000",
         12870 => x"00000000",
         12871 => x"000098f8",
         12872 => x"01510500",
         12873 => x"00000000",
         12874 => x"00000000",
         12875 => x"000098fc",
         12876 => x"01540500",
         12877 => x"00000000",
         12878 => x"00000000",
         12879 => x"00009900",
         12880 => x"01550500",
         12881 => x"00000000",
         12882 => x"00000000",
         12883 => x"00009904",
         12884 => x"01790700",
         12885 => x"00000000",
         12886 => x"00000000",
         12887 => x"0000990c",
         12888 => x"01780700",
         12889 => x"00000000",
         12890 => x"00000000",
         12891 => x"00009910",
         12892 => x"01820800",
         12893 => x"00000000",
         12894 => x"00000000",
         12895 => x"00009918",
         12896 => x"01830800",
         12897 => x"00000000",
         12898 => x"00000000",
         12899 => x"00009920",
         12900 => x"01850800",
         12901 => x"00000000",
         12902 => x"00000000",
         12903 => x"00009928",
         12904 => x"01870800",
         12905 => x"00000000",
         12906 => x"00000000",
         12907 => x"00009930",
         12908 => x"018c0900",
         12909 => x"00000000",
         12910 => x"00000000",
         12911 => x"00009938",
         12912 => x"018d0900",
         12913 => x"00000000",
         12914 => x"00000000",
         12915 => x"00009940",
         12916 => x"018e0900",
         12917 => x"00000000",
         12918 => x"00000000",
         12919 => x"00009948",
         12920 => x"018f0900",
         12921 => x"00000000",
         12922 => x"00000000",
         12923 => x"00000000",
         12924 => x"00000000",
         12925 => x"00007fff",
         12926 => x"00000000",
         12927 => x"00007fff",
         12928 => x"00010000",
         12929 => x"00007fff",
         12930 => x"00010000",
         12931 => x"00810000",
         12932 => x"01000000",
         12933 => x"017fffff",
         12934 => x"00000000",
         12935 => x"00000000",
         12936 => x"00007800",
         12937 => x"00000000",
         12938 => x"05f5e100",
         12939 => x"05f5e100",
         12940 => x"05f5e100",
         12941 => x"00000000",
         12942 => x"01010101",
         12943 => x"01010101",
         12944 => x"01011001",
         12945 => x"01000000",
         12946 => x"00000000",
         12947 => x"00000000",
         12948 => x"00000000",
         12949 => x"00000000",
         12950 => x"00000000",
         12951 => x"00000000",
         12952 => x"00000000",
         12953 => x"00000000",
         12954 => x"00000000",
         12955 => x"00000000",
         12956 => x"00000000",
         12957 => x"00000000",
         12958 => x"00000000",
         12959 => x"00000000",
         12960 => x"00000000",
         12961 => x"00000000",
         12962 => x"00000000",
         12963 => x"00000000",
         12964 => x"00000000",
         12965 => x"00000000",
         12966 => x"00000000",
         12967 => x"00000000",
         12968 => x"00000000",
         12969 => x"00000000",
         12970 => x"0000a2f4",
         12971 => x"01000000",
         12972 => x"0000a2fc",
         12973 => x"01000000",
         12974 => x"0000a304",
         12975 => x"02000000",
         12976 => x"cce0f2f3",
         12977 => x"cecff6f7",
         12978 => x"f8f9fafb",
         12979 => x"fcfdfeff",
         12980 => x"e1c1c2c3",
         12981 => x"c4c5c6e2",
         12982 => x"e3e4e5e6",
         12983 => x"ebeeeff4",
         12984 => x"00616263",
         12985 => x"64656667",
         12986 => x"68696b6a",
         12987 => x"2f2a2e2d",
         12988 => x"20212223",
         12989 => x"24252627",
         12990 => x"28294f2c",
         12991 => x"512b5749",
         12992 => x"55010203",
         12993 => x"04050607",
         12994 => x"08090a0b",
         12995 => x"0c0d0e0f",
         12996 => x"10111213",
         12997 => x"14151617",
         12998 => x"18191a52",
         12999 => x"5954be3c",
         13000 => x"c7818283",
         13001 => x"84858687",
         13002 => x"88898a8b",
         13003 => x"8c8d8e8f",
         13004 => x"90919293",
         13005 => x"94959697",
         13006 => x"98999abc",
         13007 => x"8040a5c0",
         13008 => x"00e80000",
         13009 => x"00000000",
         13010 => x"00000000",
         13011 => x"00000000",
         13012 => x"00000000",
         13013 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

